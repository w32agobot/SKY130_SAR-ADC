VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO adc_comp_latch
  CLASS BLOCK ;
  FOREIGN adc_comp_latch ;
  ORIGIN 0.000 0.000 ;
  SIZE 30.050 BY 27.980 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 17.700 0.320 18.850 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 9.100 1.720 10.260 ;
    END
  END VSS
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 11.890 4.180 12.030 ;
    END
  END clk
  PIN inp
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 15.410 9.710 15.550 ;
    END
  END inp
  PIN inn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 15.130 7.750 15.270 ;
    END
  END inn
  PIN comp_trig
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 25.310 12.590 30.050 12.730 ;
    END
  END comp_trig
  PIN latch_qn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 26.110 15.540 30.050 15.680 ;
    END
  END latch_qn
  PIN latch_q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 24.790 15.880 30.050 16.020 ;
    END
  END latch_q
  OBS
      LAYER li1 ;
        RECT 2.940 0.000 27.330 27.980 ;
      LAYER met1 ;
        RECT 0.320 19.130 29.920 26.890 ;
        RECT 0.600 17.420 29.920 19.130 ;
        RECT 0.320 16.300 29.920 17.420 ;
        RECT 0.320 15.830 24.510 16.300 ;
        RECT 9.990 15.600 24.510 15.830 ;
        RECT 9.990 15.260 25.830 15.600 ;
        RECT 9.990 15.130 29.920 15.260 ;
        RECT 8.030 14.850 29.920 15.130 ;
        RECT 0.320 13.010 29.920 14.850 ;
        RECT 0.320 12.310 25.030 13.010 ;
        RECT 4.460 11.610 29.920 12.310 ;
        RECT 0.320 10.540 29.920 11.610 ;
        RECT 2.000 8.820 29.920 10.540 ;
        RECT 0.320 1.040 29.920 8.820 ;
      LAYER met2 ;
        RECT 0.230 1.040 29.920 26.890 ;
      LAYER met3 ;
        RECT 0.230 1.040 29.920 26.890 ;
      LAYER met4 ;
        RECT 0.230 0.000 29.920 27.980 ;
  END
END adc_comp_latch
END LIBRARY

