VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_mm_sc_hd_dly5ns
  CLASS CORE ;
  FOREIGN sky130_mm_sc_hd_dly5ns ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.200 BY 2.720 ;
  SITE unithd ;
  PIN in
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.880000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 0.990 0.365 1.320 ;
    END
  END in
  PIN out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.366000 ;
    ANTENNADIFFAREA 0.361800 ;
    PORT
      LAYER li1 ;
        RECT 6.370 1.460 6.540 2.300 ;
        RECT 6.780 1.010 6.950 1.340 ;
        RECT 8.660 0.980 8.890 1.290 ;
        RECT 6.480 0.380 6.650 0.890 ;
      LAYER mcon ;
        RECT 6.370 1.540 6.540 1.820 ;
        RECT 6.780 1.090 6.950 1.260 ;
        RECT 8.690 1.100 8.860 1.270 ;
        RECT 6.480 0.720 6.650 0.890 ;
      LAYER met1 ;
        RECT 6.340 1.240 6.570 1.970 ;
        RECT 6.750 1.240 6.980 1.320 ;
        RECT 8.630 1.240 8.920 1.300 ;
        RECT 6.340 1.100 8.920 1.240 ;
        RECT 6.450 1.030 6.980 1.100 ;
        RECT 8.630 1.070 8.920 1.100 ;
        RECT 6.450 0.660 6.680 1.030 ;
    END
  END out
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.635 9.200 2.805 ;
        RECT 0.570 1.395 0.740 2.235 ;
        RECT 5.410 1.460 5.580 2.635 ;
        RECT 7.120 1.290 7.290 2.635 ;
        RECT 7.120 1.120 7.670 1.290 ;
        RECT 7.500 0.380 7.670 1.120 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 0.570 1.475 0.740 2.155 ;
      LAYER met1 ;
        RECT 0.000 2.480 9.200 2.960 ;
        RECT 0.540 1.415 0.770 2.480 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 7.970 1.180 8.140 2.300 ;
        RECT 7.970 1.010 8.490 1.180 ;
        RECT 0.570 0.455 0.740 0.915 ;
        RECT 5.520 0.085 5.690 0.840 ;
        RECT 8.320 0.085 8.490 1.010 ;
        RECT 0.000 -0.085 9.200 0.085 ;
      LAYER mcon ;
        RECT 0.570 0.535 0.740 0.835 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
      LAYER met1 ;
        RECT 0.540 0.240 0.770 0.910 ;
        RECT 4.840 0.240 5.360 0.770 ;
        RECT 0.000 -0.240 9.200 0.240 ;
      LAYER via ;
        RECT 4.940 0.420 5.260 0.770 ;
      LAYER met2 ;
        RECT 4.840 0.370 5.360 0.910 ;
      LAYER via2 ;
        RECT 4.940 0.630 5.220 0.910 ;
      LAYER met3 ;
        RECT 0.735 0.940 4.710 2.120 ;
        RECT 5.910 0.940 8.570 2.120 ;
        RECT 0.735 0.600 8.570 0.940 ;
    END
  END VGND
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.235 9.390 2.910 ;
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 -0.085 9.195 1.070 ;
    END
  END VNB
  OBS
      LAYER li1 ;
        RECT 4.860 1.180 5.030 2.235 ;
        RECT 5.890 1.460 6.060 2.300 ;
        RECT 7.460 1.460 7.660 2.300 ;
        RECT 8.450 1.460 8.650 2.300 ;
        RECT 5.450 1.180 5.810 1.290 ;
        RECT 4.860 1.010 5.810 1.180 ;
        RECT 4.860 0.365 5.030 1.010 ;
        RECT 6.000 0.380 6.170 0.840 ;
        RECT 7.020 0.380 7.190 0.840 ;
        RECT 7.980 0.380 8.150 0.840 ;
      LAYER mcon ;
        RECT 4.860 1.475 5.030 2.085 ;
        RECT 5.890 1.540 6.060 2.220 ;
        RECT 7.490 1.640 7.660 2.220 ;
        RECT 8.450 1.640 8.620 2.220 ;
        RECT 5.450 1.070 5.730 1.240 ;
        RECT 6.000 0.460 6.170 0.760 ;
        RECT 7.020 0.460 7.190 0.660 ;
        RECT 7.980 0.460 8.150 0.660 ;
      LAYER met1 ;
        RECT 4.830 1.330 5.060 2.195 ;
        RECT 5.860 2.110 8.650 2.280 ;
        RECT 5.860 1.480 6.090 2.110 ;
        RECT 7.460 1.580 7.690 2.110 ;
        RECT 8.420 1.580 8.650 2.110 ;
        RECT 4.830 1.010 5.810 1.330 ;
        RECT 5.970 0.520 6.200 0.820 ;
        RECT 6.990 0.520 7.220 0.720 ;
        RECT 7.950 0.520 8.180 0.720 ;
        RECT 5.970 0.380 8.180 0.520 ;
      LAYER via ;
        RECT 5.450 1.070 5.730 1.330 ;
      LAYER met2 ;
        RECT 5.070 1.050 5.810 1.580 ;
      LAYER via2 ;
        RECT 5.120 1.270 5.400 1.550 ;
      LAYER met3 ;
        RECT 5.070 1.240 5.480 1.960 ;
      LAYER via3 ;
        RECT 5.120 1.270 5.440 1.590 ;
      LAYER met4 ;
        RECT 5.070 1.450 5.480 1.650 ;
        RECT 4.160 1.130 6.470 1.450 ;
  END
END sky130_mm_sc_hd_dly5ns
END LIBRARY

