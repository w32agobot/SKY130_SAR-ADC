magic
tech sky130A
magscale 1 2
timestamp 1661502601
<< nwell >>
rect -10 48 408 452
<< nmos >>
rect 88 -218 118 -118
rect 184 -218 214 -118
rect 280 -218 310 -118
<< pmos >>
rect 88 110 118 310
rect 184 110 214 310
rect 280 110 310 310
<< ndiff >>
rect 26 -130 88 -118
rect 26 -206 38 -130
rect 72 -206 88 -130
rect 26 -218 88 -206
rect 118 -130 184 -118
rect 118 -206 134 -130
rect 168 -206 184 -130
rect 118 -218 184 -206
rect 214 -130 280 -118
rect 214 -206 230 -130
rect 264 -206 280 -130
rect 214 -218 280 -206
rect 310 -130 372 -118
rect 310 -206 326 -130
rect 360 -206 372 -130
rect 310 -218 372 -206
<< pdiff >>
rect 26 298 88 310
rect 26 122 38 298
rect 72 122 88 298
rect 26 110 88 122
rect 118 298 184 310
rect 118 122 134 298
rect 168 122 184 298
rect 118 110 184 122
rect 214 298 280 310
rect 214 122 230 298
rect 264 122 280 298
rect 214 110 280 122
rect 310 298 372 310
rect 310 122 326 298
rect 360 122 372 298
rect 310 110 372 122
<< ndiffc >>
rect 38 -206 72 -130
rect 134 -206 168 -130
rect 230 -206 264 -130
rect 326 -206 360 -130
<< pdiffc >>
rect 38 122 72 298
rect 134 122 168 298
rect 230 122 264 298
rect 326 122 360 298
<< psubdiff >>
rect 26 -326 360 -288
<< nsubdiff >>
rect 26 378 50 416
rect 88 378 126 416
rect 164 378 202 416
rect 240 378 278 416
rect 316 378 372 416
<< nsubdiffcont >>
rect 50 378 88 416
rect 126 378 164 416
rect 202 378 240 416
rect 278 378 316 416
<< poly >>
rect 184 336 310 366
rect 88 310 118 336
rect 184 310 214 336
rect 280 310 310 336
rect 88 84 118 110
rect 76 60 118 84
rect -42 -30 22 -18
rect 76 -30 108 60
rect 184 28 214 110
rect 280 84 310 110
rect -42 -66 108 -30
rect 150 11 214 28
rect 150 -23 160 11
rect 194 -23 214 11
rect 150 -40 214 -23
rect -42 -74 22 -66
rect 76 -68 108 -66
rect 76 -92 118 -68
rect 88 -118 118 -92
rect 184 -118 214 -40
rect 280 -118 310 -92
rect 88 -244 118 -218
rect 184 -244 214 -218
rect 280 -244 310 -218
rect 184 -274 310 -244
<< polycont >>
rect 160 -23 194 11
<< locali >>
rect -42 378 50 416
rect 88 378 126 416
rect 164 378 202 416
rect 240 378 278 416
rect 316 378 408 416
rect 38 298 72 314
rect 38 28 72 122
rect 134 298 168 378
rect 134 106 168 122
rect 230 298 264 314
rect 38 11 196 28
rect 38 -23 160 11
rect 194 -23 196 11
rect 38 -40 196 -23
rect 230 -8 264 122
rect 326 298 360 378
rect 326 106 360 122
rect 38 -130 72 -40
rect 230 -46 408 -8
rect 38 -222 72 -206
rect 134 -130 168 -114
rect 134 -288 168 -206
rect 230 -130 264 -46
rect 230 -222 264 -206
rect 326 -130 360 -114
rect 326 -288 360 -206
rect -42 -326 408 -288
<< comment >>
rect 134 88 168 102
rect 326 90 360 104
rect 134 -110 168 -96
rect 326 -110 360 -96
<< labels >>
rlabel locali -42 -326 -42 -288 7 VSS
port 2 w
rlabel locali -42 378 -42 416 7 VDD
port 1 w
rlabel locali 408 -46 408 -8 3 out
port 4 e
rlabel poly -42 -74 -42 -18 7 in
port 5 w
<< end >>
