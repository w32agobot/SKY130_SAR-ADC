magic
tech sky130A
timestamp 1663849571
<< pwell >>
rect 440 1910 680 2000
rect 1320 1910 1560 2000
rect 115 1890 1910 1910
rect 110 1880 1910 1890
rect 95 1560 1910 1880
rect 0 1320 2000 1560
rect 90 680 1910 1320
rect 0 440 2000 680
rect 90 90 1910 440
rect 440 0 680 90
rect 1320 0 1560 90
<< nmos >>
rect 180 200 1820 1800
<< ndiff >>
rect 180 1860 1820 1870
rect 180 1810 210 1860
rect 270 1810 290 1860
rect 350 1810 370 1860
rect 430 1810 450 1860
rect 510 1810 530 1860
rect 590 1810 610 1860
rect 670 1810 690 1860
rect 750 1810 770 1860
rect 830 1810 850 1860
rect 910 1810 930 1860
rect 990 1810 1010 1860
rect 1070 1810 1090 1860
rect 1150 1810 1170 1860
rect 1230 1810 1250 1860
rect 1310 1810 1330 1860
rect 1390 1810 1410 1860
rect 1470 1810 1490 1860
rect 1550 1810 1570 1860
rect 1630 1810 1650 1860
rect 1710 1810 1730 1860
rect 1785 1810 1820 1860
rect 180 1800 1820 1810
rect 180 190 1820 200
rect 180 140 210 190
rect 270 140 290 190
rect 350 140 370 190
rect 430 140 450 190
rect 510 140 530 190
rect 590 140 610 190
rect 670 140 690 190
rect 750 140 770 190
rect 830 140 850 190
rect 910 140 930 190
rect 990 140 1010 190
rect 1070 140 1090 190
rect 1150 140 1170 190
rect 1230 140 1250 190
rect 1310 140 1330 190
rect 1390 140 1410 190
rect 1470 140 1490 190
rect 1550 140 1570 190
rect 1630 140 1650 190
rect 1710 140 1730 190
rect 1785 140 1820 190
rect 180 130 1820 140
<< ndiffc >>
rect 210 1810 270 1860
rect 290 1810 350 1860
rect 370 1810 430 1860
rect 450 1810 510 1860
rect 530 1810 590 1860
rect 610 1810 670 1860
rect 690 1810 750 1860
rect 770 1810 830 1860
rect 850 1810 910 1860
rect 930 1810 990 1860
rect 1010 1810 1070 1860
rect 1090 1810 1150 1860
rect 1170 1810 1230 1860
rect 1250 1810 1310 1860
rect 1330 1810 1390 1860
rect 1410 1810 1470 1860
rect 1490 1810 1550 1860
rect 1570 1810 1630 1860
rect 1650 1810 1710 1860
rect 1730 1810 1785 1860
rect 210 140 270 190
rect 290 140 350 190
rect 370 140 430 190
rect 450 140 510 190
rect 530 140 590 190
rect 610 140 670 190
rect 690 140 750 190
rect 770 140 830 190
rect 850 140 910 190
rect 930 140 990 190
rect 1010 140 1070 190
rect 1090 140 1150 190
rect 1170 140 1230 190
rect 1250 140 1310 190
rect 1330 140 1390 190
rect 1410 140 1470 190
rect 1490 140 1550 190
rect 1570 140 1630 190
rect 1650 140 1710 190
rect 1730 140 1785 190
<< psubdiff >>
rect 445 1950 675 1960
rect 445 1925 460 1950
rect 660 1925 675 1950
rect 445 1915 675 1925
rect 1325 1950 1555 1960
rect 1325 1925 1340 1950
rect 1540 1925 1555 1950
rect 1325 1915 1555 1925
rect 40 1540 85 1555
rect 40 1340 50 1540
rect 75 1340 85 1540
rect 40 1325 85 1340
rect 40 660 85 675
rect 40 460 50 660
rect 75 460 85 660
rect 40 445 85 460
rect 1915 1540 1960 1555
rect 1915 1340 1925 1540
rect 1950 1340 1960 1540
rect 1915 1325 1960 1340
rect 1915 660 1960 675
rect 1915 460 1925 660
rect 1950 460 1960 660
rect 1915 445 1960 460
rect 445 75 675 85
rect 445 50 460 75
rect 660 50 675 75
rect 445 40 675 50
rect 1325 75 1555 85
rect 1325 50 1340 75
rect 1540 50 1555 75
rect 1325 40 1555 50
<< psubdiffcont >>
rect 460 1925 660 1950
rect 1340 1925 1540 1950
rect 50 1340 75 1540
rect 50 460 75 660
rect 1925 1340 1950 1540
rect 1925 460 1950 660
rect 460 50 660 75
rect 1340 50 1540 75
<< poly >>
rect 160 1575 180 1800
rect 105 1480 180 1575
rect 105 1425 120 1480
rect 160 1425 180 1480
rect 105 1405 180 1425
rect 105 1350 120 1405
rect 160 1350 180 1405
rect 105 1330 180 1350
rect 105 1275 120 1330
rect 160 1275 180 1330
rect 105 1255 180 1275
rect 105 1200 120 1255
rect 160 1200 180 1255
rect 105 1180 180 1200
rect 105 1125 120 1180
rect 160 1125 180 1180
rect 105 1105 180 1125
rect 105 1050 120 1105
rect 160 1050 180 1105
rect 105 1030 180 1050
rect 105 975 120 1030
rect 160 975 180 1030
rect 105 955 180 975
rect 105 900 120 955
rect 160 900 180 955
rect 105 880 180 900
rect 105 825 120 880
rect 160 825 180 880
rect 105 805 180 825
rect 105 750 120 805
rect 160 750 180 805
rect 105 730 180 750
rect 105 675 120 730
rect 160 675 180 730
rect 105 655 180 675
rect 105 600 120 655
rect 160 600 180 655
rect 105 580 180 600
rect 105 525 120 580
rect 160 525 180 580
rect 105 420 180 525
rect 160 200 180 420
rect 1820 1575 1840 1800
rect 1820 1480 1895 1575
rect 1820 1425 1840 1480
rect 1880 1425 1895 1480
rect 1820 1405 1895 1425
rect 1820 1350 1840 1405
rect 1880 1350 1895 1405
rect 1820 1330 1895 1350
rect 1820 1275 1840 1330
rect 1880 1275 1895 1330
rect 1820 1255 1895 1275
rect 1820 1200 1840 1255
rect 1880 1200 1895 1255
rect 1820 1180 1895 1200
rect 1820 1125 1840 1180
rect 1880 1125 1895 1180
rect 1820 1105 1895 1125
rect 1820 1050 1840 1105
rect 1880 1050 1895 1105
rect 1820 1030 1895 1050
rect 1820 975 1840 1030
rect 1880 975 1895 1030
rect 1820 955 1895 975
rect 1820 900 1840 955
rect 1880 900 1895 955
rect 1820 880 1895 900
rect 1820 825 1840 880
rect 1880 825 1895 880
rect 1820 805 1895 825
rect 1820 750 1840 805
rect 1880 750 1895 805
rect 1820 730 1895 750
rect 1820 675 1840 730
rect 1880 675 1895 730
rect 1820 655 1895 675
rect 1820 600 1840 655
rect 1880 600 1895 655
rect 1820 580 1895 600
rect 1820 525 1840 580
rect 1880 525 1895 580
rect 1820 420 1895 525
rect 1820 200 1840 420
<< polycont >>
rect 120 1425 160 1480
rect 120 1350 160 1405
rect 120 1275 160 1330
rect 120 1200 160 1255
rect 120 1125 160 1180
rect 120 1050 160 1105
rect 120 975 160 1030
rect 120 900 160 955
rect 120 825 160 880
rect 120 750 160 805
rect 120 675 160 730
rect 120 600 160 655
rect 120 525 160 580
rect 1840 1425 1880 1480
rect 1840 1350 1880 1405
rect 1840 1275 1880 1330
rect 1840 1200 1880 1255
rect 1840 1125 1880 1180
rect 1840 1050 1880 1105
rect 1840 975 1880 1030
rect 1840 900 1880 955
rect 1840 825 1880 880
rect 1840 750 1880 805
rect 1840 675 1880 730
rect 1840 600 1880 655
rect 1840 525 1880 580
<< locali >>
rect 445 1960 675 2000
rect 1325 1960 1555 2000
rect 40 1950 1960 1960
rect 40 1925 460 1950
rect 660 1925 1340 1950
rect 1540 1925 1960 1950
rect 40 1920 1960 1925
rect 40 1555 80 1920
rect 445 1915 675 1920
rect 1325 1915 1555 1920
rect 180 1810 210 1860
rect 270 1810 290 1860
rect 350 1810 370 1860
rect 430 1810 450 1860
rect 510 1810 530 1860
rect 590 1810 610 1860
rect 670 1810 690 1860
rect 750 1810 770 1860
rect 830 1810 850 1860
rect 910 1810 930 1860
rect 990 1810 1010 1860
rect 1070 1810 1090 1860
rect 1150 1810 1170 1860
rect 1230 1810 1250 1860
rect 1310 1810 1330 1860
rect 1390 1810 1410 1860
rect 1470 1810 1490 1860
rect 1550 1810 1570 1860
rect 1630 1810 1650 1860
rect 1710 1810 1730 1860
rect 1785 1810 1820 1860
rect 180 1800 1820 1810
rect 120 1760 520 1780
rect 120 1700 160 1760
rect 540 1740 575 1800
rect 180 1720 575 1740
rect 120 1680 520 1700
rect 120 1620 160 1680
rect 540 1660 575 1720
rect 180 1640 575 1660
rect 120 1600 520 1620
rect 0 1540 85 1555
rect 0 1340 50 1540
rect 75 1340 85 1540
rect 0 1325 85 1340
rect 120 1540 160 1600
rect 540 1580 575 1640
rect 180 1560 575 1580
rect 120 1520 520 1540
rect 120 1480 160 1520
rect 540 1500 575 1560
rect 180 1480 575 1500
rect 160 1440 520 1460
rect 120 1405 160 1425
rect 540 1420 575 1480
rect 180 1400 575 1420
rect 160 1360 520 1380
rect 120 1330 160 1350
rect 540 1340 575 1400
rect 40 675 80 1325
rect 180 1320 575 1340
rect 160 1280 520 1300
rect 120 1255 160 1275
rect 540 1260 575 1320
rect 180 1240 575 1260
rect 160 1200 520 1220
rect 120 1180 160 1200
rect 540 1180 575 1240
rect 180 1160 575 1180
rect 160 1125 520 1140
rect 120 1120 520 1125
rect 120 1105 160 1120
rect 540 1100 575 1160
rect 180 1080 575 1100
rect 160 1050 520 1060
rect 120 1040 520 1050
rect 540 1040 575 1080
rect 120 1030 160 1040
rect 595 1020 615 1780
rect 635 1040 655 1800
rect 675 1020 695 1780
rect 715 1040 735 1800
rect 755 1020 775 1780
rect 795 1040 815 1800
rect 835 1020 855 1780
rect 875 1040 895 1800
rect 915 1020 935 1780
rect 160 980 935 1020
rect 120 960 160 975
rect 120 955 520 960
rect 160 940 520 955
rect 540 920 575 960
rect 180 900 575 920
rect 120 880 160 900
rect 160 860 520 880
rect 540 840 575 900
rect 120 805 160 825
rect 180 820 575 840
rect 160 780 520 800
rect 540 760 575 820
rect 120 730 160 750
rect 180 740 575 760
rect 160 700 520 720
rect 540 680 575 740
rect 0 660 85 675
rect 0 460 50 660
rect 75 460 85 660
rect 0 445 85 460
rect 120 655 160 675
rect 180 660 575 680
rect 160 620 520 640
rect 540 600 575 660
rect 120 580 160 600
rect 180 580 575 600
rect 160 540 520 560
rect 120 480 160 525
rect 540 520 575 580
rect 180 500 575 520
rect 120 460 520 480
rect 40 80 80 445
rect 120 400 160 460
rect 540 440 575 500
rect 180 420 575 440
rect 120 380 520 400
rect 120 320 160 380
rect 540 360 575 420
rect 180 340 575 360
rect 120 300 520 320
rect 120 240 160 300
rect 540 280 575 340
rect 180 260 575 280
rect 120 220 520 240
rect 540 200 575 260
rect 595 220 615 980
rect 635 200 655 960
rect 675 220 695 980
rect 715 200 735 960
rect 755 220 775 980
rect 795 200 815 960
rect 835 220 855 980
rect 875 200 895 960
rect 915 220 935 980
rect 955 200 1045 1800
rect 1065 1020 1085 1780
rect 1105 1040 1125 1800
rect 1145 1020 1165 1780
rect 1185 1040 1205 1800
rect 1225 1020 1245 1780
rect 1265 1040 1285 1800
rect 1305 1020 1325 1780
rect 1345 1040 1365 1800
rect 1385 1020 1405 1780
rect 1425 1740 1460 1800
rect 1480 1760 1880 1780
rect 1425 1720 1820 1740
rect 1425 1660 1460 1720
rect 1840 1700 1880 1760
rect 1480 1680 1880 1700
rect 1425 1640 1820 1660
rect 1425 1580 1460 1640
rect 1840 1620 1880 1680
rect 1480 1600 1880 1620
rect 1425 1560 1820 1580
rect 1425 1500 1460 1560
rect 1840 1540 1880 1600
rect 1920 1555 1960 1920
rect 1480 1520 1880 1540
rect 1425 1480 1820 1500
rect 1840 1480 1880 1520
rect 1425 1420 1460 1480
rect 1480 1440 1840 1460
rect 1425 1400 1820 1420
rect 1840 1405 1880 1425
rect 1425 1340 1460 1400
rect 1480 1360 1840 1380
rect 1425 1320 1820 1340
rect 1840 1330 1880 1350
rect 1915 1540 2000 1555
rect 1915 1340 1925 1540
rect 1950 1340 2000 1540
rect 1915 1325 2000 1340
rect 1425 1260 1460 1320
rect 1480 1280 1840 1300
rect 1425 1240 1820 1260
rect 1840 1255 1880 1275
rect 1425 1180 1460 1240
rect 1480 1200 1840 1220
rect 1840 1180 1880 1200
rect 1425 1160 1820 1180
rect 1425 1100 1460 1160
rect 1480 1125 1840 1140
rect 1480 1120 1880 1125
rect 1840 1105 1880 1120
rect 1425 1080 1820 1100
rect 1425 1040 1460 1080
rect 1480 1050 1840 1060
rect 1480 1040 1880 1050
rect 1840 1030 1880 1040
rect 1065 980 1840 1020
rect 1065 220 1085 980
rect 1105 200 1125 960
rect 1145 220 1165 980
rect 1185 200 1205 960
rect 1225 220 1245 980
rect 1265 200 1285 960
rect 1305 220 1325 980
rect 1345 200 1365 960
rect 1385 220 1405 980
rect 1840 960 1880 975
rect 1425 920 1460 960
rect 1480 955 1880 960
rect 1480 940 1840 955
rect 1425 900 1820 920
rect 1425 840 1460 900
rect 1840 880 1880 900
rect 1480 860 1840 880
rect 1425 820 1820 840
rect 1425 760 1460 820
rect 1840 805 1880 825
rect 1480 780 1840 800
rect 1425 740 1820 760
rect 1425 680 1460 740
rect 1840 730 1880 750
rect 1480 700 1840 720
rect 1425 660 1820 680
rect 1920 675 1960 1325
rect 1425 600 1460 660
rect 1840 655 1880 675
rect 1480 620 1840 640
rect 1425 580 1820 600
rect 1840 580 1880 600
rect 1425 520 1460 580
rect 1480 540 1840 560
rect 1425 500 1820 520
rect 1425 440 1460 500
rect 1840 480 1880 525
rect 1480 460 1880 480
rect 1425 420 1820 440
rect 1425 360 1460 420
rect 1840 400 1880 460
rect 1915 660 2000 675
rect 1915 460 1925 660
rect 1950 460 2000 660
rect 1915 445 2000 460
rect 1480 380 1880 400
rect 1425 340 1820 360
rect 1425 280 1460 340
rect 1840 320 1880 380
rect 1480 300 1880 320
rect 1425 260 1820 280
rect 1425 200 1460 260
rect 1840 240 1880 300
rect 1480 220 1880 240
rect 180 190 1820 200
rect 180 140 210 190
rect 270 140 290 190
rect 350 140 370 190
rect 430 140 450 190
rect 510 140 530 190
rect 590 140 610 190
rect 670 140 690 190
rect 750 140 770 190
rect 830 140 850 190
rect 910 140 930 190
rect 990 140 1010 190
rect 1070 140 1090 190
rect 1150 140 1170 190
rect 1230 140 1250 190
rect 1310 140 1330 190
rect 1390 140 1410 190
rect 1470 140 1490 190
rect 1550 140 1570 190
rect 1630 140 1650 190
rect 1710 140 1730 190
rect 1785 140 1820 190
rect 445 80 675 85
rect 1325 80 1555 85
rect 1920 80 1960 445
rect 40 75 1960 80
rect 40 50 460 75
rect 660 50 1340 75
rect 1540 50 1960 75
rect 40 40 1960 50
rect 445 0 675 40
rect 1325 0 1555 40
<< viali >>
rect 210 1810 270 1860
rect 290 1810 350 1860
rect 370 1810 430 1860
rect 450 1810 510 1860
rect 530 1810 590 1860
rect 1410 1810 1470 1860
rect 1490 1810 1550 1860
rect 1570 1810 1630 1860
rect 1650 1810 1710 1860
rect 1730 1810 1785 1860
rect 125 1430 155 1475
rect 125 1355 155 1400
rect 125 1280 155 1325
rect 125 1205 155 1250
rect 125 1130 155 1175
rect 125 1055 155 1100
rect 125 980 155 1025
rect 125 905 155 950
rect 125 830 155 875
rect 125 755 155 800
rect 125 680 155 725
rect 125 605 155 650
rect 125 530 155 575
rect 1845 1430 1875 1475
rect 1845 1355 1875 1400
rect 1845 1280 1875 1325
rect 1845 1205 1875 1250
rect 1845 1130 1875 1175
rect 1845 1055 1875 1100
rect 1845 980 1875 1025
rect 1845 905 1875 950
rect 1845 830 1875 875
rect 1845 755 1875 800
rect 1845 680 1875 725
rect 1845 605 1875 650
rect 1845 530 1875 575
rect 210 140 270 190
rect 290 140 350 190
rect 370 140 430 190
rect 450 140 510 190
rect 530 140 590 190
rect 1410 140 1470 190
rect 1490 140 1550 190
rect 1570 140 1630 190
rect 1650 140 1710 190
rect 1730 140 1785 190
<< metal1 >>
rect 0 1990 440 2000
rect 0 1890 10 1990
rect 110 1890 170 1990
rect 270 1890 330 1990
rect 430 1985 440 1990
rect 680 1990 1320 2000
rect 430 1895 600 1985
rect 430 1890 440 1895
rect 0 1880 440 1890
rect 0 1830 120 1880
rect 455 1865 600 1895
rect 680 1890 690 1990
rect 790 1890 805 1990
rect 905 1890 920 1990
rect 1080 1890 1095 1990
rect 1195 1890 1210 1990
rect 1310 1890 1320 1990
rect 1560 1990 2000 2000
rect 1560 1980 1570 1990
rect 680 1880 1320 1890
rect 1400 1890 1570 1980
rect 1670 1890 1730 1990
rect 1830 1890 1890 1990
rect 1990 1890 2000 1990
rect 0 1730 10 1830
rect 110 1730 120 1830
rect 0 1670 120 1730
rect 0 1570 10 1670
rect 110 1570 120 1670
rect 0 1560 120 1570
rect 180 1860 600 1865
rect 180 1810 210 1860
rect 270 1810 290 1860
rect 350 1810 370 1860
rect 430 1810 450 1860
rect 510 1810 530 1860
rect 590 1845 600 1860
rect 590 1830 935 1845
rect 590 1810 600 1830
rect 950 1815 1050 1880
rect 1400 1865 1545 1890
rect 1560 1880 2000 1890
rect 1400 1860 1820 1865
rect 1400 1845 1410 1860
rect 1070 1830 1410 1845
rect 180 1800 600 1810
rect 615 1800 1385 1815
rect 1400 1810 1410 1830
rect 1470 1810 1490 1860
rect 1550 1810 1570 1860
rect 1630 1810 1650 1860
rect 1710 1810 1730 1860
rect 1785 1810 1820 1860
rect 1400 1800 1820 1810
rect 180 1515 195 1800
rect 120 1475 195 1500
rect 120 1430 125 1475
rect 155 1430 195 1475
rect 120 1400 195 1430
rect 120 1355 125 1400
rect 155 1355 195 1400
rect 120 1325 195 1355
rect 120 1320 125 1325
rect 0 1310 125 1320
rect 0 1240 10 1310
rect 80 1280 125 1310
rect 155 1280 195 1325
rect 80 1250 195 1280
rect 80 1240 125 1250
rect 0 1225 125 1240
rect 0 1155 10 1225
rect 80 1205 125 1225
rect 155 1205 195 1250
rect 80 1175 195 1205
rect 80 1155 125 1175
rect 0 1140 125 1155
rect 0 1070 10 1140
rect 80 1130 125 1140
rect 155 1130 195 1175
rect 80 1100 195 1130
rect 80 1070 125 1100
rect 0 1055 125 1070
rect 155 1055 195 1100
rect 0 1045 195 1055
rect 0 955 15 1045
rect 80 1030 195 1045
rect 210 1030 225 1785
rect 240 1045 255 1800
rect 270 1030 285 1785
rect 300 1045 315 1800
rect 330 1030 345 1785
rect 360 1045 375 1800
rect 390 1030 405 1785
rect 420 1045 435 1800
rect 450 1030 465 1785
rect 480 1045 495 1800
rect 540 1785 600 1800
rect 510 1030 525 1785
rect 540 1770 935 1785
rect 540 1725 600 1770
rect 950 1755 1050 1800
rect 1400 1785 1460 1800
rect 1065 1770 1460 1785
rect 615 1740 1385 1755
rect 540 1710 935 1725
rect 540 1665 600 1710
rect 950 1695 1050 1740
rect 1400 1725 1460 1770
rect 1065 1710 1460 1725
rect 615 1680 1385 1695
rect 540 1650 935 1665
rect 540 1605 600 1650
rect 950 1635 1050 1680
rect 1400 1665 1460 1710
rect 1065 1650 1460 1665
rect 615 1620 1385 1635
rect 540 1590 935 1605
rect 540 1545 600 1590
rect 950 1575 1050 1620
rect 1400 1605 1460 1650
rect 1065 1590 1460 1605
rect 615 1560 1385 1575
rect 540 1530 935 1545
rect 540 1485 600 1530
rect 950 1515 1050 1560
rect 1400 1545 1460 1590
rect 1065 1530 1460 1545
rect 615 1500 1385 1515
rect 540 1470 935 1485
rect 540 1425 600 1470
rect 950 1455 1050 1500
rect 1400 1485 1460 1530
rect 1065 1470 1460 1485
rect 615 1440 1385 1455
rect 540 1410 935 1425
rect 540 1365 600 1410
rect 950 1395 1050 1440
rect 1400 1425 1460 1470
rect 1065 1410 1460 1425
rect 615 1380 1385 1395
rect 540 1350 935 1365
rect 540 1305 600 1350
rect 950 1335 1050 1380
rect 1400 1365 1460 1410
rect 1065 1350 1460 1365
rect 615 1320 1385 1335
rect 540 1290 935 1305
rect 540 1245 600 1290
rect 950 1275 1050 1320
rect 1400 1305 1460 1350
rect 1065 1290 1460 1305
rect 615 1260 1385 1275
rect 540 1230 935 1245
rect 540 1185 600 1230
rect 950 1215 1050 1260
rect 1400 1245 1460 1290
rect 1065 1230 1460 1245
rect 615 1200 1385 1215
rect 540 1170 935 1185
rect 540 1125 600 1170
rect 950 1155 1050 1200
rect 1400 1185 1460 1230
rect 1065 1170 1460 1185
rect 615 1140 1385 1155
rect 540 1110 935 1125
rect 540 1065 600 1110
rect 950 1095 1050 1140
rect 1400 1125 1460 1170
rect 1065 1110 1460 1125
rect 615 1080 1385 1095
rect 540 1045 935 1065
rect 950 1030 1050 1080
rect 1400 1065 1460 1110
rect 1065 1045 1460 1065
rect 1475 1030 1490 1785
rect 1505 1045 1520 1800
rect 1535 1030 1550 1785
rect 1565 1045 1580 1800
rect 1595 1030 1610 1785
rect 1625 1045 1640 1800
rect 1655 1030 1670 1785
rect 1685 1045 1700 1800
rect 1715 1030 1730 1785
rect 1745 1045 1760 1800
rect 1775 1030 1790 1785
rect 1805 1515 1820 1800
rect 1880 1830 2000 1880
rect 1880 1730 1890 1830
rect 1990 1730 2000 1830
rect 1880 1670 2000 1730
rect 1880 1570 1890 1670
rect 1990 1570 2000 1670
rect 1880 1560 2000 1570
rect 1805 1475 1880 1500
rect 1805 1430 1845 1475
rect 1875 1430 1880 1475
rect 1805 1400 1880 1430
rect 1805 1355 1845 1400
rect 1875 1355 1880 1400
rect 1805 1325 1880 1355
rect 1805 1280 1845 1325
rect 1875 1320 1880 1325
rect 1875 1310 2000 1320
rect 1875 1280 1920 1310
rect 1805 1250 1920 1280
rect 1805 1205 1845 1250
rect 1875 1240 1920 1250
rect 1990 1240 2000 1310
rect 1875 1225 2000 1240
rect 1875 1205 1920 1225
rect 1805 1175 1920 1205
rect 1805 1130 1845 1175
rect 1875 1155 1920 1175
rect 1990 1155 2000 1225
rect 1875 1140 2000 1155
rect 1875 1130 1920 1140
rect 1805 1100 1920 1130
rect 1805 1055 1845 1100
rect 1875 1070 1920 1100
rect 1990 1070 2000 1140
rect 1875 1055 2000 1070
rect 1805 1045 2000 1055
rect 1805 1030 1920 1045
rect 80 1025 1920 1030
rect 80 980 125 1025
rect 155 980 1845 1025
rect 1875 980 1920 1025
rect 80 970 1920 980
rect 80 955 195 970
rect 0 950 195 955
rect 0 930 125 950
rect 0 860 10 930
rect 80 905 125 930
rect 155 905 195 950
rect 80 875 195 905
rect 80 860 125 875
rect 0 845 125 860
rect 0 775 10 845
rect 80 830 125 845
rect 155 830 195 875
rect 80 800 195 830
rect 80 775 125 800
rect 0 760 125 775
rect 0 690 10 760
rect 80 755 125 760
rect 155 755 195 800
rect 80 725 195 755
rect 80 690 125 725
rect 0 680 125 690
rect 155 680 195 725
rect 120 650 195 680
rect 120 605 125 650
rect 155 605 195 650
rect 120 575 195 605
rect 120 530 125 575
rect 155 530 195 575
rect 120 505 195 530
rect 0 430 120 440
rect 0 330 10 430
rect 110 330 120 430
rect 0 270 120 330
rect 0 170 10 270
rect 110 170 120 270
rect 0 120 120 170
rect 180 200 195 490
rect 210 215 225 970
rect 240 200 255 955
rect 270 215 285 970
rect 300 200 315 955
rect 330 215 345 970
rect 360 200 375 955
rect 390 215 405 970
rect 420 200 435 955
rect 450 215 465 970
rect 480 200 495 955
rect 510 215 525 970
rect 540 935 935 955
rect 540 890 600 935
rect 950 920 1050 970
rect 1065 935 1460 955
rect 615 905 1385 920
rect 540 875 935 890
rect 540 830 600 875
rect 950 860 1050 905
rect 1400 890 1460 935
rect 1065 875 1460 890
rect 615 845 1385 860
rect 540 815 935 830
rect 540 770 600 815
rect 950 800 1050 845
rect 1400 830 1460 875
rect 1065 815 1460 830
rect 615 785 1385 800
rect 540 755 935 770
rect 540 710 600 755
rect 950 740 1050 785
rect 1400 770 1460 815
rect 1065 755 1460 770
rect 615 725 1385 740
rect 540 695 935 710
rect 540 650 600 695
rect 950 680 1050 725
rect 1400 710 1460 755
rect 1065 695 1460 710
rect 615 665 1385 680
rect 540 635 935 650
rect 540 590 600 635
rect 950 620 1050 665
rect 1400 650 1460 695
rect 1065 635 1460 650
rect 615 605 1385 620
rect 540 575 935 590
rect 540 530 600 575
rect 950 560 1050 605
rect 1400 590 1460 635
rect 1065 575 1460 590
rect 615 545 1385 560
rect 540 515 935 530
rect 540 470 600 515
rect 950 500 1050 545
rect 1400 530 1460 575
rect 1065 515 1460 530
rect 615 485 1385 500
rect 540 455 935 470
rect 540 410 600 455
rect 950 440 1050 485
rect 1400 470 1460 515
rect 1065 455 1460 470
rect 615 425 1385 440
rect 540 395 935 410
rect 540 350 600 395
rect 950 380 1050 425
rect 1400 410 1460 455
rect 1065 395 1460 410
rect 615 365 1385 380
rect 540 335 935 350
rect 540 290 600 335
rect 950 320 1050 365
rect 1400 350 1460 395
rect 1065 335 1460 350
rect 615 305 1385 320
rect 540 275 935 290
rect 540 230 600 275
rect 950 260 1050 305
rect 1400 290 1460 335
rect 1065 275 1460 290
rect 615 245 1385 260
rect 540 215 935 230
rect 540 200 600 215
rect 950 200 1050 245
rect 1400 230 1460 275
rect 1065 215 1460 230
rect 1475 215 1490 970
rect 1400 200 1460 215
rect 1505 200 1520 955
rect 1535 215 1550 970
rect 1565 200 1580 955
rect 1595 215 1610 970
rect 1625 200 1640 955
rect 1655 215 1670 970
rect 1685 200 1700 955
rect 1715 215 1730 970
rect 1745 200 1760 955
rect 1775 215 1790 970
rect 1805 955 1920 970
rect 1985 955 2000 1045
rect 1805 950 2000 955
rect 1805 905 1845 950
rect 1875 930 2000 950
rect 1875 905 1920 930
rect 1805 875 1920 905
rect 1805 830 1845 875
rect 1875 860 1920 875
rect 1990 860 2000 930
rect 1875 845 2000 860
rect 1875 830 1920 845
rect 1805 800 1920 830
rect 1805 755 1845 800
rect 1875 775 1920 800
rect 1990 775 2000 845
rect 1875 760 2000 775
rect 1875 755 1920 760
rect 1805 725 1920 755
rect 1805 680 1845 725
rect 1875 690 1920 725
rect 1990 690 2000 760
rect 1875 680 2000 690
rect 1805 650 1880 680
rect 1805 605 1845 650
rect 1875 605 1880 650
rect 1805 575 1880 605
rect 1805 530 1845 575
rect 1875 530 1880 575
rect 1805 505 1880 530
rect 1805 200 1820 490
rect 180 190 600 200
rect 180 140 210 190
rect 270 140 290 190
rect 350 140 370 190
rect 430 140 450 190
rect 510 140 530 190
rect 590 170 600 190
rect 615 185 1385 200
rect 1400 190 1820 200
rect 590 155 935 170
rect 590 140 600 155
rect 180 135 600 140
rect 0 110 440 120
rect 0 10 10 110
rect 110 10 170 110
rect 270 10 330 110
rect 430 105 440 110
rect 455 105 600 135
rect 950 120 1050 185
rect 1400 170 1410 190
rect 1065 155 1410 170
rect 1400 140 1410 155
rect 1470 140 1490 190
rect 1550 140 1570 190
rect 1630 140 1650 190
rect 1710 140 1730 190
rect 1785 140 1820 190
rect 1400 135 1820 140
rect 1880 430 2000 440
rect 1880 330 1890 430
rect 1990 330 2000 430
rect 1880 270 2000 330
rect 1880 170 1890 270
rect 1990 170 2000 270
rect 430 15 600 105
rect 680 110 1320 120
rect 430 10 440 15
rect 0 0 440 10
rect 680 10 690 110
rect 790 10 800 110
rect 900 10 915 110
rect 1075 10 1095 110
rect 1195 10 1210 110
rect 1310 10 1320 110
rect 1400 105 1545 135
rect 1880 120 2000 170
rect 1560 110 2000 120
rect 1560 105 1570 110
rect 1400 15 1570 105
rect 680 0 1320 10
rect 1560 10 1570 15
rect 1670 10 1730 110
rect 1830 10 1890 110
rect 1990 10 2000 110
rect 1560 0 2000 10
<< via1 >>
rect 10 1890 110 1990
rect 170 1890 270 1990
rect 330 1890 430 1990
rect 690 1890 790 1990
rect 805 1890 905 1990
rect 920 1890 1080 1990
rect 1095 1890 1195 1990
rect 1210 1890 1310 1990
rect 1570 1890 1670 1990
rect 1730 1890 1830 1990
rect 1890 1890 1990 1990
rect 10 1730 110 1830
rect 10 1570 110 1670
rect 10 1240 80 1310
rect 10 1155 80 1225
rect 10 1070 80 1140
rect 1890 1730 1990 1830
rect 1890 1570 1990 1670
rect 1920 1240 1990 1310
rect 1920 1155 1990 1225
rect 1920 1070 1990 1140
rect 10 860 80 930
rect 10 775 80 845
rect 10 690 80 760
rect 10 330 110 430
rect 10 170 110 270
rect 1920 860 1990 930
rect 1920 775 1990 845
rect 1920 690 1990 760
rect 10 10 110 110
rect 170 10 270 110
rect 330 10 430 110
rect 1890 330 1990 430
rect 1890 170 1990 270
rect 690 10 790 110
rect 800 10 900 110
rect 915 10 1075 110
rect 1095 10 1195 110
rect 1210 10 1310 110
rect 1570 10 1670 110
rect 1730 10 1830 110
rect 1890 10 1990 110
<< metal2 >>
rect 0 1990 440 2000
rect 0 1890 10 1990
rect 110 1890 170 1990
rect 270 1890 330 1990
rect 430 1890 440 1990
rect 680 1990 1320 2000
rect 680 1910 690 1990
rect 0 1880 440 1890
rect 490 1890 690 1910
rect 790 1890 805 1990
rect 905 1890 920 1990
rect 1080 1890 1095 1990
rect 1195 1890 1210 1990
rect 1310 1910 1320 1990
rect 1560 1990 2000 2000
rect 1310 1890 1510 1910
rect 0 1830 121 1880
rect 490 1860 1510 1890
rect 1560 1890 1570 1990
rect 1670 1890 1730 1990
rect 1830 1890 1890 1990
rect 1990 1890 2000 1990
rect 1560 1880 2000 1890
rect 0 1730 10 1830
rect 110 1785 121 1830
rect 180 1855 1820 1860
rect 180 1800 560 1855
rect 110 1770 515 1785
rect 110 1730 160 1770
rect 530 1755 560 1800
rect 175 1740 560 1755
rect 0 1725 160 1730
rect 0 1710 515 1725
rect 0 1670 160 1710
rect 530 1695 560 1740
rect 175 1680 560 1695
rect 0 1570 10 1670
rect 110 1665 160 1670
rect 110 1650 515 1665
rect 110 1605 160 1650
rect 530 1635 560 1680
rect 175 1620 560 1635
rect 110 1590 515 1605
rect 110 1570 160 1590
rect 530 1575 560 1620
rect 0 1560 160 1570
rect 175 1560 560 1575
rect 120 1545 160 1560
rect 120 1530 515 1545
rect 120 1485 160 1530
rect 530 1515 560 1560
rect 175 1500 560 1515
rect 120 1470 515 1485
rect 120 1425 160 1470
rect 530 1455 560 1500
rect 175 1440 560 1455
rect 120 1410 515 1425
rect 120 1365 160 1410
rect 530 1395 560 1440
rect 175 1380 560 1395
rect 120 1350 515 1365
rect 0 1310 90 1320
rect 0 1240 10 1310
rect 80 1240 90 1310
rect 0 1225 90 1240
rect 0 1155 10 1225
rect 80 1155 90 1225
rect 0 1140 90 1155
rect 0 1070 10 1140
rect 80 1070 90 1140
rect 0 930 90 1070
rect 0 860 10 930
rect 80 860 90 930
rect 0 845 90 860
rect 0 775 10 845
rect 80 775 90 845
rect 0 760 90 775
rect 0 690 10 760
rect 80 690 90 760
rect 0 680 90 690
rect 120 1305 160 1350
rect 530 1335 560 1380
rect 175 1320 560 1335
rect 120 1290 515 1305
rect 120 1245 160 1290
rect 530 1275 560 1320
rect 175 1260 560 1275
rect 120 1230 515 1245
rect 120 1185 160 1230
rect 530 1215 560 1260
rect 175 1200 560 1215
rect 120 1170 515 1185
rect 120 1125 160 1170
rect 530 1155 560 1200
rect 175 1140 560 1155
rect 120 1110 515 1125
rect 120 1065 160 1110
rect 530 1095 560 1140
rect 175 1080 560 1095
rect 120 1050 515 1065
rect 120 1020 160 1050
rect 530 1035 560 1080
rect 575 1020 590 1840
rect 605 1035 620 1855
rect 635 1020 650 1840
rect 665 1035 680 1855
rect 695 1020 710 1840
rect 725 1035 740 1855
rect 755 1020 770 1840
rect 785 1035 800 1855
rect 815 1020 830 1840
rect 845 1035 860 1855
rect 875 1020 890 1840
rect 905 1035 920 1855
rect 935 1020 950 1840
rect 120 980 950 1020
rect 120 950 160 980
rect 120 935 515 950
rect 120 890 160 935
rect 530 920 560 965
rect 175 905 560 920
rect 120 875 515 890
rect 120 830 160 875
rect 530 860 560 905
rect 175 845 560 860
rect 120 815 515 830
rect 120 770 160 815
rect 530 800 560 845
rect 175 785 560 800
rect 120 755 515 770
rect 120 710 160 755
rect 530 740 560 785
rect 175 725 560 740
rect 120 695 515 710
rect 120 650 160 695
rect 530 680 560 725
rect 175 665 560 680
rect 120 635 515 650
rect 120 590 160 635
rect 530 620 560 665
rect 175 605 560 620
rect 120 575 515 590
rect 120 530 160 575
rect 530 560 560 605
rect 175 545 560 560
rect 120 515 515 530
rect 120 470 160 515
rect 530 500 560 545
rect 175 485 560 500
rect 120 455 515 470
rect 120 440 160 455
rect 530 440 560 485
rect 0 430 160 440
rect 0 330 10 430
rect 110 410 160 430
rect 175 425 560 440
rect 110 395 515 410
rect 110 350 160 395
rect 530 380 560 425
rect 175 365 560 380
rect 110 335 515 350
rect 110 330 160 335
rect 0 290 160 330
rect 530 320 560 365
rect 175 305 560 320
rect 0 275 515 290
rect 0 270 160 275
rect 0 170 10 270
rect 110 230 160 270
rect 530 260 560 305
rect 175 245 560 260
rect 110 215 515 230
rect 110 170 120 215
rect 530 200 560 245
rect 0 120 120 170
rect 180 145 560 200
rect 575 160 590 980
rect 605 145 620 965
rect 635 160 650 980
rect 665 145 680 965
rect 695 160 710 980
rect 725 145 740 965
rect 755 160 770 980
rect 785 145 800 965
rect 815 160 830 980
rect 845 145 860 965
rect 875 160 890 980
rect 905 145 920 965
rect 935 160 950 980
rect 965 145 1035 1855
rect 1050 1020 1065 1840
rect 1080 1035 1095 1855
rect 1110 1020 1125 1840
rect 1140 1035 1155 1855
rect 1170 1020 1185 1840
rect 1200 1035 1215 1855
rect 1230 1020 1245 1840
rect 1260 1035 1275 1855
rect 1290 1020 1305 1840
rect 1320 1035 1335 1855
rect 1350 1020 1365 1840
rect 1380 1035 1395 1855
rect 1410 1020 1425 1840
rect 1440 1800 1820 1855
rect 1880 1830 2000 1880
rect 1440 1755 1470 1800
rect 1880 1785 1890 1830
rect 1485 1770 1890 1785
rect 1440 1740 1825 1755
rect 1440 1695 1470 1740
rect 1840 1730 1890 1770
rect 1990 1730 2000 1830
rect 1840 1725 2000 1730
rect 1485 1710 2000 1725
rect 1440 1680 1825 1695
rect 1440 1635 1470 1680
rect 1840 1670 2000 1710
rect 1840 1665 1890 1670
rect 1485 1650 1890 1665
rect 1440 1620 1825 1635
rect 1440 1575 1470 1620
rect 1840 1605 1890 1650
rect 1485 1590 1890 1605
rect 1440 1560 1825 1575
rect 1840 1570 1890 1590
rect 1990 1570 2000 1670
rect 1840 1560 2000 1570
rect 1440 1515 1470 1560
rect 1840 1545 1880 1560
rect 1485 1530 1880 1545
rect 1440 1500 1825 1515
rect 1440 1455 1470 1500
rect 1840 1485 1880 1530
rect 1485 1470 1880 1485
rect 1440 1440 1825 1455
rect 1440 1395 1470 1440
rect 1840 1425 1880 1470
rect 1485 1410 1880 1425
rect 1440 1380 1825 1395
rect 1440 1335 1470 1380
rect 1840 1365 1880 1410
rect 1485 1350 1880 1365
rect 1440 1320 1825 1335
rect 1440 1275 1470 1320
rect 1840 1305 1880 1350
rect 1485 1290 1880 1305
rect 1440 1260 1825 1275
rect 1440 1215 1470 1260
rect 1840 1245 1880 1290
rect 1485 1230 1880 1245
rect 1440 1200 1825 1215
rect 1440 1155 1470 1200
rect 1840 1185 1880 1230
rect 1485 1170 1880 1185
rect 1440 1140 1825 1155
rect 1440 1095 1470 1140
rect 1840 1125 1880 1170
rect 1485 1110 1880 1125
rect 1440 1080 1825 1095
rect 1440 1035 1470 1080
rect 1840 1065 1880 1110
rect 1485 1050 1880 1065
rect 1840 1020 1880 1050
rect 1050 980 1880 1020
rect 1050 160 1065 980
rect 1080 145 1095 965
rect 1110 160 1125 980
rect 1140 145 1155 965
rect 1170 160 1185 980
rect 1200 145 1215 965
rect 1230 160 1245 980
rect 1260 145 1275 965
rect 1290 160 1305 980
rect 1320 145 1335 965
rect 1350 160 1365 980
rect 1380 145 1395 965
rect 1410 160 1425 980
rect 1440 920 1470 965
rect 1840 950 1880 980
rect 1485 935 1880 950
rect 1440 905 1825 920
rect 1440 860 1470 905
rect 1840 890 1880 935
rect 1485 875 1880 890
rect 1440 845 1825 860
rect 1440 800 1470 845
rect 1840 830 1880 875
rect 1485 815 1880 830
rect 1440 785 1825 800
rect 1440 740 1470 785
rect 1840 770 1880 815
rect 1485 755 1880 770
rect 1440 725 1825 740
rect 1440 680 1470 725
rect 1840 710 1880 755
rect 1485 695 1880 710
rect 1440 665 1825 680
rect 1440 620 1470 665
rect 1840 650 1880 695
rect 1910 1310 2000 1320
rect 1910 1240 1920 1310
rect 1990 1240 2000 1310
rect 1910 1225 2000 1240
rect 1910 1155 1920 1225
rect 1990 1155 2000 1225
rect 1910 1140 2000 1155
rect 1910 1070 1920 1140
rect 1990 1070 2000 1140
rect 1910 930 2000 1070
rect 1910 860 1920 930
rect 1990 860 2000 930
rect 1910 845 2000 860
rect 1910 775 1920 845
rect 1990 775 2000 845
rect 1910 760 2000 775
rect 1910 690 1920 760
rect 1990 690 2000 760
rect 1910 680 2000 690
rect 1485 635 1880 650
rect 1440 605 1825 620
rect 1440 560 1470 605
rect 1840 590 1880 635
rect 1485 575 1880 590
rect 1440 545 1825 560
rect 1440 500 1470 545
rect 1840 530 1880 575
rect 1485 515 1880 530
rect 1440 485 1825 500
rect 1440 440 1470 485
rect 1840 470 1880 515
rect 1485 455 1880 470
rect 1840 440 1880 455
rect 1440 425 1825 440
rect 1840 430 2000 440
rect 1440 380 1470 425
rect 1840 410 1890 430
rect 1485 395 1890 410
rect 1440 365 1825 380
rect 1440 320 1470 365
rect 1840 350 1890 395
rect 1485 335 1890 350
rect 1840 330 1890 335
rect 1990 330 2000 430
rect 1440 305 1825 320
rect 1440 260 1470 305
rect 1840 290 2000 330
rect 1485 275 2000 290
rect 1840 270 2000 275
rect 1440 245 1825 260
rect 1440 200 1470 245
rect 1840 230 1890 270
rect 1485 215 1890 230
rect 1440 145 1820 200
rect 180 140 1820 145
rect 1880 170 1890 215
rect 1990 170 2000 270
rect 0 110 440 120
rect 0 10 10 110
rect 110 10 170 110
rect 270 10 330 110
rect 430 10 440 110
rect 490 110 1510 140
rect 1880 120 2000 170
rect 490 90 690 110
rect 0 0 440 10
rect 680 10 690 90
rect 790 10 800 110
rect 900 10 915 110
rect 1075 10 1095 110
rect 1195 10 1210 110
rect 1310 90 1510 110
rect 1560 110 2000 120
rect 1310 10 1320 90
rect 680 0 1320 10
rect 1560 10 1570 110
rect 1670 10 1730 110
rect 1830 10 1890 110
rect 1990 10 2000 110
rect 1560 0 2000 10
<< metal3 >>
rect 0 1990 440 2000
rect 0 1905 10 1990
rect 95 1905 105 1990
rect 190 1905 250 1990
rect 335 1905 345 1990
rect 430 1905 440 1990
rect 680 1990 1320 2000
rect 680 1925 690 1990
rect 755 1925 770 1990
rect 835 1925 850 1990
rect 915 1925 1085 1990
rect 1150 1925 1165 1990
rect 1230 1925 1245 1990
rect 1310 1925 1320 1990
rect 680 1915 1320 1925
rect 1560 1990 2000 2000
rect 0 1895 440 1905
rect 0 1810 10 1895
rect 95 1875 440 1895
rect 1560 1905 1570 1990
rect 1655 1905 1665 1990
rect 1750 1905 1810 1990
rect 1895 1905 1905 1990
rect 1990 1905 2000 1990
rect 1560 1895 2000 1905
rect 1560 1875 1905 1895
rect 95 1810 1905 1875
rect 1990 1810 2000 1895
rect 0 1750 2000 1810
rect 0 1665 10 1750
rect 95 1665 1905 1750
rect 1990 1665 2000 1750
rect 0 1655 2000 1665
rect 0 1570 10 1655
rect 95 1570 1905 1655
rect 1990 1570 2000 1655
rect 0 1560 2000 1570
rect 0 1310 85 1320
rect 0 1245 10 1310
rect 75 1245 85 1310
rect 0 1230 85 1245
rect 0 1165 10 1230
rect 75 1165 85 1230
rect 0 1150 85 1165
rect 0 1085 10 1150
rect 75 1085 85 1150
rect 0 915 85 1085
rect 0 850 10 915
rect 75 850 85 915
rect 0 835 85 850
rect 0 770 10 835
rect 75 770 85 835
rect 0 755 85 770
rect 0 690 10 755
rect 75 690 85 755
rect 0 680 85 690
rect 125 440 1875 1560
rect 1915 1310 2000 1320
rect 1915 1245 1925 1310
rect 1990 1245 2000 1310
rect 1915 1230 2000 1245
rect 1915 1165 1925 1230
rect 1990 1165 2000 1230
rect 1915 1150 2000 1165
rect 1915 1085 1925 1150
rect 1990 1085 2000 1150
rect 1915 915 2000 1085
rect 1915 850 1925 915
rect 1990 850 2000 915
rect 1915 835 2000 850
rect 1915 770 1925 835
rect 1990 770 2000 835
rect 1915 755 2000 770
rect 1915 690 1925 755
rect 1990 690 2000 755
rect 1915 680 2000 690
rect 0 430 2000 440
rect 0 345 10 430
rect 95 345 1905 430
rect 1990 345 2000 430
rect 0 335 2000 345
rect 0 250 10 335
rect 95 250 1905 335
rect 1990 250 2000 335
rect 0 190 2000 250
rect 0 105 10 190
rect 95 125 1905 190
rect 95 105 440 125
rect 0 95 440 105
rect 0 10 10 95
rect 95 10 105 95
rect 190 10 250 95
rect 335 10 345 95
rect 430 10 440 95
rect 1560 105 1905 125
rect 1990 105 2000 190
rect 1560 95 2000 105
rect 0 0 440 10
rect 680 75 1320 85
rect 680 10 690 75
rect 755 10 770 75
rect 835 10 850 75
rect 915 10 1085 75
rect 1150 10 1165 75
rect 1230 10 1245 75
rect 1310 10 1320 75
rect 680 0 1320 10
rect 1560 10 1570 95
rect 1655 10 1665 95
rect 1750 10 1810 95
rect 1895 10 1905 95
rect 1990 10 2000 95
rect 1560 0 2000 10
<< via3 >>
rect 10 1905 95 1990
rect 105 1905 190 1990
rect 250 1905 335 1990
rect 345 1905 430 1990
rect 690 1925 755 1990
rect 770 1925 835 1990
rect 850 1925 915 1990
rect 1085 1925 1150 1990
rect 1165 1925 1230 1990
rect 1245 1925 1310 1990
rect 10 1810 95 1895
rect 1570 1905 1655 1990
rect 1665 1905 1750 1990
rect 1810 1905 1895 1990
rect 1905 1905 1990 1990
rect 1905 1810 1990 1895
rect 10 1665 95 1750
rect 1905 1665 1990 1750
rect 10 1570 95 1655
rect 1905 1570 1990 1655
rect 10 1245 75 1310
rect 10 1165 75 1230
rect 10 1085 75 1150
rect 10 850 75 915
rect 10 770 75 835
rect 10 690 75 755
rect 1925 1245 1990 1310
rect 1925 1165 1990 1230
rect 1925 1085 1990 1150
rect 1925 850 1990 915
rect 1925 770 1990 835
rect 1925 690 1990 755
rect 10 345 95 430
rect 1905 345 1990 430
rect 10 250 95 335
rect 1905 250 1990 335
rect 10 105 95 190
rect 10 10 95 95
rect 105 10 190 95
rect 250 10 335 95
rect 345 10 430 95
rect 1905 105 1990 190
rect 690 10 755 75
rect 770 10 835 75
rect 850 10 915 75
rect 1085 10 1150 75
rect 1165 10 1230 75
rect 1245 10 1310 75
rect 1570 10 1655 95
rect 1665 10 1750 95
rect 1810 10 1895 95
rect 1905 10 1990 95
<< mimcap >>
rect 140 1845 1860 1860
rect 140 155 155 1845
rect 1845 155 1860 1845
rect 140 140 1860 155
<< mimcapcontact >>
rect 155 155 1845 1845
<< metal4 >>
rect 0 1990 440 2000
rect 0 1905 10 1990
rect 95 1905 105 1990
rect 190 1905 250 1990
rect 335 1905 345 1990
rect 430 1905 440 1990
rect 0 1895 440 1905
rect 680 1990 1320 2000
rect 680 1925 690 1990
rect 755 1925 770 1990
rect 835 1925 850 1990
rect 915 1925 1085 1990
rect 1150 1925 1165 1990
rect 1230 1925 1245 1990
rect 1310 1925 1320 1990
rect 0 1810 10 1895
rect 95 1810 105 1895
rect 680 1855 1320 1925
rect 1560 1990 2000 2000
rect 1560 1905 1570 1990
rect 1655 1905 1665 1990
rect 1750 1905 1810 1990
rect 1895 1905 1905 1990
rect 1990 1905 2000 1990
rect 1560 1895 2000 1905
rect 0 1750 105 1810
rect 0 1665 10 1750
rect 95 1665 105 1750
rect 0 1655 105 1665
rect 0 1570 10 1655
rect 95 1570 105 1655
rect 0 1560 105 1570
rect 145 1845 1855 1855
rect 145 1320 155 1845
rect 0 1310 155 1320
rect 0 1245 10 1310
rect 75 1245 155 1310
rect 0 1230 155 1245
rect 0 1165 10 1230
rect 75 1165 155 1230
rect 0 1150 155 1165
rect 0 1085 10 1150
rect 75 1085 155 1150
rect 0 915 155 1085
rect 0 850 10 915
rect 75 850 155 915
rect 0 835 155 850
rect 0 770 10 835
rect 75 770 155 835
rect 0 755 155 770
rect 0 690 10 755
rect 75 690 155 755
rect 0 680 155 690
rect 0 430 105 440
rect 0 345 10 430
rect 95 345 105 430
rect 0 335 105 345
rect 0 250 10 335
rect 95 250 105 335
rect 0 190 105 250
rect 0 105 10 190
rect 95 105 105 190
rect 145 155 155 680
rect 1845 1320 1855 1845
rect 1895 1810 1905 1895
rect 1990 1810 2000 1895
rect 1895 1750 2000 1810
rect 1895 1665 1905 1750
rect 1990 1665 2000 1750
rect 1895 1655 2000 1665
rect 1895 1570 1905 1655
rect 1990 1570 2000 1655
rect 1895 1560 2000 1570
rect 1845 1310 2000 1320
rect 1845 1245 1925 1310
rect 1990 1245 2000 1310
rect 1845 1230 2000 1245
rect 1845 1165 1925 1230
rect 1990 1165 2000 1230
rect 1845 1150 2000 1165
rect 1845 1085 1925 1150
rect 1990 1085 2000 1150
rect 1845 915 2000 1085
rect 1845 850 1925 915
rect 1990 850 2000 915
rect 1845 835 2000 850
rect 1845 770 1925 835
rect 1990 770 2000 835
rect 1845 755 2000 770
rect 1845 690 1925 755
rect 1990 690 2000 755
rect 1845 680 2000 690
rect 1845 155 1855 680
rect 145 145 1855 155
rect 1895 430 2000 440
rect 1895 345 1905 430
rect 1990 345 2000 430
rect 1895 335 2000 345
rect 1895 250 1905 335
rect 1990 250 2000 335
rect 1895 190 2000 250
rect 0 95 440 105
rect 0 10 10 95
rect 95 10 105 95
rect 190 10 250 95
rect 335 10 345 95
rect 430 10 440 95
rect 0 0 440 10
rect 680 75 1320 145
rect 1895 105 1905 190
rect 1990 105 2000 190
rect 680 10 690 75
rect 755 10 770 75
rect 835 10 850 75
rect 915 10 1085 75
rect 1150 10 1165 75
rect 1230 10 1245 75
rect 1310 10 1320 75
rect 680 0 1320 10
rect 1560 95 2000 105
rect 1560 10 1570 95
rect 1655 10 1665 95
rect 1750 10 1810 95
rect 1895 10 1905 95
rect 1990 10 2000 95
rect 1560 0 2000 10
<< labels >>
flabel metal1 s 680 0 1320 90 5 FreeSans 160 0 0 0 nmoscap_top
port 1 s
flabel metal1 s 680 1910 1320 2000 1 FreeSans 160 0 0 0 nmoscap_top
port 1 n
flabel metal1 s 1910 680 2000 1320 3 FreeSans 160 90 0 0 nmoscap_top
port 1 e
flabel metal1 s 0 680 90 1320 7 FreeSans 160 90 0 0 nmoscap_top
port 1 w
flabel metal1 s 0 1560 120 2000 7 FreeSans 160 90 0 0 nmoscap_bot
port 2 w
flabel metal1 s 0 0 120 440 7 FreeSans 160 90 0 0 nmoscap_bot
port 2 w
flabel metal1 s 1880 0 2000 440 3 FreeSans 160 90 0 0 nmoscap_bot
port 2 e
flabel metal1 s 1880 1560 2000 2000 3 FreeSans 160 90 0 0 nmoscap_bot
port 2 e
flabel metal1 s 1560 1880 2000 2000 1 FreeSans 160 0 0 0 nmoscap_bot
port 2 n
flabel metal1 s 0 1880 440 2000 1 FreeSans 160 0 0 0 nmoscap_bot
port 2 n
flabel metal1 s 0 0 440 120 5 FreeSans 160 0 0 0 nmoscap_bot
port 2 s
flabel metal1 s 1560 0 2000 120 5 FreeSans 160 0 0 0 nmoscap_bot
port 2 s
flabel locali s 445 0 675 40 5 FreeSans 160 0 0 0 pwell
port 3 s
flabel locali s 1325 0 1555 40 5 FreeSans 160 0 0 0 pwell
port 3 s
flabel locali s 1325 1960 1555 2000 1 FreeSans 160 0 0 0 pwell
port 3 n
flabel locali s 445 1960 675 2000 1 FreeSans 160 0 0 0 pwell
port 3 n
flabel locali s 1960 1325 2000 1555 3 FreeSans 160 90 0 0 pwell
port 3 e
flabel locali s 1960 445 2000 675 3 FreeSans 160 90 0 0 pwell
port 3 e
flabel locali s 0 445 40 675 7 FreeSans 160 90 0 0 pwell
port 3 w
flabel locali s 0 1325 40 1555 7 FreeSans 160 90 0 0 pwell
port 3 w
flabel metal3 680 1915 1320 2000 1 FreeSans 160 0 0 0 mimcap_top
port 4 n
flabel metal3 680 0 1320 85 5 FreeSans 160 0 0 0 mimcap_top
port 4 s
flabel metal3 1915 680 2000 1320 3 FreeSans 160 90 0 0 mimcap_top
port 4 e
flabel metal3 0 680 85 1320 7 FreeSans 160 90 0 0 mimcap_top
port 4 w
flabel metal3 1560 0 2000 125 5 FreeSans 160 0 0 0 mimcap_bot
port 5 s
flabel metal3 0 0 440 125 5 FreeSans 160 0 0 0 mimcap_bot
port 5 s
flabel metal3 0 1875 440 2000 1 FreeSans 160 0 0 0 mimcap_bot
port 5 n
flabel metal3 1560 1875 2000 2000 1 FreeSans 160 0 0 0 mimcap_bot
port 5 n
flabel metal3 1875 1560 2000 2000 3 FreeSans 160 90 0 0 mimcap_bot
port 5 e
flabel metal3 1875 0 2000 440 3 FreeSans 160 90 0 0 mimcap_bot
port 5 e
flabel metal3 0 0 125 440 7 FreeSans 160 90 0 0 mimcap_bot
port 5 w
flabel metal3 0 1560 125 2000 7 FreeSans 160 90 0 0 mimcap_bot
port 5 w
<< properties >>
string FIXED_BBOX 0 0 2000 2000
<< end >>
