magic
tech sky130A
magscale 1 2
timestamp 1661178173
<< error_p >>
rect -9 1873 2191 1933
rect 2291 1873 4491 1933
rect -9 1793 2191 1853
rect 2291 1793 4491 1853
<< nwell >>
rect -50 -196 848 144
<< nmos >>
rect 48 -910 78 -510
rect 144 -910 174 -510
rect 240 -910 270 -510
rect 336 -910 366 -510
rect 432 -910 462 -510
rect 528 -910 558 -510
rect 624 -910 654 -510
rect 720 -910 750 -510
rect 48 -1170 78 -1070
rect 144 -1170 174 -1070
rect 240 -1170 270 -1070
rect 336 -1170 366 -1070
rect 432 -1170 462 -1070
rect 528 -1170 558 -1070
rect 624 -1170 654 -1070
rect 720 -1170 750 -1070
<< pmos >>
rect 48 -96 78 4
rect 144 -96 174 4
rect 240 -96 270 4
rect 336 -96 366 4
rect 432 -96 462 4
rect 528 -96 558 4
rect 624 -96 654 4
rect 720 -96 750 4
<< ndiff >>
rect -14 -522 48 -510
rect -14 -898 -2 -522
rect 32 -898 48 -522
rect -14 -910 48 -898
rect 78 -522 144 -510
rect 78 -898 94 -522
rect 128 -898 144 -522
rect 78 -910 144 -898
rect 174 -522 240 -510
rect 174 -898 190 -522
rect 224 -898 240 -522
rect 174 -910 240 -898
rect 270 -522 336 -510
rect 270 -898 286 -522
rect 320 -898 336 -522
rect 270 -910 336 -898
rect 366 -522 432 -510
rect 366 -898 382 -522
rect 416 -898 432 -522
rect 366 -910 432 -898
rect 462 -522 528 -510
rect 462 -898 478 -522
rect 512 -898 528 -522
rect 462 -910 528 -898
rect 558 -522 624 -510
rect 558 -898 574 -522
rect 608 -898 624 -522
rect 558 -910 624 -898
rect 654 -522 720 -510
rect 654 -898 670 -522
rect 704 -898 720 -522
rect 654 -910 720 -898
rect 750 -522 812 -510
rect 750 -898 766 -522
rect 800 -898 812 -522
rect 750 -910 812 -898
rect -14 -1082 48 -1070
rect -14 -1158 -2 -1082
rect 32 -1158 48 -1082
rect -14 -1170 48 -1158
rect 78 -1082 144 -1070
rect 78 -1158 94 -1082
rect 128 -1158 144 -1082
rect 78 -1170 144 -1158
rect 174 -1082 240 -1070
rect 174 -1158 190 -1082
rect 224 -1158 240 -1082
rect 174 -1170 240 -1158
rect 270 -1082 336 -1070
rect 270 -1158 286 -1082
rect 320 -1158 336 -1082
rect 270 -1170 336 -1158
rect 366 -1082 432 -1070
rect 366 -1158 382 -1082
rect 416 -1158 432 -1082
rect 366 -1170 432 -1158
rect 462 -1082 528 -1070
rect 462 -1158 478 -1082
rect 512 -1158 528 -1082
rect 462 -1170 528 -1158
rect 558 -1082 624 -1070
rect 558 -1158 574 -1082
rect 608 -1158 624 -1082
rect 558 -1170 624 -1158
rect 654 -1082 720 -1070
rect 654 -1158 670 -1082
rect 704 -1158 720 -1082
rect 654 -1170 720 -1158
rect 750 -1082 812 -1070
rect 750 -1158 766 -1082
rect 800 -1158 812 -1082
rect 750 -1170 812 -1158
<< pdiff >>
rect -14 -8 48 4
rect -14 -84 -2 -8
rect 32 -84 48 -8
rect -14 -96 48 -84
rect 78 -8 144 4
rect 78 -84 94 -8
rect 128 -84 144 -8
rect 78 -96 144 -84
rect 174 -8 240 4
rect 174 -84 190 -8
rect 224 -84 240 -8
rect 174 -96 240 -84
rect 270 -8 336 4
rect 270 -84 286 -8
rect 320 -84 336 -8
rect 270 -96 336 -84
rect 366 -8 432 4
rect 366 -84 382 -8
rect 416 -84 432 -8
rect 366 -96 432 -84
rect 462 -8 528 4
rect 462 -84 478 -8
rect 512 -84 528 -8
rect 462 -96 528 -84
rect 558 -8 624 4
rect 558 -84 574 -8
rect 608 -84 624 -8
rect 558 -96 624 -84
rect 654 -8 720 4
rect 654 -84 670 -8
rect 704 -84 720 -8
rect 654 -96 720 -84
rect 750 -8 812 4
rect 750 -84 766 -8
rect 800 -84 812 -8
rect 750 -96 812 -84
<< ndiffc >>
rect -2 -898 32 -522
rect 94 -898 128 -522
rect 190 -898 224 -522
rect 286 -898 320 -522
rect 382 -898 416 -522
rect 478 -898 512 -522
rect 574 -898 608 -522
rect 670 -898 704 -522
rect 766 -898 800 -522
rect -2 -1158 32 -1082
rect 94 -1158 128 -1082
rect 190 -1158 224 -1082
rect 286 -1158 320 -1082
rect 382 -1158 416 -1082
rect 478 -1158 512 -1082
rect 574 -1158 608 -1082
rect 670 -1158 704 -1082
rect 766 -1158 800 -1082
<< pdiffc >>
rect -2 -84 32 -8
rect 94 -84 128 -8
rect 190 -84 224 -8
rect 286 -84 320 -8
rect 382 -84 416 -8
rect 478 -84 512 -8
rect 574 -84 608 -8
rect 670 -84 704 -8
rect 766 -84 800 -8
<< psubdiff >>
rect -26 -1228 830 -1226
rect -26 -1264 4 -1228
rect 40 -1264 122 -1228
rect 158 -1264 240 -1228
rect 276 -1264 358 -1228
rect 394 -1264 476 -1228
rect 512 -1264 594 -1228
rect 630 -1264 712 -1228
rect 748 -1264 830 -1228
rect -26 -1268 830 -1264
<< nsubdiff >>
rect -14 100 812 108
rect -14 66 16 100
rect 50 66 100 100
rect 134 66 184 100
rect 218 66 268 100
rect 302 66 352 100
rect 386 66 436 100
rect 470 66 520 100
rect 554 66 604 100
rect 638 66 688 100
rect 722 66 812 100
rect -14 60 812 66
<< psubdiffcont >>
rect 4 -1264 40 -1228
rect 122 -1264 158 -1228
rect 240 -1264 276 -1228
rect 358 -1264 394 -1228
rect 476 -1264 512 -1228
rect 594 -1264 630 -1228
rect 712 -1264 748 -1228
<< nsubdiffcont >>
rect 16 66 50 100
rect 100 66 134 100
rect 184 66 218 100
rect 268 66 302 100
rect 352 66 386 100
rect 436 66 470 100
rect 520 66 554 100
rect 604 66 638 100
rect 688 66 722 100
<< poly >>
rect 48 4 78 30
rect 144 4 174 30
rect 240 4 270 30
rect 336 4 366 30
rect 432 4 462 30
rect 528 4 558 30
rect 624 4 654 30
rect 720 4 750 30
rect 48 -122 78 -96
rect 144 -122 174 -96
rect 240 -122 270 -96
rect 336 -122 366 -96
rect 432 -122 462 -96
rect 528 -122 558 -96
rect 624 -122 654 -96
rect 720 -122 750 -96
rect 48 -154 750 -122
rect 174 -316 226 -260
rect 188 -454 226 -316
rect 566 -382 618 -326
rect 572 -454 610 -382
rect 48 -484 366 -454
rect 48 -510 78 -484
rect 144 -510 174 -484
rect 240 -510 270 -484
rect 336 -510 366 -484
rect 432 -484 750 -454
rect 432 -510 462 -484
rect 528 -510 558 -484
rect 624 -510 654 -484
rect 720 -510 750 -484
rect 48 -938 78 -910
rect 144 -938 174 -910
rect 240 -938 270 -910
rect 336 -938 366 -910
rect 432 -938 462 -910
rect 528 -938 558 -910
rect 624 -938 654 -910
rect 720 -938 750 -910
rect 48 -1044 750 -1014
rect 48 -1070 78 -1044
rect 144 -1070 174 -1044
rect 240 -1070 270 -1044
rect 336 -1070 366 -1044
rect 432 -1070 462 -1044
rect 528 -1070 558 -1044
rect 624 -1070 654 -1044
rect 720 -1070 750 -1044
rect 48 -1196 78 -1170
rect 144 -1196 174 -1170
rect 240 -1196 270 -1170
rect 336 -1196 366 -1170
rect 432 -1196 462 -1170
rect 528 -1196 558 -1170
rect 624 -1196 654 -1170
rect 720 -1196 750 -1170
<< locali >>
rect -14 100 812 108
rect -14 66 16 100
rect 50 66 100 100
rect 134 66 184 100
rect 218 66 268 100
rect 302 66 352 100
rect 386 66 436 100
rect 470 66 520 100
rect 554 66 604 100
rect 638 66 688 100
rect 722 66 812 100
rect -14 60 812 66
rect -2 42 800 60
rect -2 -8 32 42
rect -2 -100 32 -84
rect 94 -8 128 8
rect 94 -160 128 -84
rect 190 -8 224 42
rect 190 -100 224 -84
rect 286 -8 320 8
rect 286 -160 320 -84
rect 382 -8 416 42
rect 382 -100 416 -84
rect 478 -8 512 8
rect 94 -194 320 -160
rect 174 -266 226 -260
rect 174 -306 180 -266
rect 220 -306 226 -266
rect 174 -316 226 -306
rect 286 -418 320 -194
rect 94 -452 320 -418
rect -2 -522 32 -506
rect -2 -948 32 -898
rect 94 -522 128 -452
rect 94 -914 128 -898
rect 190 -522 224 -506
rect 190 -948 224 -898
rect 286 -522 320 -452
rect 478 -156 512 -84
rect 574 -8 608 42
rect 574 -100 608 -84
rect 670 -8 704 8
rect 670 -156 704 -84
rect 766 -8 800 42
rect 766 -100 800 -84
rect 478 -190 704 -156
rect 478 -416 512 -190
rect 566 -332 618 -326
rect 566 -372 572 -332
rect 612 -372 618 -332
rect 566 -382 618 -372
rect 478 -450 704 -416
rect 286 -914 320 -898
rect 382 -522 416 -506
rect 382 -948 416 -898
rect 478 -522 512 -450
rect 478 -914 512 -898
rect 574 -522 608 -506
rect 574 -948 608 -898
rect 670 -522 704 -450
rect 670 -914 704 -898
rect 766 -522 800 -506
rect 766 -948 800 -898
rect -2 -984 800 -948
rect -2 -1082 32 -984
rect -2 -1174 32 -1158
rect 94 -1082 128 -1064
rect 94 -1212 128 -1158
rect 190 -1082 224 -984
rect 190 -1174 224 -1158
rect 286 -1082 320 -1066
rect 286 -1212 320 -1158
rect 382 -1082 416 -984
rect 382 -1174 416 -1158
rect 478 -1082 512 -1066
rect 478 -1212 512 -1158
rect 574 -1082 608 -984
rect 574 -1174 608 -1158
rect 670 -1082 704 -1066
rect 670 -1212 704 -1158
rect 766 -1082 800 -984
rect 766 -1174 800 -1158
rect 94 -1226 704 -1212
rect -26 -1228 830 -1226
rect -26 -1264 4 -1228
rect 40 -1264 122 -1228
rect 158 -1264 240 -1228
rect 276 -1264 358 -1228
rect 394 -1264 476 -1228
rect 512 -1264 594 -1228
rect 630 -1264 712 -1228
rect 748 -1264 830 -1228
rect -26 -1268 830 -1264
<< viali >>
rect -2 -84 32 -8
rect 94 -84 128 -8
rect 190 -84 224 -8
rect 286 -84 320 -8
rect 382 -84 416 -8
rect 478 -84 512 -8
rect 180 -306 220 -266
rect -2 -898 32 -522
rect 94 -898 128 -522
rect 190 -898 224 -522
rect 574 -84 608 -8
rect 670 -84 704 -8
rect 766 -84 800 -8
rect 572 -372 612 -332
rect 286 -898 320 -522
rect 382 -898 416 -522
rect 478 -898 512 -522
rect 574 -898 608 -522
rect 670 -898 704 -522
rect 766 -898 800 -522
rect -2 -1158 32 -1082
rect 94 -1158 128 -1082
rect 190 -1158 224 -1082
rect 286 -1158 320 -1082
rect 382 -1158 416 -1082
rect 478 -1158 512 -1082
rect 574 -1158 608 -1082
rect 670 -1158 704 -1082
rect 766 -1158 800 -1082
rect 4 -1264 40 -1228
rect 122 -1264 158 -1228
rect 240 -1264 276 -1228
rect 358 -1264 394 -1228
rect 476 -1264 512 -1228
rect 594 -1264 630 -1228
rect 712 -1264 748 -1228
<< metal1 >>
rect -14 60 812 108
rect -8 -8 38 4
rect -8 -84 -2 -8
rect 32 -84 38 -8
rect -8 -96 38 -84
rect 88 -8 134 4
rect 88 -84 94 -8
rect 128 -84 134 -8
rect 88 -96 134 -84
rect 184 -8 230 4
rect 184 -84 190 -8
rect 224 -84 230 -8
rect 184 -96 230 -84
rect 280 -8 326 4
rect 280 -84 286 -8
rect 320 -84 326 -8
rect 280 -96 326 -84
rect 376 -8 422 4
rect 376 -84 382 -8
rect 416 -84 422 -8
rect 376 -96 422 -84
rect 472 -8 518 4
rect 472 -84 478 -8
rect 512 -84 518 -8
rect 472 -96 518 -84
rect 568 -8 614 4
rect 568 -84 574 -8
rect 608 -84 614 -8
rect 568 -96 614 -84
rect 664 -8 710 4
rect 664 -84 670 -8
rect 704 -84 710 -8
rect 664 -96 710 -84
rect 760 -8 806 4
rect 760 -84 766 -8
rect 800 -84 806 -8
rect 760 -96 806 -84
rect 94 -230 296 -202
rect 88 -266 232 -258
rect 88 -286 180 -266
rect 168 -306 180 -286
rect 220 -306 232 -266
rect 168 -316 232 -306
rect 268 -378 296 -230
rect 560 -332 624 -326
rect 560 -372 572 -332
rect 612 -372 624 -332
rect 560 -378 624 -372
rect 268 -406 624 -378
rect -8 -522 38 -510
rect -8 -898 -2 -522
rect 32 -898 38 -522
rect -8 -910 38 -898
rect 88 -522 134 -510
rect 88 -898 94 -522
rect 128 -898 134 -522
rect 88 -910 134 -898
rect 184 -522 230 -510
rect 184 -898 190 -522
rect 224 -898 230 -522
rect 184 -910 230 -898
rect 280 -522 326 -510
rect 280 -898 286 -522
rect 320 -898 326 -522
rect 280 -910 326 -898
rect 376 -522 422 -510
rect 376 -898 382 -522
rect 416 -898 422 -522
rect 376 -910 422 -898
rect 472 -522 518 -510
rect 472 -898 478 -522
rect 512 -898 518 -522
rect 472 -910 518 -898
rect 568 -522 614 -510
rect 568 -898 574 -522
rect 608 -898 614 -522
rect 568 -910 614 -898
rect 664 -522 710 -510
rect 664 -898 670 -522
rect 704 -898 710 -522
rect 664 -910 710 -898
rect 760 -522 806 -510
rect 760 -898 766 -522
rect 800 -898 806 -522
rect 760 -910 806 -898
rect -8 -1082 38 -1070
rect -8 -1158 -2 -1082
rect 32 -1158 38 -1082
rect -8 -1170 38 -1158
rect 88 -1082 134 -1070
rect 88 -1158 94 -1082
rect 128 -1158 134 -1082
rect 88 -1170 134 -1158
rect 184 -1082 230 -1070
rect 184 -1158 190 -1082
rect 224 -1158 230 -1082
rect 184 -1170 230 -1158
rect 280 -1082 326 -1070
rect 280 -1158 286 -1082
rect 320 -1158 326 -1082
rect 280 -1170 326 -1158
rect 376 -1082 422 -1070
rect 376 -1158 382 -1082
rect 416 -1158 422 -1082
rect 376 -1170 422 -1158
rect 472 -1082 518 -1070
rect 472 -1158 478 -1082
rect 512 -1158 518 -1082
rect 472 -1170 518 -1158
rect 568 -1082 614 -1070
rect 568 -1158 574 -1082
rect 608 -1158 614 -1082
rect 568 -1170 614 -1158
rect 664 -1082 710 -1070
rect 664 -1158 670 -1082
rect 704 -1158 710 -1082
rect 664 -1170 710 -1158
rect 760 -1082 806 -1070
rect 760 -1158 766 -1082
rect 800 -1158 806 -1082
rect 760 -1170 806 -1158
rect -26 -1228 830 -1222
rect -26 -1264 4 -1228
rect 40 -1264 122 -1228
rect 158 -1264 240 -1228
rect 276 -1264 358 -1228
rect 394 -1264 476 -1228
rect 512 -1264 594 -1228
rect 630 -1264 712 -1228
rect 748 -1264 830 -1228
rect -26 -1270 830 -1264
use sky130_fd_pr__cap_mim_m3_1_55Z62P  sky130_fd_pr__cap_mim_m3_1_55Z62P_0
timestamp 1661178173
transform 0 1 2241 -1 0 1863
box -1509 -2300 1509 2300
<< end >>
