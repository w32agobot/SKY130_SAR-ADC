magic
tech sky130A
timestamp 1662907922
<< nwell >>
rect 117 474 521 661
<< nmos >>
rect 186 347 201 389
rect 234 347 249 389
rect 338 347 353 389
rect 386 347 401 389
rect 434 347 449 389
<< pmos >>
rect 186 492 201 572
rect 234 492 249 572
rect 338 508 353 588
rect 386 508 401 588
rect 434 508 449 588
<< ndiff >>
rect 155 383 186 389
rect 155 353 161 383
rect 178 353 186 383
rect 155 347 186 353
rect 201 383 234 389
rect 201 353 209 383
rect 226 353 234 383
rect 201 347 234 353
rect 249 383 280 389
rect 249 353 257 383
rect 274 353 280 383
rect 249 347 280 353
rect 307 383 338 389
rect 307 353 313 383
rect 330 353 338 383
rect 307 347 338 353
rect 353 383 386 389
rect 353 353 361 383
rect 378 353 386 383
rect 353 347 386 353
rect 401 383 434 389
rect 401 353 409 383
rect 426 353 434 383
rect 401 347 434 353
rect 449 383 480 389
rect 449 353 457 383
rect 474 353 480 383
rect 449 347 480 353
<< pdiff >>
rect 307 582 338 588
rect 155 566 186 572
rect 155 498 161 566
rect 178 498 186 566
rect 155 492 186 498
rect 201 566 234 572
rect 201 498 209 566
rect 226 498 234 566
rect 201 492 234 498
rect 249 566 280 572
rect 249 498 257 566
rect 274 498 280 566
rect 307 514 313 582
rect 330 514 338 582
rect 307 508 338 514
rect 353 582 386 588
rect 353 514 361 582
rect 378 514 386 582
rect 353 508 386 514
rect 401 582 434 588
rect 401 514 409 582
rect 426 514 434 582
rect 401 508 434 514
rect 449 582 480 588
rect 449 514 457 582
rect 474 514 480 582
rect 449 508 480 514
rect 249 492 280 498
<< ndiffc >>
rect 161 353 178 383
rect 209 353 226 383
rect 257 353 274 383
rect 313 353 330 383
rect 361 353 378 383
rect 409 353 426 383
rect 457 353 474 383
<< pdiffc >>
rect 161 498 178 566
rect 209 498 226 566
rect 257 498 274 566
rect 313 514 330 582
rect 361 514 378 582
rect 409 514 426 582
rect 457 514 474 582
<< psubdiff >>
rect 161 295 185 312
rect 202 295 233 312
rect 250 295 262 312
rect 409 295 433 312
rect 450 295 466 312
<< nsubdiff >>
rect 221 640 473 643
rect 221 623 233 640
rect 250 623 285 640
rect 302 623 337 640
rect 354 623 385 640
rect 402 623 432 640
rect 449 623 473 640
rect 221 620 473 623
<< psubdiffcont >>
rect 185 295 202 312
rect 233 295 250 312
rect 433 295 450 312
<< nsubdiffcont >>
rect 233 623 250 640
rect 285 623 302 640
rect 337 623 354 640
rect 385 623 402 640
rect 432 623 449 640
<< poly >>
rect 176 630 210 635
rect 176 612 184 630
rect 202 612 210 630
rect 176 580 210 612
rect 338 588 353 601
rect 386 588 401 601
rect 434 588 449 601
rect 186 572 201 580
rect 234 572 249 585
rect 186 389 201 492
rect 234 475 249 492
rect 338 489 353 508
rect 386 495 401 508
rect 434 500 449 508
rect 434 495 487 500
rect 234 465 268 475
rect 234 446 243 465
rect 260 446 268 465
rect 234 397 268 446
rect 317 420 353 489
rect 374 479 487 495
rect 374 461 408 479
rect 382 436 400 461
rect 453 459 487 479
rect 382 434 408 436
rect 338 417 353 420
rect 374 417 408 434
rect 338 402 449 417
rect 234 389 249 397
rect 338 389 353 402
rect 386 389 401 402
rect 434 389 449 402
rect 186 334 201 347
rect 234 334 249 347
rect 338 334 353 347
rect 386 334 401 347
rect 434 334 449 347
rect 338 324 401 334
rect 325 319 401 324
rect 323 302 331 319
rect 348 302 365 319
rect 382 302 390 319
rect 323 296 390 302
<< polycont >>
rect 184 612 202 630
rect 243 446 260 465
rect 331 302 348 319
rect 365 302 382 319
<< locali >>
rect 127 574 144 664
rect 221 640 473 643
rect 184 630 202 638
rect 221 623 233 640
rect 250 623 285 640
rect 302 623 337 640
rect 354 623 385 640
rect 402 623 432 640
rect 449 623 473 640
rect 221 620 473 623
rect 184 607 202 612
rect 184 590 185 607
rect 257 582 330 590
rect 127 566 178 574
rect 127 498 161 566
rect 127 491 178 498
rect 127 354 144 491
rect 161 490 178 491
rect 209 566 226 574
rect 161 389 184 391
rect 161 383 167 389
rect 178 367 184 372
rect 209 383 226 498
rect 257 571 313 582
rect 257 566 286 571
rect 274 553 286 566
rect 303 553 313 571
rect 274 532 313 553
rect 274 514 286 532
rect 303 514 313 532
rect 274 506 330 514
rect 361 582 378 620
rect 361 506 378 514
rect 409 582 426 602
rect 274 498 294 506
rect 409 501 426 514
rect 457 582 474 590
rect 457 506 474 514
rect 257 490 294 498
rect 243 465 260 473
rect 243 428 260 446
rect 243 408 260 411
rect 277 425 294 490
rect 277 408 308 425
rect 291 391 308 408
rect 161 345 178 353
rect 209 345 226 353
rect 257 383 274 391
rect 291 389 330 391
rect 291 372 299 389
rect 316 383 330 389
rect 291 371 313 372
rect 257 351 274 353
rect 127 285 144 337
rect 313 345 330 353
rect 361 383 378 391
rect 361 345 378 353
rect 409 383 426 391
rect 257 331 274 334
rect 331 319 348 324
rect 365 319 382 324
rect 161 295 185 312
rect 202 295 233 312
rect 250 295 262 312
rect 323 302 331 319
rect 348 302 365 319
rect 382 302 390 319
rect 409 312 426 353
rect 457 383 474 391
rect 457 345 474 353
rect 331 285 348 302
rect 365 296 382 302
rect 409 295 433 312
rect 450 295 466 312
rect 497 285 514 664
<< viali >>
rect 233 623 250 640
rect 285 623 302 640
rect 337 623 354 640
rect 385 623 402 640
rect 432 623 449 640
rect 185 590 202 607
rect 209 547 226 565
rect 209 508 226 526
rect 127 337 144 354
rect 167 383 184 389
rect 167 372 178 383
rect 178 372 184 383
rect 286 553 303 571
rect 286 514 303 532
rect 457 553 474 571
rect 457 514 474 532
rect 243 411 260 428
rect 299 383 316 389
rect 299 372 313 383
rect 313 372 316 383
rect 257 334 274 351
rect 361 366 378 383
rect 185 295 202 312
rect 233 295 250 312
rect 457 366 474 383
rect 433 295 450 312
<< metal1 >>
rect 117 640 521 648
rect 117 624 233 640
rect 117 620 168 624
rect 219 623 233 624
rect 250 623 285 640
rect 302 623 337 640
rect 354 623 385 640
rect 402 623 432 640
rect 449 623 521 640
rect 219 620 521 623
rect 179 607 208 610
rect 179 606 185 607
rect 117 591 185 606
rect 179 590 185 591
rect 202 606 208 607
rect 202 591 521 606
rect 202 590 208 591
rect 179 587 208 590
rect 203 570 232 572
rect 283 571 306 577
rect 202 544 205 570
rect 231 544 234 570
rect 202 531 234 544
rect 202 505 205 531
rect 231 505 234 531
rect 283 553 286 571
rect 303 554 306 571
rect 454 571 477 577
rect 454 554 457 571
rect 303 553 457 554
rect 474 553 477 571
rect 283 540 477 553
rect 283 532 306 540
rect 283 514 286 532
rect 303 514 306 532
rect 283 508 306 514
rect 454 532 477 540
rect 454 514 457 532
rect 474 514 477 532
rect 454 508 477 514
rect 457 505 474 508
rect 117 477 521 491
rect 318 464 347 477
rect 153 450 295 460
rect 367 450 398 453
rect 455 450 485 463
rect 117 445 521 450
rect 117 436 167 445
rect 281 436 521 445
rect 237 428 266 431
rect 367 430 398 436
rect 237 422 243 428
rect 117 411 243 422
rect 260 422 266 428
rect 260 416 353 422
rect 438 416 521 422
rect 260 411 521 416
rect 117 408 521 411
rect 237 405 266 408
rect 335 402 478 408
rect 161 389 190 394
rect 161 372 167 389
rect 184 385 190 389
rect 293 389 322 394
rect 293 385 299 389
rect 184 372 299 385
rect 316 372 322 389
rect 161 371 322 372
rect 161 367 190 371
rect 293 367 322 371
rect 355 383 480 387
rect 355 366 361 383
rect 378 366 457 383
rect 474 366 480 383
rect 355 363 480 366
rect 124 354 147 360
rect 124 345 127 354
rect 117 337 127 345
rect 144 345 147 354
rect 254 351 278 357
rect 254 345 257 351
rect 144 337 257 345
rect 117 334 257 337
rect 274 345 278 351
rect 274 334 521 345
rect 117 331 521 334
rect 117 312 521 317
rect 117 295 185 312
rect 202 295 233 312
rect 250 295 433 312
rect 450 295 521 312
rect 117 289 521 295
<< via1 >>
rect 205 565 231 570
rect 205 547 209 565
rect 209 547 226 565
rect 226 547 231 565
rect 205 544 231 547
rect 205 526 231 531
rect 205 508 209 526
rect 209 508 226 526
rect 226 508 231 526
rect 205 505 231 508
<< metal2 >>
rect 202 570 234 572
rect 202 544 205 570
rect 231 544 234 570
rect 202 531 234 544
rect 202 505 205 531
rect 231 505 234 531
rect 202 500 234 505
<< labels >>
rlabel metal1 117 436 117 450 7 col_n
port 6 w
rlabel metal1 117 477 117 491 7 colon_n
port 7 w
rlabel metal1 117 331 117 345 7 vcom
port 3 w
rlabel metal1 117 591 117 606 7 sample_n
port 5 w
rlabel metal1 117 408 117 422 7 sample
port 4 w
rlabel metal1 117 289 117 317 7 VSS
port 2 w
rlabel metal1 117 620 117 648 7 VDD
port 1 w
rlabel locali 409 501 426 501 5 vint1
rlabel locali 497 285 514 285 5 row_n
port 8 s
rlabel locali 457 391 474 391 1 vint2
rlabel locali 291 390 291 405 7 vdrv
rlabel metal2 202 500 234 500 5 cbot
port 9 s
rlabel locali 331 285 348 285 1 en_n
port 10 n
<< end >>
