magic
tech sky130A
magscale 1 2
timestamp 1661174129
<< nwell >>
rect -353 112 449 150
rect -449 -112 449 112
rect -449 -150 353 -112
<< pmos >>
rect -351 -50 -321 50
rect -255 -50 -225 50
rect -159 -50 -129 50
rect -63 -50 -33 50
rect 33 -50 63 50
rect 129 -50 159 50
rect 225 -50 255 50
rect 321 -50 351 50
<< pdiff >>
rect -413 38 -351 50
rect -413 -38 -401 38
rect -367 -38 -351 38
rect -413 -50 -351 -38
rect -321 38 -255 50
rect -321 -38 -305 38
rect -271 -38 -255 38
rect -321 -50 -255 -38
rect -225 38 -159 50
rect -225 -38 -209 38
rect -175 -38 -159 38
rect -225 -50 -159 -38
rect -129 38 -63 50
rect -129 -38 -113 38
rect -79 -38 -63 38
rect -129 -50 -63 -38
rect -33 38 33 50
rect -33 -38 -17 38
rect 17 -38 33 38
rect -33 -50 33 -38
rect 63 38 129 50
rect 63 -38 79 38
rect 113 -38 129 38
rect 63 -50 129 -38
rect 159 38 225 50
rect 159 -38 175 38
rect 209 -38 225 38
rect 159 -50 225 -38
rect 255 38 321 50
rect 255 -38 271 38
rect 305 -38 321 38
rect 255 -50 321 -38
rect 351 38 413 50
rect 351 -38 367 38
rect 401 -38 413 38
rect 351 -50 413 -38
<< pdiffc >>
rect -401 -38 -367 38
rect -305 -38 -271 38
rect -209 -38 -175 38
rect -113 -38 -79 38
rect -17 -38 17 38
rect 79 -38 113 38
rect 175 -38 209 38
rect 271 -38 305 38
rect 367 -38 401 38
<< poly >>
rect -273 131 -207 147
rect -273 97 -257 131
rect -223 97 -207 131
rect -273 81 -207 97
rect -81 131 -15 147
rect -81 97 -65 131
rect -31 97 -15 131
rect -81 81 -15 97
rect 111 131 177 147
rect 111 97 127 131
rect 161 97 177 131
rect 111 81 177 97
rect 303 131 369 147
rect 303 97 319 131
rect 353 97 369 131
rect 303 81 369 97
rect -351 50 -321 76
rect -255 50 -225 81
rect -159 50 -129 76
rect -63 50 -33 81
rect 33 50 63 76
rect 129 50 159 81
rect 225 50 255 76
rect 321 50 351 81
rect -351 -81 -321 -50
rect -255 -76 -225 -50
rect -159 -81 -129 -50
rect -63 -76 -33 -50
rect 33 -81 63 -50
rect 129 -76 159 -50
rect 225 -81 255 -50
rect 321 -76 351 -50
rect -369 -97 -303 -81
rect -369 -131 -353 -97
rect -319 -131 -303 -97
rect -369 -147 -303 -131
rect -177 -97 -111 -81
rect -177 -131 -161 -97
rect -127 -131 -111 -97
rect -177 -147 -111 -131
rect 15 -97 81 -81
rect 15 -131 31 -97
rect 65 -131 81 -97
rect 15 -147 81 -131
rect 207 -97 273 -81
rect 207 -131 223 -97
rect 257 -131 273 -97
rect 207 -147 273 -131
<< polycont >>
rect -257 97 -223 131
rect -65 97 -31 131
rect 127 97 161 131
rect 319 97 353 131
rect -353 -131 -319 -97
rect -161 -131 -127 -97
rect 31 -131 65 -97
rect 223 -131 257 -97
<< locali >>
rect -273 97 -257 131
rect -223 97 -207 131
rect -81 97 -65 131
rect -31 97 -15 131
rect 111 97 127 131
rect 161 97 177 131
rect 303 97 319 131
rect 353 97 369 131
rect -401 38 -367 54
rect -401 -54 -367 -38
rect -305 38 -271 54
rect -305 -54 -271 -38
rect -209 38 -175 54
rect -209 -54 -175 -38
rect -113 38 -79 54
rect -113 -54 -79 -38
rect -17 38 17 54
rect -17 -54 17 -38
rect 79 38 113 54
rect 79 -54 113 -38
rect 175 38 209 54
rect 175 -54 209 -38
rect 271 38 305 54
rect 271 -54 305 -38
rect 367 38 401 54
rect 367 -54 401 -38
rect -369 -131 -353 -97
rect -319 -131 -303 -97
rect -177 -131 -161 -97
rect -127 -131 -111 -97
rect 15 -131 31 -97
rect 65 -131 81 -97
rect 207 -131 223 -97
rect 257 -131 273 -97
<< viali >>
rect -257 97 -223 131
rect -65 97 -31 131
rect 127 97 161 131
rect 319 97 353 131
rect -401 -38 -367 38
rect -305 -38 -271 38
rect -209 -38 -175 38
rect -113 -38 -79 38
rect -17 -38 17 38
rect 79 -38 113 38
rect 175 -38 209 38
rect 271 -38 305 38
rect 367 -38 401 38
rect -353 -131 -319 -97
rect -161 -131 -127 -97
rect 31 -131 65 -97
rect 223 -131 257 -97
<< metal1 >>
rect -269 131 -211 137
rect -269 97 -257 131
rect -223 97 -211 131
rect -269 91 -211 97
rect -77 131 -19 137
rect -77 97 -65 131
rect -31 97 -19 131
rect -77 91 -19 97
rect 115 131 173 137
rect 115 97 127 131
rect 161 97 173 131
rect 115 91 173 97
rect 307 131 365 137
rect 307 97 319 131
rect 353 97 365 131
rect 307 91 365 97
rect -407 38 -361 50
rect -407 -38 -401 38
rect -367 -38 -361 38
rect -407 -50 -361 -38
rect -311 38 -265 50
rect -311 -38 -305 38
rect -271 -38 -265 38
rect -311 -50 -265 -38
rect -215 38 -169 50
rect -215 -38 -209 38
rect -175 -38 -169 38
rect -215 -50 -169 -38
rect -119 38 -73 50
rect -119 -38 -113 38
rect -79 -38 -73 38
rect -119 -50 -73 -38
rect -23 38 23 50
rect -23 -38 -17 38
rect 17 -38 23 38
rect -23 -50 23 -38
rect 73 38 119 50
rect 73 -38 79 38
rect 113 -38 119 38
rect 73 -50 119 -38
rect 169 38 215 50
rect 169 -38 175 38
rect 209 -38 215 38
rect 169 -50 215 -38
rect 265 38 311 50
rect 265 -38 271 38
rect 305 -38 311 38
rect 265 -50 311 -38
rect 361 38 407 50
rect 361 -38 367 38
rect 401 -38 407 38
rect 361 -50 407 -38
rect -365 -97 -307 -91
rect -365 -131 -353 -97
rect -319 -131 -307 -97
rect -365 -137 -307 -131
rect -173 -97 -115 -91
rect -173 -131 -161 -97
rect -127 -131 -115 -97
rect -173 -137 -115 -131
rect 19 -97 77 -91
rect 19 -131 31 -97
rect 65 -131 77 -97
rect 19 -137 77 -131
rect 211 -97 269 -91
rect 211 -131 223 -97
rect 257 -131 269 -97
rect 211 -137 269 -131
<< end >>
