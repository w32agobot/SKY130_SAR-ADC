magic
tech sky130A
timestamp 1659694242
<< metal2 >>
rect 154 2402 184 2538
rect 33 2372 2535 2402
rect 1 139 72 169
rect 154 36 184 2372
rect 1244 1249 1314 1323
rect 1888 1252 1958 1326
rect 656 656 698 707
rect 2529 304 2595 334
rect 605 159 671 189
rect 1254 164 1316 195
rect 1892 166 1954 197
rect 3013 32 3043 2534
rect 3364 2402 3394 2538
rect 6223 2402 6253 2534
rect 6574 2402 6604 2538
rect 9433 2402 9463 2534
rect 9784 2402 9814 2538
rect 12643 2402 12673 2534
rect 12994 2402 13024 2538
rect 15853 2410 15883 2534
rect 15354 2402 16043 2410
rect 3243 2380 16043 2402
rect 3243 2372 15375 2380
rect 3177 159 3246 189
rect 3364 36 3394 2372
rect 4459 1249 4529 1323
rect 5095 1247 5165 1321
rect 4508 656 4550 707
rect 4949 628 4966 657
rect 5739 304 5805 334
rect 3815 159 3881 189
rect 6223 32 6253 2372
rect 6399 189 6470 190
rect 6387 160 6470 189
rect 6387 159 6464 160
rect 6393 157 6464 159
rect 6574 36 6604 2372
rect 7665 1254 7735 1328
rect 8309 1256 8379 1330
rect 7718 656 7760 707
rect 8159 628 8176 657
rect 8949 304 9015 334
rect 7025 159 7091 189
rect 9433 32 9463 2372
rect 9602 189 9673 192
rect 9597 162 9673 189
rect 9597 159 9669 162
rect 9784 36 9814 2372
rect 10882 1256 10952 1330
rect 11490 1232 11607 1336
rect 10928 656 10970 707
rect 11369 627 11386 656
rect 12159 304 12225 334
rect 10235 159 10301 189
rect 12643 32 12673 2372
rect 12816 189 12887 190
rect 12807 160 12887 189
rect 12807 159 12882 160
rect 12994 36 13024 2372
rect 14089 1256 14159 1330
rect 14734 1249 14804 1323
rect 14138 656 14180 707
rect 14583 627 14600 656
rect 15369 304 15435 334
rect 13445 159 13511 189
rect 15853 32 15883 2380
rect 16017 159 16050 189
<< metal4 >>
rect 90 2478 120 2535
rect 234 2478 264 2535
rect 378 2478 408 2535
rect 522 2478 552 2535
rect 33 2448 2535 2478
rect 90 2334 120 2448
rect 234 2334 264 2448
rect 378 2334 408 2448
rect 522 2334 552 2448
rect 33 2304 2535 2334
rect 90 2190 120 2304
rect 234 2190 264 2304
rect 378 2190 408 2304
rect 522 2190 552 2304
rect 33 2160 2535 2190
rect 90 2046 120 2160
rect 234 2046 264 2160
rect 378 2046 408 2160
rect 522 2046 552 2160
rect 33 2016 2535 2046
rect 2 90 73 120
rect 90 33 120 2016
rect 234 33 264 2016
rect 378 33 408 2016
rect 522 33 552 2016
rect 732 1836 762 1926
rect 876 1836 906 1926
rect 1020 1836 1050 1926
rect 1164 1836 1194 1926
rect 1374 1836 1404 1926
rect 1518 1836 1548 1926
rect 1662 1836 1692 1926
rect 1806 1836 1836 1926
rect 2016 1836 2046 1926
rect 2160 1836 2190 1926
rect 2304 1836 2334 1926
rect 2448 1836 2478 1926
rect 642 1806 2568 1836
rect 732 1692 762 1806
rect 876 1692 906 1806
rect 1020 1692 1050 1806
rect 1164 1692 1194 1806
rect 1374 1692 1404 1806
rect 1518 1692 1548 1806
rect 1662 1692 1692 1806
rect 1806 1692 1836 1806
rect 2016 1692 2046 1806
rect 2160 1692 2190 1806
rect 2304 1692 2334 1806
rect 2448 1692 2478 1806
rect 642 1662 2568 1692
rect 732 1548 762 1662
rect 876 1548 906 1662
rect 1020 1548 1050 1662
rect 1164 1548 1194 1662
rect 1374 1548 1404 1662
rect 1518 1548 1548 1662
rect 1662 1548 1692 1662
rect 1806 1548 1836 1662
rect 2016 1548 2046 1662
rect 2160 1548 2190 1662
rect 2304 1548 2334 1662
rect 2448 1548 2478 1662
rect 642 1518 2568 1548
rect 732 1404 762 1518
rect 876 1404 906 1518
rect 1020 1404 1050 1518
rect 1164 1404 1194 1518
rect 1374 1404 1404 1518
rect 1518 1404 1548 1518
rect 1662 1404 1692 1518
rect 1806 1404 1836 1518
rect 2016 1404 2046 1518
rect 2160 1404 2190 1518
rect 2304 1404 2334 1518
rect 2448 1404 2478 1518
rect 642 1374 2568 1404
rect 732 1194 762 1374
rect 876 1194 906 1374
rect 1020 1194 1050 1374
rect 1164 1194 1194 1374
rect 1374 1194 1404 1374
rect 1518 1194 1548 1374
rect 1662 1194 1692 1374
rect 1806 1194 1836 1374
rect 2016 1194 2046 1374
rect 2160 1194 2190 1374
rect 2304 1194 2334 1374
rect 2448 1194 2478 1374
rect 642 1164 2568 1194
rect 732 1050 762 1164
rect 876 1050 906 1164
rect 1020 1050 1050 1164
rect 1164 1050 1194 1164
rect 1374 1050 1404 1164
rect 1518 1050 1548 1164
rect 1662 1050 1692 1164
rect 1806 1050 1836 1164
rect 2016 1050 2046 1164
rect 2160 1050 2190 1164
rect 2304 1050 2334 1164
rect 2448 1050 2478 1164
rect 642 1020 2568 1050
rect 732 906 762 1020
rect 876 906 906 1020
rect 1020 906 1050 1020
rect 1164 906 1194 1020
rect 1374 906 1404 1020
rect 1518 906 1548 1020
rect 1662 906 1692 1020
rect 1806 906 1836 1020
rect 2016 906 2046 1020
rect 2160 906 2190 1020
rect 2304 906 2334 1020
rect 2448 906 2478 1020
rect 642 876 2568 906
rect 732 762 762 876
rect 876 762 906 876
rect 1020 762 1050 876
rect 1164 762 1194 876
rect 1374 762 1404 876
rect 1518 762 1548 876
rect 1662 762 1692 876
rect 1806 762 1836 876
rect 2016 762 2046 876
rect 2160 762 2190 876
rect 2304 762 2334 876
rect 2448 762 2478 876
rect 642 732 2568 762
rect 732 642 762 732
rect 876 643 906 732
rect 1020 642 1050 732
rect 1164 643 1194 732
rect 1374 642 1404 732
rect 1518 642 1548 732
rect 1662 642 1692 732
rect 1806 642 1836 732
rect 2016 642 2046 732
rect 2160 642 2190 732
rect 2304 642 2334 732
rect 2448 643 2478 732
rect 609 522 675 552
rect 1178 521 2049 552
rect 2535 522 2604 552
rect 609 378 675 408
rect 1178 377 2049 408
rect 2535 378 2604 408
rect 609 234 675 264
rect 1181 232 2052 263
rect 2535 234 2604 264
rect 609 90 675 120
rect 1141 90 2012 121
rect 2535 90 2604 120
rect 2658 33 2688 2535
rect 2802 33 2832 2535
rect 2946 33 2976 2535
rect 3090 33 3120 2535
rect 3300 2478 3330 2535
rect 3444 2478 3474 2535
rect 3588 2478 3618 2535
rect 3732 2478 3762 2535
rect 5868 2478 5898 2535
rect 6012 2478 6042 2535
rect 6156 2478 6186 2535
rect 6300 2478 6330 2535
rect 6510 2478 6540 2535
rect 6654 2478 6684 2535
rect 6798 2478 6828 2535
rect 6942 2478 6972 2535
rect 9078 2478 9108 2535
rect 9222 2478 9252 2535
rect 9366 2478 9396 2535
rect 9510 2478 9540 2535
rect 9720 2478 9750 2535
rect 9864 2478 9894 2535
rect 10008 2478 10038 2535
rect 10152 2478 10182 2535
rect 12288 2478 12318 2535
rect 12432 2478 12462 2535
rect 12576 2478 12606 2535
rect 12720 2478 12750 2535
rect 12930 2478 12960 2535
rect 13074 2478 13104 2535
rect 13218 2478 13248 2535
rect 13362 2478 13392 2535
rect 15498 2478 15528 2535
rect 15642 2478 15672 2535
rect 15786 2478 15816 2535
rect 15930 2478 15960 2535
rect 3243 2448 16031 2478
rect 3300 2334 3330 2448
rect 3444 2334 3474 2448
rect 3588 2334 3618 2448
rect 3732 2334 3762 2448
rect 5868 2334 5898 2448
rect 6012 2334 6042 2448
rect 6156 2334 6186 2448
rect 6300 2334 6330 2448
rect 6510 2334 6540 2448
rect 6654 2334 6684 2448
rect 6798 2334 6828 2448
rect 6942 2334 6972 2448
rect 9078 2334 9108 2448
rect 9222 2334 9252 2448
rect 9366 2334 9396 2448
rect 9510 2334 9540 2448
rect 9720 2334 9750 2448
rect 9864 2334 9894 2448
rect 10008 2334 10038 2448
rect 10152 2334 10182 2448
rect 12288 2334 12318 2448
rect 12432 2334 12462 2448
rect 12576 2334 12606 2448
rect 12720 2334 12750 2448
rect 12930 2334 12960 2448
rect 13074 2334 13104 2448
rect 13218 2334 13248 2448
rect 13362 2334 13392 2448
rect 15498 2334 15528 2448
rect 15642 2334 15672 2448
rect 15786 2334 15816 2448
rect 15930 2334 15960 2448
rect 3243 2304 16035 2334
rect 3300 2190 3330 2304
rect 3444 2190 3474 2304
rect 3588 2190 3618 2304
rect 3732 2190 3762 2304
rect 5868 2190 5898 2304
rect 6012 2190 6042 2304
rect 6156 2190 6186 2304
rect 6300 2190 6330 2304
rect 6510 2190 6540 2304
rect 6654 2190 6684 2304
rect 6798 2190 6828 2304
rect 6942 2190 6972 2304
rect 9078 2190 9108 2304
rect 9222 2190 9252 2304
rect 9366 2190 9396 2304
rect 9510 2190 9540 2304
rect 9720 2190 9750 2304
rect 9864 2190 9894 2304
rect 10008 2190 10038 2304
rect 10152 2190 10182 2304
rect 12288 2190 12318 2304
rect 12432 2190 12462 2304
rect 12576 2190 12606 2304
rect 12720 2190 12750 2304
rect 12930 2190 12960 2304
rect 13074 2190 13104 2304
rect 13218 2190 13248 2304
rect 13362 2190 13392 2304
rect 15498 2190 15528 2304
rect 15642 2190 15672 2304
rect 15786 2190 15816 2304
rect 15930 2190 15960 2304
rect 3243 2160 16031 2190
rect 3300 2046 3330 2160
rect 3444 2046 3474 2160
rect 3588 2046 3618 2160
rect 3732 2046 3762 2160
rect 5868 2046 5898 2160
rect 6012 2046 6042 2160
rect 6156 2046 6186 2160
rect 6300 2046 6330 2160
rect 6510 2046 6540 2160
rect 6654 2046 6684 2160
rect 6798 2046 6828 2160
rect 6942 2046 6972 2160
rect 9078 2046 9108 2160
rect 9222 2046 9252 2160
rect 9366 2046 9396 2160
rect 9510 2046 9540 2160
rect 9720 2046 9750 2160
rect 9864 2046 9894 2160
rect 10008 2046 10038 2160
rect 10152 2046 10182 2160
rect 12288 2046 12318 2160
rect 12432 2046 12462 2160
rect 12576 2046 12606 2160
rect 12720 2046 12750 2160
rect 12930 2046 12960 2160
rect 13074 2046 13104 2160
rect 13218 2046 13248 2160
rect 13362 2046 13392 2160
rect 15498 2046 15528 2160
rect 15642 2046 15672 2160
rect 15786 2046 15816 2160
rect 15930 2046 15960 2160
rect 3243 2016 16029 2046
rect 3177 90 3253 120
rect 3300 33 3330 2016
rect 3444 33 3474 2016
rect 3588 33 3618 2016
rect 3732 33 3762 2016
rect 3942 1836 3972 1926
rect 4086 1836 4116 1926
rect 4230 1836 4260 1926
rect 4374 1836 4404 1926
rect 4584 1836 4614 1926
rect 4728 1836 4758 1926
rect 4872 1836 4902 1926
rect 5016 1836 5046 1926
rect 5226 1836 5256 1926
rect 5370 1836 5400 1926
rect 5514 1836 5544 1926
rect 5658 1836 5688 1926
rect 3852 1806 5778 1836
rect 3942 1692 3972 1806
rect 4086 1692 4116 1806
rect 4230 1692 4260 1806
rect 4374 1692 4404 1806
rect 4584 1692 4614 1806
rect 4728 1692 4758 1806
rect 4872 1692 4902 1806
rect 5016 1692 5046 1806
rect 5226 1692 5256 1806
rect 5370 1692 5400 1806
rect 5514 1692 5544 1806
rect 5658 1692 5688 1806
rect 3852 1662 5778 1692
rect 3942 1548 3972 1662
rect 4086 1548 4116 1662
rect 4230 1548 4260 1662
rect 4374 1548 4404 1662
rect 4584 1548 4614 1662
rect 4728 1548 4758 1662
rect 4872 1548 4902 1662
rect 5016 1548 5046 1662
rect 5226 1548 5256 1662
rect 5370 1548 5400 1662
rect 5514 1548 5544 1662
rect 5658 1548 5688 1662
rect 3852 1518 5778 1548
rect 3942 1404 3972 1518
rect 4086 1404 4116 1518
rect 4230 1404 4260 1518
rect 4374 1404 4404 1518
rect 4584 1404 4614 1518
rect 4728 1404 4758 1518
rect 4872 1404 4902 1518
rect 5016 1404 5046 1518
rect 5226 1404 5256 1518
rect 5370 1404 5400 1518
rect 5514 1404 5544 1518
rect 5658 1404 5688 1518
rect 3852 1374 5778 1404
rect 3942 1194 3972 1374
rect 4086 1194 4116 1374
rect 4230 1194 4260 1374
rect 4374 1194 4404 1374
rect 4584 1194 4614 1374
rect 4728 1194 4758 1374
rect 4872 1194 4902 1374
rect 5016 1194 5046 1374
rect 5226 1194 5256 1374
rect 5370 1194 5400 1374
rect 5514 1194 5544 1374
rect 5658 1194 5688 1374
rect 3852 1164 5778 1194
rect 3942 1050 3972 1164
rect 4086 1050 4116 1164
rect 4230 1050 4260 1164
rect 4374 1050 4404 1164
rect 4584 1050 4614 1164
rect 4728 1050 4758 1164
rect 4872 1050 4902 1164
rect 5016 1050 5046 1164
rect 5226 1050 5256 1164
rect 5370 1050 5400 1164
rect 5514 1050 5544 1164
rect 5658 1050 5688 1164
rect 3852 1020 5778 1050
rect 3942 906 3972 1020
rect 4086 906 4116 1020
rect 4230 906 4260 1020
rect 4374 906 4404 1020
rect 4584 906 4614 1020
rect 4728 906 4758 1020
rect 4872 906 4902 1020
rect 5016 906 5046 1020
rect 5226 906 5256 1020
rect 5370 906 5400 1020
rect 5514 906 5544 1020
rect 5658 906 5688 1020
rect 3852 876 5778 906
rect 3942 762 3972 876
rect 4086 762 4116 876
rect 4230 762 4260 876
rect 4374 762 4404 876
rect 4584 762 4614 876
rect 4728 762 4758 876
rect 4872 762 4902 876
rect 5016 762 5046 876
rect 5226 762 5256 876
rect 5370 762 5400 876
rect 5514 762 5544 876
rect 5658 762 5688 876
rect 3852 732 5778 762
rect 3942 642 3972 732
rect 4086 643 4116 732
rect 4230 642 4260 732
rect 4374 643 4404 732
rect 4584 609 4614 732
rect 4728 609 4758 732
rect 4872 609 4902 732
rect 5016 609 5046 732
rect 5226 642 5256 732
rect 5370 642 5400 732
rect 5514 642 5544 732
rect 5658 643 5688 732
rect 3819 522 3885 552
rect 4494 522 4527 552
rect 5103 522 5136 552
rect 5745 522 5814 552
rect 3819 378 3885 408
rect 4494 378 4527 408
rect 5103 378 5136 408
rect 5745 378 5814 408
rect 3819 234 3885 264
rect 5745 234 5814 264
rect 3819 90 3885 120
rect 5745 90 5814 120
rect 4584 51 4611 74
rect 5868 33 5898 2016
rect 6012 33 6042 2016
rect 6156 33 6186 2016
rect 6300 33 6330 2016
rect 6387 90 6470 120
rect 6510 33 6540 2016
rect 6654 33 6684 2016
rect 6798 33 6828 2016
rect 6942 33 6972 2016
rect 7152 1836 7182 1926
rect 7296 1836 7326 1926
rect 7440 1836 7470 1926
rect 7584 1836 7614 1926
rect 7794 1836 7824 1926
rect 7938 1836 7968 1926
rect 8082 1836 8112 1926
rect 8226 1836 8256 1926
rect 8436 1836 8466 1926
rect 8580 1836 8610 1926
rect 8724 1836 8754 1926
rect 8868 1836 8898 1926
rect 7062 1806 8988 1836
rect 7152 1692 7182 1806
rect 7296 1692 7326 1806
rect 7440 1692 7470 1806
rect 7584 1692 7614 1806
rect 7794 1692 7824 1806
rect 7938 1692 7968 1806
rect 8082 1692 8112 1806
rect 8226 1692 8256 1806
rect 8436 1692 8466 1806
rect 8580 1692 8610 1806
rect 8724 1692 8754 1806
rect 8868 1692 8898 1806
rect 7062 1662 8988 1692
rect 7152 1548 7182 1662
rect 7296 1548 7326 1662
rect 7440 1548 7470 1662
rect 7584 1548 7614 1662
rect 7794 1548 7824 1662
rect 7938 1548 7968 1662
rect 8082 1548 8112 1662
rect 8226 1548 8256 1662
rect 8436 1548 8466 1662
rect 8580 1548 8610 1662
rect 8724 1548 8754 1662
rect 8868 1548 8898 1662
rect 7062 1518 8988 1548
rect 7152 1404 7182 1518
rect 7296 1404 7326 1518
rect 7440 1404 7470 1518
rect 7584 1404 7614 1518
rect 7794 1404 7824 1518
rect 7938 1404 7968 1518
rect 8082 1404 8112 1518
rect 8226 1404 8256 1518
rect 8436 1404 8466 1518
rect 8580 1404 8610 1518
rect 8724 1404 8754 1518
rect 8868 1404 8898 1518
rect 7062 1374 8988 1404
rect 7152 1194 7182 1374
rect 7296 1194 7326 1374
rect 7440 1194 7470 1374
rect 7584 1194 7614 1374
rect 7794 1194 7824 1374
rect 7938 1194 7968 1374
rect 8082 1194 8112 1374
rect 8226 1194 8256 1374
rect 8436 1194 8466 1374
rect 8580 1194 8610 1374
rect 8724 1194 8754 1374
rect 8868 1194 8898 1374
rect 7062 1164 8988 1194
rect 7152 1050 7182 1164
rect 7296 1050 7326 1164
rect 7440 1050 7470 1164
rect 7584 1050 7614 1164
rect 7794 1050 7824 1164
rect 7938 1050 7968 1164
rect 8082 1050 8112 1164
rect 8226 1050 8256 1164
rect 8436 1050 8466 1164
rect 8580 1050 8610 1164
rect 8724 1050 8754 1164
rect 8868 1050 8898 1164
rect 7062 1020 8988 1050
rect 7152 906 7182 1020
rect 7296 906 7326 1020
rect 7440 906 7470 1020
rect 7584 906 7614 1020
rect 7794 906 7824 1020
rect 7938 906 7968 1020
rect 8082 906 8112 1020
rect 8226 906 8256 1020
rect 8436 906 8466 1020
rect 8580 906 8610 1020
rect 8724 906 8754 1020
rect 8868 906 8898 1020
rect 7062 876 8988 906
rect 7152 762 7182 876
rect 7296 762 7326 876
rect 7440 762 7470 876
rect 7584 762 7614 876
rect 7794 762 7824 876
rect 7938 762 7968 876
rect 8082 762 8112 876
rect 8226 762 8256 876
rect 8436 762 8466 876
rect 8580 762 8610 876
rect 8724 762 8754 876
rect 8868 762 8898 876
rect 7062 732 8988 762
rect 7152 642 7182 732
rect 7296 643 7326 732
rect 7440 642 7470 732
rect 7584 643 7614 732
rect 7794 590 7824 732
rect 7938 593 7968 732
rect 8082 642 8112 732
rect 8226 642 8256 732
rect 8436 642 8466 732
rect 8580 642 8610 732
rect 8724 642 8754 732
rect 8868 643 8898 732
rect 7029 522 7095 552
rect 7704 522 7737 552
rect 8955 522 9024 552
rect 7029 378 7095 408
rect 7704 378 7737 408
rect 8955 378 9024 408
rect 7029 234 7095 264
rect 8955 234 9024 264
rect 7029 90 7095 120
rect 8955 90 9024 120
rect 7794 52 7812 76
rect 9078 33 9108 2016
rect 9222 33 9252 2016
rect 9366 33 9396 2016
rect 9510 33 9540 2016
rect 9597 90 9674 120
rect 9720 33 9750 2016
rect 9864 33 9894 2016
rect 10008 33 10038 2016
rect 10152 33 10182 2016
rect 10362 1836 10392 1926
rect 10506 1836 10536 1926
rect 10650 1836 10680 1926
rect 10794 1836 10824 1926
rect 11004 1836 11034 1926
rect 11148 1836 11178 1926
rect 11292 1836 11322 1926
rect 11436 1836 11466 1926
rect 11646 1836 11676 1926
rect 11790 1836 11820 1926
rect 11934 1836 11964 1926
rect 12078 1836 12108 1926
rect 10272 1806 12198 1836
rect 10362 1692 10392 1806
rect 10506 1692 10536 1806
rect 10650 1692 10680 1806
rect 10794 1692 10824 1806
rect 11004 1692 11034 1806
rect 11148 1692 11178 1806
rect 11292 1692 11322 1806
rect 11436 1692 11466 1806
rect 11646 1692 11676 1806
rect 11790 1692 11820 1806
rect 11934 1692 11964 1806
rect 12078 1692 12108 1806
rect 10272 1662 12198 1692
rect 10362 1548 10392 1662
rect 10506 1548 10536 1662
rect 10650 1548 10680 1662
rect 10794 1548 10824 1662
rect 11004 1548 11034 1662
rect 11148 1548 11178 1662
rect 11292 1548 11322 1662
rect 11436 1548 11466 1662
rect 11646 1548 11676 1662
rect 11790 1548 11820 1662
rect 11934 1548 11964 1662
rect 12078 1548 12108 1662
rect 10272 1518 12198 1548
rect 10362 1404 10392 1518
rect 10506 1404 10536 1518
rect 10650 1404 10680 1518
rect 10794 1404 10824 1518
rect 11004 1404 11034 1518
rect 11148 1404 11178 1518
rect 11292 1404 11322 1518
rect 11436 1404 11466 1518
rect 11646 1404 11676 1518
rect 11790 1404 11820 1518
rect 11934 1404 11964 1518
rect 12078 1404 12108 1518
rect 10272 1374 12198 1404
rect 10362 1194 10392 1374
rect 10506 1194 10536 1374
rect 10650 1194 10680 1374
rect 10794 1194 10824 1374
rect 11004 1194 11034 1374
rect 11148 1194 11178 1374
rect 11292 1194 11322 1374
rect 11436 1194 11466 1374
rect 11646 1194 11676 1374
rect 11790 1194 11820 1374
rect 11934 1194 11964 1374
rect 12078 1194 12108 1374
rect 10272 1164 12198 1194
rect 10362 1050 10392 1164
rect 10506 1050 10536 1164
rect 10650 1050 10680 1164
rect 10794 1050 10824 1164
rect 11004 1050 11034 1164
rect 11148 1050 11178 1164
rect 11292 1050 11322 1164
rect 11436 1050 11466 1164
rect 11646 1050 11676 1164
rect 11790 1050 11820 1164
rect 11934 1050 11964 1164
rect 12078 1050 12108 1164
rect 10272 1020 12198 1050
rect 10362 906 10392 1020
rect 10506 906 10536 1020
rect 10650 906 10680 1020
rect 10794 906 10824 1020
rect 11004 906 11034 1020
rect 11148 906 11178 1020
rect 11292 906 11322 1020
rect 11436 906 11466 1020
rect 11646 906 11676 1020
rect 11790 906 11820 1020
rect 11934 906 11964 1020
rect 12078 906 12108 1020
rect 10272 876 12198 906
rect 10362 762 10392 876
rect 10506 762 10536 876
rect 10650 762 10680 876
rect 10794 762 10824 876
rect 11004 762 11034 876
rect 11148 762 11178 876
rect 11292 762 11322 876
rect 11436 762 11466 876
rect 11646 762 11676 876
rect 11790 762 11820 876
rect 11934 762 11964 876
rect 12078 762 12108 876
rect 10272 732 12198 762
rect 10362 642 10392 732
rect 10506 643 10536 732
rect 10650 642 10680 732
rect 10794 643 10824 732
rect 11004 642 11034 732
rect 11148 586 11178 732
rect 11292 596 11322 732
rect 11436 642 11466 732
rect 11646 642 11676 732
rect 11790 642 11820 732
rect 11934 642 11964 732
rect 12078 643 12108 732
rect 10239 522 10305 552
rect 12165 522 12234 552
rect 10239 378 10305 408
rect 12165 378 12234 408
rect 10239 234 10305 264
rect 12165 234 12234 264
rect 10239 90 10305 120
rect 12165 90 12234 120
rect 11004 55 11026 78
rect 12288 33 12318 2016
rect 12432 33 12462 2016
rect 12576 33 12606 2016
rect 12720 33 12750 2016
rect 12807 90 12890 120
rect 12930 33 12960 2016
rect 13074 33 13104 2016
rect 13218 33 13248 2016
rect 13362 33 13392 2016
rect 13572 1836 13602 1926
rect 13716 1836 13746 1926
rect 13860 1836 13890 1926
rect 14004 1836 14034 1926
rect 14214 1836 14244 1926
rect 14358 1836 14388 1926
rect 14502 1836 14532 1926
rect 14646 1836 14676 1926
rect 14856 1836 14886 1926
rect 15000 1836 15030 1926
rect 15144 1836 15174 1926
rect 15288 1836 15318 1926
rect 13482 1806 15408 1836
rect 13572 1692 13602 1806
rect 13716 1692 13746 1806
rect 13860 1692 13890 1806
rect 14004 1692 14034 1806
rect 14214 1692 14244 1806
rect 14358 1692 14388 1806
rect 14502 1692 14532 1806
rect 14646 1692 14676 1806
rect 14856 1692 14886 1806
rect 15000 1692 15030 1806
rect 15144 1692 15174 1806
rect 15288 1692 15318 1806
rect 13482 1662 15408 1692
rect 13572 1548 13602 1662
rect 13716 1548 13746 1662
rect 13860 1548 13890 1662
rect 14004 1548 14034 1662
rect 14214 1548 14244 1662
rect 14358 1548 14388 1662
rect 14502 1548 14532 1662
rect 14646 1548 14676 1662
rect 14856 1548 14886 1662
rect 15000 1548 15030 1662
rect 15144 1548 15174 1662
rect 15288 1548 15318 1662
rect 13482 1518 15408 1548
rect 13572 1404 13602 1518
rect 13716 1404 13746 1518
rect 13860 1404 13890 1518
rect 14004 1404 14034 1518
rect 14214 1404 14244 1518
rect 14358 1404 14388 1518
rect 14502 1404 14532 1518
rect 14646 1404 14676 1518
rect 14856 1404 14886 1518
rect 15000 1404 15030 1518
rect 15144 1404 15174 1518
rect 15288 1404 15318 1518
rect 13482 1374 15408 1404
rect 13572 1194 13602 1374
rect 13716 1194 13746 1374
rect 13860 1194 13890 1374
rect 14004 1194 14034 1374
rect 14214 1194 14244 1374
rect 14358 1194 14388 1374
rect 14502 1194 14532 1374
rect 14646 1194 14676 1374
rect 14856 1194 14886 1374
rect 15000 1194 15030 1374
rect 15144 1194 15174 1374
rect 15288 1194 15318 1374
rect 13482 1164 15408 1194
rect 13572 1050 13602 1164
rect 13716 1050 13746 1164
rect 13860 1050 13890 1164
rect 14004 1050 14034 1164
rect 14214 1050 14244 1164
rect 14358 1050 14388 1164
rect 14502 1050 14532 1164
rect 14646 1050 14676 1164
rect 14856 1050 14886 1164
rect 15000 1050 15030 1164
rect 15144 1050 15174 1164
rect 15288 1050 15318 1164
rect 13482 1020 15408 1050
rect 13572 906 13602 1020
rect 13716 906 13746 1020
rect 13860 906 13890 1020
rect 14004 906 14034 1020
rect 14214 906 14244 1020
rect 14358 906 14388 1020
rect 14502 906 14532 1020
rect 14646 906 14676 1020
rect 14856 906 14886 1020
rect 15000 906 15030 1020
rect 15144 906 15174 1020
rect 15288 906 15318 1020
rect 13482 876 15408 906
rect 13572 762 13602 876
rect 13716 762 13746 876
rect 13860 762 13890 876
rect 14004 762 14034 876
rect 14214 762 14244 876
rect 14358 762 14388 876
rect 14502 762 14532 876
rect 14646 762 14676 876
rect 14856 762 14886 876
rect 15000 762 15030 876
rect 15144 762 15174 876
rect 15288 762 15318 876
rect 13482 732 15408 762
rect 13572 642 13602 732
rect 13716 643 13746 732
rect 13860 642 13890 732
rect 14004 643 14034 732
rect 14214 642 14244 732
rect 14358 587 14388 732
rect 14502 642 14532 732
rect 14646 642 14676 732
rect 14856 642 14886 732
rect 15000 642 15030 732
rect 15144 642 15174 732
rect 15288 643 15318 732
rect 13449 522 13515 552
rect 15375 522 15444 552
rect 13449 378 13515 408
rect 15375 378 15444 408
rect 13449 234 13515 264
rect 15375 234 15444 264
rect 13449 90 13515 120
rect 15375 90 15444 120
rect 14214 55 14242 78
rect 15498 33 15528 2016
rect 15642 33 15672 2016
rect 15786 33 15816 2016
rect 15930 33 15960 2016
rect 16017 90 16050 120
use adc_array_wafflecap_16(1)_41um2  adc_array_wafflecap_16(1)_41um2_0
timestamp 1659692885
transform 1 0 14124 0 1 0
box 0 0 642 642
use adc_array_wafflecap_16(2)_41um2  adc_array_wafflecap_16(2)_41um2_0
timestamp 1659692910
transform 1 0 10914 0 1 0
box 0 0 642 642
use adc_array_wafflecap_16(4)_41um2  adc_array_wafflecap_16(4)_41um2_0
timestamp 1659692964
transform 1 0 7704 0 1 0
box 0 0 642 642
use adc_array_wafflecap_16(8)_41um2  adc_array_wafflecap_16(8)_41um2_0
timestamp 1659692976
transform 1 0 4494 0 1 0
box 0 0 642 642
use adc_array_wafflecap_16(16)_41um2  adc_array_wafflecap_16(16)_41um2_0
array 0 4 3210 0 0 2568
timestamp 1659692990
transform 1 0 0 0 1 0
box 0 0 642 642
use adc_array_wafflecap_16(16)_41um2  adc_array_wafflecap_16(16)_41um2_1
array 0 4 3210 0 0 2568
timestamp 1659692990
transform 1 0 0 0 1 642
box 0 0 642 642
use adc_array_wafflecap_16(16)_41um2  adc_array_wafflecap_16(16)_41um2_2
array 0 4 3210 0 0 2568
timestamp 1659692990
transform 1 0 0 0 1 1284
box 0 0 642 642
use adc_array_wafflecap_16(16)_41um2  adc_array_wafflecap_16(16)_41um2_3
array 0 4 3210 0 0 2568
timestamp 1659692990
transform 1 0 0 0 1 1926
box 0 0 642 642
use adc_array_wafflecap_16(16)_41um2  adc_array_wafflecap_16(16)_41um2_4
array 0 4 3210 0 0 2568
timestamp 1659692990
transform 1 0 642 0 1 1926
box 0 0 642 642
use adc_array_wafflecap_16(16)_41um2  adc_array_wafflecap_16(16)_41um2_5
array 0 4 3210 0 0 2568
timestamp 1659692990
transform 1 0 1284 0 1 1926
box 0 0 642 642
use adc_array_wafflecap_16(16)_41um2  adc_array_wafflecap_16(16)_41um2_6
array 0 4 3210 0 0 2568
timestamp 1659692990
transform 1 0 1926 0 1 1926
box 0 0 642 642
use adc_array_wafflecap_16(16)_41um2  adc_array_wafflecap_16(16)_41um2_7
array 0 4 3210 0 0 2568
timestamp 1659692990
transform 1 0 2568 0 1 1926
box 0 0 642 642
use adc_array_wafflecap_16(16)_41um2  adc_array_wafflecap_16(16)_41um2_8
array 0 4 3210 0 0 2568
timestamp 1659692990
transform 1 0 2568 0 1 1284
box 0 0 642 642
use adc_array_wafflecap_16(16)_41um2  adc_array_wafflecap_16(16)_41um2_9
array 0 4 3210 0 0 2568
timestamp 1659692990
transform 1 0 2568 0 1 642
box 0 0 642 642
use adc_array_wafflecap_16(16)_41um2  adc_array_wafflecap_16(16)_41um2_10
array 0 4 3210 0 0 2568
timestamp 1659692990
transform 1 0 2568 0 1 0
box 0 0 642 642
use adc_array_wafflecap_16(16)_41um2  adc_array_wafflecap_16(16)_41um2_11
array 0 4 3210 0 0 2568
timestamp 1659692990
transform 1 0 642 0 1 1284
box 0 0 642 642
use adc_array_wafflecap_16(16)_41um2  adc_array_wafflecap_16(16)_41um2_12
array 0 4 3210 0 0 2568
timestamp 1659692990
transform 1 0 1284 0 1 1284
box 0 0 642 642
use adc_array_wafflecap_16(16)_41um2  adc_array_wafflecap_16(16)_41um2_13
array 0 4 3210 0 0 2568
timestamp 1659692990
transform 1 0 1926 0 1 1284
box 0 0 642 642
use adc_array_wafflecap_16(16)_41um2  adc_array_wafflecap_16(16)_41um2_14
array 0 4 3210 0 0 2568
timestamp 1659692990
transform 1 0 642 0 1 642
box 0 0 642 642
use adc_array_wafflecap_16(16)_41um2  adc_array_wafflecap_16(16)_41um2_15
array 0 4 3210 0 0 2568
timestamp 1659692990
transform 1 0 1284 0 1 642
box 0 0 642 642
use adc_array_wafflecap_16(16)_41um2  adc_array_wafflecap_16(16)_41um2_16
array 0 4 3210 0 0 2568
timestamp 1659692990
transform 1 0 1926 0 1 642
box 0 0 642 642
use adc_array_wafflecap_16(16)_41um2  adc_array_wafflecap_16(16)_41um2_17
array 0 4 3210 0 0 2568
timestamp 1659692990
transform 1 0 642 0 1 0
box 0 0 642 642
use adc_array_wafflecap_16(16)_41um2  adc_array_wafflecap_16(16)_41um2_18
array 0 4 3210 0 0 2568
timestamp 1659692990
transform 1 0 1926 0 1 0
box 0 0 642 642
use adc_array_wafflecap_16(16)_41um2  adc_array_wafflecap_16(16)_41um2_19
timestamp 1659692990
transform 1 0 1284 0 1 0
box 0 0 642 642
<< labels >>
rlabel metal4 2 90 2 120 7 ctop_dummy
rlabel metal2 1 139 1 169 7 cdummy_bot
rlabel metal4 14358 632 14358 650 7 ctop_1
rlabel metal2 14138 662 14138 680 7 cbot_1
rlabel metal4 11148 634 11148 652 7 ctop_2
rlabel metal2 10928 667 10928 685 7 cbot_2
rlabel metal4 7938 633 7938 651 7 ctop_4
rlabel metal2 7718 671 7718 689 7 cbot_4
rlabel metal4 4584 633 4584 651 7 ctop_8
rlabel metal4 876 646 876 664 7 ctop_16
rlabel metal2 656 676 656 694 7 cbot_16
rlabel metal4 14214 55 14214 75 7 ctop_1_floating
rlabel metal4 11004 57 11004 75 7 ctop_2_floating
rlabel metal4 7794 56 7794 74 7 ctop_4_floating
rlabel metal4 4584 53 4584 71 7 ctop_8_floating
rlabel metal2 4508 670 4508 695 7 cbot_8
<< end >>
