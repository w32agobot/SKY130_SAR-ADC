* NGSPICE file created from adc_array_wafflecap_8_Gate_25um2.ext - technology: sky130A


* Top level circuit adc_array_wafflecap_8_Gate_25um2

.end

