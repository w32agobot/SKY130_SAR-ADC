magic
tech sky130A
timestamp 1661165658
<< checkpaint >>
rect -564 -660 1250 1322
<< metal2 >>
rect 163 590 579 608
rect 163 559 348 590
rect 394 559 579 590
rect 163 465 579 559
rect 163 434 348 465
rect 394 434 579 465
rect 163 341 579 434
rect 163 310 348 341
rect 394 310 579 341
rect 163 217 579 310
rect 163 186 348 217
rect 394 186 579 217
rect 163 93 579 186
rect 163 62 348 93
rect 394 62 579 93
rect 163 43 579 62
<< via2 >>
rect 348 559 394 590
rect 348 434 394 465
rect 348 310 394 341
rect 348 186 394 217
rect 348 62 394 93
<< metal3 >>
rect 343 590 399 593
rect 343 589 348 590
rect 182 559 348 589
rect 394 589 399 590
rect 394 559 560 589
rect 343 555 399 559
rect 246 527 284 528
rect 246 526 249 527
rect 201 496 249 526
rect 246 495 249 496
rect 281 526 284 527
rect 458 527 496 528
rect 458 526 461 527
rect 281 496 328 526
rect 414 496 461 526
rect 281 495 284 496
rect 246 494 284 495
rect 458 495 461 496
rect 493 526 496 527
rect 493 496 541 526
rect 493 495 496 496
rect 458 494 496 495
rect 343 465 399 468
rect 343 464 348 465
rect 182 434 348 464
rect 394 464 399 465
rect 394 434 560 464
rect 343 430 399 434
rect 246 403 284 404
rect 246 402 249 403
rect 201 372 249 402
rect 246 371 249 372
rect 281 402 284 403
rect 458 403 496 404
rect 458 402 461 403
rect 281 372 328 402
rect 414 372 461 402
rect 281 371 284 372
rect 246 370 284 371
rect 458 371 461 372
rect 493 402 496 403
rect 493 372 541 402
rect 493 371 496 372
rect 458 370 496 371
rect 343 341 399 344
rect 343 340 348 341
rect 182 310 348 340
rect 394 340 399 341
rect 394 310 560 340
rect 343 306 399 310
rect 246 279 284 280
rect 246 278 249 279
rect 201 248 249 278
rect 246 247 249 248
rect 281 278 284 279
rect 458 279 496 280
rect 458 278 461 279
rect 281 248 328 278
rect 414 248 461 278
rect 281 247 284 248
rect 246 246 284 247
rect 458 247 461 248
rect 493 278 496 279
rect 493 248 541 278
rect 493 247 496 248
rect 458 246 496 247
rect 343 217 399 220
rect 343 216 348 217
rect 182 186 348 216
rect 394 216 399 217
rect 394 186 560 216
rect 343 182 399 186
rect 246 155 284 156
rect 246 154 249 155
rect 201 124 249 154
rect 246 123 249 124
rect 281 154 284 155
rect 458 155 496 156
rect 458 154 461 155
rect 281 124 328 154
rect 414 124 461 154
rect 281 123 284 124
rect 246 122 284 123
rect 458 123 461 124
rect 493 154 496 155
rect 493 124 541 154
rect 493 123 496 124
rect 458 122 496 123
rect 343 93 399 96
rect 343 92 348 93
rect 182 62 348 92
rect 394 92 399 93
rect 394 62 560 92
rect 343 58 399 62
<< via3 >>
rect 249 495 281 527
rect 461 495 493 527
rect 249 371 281 403
rect 461 371 493 403
rect 249 247 281 279
rect 461 247 493 279
rect 249 123 281 155
rect 461 123 493 155
<< metal4 >>
rect 147 619 595 635
rect 248 528 281 619
rect 461 528 494 619
rect 246 527 284 528
rect 246 526 249 527
rect 201 496 249 526
rect 246 495 249 496
rect 281 526 284 527
rect 458 527 496 528
rect 458 526 461 527
rect 281 496 328 526
rect 414 496 461 526
rect 281 495 284 496
rect 246 494 284 495
rect 458 495 461 496
rect 493 526 496 527
rect 493 496 541 526
rect 493 495 496 496
rect 458 494 496 495
rect 248 404 281 494
rect 461 404 494 494
rect 246 403 284 404
rect 246 402 249 403
rect 201 372 249 402
rect 246 371 249 372
rect 281 402 284 403
rect 458 403 496 404
rect 458 402 461 403
rect 281 372 328 402
rect 414 372 461 402
rect 281 371 284 372
rect 246 370 284 371
rect 458 371 461 372
rect 493 402 496 403
rect 493 372 541 402
rect 493 371 496 372
rect 458 370 496 371
rect 248 280 281 370
rect 461 280 494 370
rect 246 279 284 280
rect 246 278 249 279
rect 201 248 249 278
rect 246 247 249 248
rect 281 278 284 279
rect 458 279 496 280
rect 458 278 461 279
rect 281 248 328 278
rect 414 248 461 278
rect 281 247 284 248
rect 246 246 284 247
rect 458 247 461 248
rect 493 278 496 279
rect 493 248 541 278
rect 493 247 496 248
rect 458 246 496 247
rect 248 156 281 246
rect 461 156 494 246
rect 246 155 284 156
rect 246 154 249 155
rect 201 124 249 154
rect 246 123 249 124
rect 281 154 284 155
rect 458 155 496 156
rect 458 154 461 155
rect 281 124 328 154
rect 414 124 461 154
rect 281 123 284 124
rect 246 122 284 123
rect 458 123 461 124
rect 493 154 496 155
rect 493 124 541 154
rect 493 123 496 124
rect 458 122 496 123
rect 248 32 281 122
rect 461 32 494 122
rect 147 16 595 32
<< comment >>
rect 147 620 163 635
rect 579 620 595 635
rect 147 16 163 31
rect 579 16 595 31
<< end >>
