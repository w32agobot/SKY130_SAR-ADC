magic
tech sky130A
timestamp 1661171482
<< nwell >>
rect 117 152 130 306
<< poly >>
rect 0 129 4 152
<< locali >>
rect 0 129 4 152
rect 230 129 234 152
<< metal1 >>
rect 0 286 5 309
rect 0 0 5 23
use inverter  inverter_0 ../inverter
array 0 1 117 0 0 309
timestamp 1661171367
transform 1 0 13 0 1 63
box -13 -63 104 246
<< labels >>
rlabel metal1 0 286 0 309 7 VDD
port 1 w
rlabel metal1 0 0 0 23 7 VSS
port 2 w
rlabel locali 0 129 0 152 7 in
port 3 w
rlabel locali 234 129 234 152 3 out
port 4 e
<< end >>
