magic
tech sky130A
timestamp 1667211608
<< nwell >>
rect 2986 6600 3045 6804
rect 1367 6361 1549 6406
rect 1344 6349 1549 6361
rect 1344 6220 1372 6349
rect 1427 6294 1549 6349
rect 1421 6275 1549 6294
rect 1427 6220 1549 6275
rect 1344 6207 1549 6220
rect 2985 6028 3125 6230
<< poly >>
rect 3040 6556 3056 6570
rect 3040 6474 3055 6556
rect 3040 6465 3077 6474
rect 3040 6448 3055 6465
rect 3072 6448 3077 6465
rect 3040 6440 3077 6448
rect 2239 6062 2278 6067
rect 2239 6045 2247 6062
rect 2264 6045 2278 6062
rect 2239 6040 2278 6045
<< polycont >>
rect 3055 6448 3072 6465
rect 1339 6187 1356 6204
rect 2247 6045 2264 6062
<< locali >>
rect 1491 6740 1599 6743
rect 1491 6722 1497 6740
rect 1514 6722 1536 6740
rect 1553 6722 1572 6740
rect 1589 6722 1599 6740
rect 1491 6719 1599 6722
rect 1491 6406 1534 6719
rect 3471 6570 3538 6573
rect 3471 6552 3477 6570
rect 3495 6552 3514 6570
rect 3532 6552 3538 6570
rect 3471 6549 3538 6552
rect 1375 6386 1534 6406
rect 3051 6465 3075 6473
rect 3051 6448 3055 6465
rect 3072 6448 3075 6465
rect 3104 6448 3654 6474
rect 1444 6294 1466 6386
rect 1444 6275 1490 6294
rect 3051 6282 3075 6448
rect 3051 6264 3054 6282
rect 3072 6264 3075 6282
rect 1331 6204 1358 6212
rect 1331 6187 1339 6204
rect 1356 6187 1358 6204
rect 1331 6179 1358 6187
rect 1448 6204 1475 6212
rect 1448 6187 1456 6204
rect 1473 6187 1475 6204
rect 1448 6179 1475 6187
rect 3051 6106 3075 6264
rect 3092 6420 3116 6426
rect 3092 6402 3095 6420
rect 3113 6402 3116 6420
rect 3092 6252 3116 6402
rect 3185 6365 3228 6448
rect 3358 6275 3458 6278
rect 3358 6259 3396 6275
rect 3390 6257 3396 6259
rect 3414 6257 3434 6275
rect 3452 6257 3458 6275
rect 3390 6254 3458 6257
rect 3092 6234 3095 6252
rect 3113 6234 3116 6252
rect 3092 6228 3116 6234
rect 3051 6080 3180 6106
rect 2239 6062 2278 6067
rect 2239 6045 2247 6062
rect 2264 6045 2278 6062
rect 3002 6046 3170 6063
rect 2239 6040 2278 6045
<< viali >>
rect 1497 6722 1514 6740
rect 1536 6722 1553 6740
rect 1572 6722 1589 6740
rect 3477 6552 3495 6570
rect 3514 6552 3532 6570
rect 3054 6264 3072 6282
rect 1339 6187 1356 6204
rect 1456 6187 1473 6204
rect 3095 6402 3113 6420
rect 3396 6257 3414 6275
rect 3434 6257 3452 6275
rect 3095 6234 3113 6252
rect 2247 6045 2264 6062
rect 2286 6045 2303 6062
<< metal1 >>
rect 801 6770 815 6885
rect 1491 6740 1599 6770
rect 1491 6722 1497 6740
rect 1514 6722 1536 6740
rect 1553 6722 1572 6740
rect 1589 6722 1599 6740
rect 1491 6719 1599 6722
rect 2981 6738 3042 6755
rect 801 6541 808 6555
rect 801 6513 808 6527
rect 2981 6426 2999 6738
rect 3528 6588 4033 6602
rect 3471 6570 3538 6573
rect 3471 6552 3477 6570
rect 3495 6552 3514 6570
rect 3532 6568 3538 6570
rect 3532 6554 4033 6568
rect 3532 6552 3538 6554
rect 3471 6549 3538 6552
rect 2981 6420 3116 6426
rect 2981 6407 3095 6420
rect 3092 6402 3095 6407
rect 3113 6402 3116 6420
rect 3092 6396 3116 6402
rect 3051 6282 3075 6288
rect 3051 6277 3054 6282
rect 2953 6264 3054 6277
rect 3072 6264 3075 6282
rect 2953 6258 3075 6264
rect 3390 6275 3458 6278
rect 3092 6252 3116 6258
rect 3390 6257 3396 6275
rect 3414 6257 3434 6275
rect 3452 6273 3458 6275
rect 3452 6259 4033 6273
rect 3452 6257 3458 6259
rect 3390 6254 3458 6257
rect 3092 6234 3095 6252
rect 3113 6245 3116 6252
rect 3113 6234 3141 6245
rect 3092 6226 3141 6234
rect 1328 6204 1359 6212
rect 1328 6203 1339 6204
rect 801 6189 1339 6203
rect 1328 6187 1339 6189
rect 1356 6187 1359 6204
rect 1328 6179 1359 6187
rect 1448 6204 1476 6212
rect 1448 6187 1456 6204
rect 1473 6195 1476 6204
rect 1473 6187 1578 6195
rect 1448 6179 1578 6187
rect 801 5910 812 6026
rect 1314 6025 1542 6078
rect 1557 6067 1578 6179
rect 1557 6062 2311 6067
rect 1557 6045 2247 6062
rect 2264 6045 2286 6062
rect 2303 6045 2311 6062
rect 1557 6040 2311 6045
<< metal4 >>
rect 824 5000 984 7798
rect 1022 5000 1182 7798
rect 3678 5000 3838 7798
rect 3873 5000 4033 7798
use adc_comp_circuit  adc_comp_circuit_0
timestamp 1667211141
transform 1 0 1558 0 1 6689
box -757 -1689 2475 1109
use adc_inverter  adc_inverter_0
timestamp 1664803391
transform 1 0 1344 0 1 6118
box -13 -65 104 291
use adc_inverter  adc_inverter_1
timestamp 1664803391
transform 1 0 1461 0 1 6118
box -13 -65 104 291
use adc_nor  adc_nor_0
timestamp 1661513809
transform 1 0 3129 0 -1 6258
box -4 -118 253 230
use adc_nor_latch  adc_nor_latch_0
timestamp 1661515501
transform 1 0 3045 0 1 6456
box -3 0 505 348
<< labels >>
flabel metal1 s 801 6189 808 6203 7 FreeSans 80 0 0 0 clk
port 3 w signal input
flabel metal1 s 801 6541 808 6555 7 FreeSans 80 0 0 0 inp
port 4 w signal input
flabel metal1 s 801 6513 808 6527 7 FreeSans 80 0 0 0 inn
port 5 w signal input
flabel metal1 s 3952 6259 4033 6273 3 FreeSans 80 0 0 0 comp_trig
port 6 e signal output
flabel metal1 s 3952 6554 4033 6568 3 FreeSans 80 0 0 0 latch_qn
port 7 e signal output
flabel metal1 s 3952 6588 4033 6602 3 FreeSans 80 0 0 0 latch_q
port 8 e signal output
flabel metal4 3873 5000 4033 7798 0 FreeSans 800 90 0 0 VDD
port 1 nsew power bidirectional 
flabel metal4 3678 5000 3838 7798 0 FreeSans 800 90 0 0 VSS
port 2 nsew ground bidirectional
flabel metal4 1022 5000 1182 7798 0 FreeSans 800 90 0 0 VSS
port 2 nsew ground bidirectional
flabel metal4 824 5000 984 7798 0 FreeSans 800 90 0 0 VDD
port 1 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 4200 12900
string LEFclass BLOCK
string LEForigin 0 0
string LEFsource USER
<< end >>
