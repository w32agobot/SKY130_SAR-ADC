* SPICE3 file created from extract2.ext - technology: sky130A

C0 m4_21860_n30# top_1 1.27fF
C1 top_8 dummy_top 4.98fF
C2 dummy_bot bot_4 9.63fF
C3 dummy_bot bot_8 8.51fF
C4 dummy_bot top_2 1.56fF
C5 top_4 bot_4 7.12fF
C6 dummy_bot bot_1 9.63fF
C7 dummy_bot top_1 1.55fF
C8 m4_15440_n30# top_2 1.18fF
C9 top_4 dummy_bot 1.35fF
C10 top_1 bot_1 6.78fF
C11 top_8 bot_8 6.43fF
C12 top_8 dummy_bot 1.77fF
C13 dummy_bot dummy_top 55.72fF
C14 top_2 dummy_top 4.25fF
C15 top_1 dummy_top 4.24fF
C16 dummy_bot bot_2 9.64fF
C17 top_4 dummy_top 3.57fF
C18 bot_2 top_2 6.91fF
C19 dummy_top VSUBS 10.08fF
C20 bot_1 VSUBS 3.43fF
C21 bot_2 VSUBS 3.65fF
C22 bot_4 VSUBS 3.61fF
C23 bot_8 VSUBS 2.87fF
C24 dummy_bot VSUBS 38.21fF
