magic
tech sky130A
magscale 1 2
timestamp 1665042887
<< nwell >>
rect 0 506 1004 880
<< nmos >>
rect 232 252 262 336
rect 328 252 358 336
rect 536 252 566 336
rect 632 252 662 336
rect 728 252 758 336
<< pmos >>
rect 232 542 262 702
rect 328 542 358 702
rect 536 574 566 734
rect 632 574 662 734
rect 728 574 758 734
<< ndiff >>
rect 170 324 232 336
rect 170 264 182 324
rect 216 264 232 324
rect 170 252 232 264
rect 262 324 328 336
rect 262 264 278 324
rect 312 264 328 324
rect 262 252 328 264
rect 358 324 420 336
rect 358 264 374 324
rect 408 264 420 324
rect 358 252 420 264
rect 474 324 536 336
rect 474 264 486 324
rect 520 264 536 324
rect 474 252 536 264
rect 566 324 632 336
rect 566 264 582 324
rect 616 264 632 324
rect 566 252 632 264
rect 662 324 728 336
rect 662 264 678 324
rect 712 264 728 324
rect 662 252 728 264
rect 758 324 820 336
rect 758 264 774 324
rect 808 264 820 324
rect 758 252 820 264
<< pdiff >>
rect 474 722 536 734
rect 170 690 232 702
rect 170 554 182 690
rect 216 554 232 690
rect 170 542 232 554
rect 262 690 328 702
rect 262 554 278 690
rect 312 554 328 690
rect 262 542 328 554
rect 358 690 420 702
rect 358 554 374 690
rect 408 554 420 690
rect 474 586 486 722
rect 520 586 536 722
rect 474 574 536 586
rect 566 722 632 734
rect 566 586 582 722
rect 616 586 632 722
rect 566 574 632 586
rect 662 722 728 734
rect 662 586 678 722
rect 712 586 728 722
rect 662 574 728 586
rect 758 722 820 734
rect 758 586 774 722
rect 808 586 820 722
rect 758 574 820 586
rect 358 542 420 554
<< ndiffc >>
rect 182 264 216 324
rect 278 264 312 324
rect 374 264 408 324
rect 486 264 520 324
rect 582 264 616 324
rect 678 264 712 324
rect 774 264 808 324
<< pdiffc >>
rect 182 554 216 690
rect 278 554 312 690
rect 374 554 408 690
rect 486 586 520 722
rect 582 586 616 722
rect 678 586 712 722
rect 774 586 808 722
<< psubdiff >>
rect 182 148 230 182
rect 264 148 326 182
rect 360 148 384 182
rect 678 148 726 182
rect 760 148 792 182
<< nsubdiff >>
rect 302 838 806 844
rect 302 804 326 838
rect 360 804 430 838
rect 464 804 534 838
rect 568 804 630 838
rect 664 804 724 838
rect 758 804 806 838
rect 302 798 806 804
<< psubdiffcont >>
rect 230 148 264 182
rect 326 148 360 182
rect 726 148 760 182
<< nsubdiffcont >>
rect 326 804 360 838
rect 430 804 464 838
rect 534 804 568 838
rect 630 804 664 838
rect 724 804 758 838
<< poly >>
rect 212 818 280 828
rect 212 782 228 818
rect 264 782 280 818
rect 212 718 280 782
rect 536 734 566 760
rect 632 734 662 760
rect 728 734 758 760
rect 232 702 262 718
rect 328 702 358 728
rect 232 336 262 542
rect 328 508 358 542
rect 536 536 566 574
rect 632 548 662 574
rect 728 558 758 574
rect 728 548 834 558
rect 328 488 396 508
rect 328 450 346 488
rect 380 450 396 488
rect 328 352 396 450
rect 494 398 566 536
rect 608 516 834 548
rect 608 480 676 516
rect 624 430 660 480
rect 766 476 834 516
rect 624 426 676 430
rect 536 392 566 398
rect 608 392 676 426
rect 536 362 758 392
rect 328 336 358 352
rect 536 336 566 362
rect 632 336 662 362
rect 728 336 758 362
rect 232 226 262 252
rect 328 226 358 252
rect 536 226 566 252
rect 632 226 662 252
rect 728 226 758 252
rect 536 206 662 226
rect 510 196 662 206
rect 506 162 522 196
rect 556 162 590 196
rect 624 162 640 196
rect 506 150 640 162
<< polycont >>
rect 228 782 264 818
rect 346 450 380 488
rect 522 162 556 196
rect 590 162 624 196
<< locali >>
rect 34 922 148 1004
rect 34 888 46 922
rect 136 888 148 922
rect 854 922 970 1004
rect 854 920 868 922
rect 34 706 148 888
rect 844 888 868 920
rect 958 888 970 922
rect 302 838 806 844
rect 228 818 264 834
rect 302 804 326 838
rect 360 804 430 838
rect 464 804 534 838
rect 568 804 630 838
rect 664 804 724 838
rect 758 804 806 838
rect 302 798 806 804
rect 228 772 264 782
rect 228 738 230 772
rect 374 722 520 738
rect 34 672 46 706
rect 136 690 216 706
rect 136 672 182 690
rect 34 608 182 672
rect 34 574 46 608
rect 136 574 182 608
rect 34 554 182 574
rect 34 374 216 554
rect 278 690 312 706
rect 34 266 148 374
rect 34 232 114 266
rect 182 336 228 340
rect 182 324 194 336
rect 216 292 228 302
rect 278 324 312 554
rect 374 700 486 722
rect 374 690 432 700
rect 408 664 432 690
rect 466 664 486 700
rect 408 622 486 664
rect 408 586 432 622
rect 466 586 486 622
rect 408 570 520 586
rect 582 722 616 798
rect 582 570 616 586
rect 678 722 712 762
rect 408 554 476 570
rect 678 560 712 586
rect 774 722 808 738
rect 774 570 808 586
rect 844 706 970 888
rect 844 672 862 706
rect 952 672 970 706
rect 844 608 970 672
rect 844 574 862 608
rect 952 574 970 608
rect 374 538 476 554
rect 346 488 380 504
rect 346 414 380 450
rect 346 374 380 380
rect 414 374 476 538
rect 442 340 476 374
rect 844 340 970 574
rect 182 248 216 264
rect 278 248 312 264
rect 374 324 408 340
rect 442 336 520 340
rect 442 302 458 336
rect 492 324 520 336
rect 442 300 486 302
rect 374 260 408 264
rect 34 100 148 232
rect 486 248 520 264
rect 582 324 616 340
rect 582 248 616 264
rect 678 324 712 340
rect 374 220 408 226
rect 522 196 556 206
rect 590 196 624 206
rect 182 148 230 182
rect 264 148 326 182
rect 360 148 384 182
rect 506 162 522 196
rect 556 162 590 196
rect 624 162 640 196
rect 678 182 712 264
rect 774 324 808 340
rect 774 248 808 264
rect 844 282 864 340
rect 954 282 970 340
rect 34 66 46 100
rect 136 66 148 100
rect 34 0 148 66
rect 522 0 556 162
rect 590 150 624 162
rect 678 148 726 182
rect 760 148 792 182
rect 844 102 970 282
rect 844 68 864 102
rect 954 68 970 102
rect 844 56 970 68
rect 854 0 970 56
<< viali >>
rect 46 888 136 922
rect 868 888 958 922
rect 326 804 360 838
rect 430 804 464 838
rect 534 804 568 838
rect 630 804 664 838
rect 724 804 758 838
rect 230 738 264 772
rect 46 672 136 706
rect 46 574 136 608
rect 278 652 312 688
rect 278 574 312 610
rect 114 232 148 266
rect 194 324 228 336
rect 194 302 216 324
rect 216 302 228 324
rect 432 664 466 700
rect 432 586 466 622
rect 774 664 808 700
rect 774 586 808 622
rect 862 672 952 706
rect 862 574 952 608
rect 346 380 380 414
rect 458 324 492 336
rect 458 302 486 324
rect 486 302 492 324
rect 374 226 408 260
rect 582 290 616 324
rect 230 148 264 182
rect 326 148 360 182
rect 774 290 808 324
rect 864 282 954 340
rect 46 66 136 100
rect 726 148 760 182
rect 864 68 954 102
<< metal1 >>
rect 34 922 148 1004
rect 34 888 46 922
rect 136 888 148 922
rect 854 922 970 1004
rect 854 920 868 922
rect 34 882 148 888
rect 844 888 868 920
rect 958 888 970 922
rect 844 882 970 888
rect 0 838 1004 854
rect 0 806 326 838
rect 0 798 196 806
rect 298 804 326 806
rect 360 804 430 838
rect 464 804 534 838
rect 568 804 630 838
rect 664 804 724 838
rect 758 804 1004 838
rect 298 798 1004 804
rect 218 772 276 778
rect 218 770 230 772
rect 0 740 230 770
rect 218 738 230 740
rect 264 770 276 772
rect 264 740 1004 770
rect 264 738 276 740
rect 218 732 276 738
rect 34 706 148 712
rect 34 672 46 706
rect 136 672 148 706
rect 266 698 324 702
rect 426 700 472 712
rect 34 608 148 672
rect 34 574 46 608
rect 136 574 148 608
rect 34 568 148 574
rect 264 646 270 698
rect 322 646 328 698
rect 264 620 328 646
rect 264 568 270 620
rect 322 568 328 620
rect 426 664 432 700
rect 466 666 472 700
rect 768 700 814 712
rect 768 666 774 700
rect 466 664 774 666
rect 808 664 814 700
rect 426 638 814 664
rect 426 622 472 638
rect 426 586 432 622
rect 466 586 472 622
rect 426 574 472 586
rect 768 622 814 638
rect 768 586 774 622
rect 808 586 814 622
rect 768 574 814 586
rect 844 706 970 712
rect 844 672 862 706
rect 952 672 970 706
rect 844 608 970 672
rect 844 574 862 608
rect 952 574 970 608
rect 774 568 808 574
rect 844 568 970 574
rect 0 512 1004 540
rect 496 486 554 512
rect 166 458 450 478
rect 594 458 656 464
rect 770 458 830 484
rect 0 448 1004 458
rect 0 430 194 448
rect 422 430 1004 448
rect 334 414 392 420
rect 594 418 656 430
rect 334 402 346 414
rect 0 380 346 402
rect 380 402 392 414
rect 380 390 566 402
rect 736 390 1004 402
rect 380 380 1004 390
rect 0 374 1004 380
rect 334 368 392 374
rect 530 362 816 374
rect 182 336 240 346
rect 182 302 194 336
rect 228 328 240 336
rect 446 336 504 346
rect 446 328 458 336
rect 228 302 458 328
rect 492 302 504 336
rect 848 340 970 346
rect 182 300 504 302
rect 182 292 240 300
rect 446 292 504 300
rect 570 324 820 332
rect 570 290 582 324
rect 616 290 774 324
rect 808 290 820 324
rect 570 284 820 290
rect 848 282 864 340
rect 954 282 970 340
rect 108 266 154 278
rect 848 276 970 282
rect 108 248 114 266
rect 0 232 114 248
rect 148 248 154 266
rect 368 260 416 272
rect 368 248 374 260
rect 148 232 374 248
rect 0 226 374 232
rect 408 248 416 260
rect 408 226 1004 248
rect 0 220 1004 226
rect 0 182 1004 192
rect 0 148 230 182
rect 264 148 326 182
rect 360 148 726 182
rect 760 148 1004 182
rect 0 136 1004 148
rect 34 100 148 108
rect 34 66 46 100
rect 136 66 148 100
rect 34 0 148 66
rect 844 102 970 108
rect 844 68 864 102
rect 954 68 970 102
rect 844 56 970 68
rect 854 0 970 56
<< via1 >>
rect 270 688 322 698
rect 270 652 278 688
rect 278 652 312 688
rect 312 652 322 688
rect 270 646 322 652
rect 270 610 322 620
rect 270 574 278 610
rect 278 574 312 610
rect 312 574 322 610
rect 270 568 322 574
<< metal2 >>
rect 32 962 972 972
rect 32 906 42 962
rect 98 906 138 962
rect 194 906 234 962
rect 290 906 330 962
rect 386 906 426 962
rect 482 906 522 962
rect 578 906 618 962
rect 674 906 714 962
rect 770 906 810 962
rect 866 906 906 962
rect 962 906 972 962
rect 32 866 972 906
rect 32 810 42 866
rect 98 810 330 866
rect 386 810 618 866
rect 674 810 906 866
rect 962 810 972 866
rect 32 770 972 810
rect 32 714 42 770
rect 98 714 330 770
rect 386 714 618 770
rect 674 714 906 770
rect 962 714 972 770
rect 32 698 972 714
rect 32 674 270 698
rect 322 674 972 698
rect 32 618 42 674
rect 98 618 138 674
rect 194 618 234 674
rect 322 646 330 674
rect 290 620 330 646
rect 322 618 330 620
rect 386 618 426 674
rect 482 618 522 674
rect 578 618 618 674
rect 674 618 714 674
rect 770 618 810 674
rect 866 618 906 674
rect 962 618 972 674
rect 32 578 270 618
rect 32 522 42 578
rect 98 568 270 578
rect 322 608 972 618
rect 322 578 396 608
rect 322 568 330 578
rect 98 522 330 568
rect 386 522 396 578
rect 608 578 972 608
rect 32 482 396 522
rect 32 426 42 482
rect 98 426 330 482
rect 386 426 396 482
rect 460 460 544 544
rect 608 522 618 578
rect 674 522 906 578
rect 962 522 972 578
rect 608 482 972 522
rect 32 396 396 426
rect 608 426 618 482
rect 674 426 906 482
rect 962 426 972 482
rect 608 396 972 426
rect 32 386 972 396
rect 32 330 42 386
rect 98 330 138 386
rect 194 330 234 386
rect 290 330 330 386
rect 386 330 426 386
rect 482 330 522 386
rect 578 330 618 386
rect 674 330 714 386
rect 770 330 810 386
rect 866 330 906 386
rect 962 330 972 386
rect 32 290 972 330
rect 32 234 42 290
rect 98 234 330 290
rect 386 234 618 290
rect 674 234 906 290
rect 962 234 972 290
rect 32 194 972 234
rect 32 138 42 194
rect 98 138 330 194
rect 386 138 618 194
rect 674 138 906 194
rect 962 138 972 194
rect 32 98 972 138
rect 32 42 42 98
rect 98 42 138 98
rect 194 42 234 98
rect 290 42 330 98
rect 386 42 426 98
rect 482 42 522 98
rect 578 42 618 98
rect 674 42 714 98
rect 770 42 810 98
rect 866 42 906 98
rect 962 42 972 98
rect 32 32 972 42
<< via2 >>
rect 42 906 98 962
rect 138 906 194 962
rect 234 906 290 962
rect 330 906 386 962
rect 426 906 482 962
rect 522 906 578 962
rect 618 906 674 962
rect 714 906 770 962
rect 810 906 866 962
rect 906 906 962 962
rect 42 810 98 866
rect 330 810 386 866
rect 618 810 674 866
rect 906 810 962 866
rect 42 714 98 770
rect 330 714 386 770
rect 618 714 674 770
rect 906 714 962 770
rect 42 618 98 674
rect 138 618 194 674
rect 234 646 270 674
rect 270 646 290 674
rect 234 620 290 646
rect 234 618 270 620
rect 270 618 290 620
rect 330 618 386 674
rect 426 618 482 674
rect 522 618 578 674
rect 618 618 674 674
rect 714 618 770 674
rect 810 618 866 674
rect 906 618 962 674
rect 42 522 98 578
rect 330 522 386 578
rect 42 426 98 482
rect 330 426 386 482
rect 618 522 674 578
rect 906 522 962 578
rect 618 426 674 482
rect 906 426 962 482
rect 42 330 98 386
rect 138 330 194 386
rect 234 330 290 386
rect 330 330 386 386
rect 426 330 482 386
rect 522 330 578 386
rect 618 330 674 386
rect 714 330 770 386
rect 810 330 866 386
rect 906 330 962 386
rect 42 234 98 290
rect 330 234 386 290
rect 618 234 674 290
rect 906 234 962 290
rect 42 138 98 194
rect 330 138 386 194
rect 618 138 674 194
rect 906 138 962 194
rect 42 42 98 98
rect 138 42 194 98
rect 234 42 290 98
rect 330 42 386 98
rect 426 42 482 98
rect 522 42 578 98
rect 618 42 674 98
rect 714 42 770 98
rect 810 42 866 98
rect 906 42 962 98
<< metal3 >>
rect 36 962 968 968
rect 36 906 42 962
rect 98 906 138 962
rect 194 906 234 962
rect 290 906 330 962
rect 386 906 426 962
rect 482 906 522 962
rect 578 906 618 962
rect 674 906 714 962
rect 770 906 810 962
rect 866 906 906 962
rect 962 906 968 962
rect 36 900 968 906
rect 36 866 104 900
rect 36 810 42 866
rect 98 810 104 866
rect 324 866 392 900
rect 36 770 104 810
rect 36 714 42 770
rect 98 714 104 770
rect 164 824 264 840
rect 164 756 180 824
rect 248 756 264 824
rect 164 740 264 756
rect 324 810 330 866
rect 386 810 392 866
rect 612 866 680 900
rect 324 770 392 810
rect 36 680 104 714
rect 324 714 330 770
rect 386 714 392 770
rect 452 824 552 840
rect 452 756 468 824
rect 536 756 552 824
rect 452 740 552 756
rect 612 810 618 866
rect 674 810 680 866
rect 900 866 968 900
rect 612 770 680 810
rect 324 680 392 714
rect 612 714 618 770
rect 674 714 680 770
rect 740 824 840 840
rect 740 756 756 824
rect 824 756 840 824
rect 740 740 840 756
rect 900 810 906 866
rect 962 810 968 866
rect 900 770 968 810
rect 612 680 680 714
rect 900 714 906 770
rect 962 714 968 770
rect 900 680 968 714
rect 36 674 968 680
rect 36 618 42 674
rect 98 618 138 674
rect 194 618 234 674
rect 290 618 330 674
rect 386 618 426 674
rect 482 618 522 674
rect 578 618 618 674
rect 674 618 714 674
rect 770 618 810 674
rect 866 618 906 674
rect 962 618 968 674
rect 36 612 968 618
rect 36 578 104 612
rect 36 522 42 578
rect 98 522 104 578
rect 324 578 392 612
rect 36 482 104 522
rect 36 426 42 482
rect 98 426 104 482
rect 164 536 264 552
rect 164 468 180 536
rect 248 468 264 536
rect 164 452 264 468
rect 324 522 330 578
rect 386 522 392 578
rect 324 482 392 522
rect 36 392 104 426
rect 324 426 330 482
rect 386 426 392 482
rect 324 392 392 426
rect 612 578 680 612
rect 612 522 618 578
rect 674 522 680 578
rect 900 578 968 612
rect 612 482 680 522
rect 612 426 618 482
rect 674 426 680 482
rect 740 536 840 552
rect 740 468 756 536
rect 824 468 840 536
rect 740 452 840 468
rect 900 522 906 578
rect 962 522 968 578
rect 900 482 968 522
rect 612 392 680 426
rect 900 426 906 482
rect 962 426 968 482
rect 900 392 968 426
rect 36 386 968 392
rect 36 330 42 386
rect 98 330 138 386
rect 194 330 234 386
rect 290 330 330 386
rect 386 330 426 386
rect 482 330 522 386
rect 578 330 618 386
rect 674 330 714 386
rect 770 330 810 386
rect 866 330 906 386
rect 962 330 968 386
rect 36 324 968 330
rect 36 290 104 324
rect 36 234 42 290
rect 98 234 104 290
rect 324 290 392 324
rect 36 194 104 234
rect 36 138 42 194
rect 98 138 104 194
rect 164 248 264 264
rect 164 180 180 248
rect 248 180 264 248
rect 164 164 264 180
rect 324 234 330 290
rect 386 234 392 290
rect 612 290 680 324
rect 324 194 392 234
rect 36 104 104 138
rect 324 138 330 194
rect 386 138 392 194
rect 452 248 552 264
rect 452 180 468 248
rect 536 180 552 248
rect 452 164 552 180
rect 612 234 618 290
rect 674 234 680 290
rect 900 290 968 324
rect 612 194 680 234
rect 324 104 392 138
rect 612 138 618 194
rect 674 138 680 194
rect 740 248 840 264
rect 740 180 756 248
rect 824 180 840 248
rect 740 164 840 180
rect 900 234 906 290
rect 962 234 968 290
rect 900 194 968 234
rect 612 104 680 138
rect 900 138 906 194
rect 962 138 968 194
rect 900 104 968 138
rect 36 98 968 104
rect 36 42 42 98
rect 98 42 138 98
rect 194 42 234 98
rect 290 42 330 98
rect 386 42 426 98
rect 482 42 522 98
rect 578 42 618 98
rect 674 42 714 98
rect 770 42 810 98
rect 866 42 906 98
rect 962 42 968 98
rect 36 36 968 42
<< via3 >>
rect 180 756 248 824
rect 468 756 536 824
rect 756 756 824 824
rect 180 468 248 536
rect 756 468 824 536
rect 180 180 248 248
rect 468 180 536 248
rect 756 180 824 248
<< metal4 >>
rect 184 840 244 934
rect 472 840 532 934
rect 760 840 820 934
rect 164 824 264 840
rect 164 820 180 824
rect 70 760 180 820
rect 164 756 180 760
rect 248 756 264 824
rect 452 824 552 840
rect 452 820 468 824
rect 358 760 468 820
rect 164 740 264 756
rect 452 756 468 760
rect 536 820 552 824
rect 740 824 840 840
rect 740 820 756 824
rect 536 760 756 820
rect 536 756 552 760
rect 452 740 552 756
rect 740 756 756 760
rect 824 820 840 824
rect 824 760 934 820
rect 824 756 840 760
rect 740 740 840 756
rect 184 653 244 740
rect 183 552 244 653
rect 472 646 532 740
rect 760 646 820 740
rect 164 536 264 552
rect 164 532 180 536
rect 70 472 180 532
rect 164 468 180 472
rect 248 532 264 536
rect 740 536 840 552
rect 740 532 756 536
rect 248 472 358 532
rect 646 472 756 532
rect 248 468 264 472
rect 164 452 264 468
rect 740 468 756 472
rect 824 532 840 536
rect 824 472 934 532
rect 824 468 840 472
rect 740 452 840 468
rect 184 264 244 452
rect 472 264 532 358
rect 760 264 820 452
rect 164 248 264 264
rect 164 244 180 248
rect 70 184 180 244
rect 164 180 180 184
rect 248 244 264 248
rect 452 248 552 264
rect 452 244 468 248
rect 248 184 468 244
rect 248 180 264 184
rect 164 164 264 180
rect 452 180 468 184
rect 536 244 552 248
rect 740 248 840 264
rect 740 244 756 248
rect 536 184 756 244
rect 536 180 552 184
rect 452 164 552 180
rect 740 180 756 184
rect 824 244 840 248
rect 824 184 934 244
rect 824 180 840 184
rect 740 164 840 180
rect 184 70 244 164
rect 472 70 532 164
rect 760 70 820 164
<< comment >>
rect 0 972 32 1004
rect 972 972 1004 1004
rect 576 576 608 608
rect 544 544 576 576
rect 428 428 460 460
rect 396 396 428 428
rect 0 0 32 32
rect 972 0 1004 32
<< labels >>
rlabel metal1 0 798 0 854 7 VDD
port 1 w
rlabel metal1 0 740 0 770 7 sample_n
port 2 w
rlabel metal1 0 512 0 540 7 colon_n
port 3 w
rlabel metal1 0 430 0 458 7 col_n
port 4 w
rlabel metal1 0 374 0 402 7 sample
port 5 w
rlabel metal1 0 220 0 248 7 vcom
port 6 w
rlabel metal1 0 136 0 192 7 VSS
port 7 w
rlabel locali 854 0 970 0 5 row_n
port 8 s
rlabel locali 522 0 556 0 5 en_n
port 9 s
rlabel metal4 760 934 820 934 1 ctop
port 10 n
<< end >>
