** sch_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_vcm_clkgen.sch
.subckt adc_vcm_clkgen VDD VSS phi2_n phi2 phi1 phi1_n clk
*.PININFO VDD:B VSS:B phi2_n:O phi2:O phi1:O phi1_n:O clk:I
x23 clk VSS VSS VDD VDD net5 sky130_fd_sc_hd__inv_1
x2 net6 VSS VSS VDD VDD phi1 sky130_fd_sc_hd__buf_4
x5 net6 VSS VSS VDD VDD net3 sky130_fd_sc_hd__inv_1
x11 net11 VSS VSS VDD VDD net6 sky130_fd_sc_hd__inv_1
x12 net7 VSS VSS VDD VDD net4 sky130_fd_sc_hd__inv_1
x4 net3 VSS VSS VDD VDD phi1_n sky130_fd_sc_hd__buf_4
x7 net4 VSS VSS VDD VDD phi2_n sky130_fd_sc_hd__buf_4
x8 net7 VSS VSS VDD VDD phi2 sky130_fd_sc_hd__buf_4
x3 net1 VSS VSS VDD VDD net8 sky130_fd_sc_hd__dlymetal6s6s_1
x10 net2 VSS VSS VDD VDD net9 sky130_fd_sc_hd__dlymetal6s6s_1
x6 net8 VSS VSS VDD VDD net10 sky130_fd_sc_hd__dlymetal6s6s_1
x13 net9 VSS VSS VDD VDD net13 sky130_fd_sc_hd__dlymetal6s6s_1
x1 net12 VSS VSS VDD VDD net7 sky130_fd_sc_hd__inv_1
x9 net10 VSS VSS VDD VDD net11 sky130_fd_sc_hd__dlymetal6s6s_1
x14 net13 VSS VSS VDD VDD net12 sky130_fd_sc_hd__dlymetal6s6s_1
x15 clk net4 VSS VSS VDD VDD net1 sky130_fd_sc_hd__nand2_1
x16 net3 net5 VSS VSS VDD VDD net2 sky130_fd_sc_hd__nand2_1
.ends
.end
