magic
tech sky130A
magscale 1 2
timestamp 1673875808
<< nwell >>
rect 160 493 1192 814
<< nmos >>
rect 354 298 384 382
rect 450 298 480 382
rect 872 298 902 382
rect 968 298 998 382
<< pmos >>
rect 258 530 288 690
rect 354 530 384 690
rect 450 530 480 690
rect 546 530 576 690
rect 776 530 806 690
rect 872 530 902 690
rect 968 530 998 690
rect 1064 530 1094 690
<< ndiff >>
rect 292 370 354 382
rect 292 310 304 370
rect 338 310 354 370
rect 292 298 354 310
rect 384 370 450 382
rect 384 310 400 370
rect 434 310 450 370
rect 384 298 450 310
rect 480 370 542 382
rect 480 310 496 370
rect 530 310 542 370
rect 480 298 542 310
rect 810 370 872 382
rect 810 310 822 370
rect 856 310 872 370
rect 810 298 872 310
rect 902 370 968 382
rect 902 310 918 370
rect 952 310 968 370
rect 902 298 968 310
rect 998 370 1060 382
rect 998 310 1014 370
rect 1048 310 1060 370
rect 998 298 1060 310
<< pdiff >>
rect 196 678 258 690
rect 196 542 208 678
rect 242 542 258 678
rect 196 530 258 542
rect 288 678 354 690
rect 288 542 304 678
rect 338 542 354 678
rect 288 530 354 542
rect 384 678 450 690
rect 384 542 400 678
rect 434 542 450 678
rect 384 530 450 542
rect 480 678 546 690
rect 480 542 496 678
rect 530 542 546 678
rect 480 530 546 542
rect 576 678 638 690
rect 576 542 592 678
rect 626 542 638 678
rect 576 530 638 542
rect 714 678 776 690
rect 714 542 726 678
rect 760 542 776 678
rect 714 530 776 542
rect 806 678 872 690
rect 806 542 822 678
rect 856 542 872 678
rect 806 530 872 542
rect 902 678 968 690
rect 902 542 918 678
rect 952 542 968 678
rect 902 530 968 542
rect 998 678 1064 690
rect 998 542 1014 678
rect 1048 542 1064 678
rect 998 530 1064 542
rect 1094 678 1156 690
rect 1094 542 1110 678
rect 1144 542 1156 678
rect 1094 530 1156 542
<< ndiffc >>
rect 304 310 338 370
rect 400 310 434 370
rect 496 310 530 370
rect 822 310 856 370
rect 918 310 952 370
rect 1014 310 1048 370
<< pdiffc >>
rect 208 542 242 678
rect 304 542 338 678
rect 400 542 434 678
rect 496 542 530 678
rect 592 542 626 678
rect 726 542 760 678
rect 822 542 856 678
rect 918 542 952 678
rect 1014 542 1048 678
rect 1110 542 1144 678
<< psubdiff >>
rect 230 210 264 244
rect 298 210 332 244
rect 366 210 400 244
rect 434 210 468 244
rect 502 210 536 244
rect 570 210 782 244
rect 816 210 850 244
rect 884 210 918 244
rect 952 210 986 244
rect 1020 210 1054 244
rect 1088 210 1122 244
<< nsubdiff >>
rect 208 744 264 778
rect 298 744 332 778
rect 366 744 400 778
rect 434 744 468 778
rect 502 744 536 778
rect 570 744 782 778
rect 816 744 850 778
rect 884 744 918 778
rect 952 744 986 778
rect 1020 744 1054 778
rect 1088 744 1144 778
<< psubdiffcont >>
rect 264 210 298 244
rect 332 210 366 244
rect 400 210 434 244
rect 468 210 502 244
rect 536 210 570 244
rect 782 210 816 244
rect 850 210 884 244
rect 918 210 952 244
rect 986 210 1020 244
rect 1054 210 1088 244
<< nsubdiffcont >>
rect 264 744 298 778
rect 332 744 366 778
rect 400 744 434 778
rect 468 744 502 778
rect 536 744 570 778
rect 782 744 816 778
rect 850 744 884 778
rect 918 744 952 778
rect 986 744 1020 778
rect 1054 744 1088 778
<< poly >>
rect 258 690 288 717
rect 354 690 384 716
rect 450 690 480 717
rect 546 690 576 716
rect 776 690 806 717
rect 872 690 902 716
rect 968 690 998 717
rect 1064 690 1094 716
rect 258 484 288 530
rect 354 490 384 530
rect 220 468 288 484
rect 220 434 238 468
rect 272 434 288 468
rect 220 424 288 434
rect 330 480 390 490
rect 450 484 480 530
rect 546 490 576 530
rect 330 446 346 480
rect 380 446 390 480
rect 330 430 390 446
rect 444 469 504 484
rect 444 435 454 469
rect 488 435 504 469
rect 354 382 384 430
rect 444 425 504 435
rect 546 480 614 490
rect 776 484 806 530
rect 872 490 902 530
rect 546 446 564 480
rect 598 446 614 480
rect 546 430 614 446
rect 738 468 806 484
rect 738 434 756 468
rect 790 434 806 468
rect 450 382 480 425
rect 738 424 806 434
rect 848 480 908 490
rect 968 484 998 530
rect 1064 490 1094 530
rect 848 446 864 480
rect 898 446 908 480
rect 848 430 908 446
rect 962 469 1022 484
rect 962 435 972 469
rect 1006 435 1022 469
rect 872 382 902 430
rect 962 425 1022 435
rect 1064 480 1132 490
rect 1064 446 1082 480
rect 1116 446 1132 480
rect 1064 430 1132 446
rect 968 382 998 425
rect 354 272 384 298
rect 450 272 480 298
rect 872 272 902 298
rect 968 272 998 298
<< polycont >>
rect 238 434 272 468
rect 346 446 380 480
rect 454 435 488 469
rect 564 446 598 480
rect 756 434 790 468
rect 864 446 898 480
rect 972 435 1006 469
rect 1082 446 1116 480
<< locali >>
rect 208 744 264 778
rect 298 744 332 778
rect 366 744 400 778
rect 434 744 468 778
rect 502 744 536 778
rect 570 744 782 778
rect 816 744 850 778
rect 884 744 918 778
rect 952 744 986 778
rect 1020 744 1054 778
rect 1088 744 1144 778
rect 208 678 242 744
rect 208 526 242 542
rect 304 678 338 694
rect 304 526 338 542
rect 400 678 434 694
rect 400 526 434 542
rect 496 678 530 694
rect 496 526 530 542
rect 592 678 626 744
rect 592 526 626 542
rect 726 678 760 744
rect 726 526 760 542
rect 822 678 856 694
rect 822 526 856 542
rect 918 678 952 694
rect 918 526 952 542
rect 1014 678 1048 694
rect 1014 526 1048 542
rect 1110 678 1144 744
rect 1110 526 1144 542
rect 220 468 288 484
rect 220 434 238 468
rect 272 434 288 468
rect 220 424 288 434
rect 330 480 398 490
rect 330 446 346 480
rect 380 446 398 480
rect 330 430 398 446
rect 436 469 504 484
rect 436 434 454 469
rect 488 434 504 469
rect 436 425 504 434
rect 546 480 614 490
rect 546 446 564 480
rect 598 446 614 480
rect 546 430 614 446
rect 738 468 806 484
rect 738 434 756 468
rect 790 434 806 468
rect 738 424 806 434
rect 848 480 916 490
rect 848 446 864 480
rect 898 446 916 480
rect 848 430 916 446
rect 954 469 1022 484
rect 954 434 972 469
rect 1006 434 1022 469
rect 954 425 1022 434
rect 1064 480 1132 490
rect 1064 446 1082 480
rect 1116 446 1132 480
rect 1064 430 1132 446
rect 304 370 338 386
rect 304 244 338 310
rect 400 370 434 386
rect 400 294 434 302
rect 496 370 530 386
rect 496 244 530 310
rect 822 370 856 386
rect 822 244 856 310
rect 918 370 952 386
rect 918 294 952 302
rect 1014 370 1048 386
rect 1014 244 1048 310
rect 230 210 264 244
rect 298 210 332 244
rect 366 210 400 244
rect 434 210 468 244
rect 502 210 536 244
rect 570 210 782 244
rect 816 210 850 244
rect 884 210 918 244
rect 952 210 986 244
rect 1020 210 1054 244
rect 1088 210 1122 244
<< viali >>
rect 400 594 434 628
rect 918 594 952 628
rect 238 434 272 468
rect 346 446 380 480
rect 454 435 488 468
rect 454 434 488 435
rect 564 446 598 480
rect 756 434 790 468
rect 864 446 898 480
rect 972 435 1006 468
rect 972 434 1006 435
rect 1082 446 1116 480
rect 400 310 434 336
rect 400 302 434 310
rect 918 310 952 336
rect 918 302 952 310
<< metal1 >>
rect 391 637 443 643
rect 391 579 443 585
rect 909 637 961 643
rect 909 579 961 585
rect 190 508 644 536
rect 708 508 1162 536
rect 336 480 388 508
rect 554 486 618 508
rect 229 468 281 480
rect 229 434 238 468
rect 272 434 281 468
rect 336 446 346 480
rect 380 446 388 480
rect 336 434 388 446
rect 444 468 504 480
rect 444 434 454 468
rect 488 434 504 468
rect 554 434 560 486
rect 612 434 618 486
rect 854 480 906 508
rect 1072 486 1136 508
rect 747 468 799 480
rect 747 434 756 468
rect 790 434 799 468
rect 854 446 864 480
rect 898 446 906 480
rect 854 434 906 446
rect 962 468 1022 480
rect 962 434 972 468
rect 1006 434 1022 468
rect 1072 434 1078 486
rect 1130 434 1136 486
rect 229 405 281 434
rect 444 405 504 434
rect 747 406 799 434
rect 190 377 627 405
rect 391 340 443 348
rect 391 277 443 284
rect 596 305 627 377
rect 655 354 661 406
rect 713 405 799 406
rect 962 405 1022 434
rect 713 377 1162 405
rect 713 354 719 377
rect 909 340 961 348
rect 655 305 661 324
rect 596 277 661 305
rect 655 272 661 277
rect 713 305 719 324
rect 713 277 795 305
rect 909 277 961 284
rect 713 272 719 277
<< via1 >>
rect 391 628 443 637
rect 391 594 400 628
rect 400 594 434 628
rect 434 594 443 628
rect 391 585 443 594
rect 909 628 961 637
rect 909 594 918 628
rect 918 594 952 628
rect 952 594 961 628
rect 909 585 961 594
rect 560 480 612 486
rect 560 446 564 480
rect 564 446 598 480
rect 598 446 612 480
rect 560 434 612 446
rect 1078 480 1130 486
rect 1078 446 1082 480
rect 1082 446 1116 480
rect 1116 446 1130 480
rect 1078 434 1130 446
rect 391 336 443 340
rect 391 302 400 336
rect 400 302 434 336
rect 434 302 443 336
rect 391 284 443 302
rect 661 354 713 406
rect 909 336 961 340
rect 661 272 713 324
rect 909 302 918 336
rect 918 302 952 336
rect 952 302 961 336
rect 909 284 961 302
<< metal2 >>
rect 389 637 445 648
rect 389 585 391 637
rect 443 585 445 637
rect 389 574 445 585
rect 391 340 443 574
rect 618 499 682 638
rect 907 637 963 648
rect 907 585 909 637
rect 961 585 963 637
rect 907 574 963 585
rect 1136 630 1200 639
rect 1136 574 1139 630
rect 1197 574 1200 630
rect 618 486 621 499
rect 554 434 560 486
rect 612 443 621 486
rect 679 443 682 499
rect 612 434 682 443
rect 655 405 661 406
rect 190 284 391 305
rect 596 377 661 405
rect 596 305 627 377
rect 655 354 661 377
rect 713 354 719 406
rect 909 340 961 574
rect 1136 486 1200 574
rect 1072 434 1078 486
rect 1130 434 1200 486
rect 443 284 627 305
rect 190 277 627 284
rect 655 272 661 324
rect 713 305 719 324
rect 713 284 909 305
rect 961 284 1162 305
rect 713 277 1162 284
rect 713 272 719 277
<< via2 >>
rect 1139 574 1197 630
rect 621 443 679 499
<< metal3 >>
rect 618 629 684 642
rect 1134 630 1202 642
rect 1134 629 1139 630
rect 190 574 1139 629
rect 1197 574 1202 630
rect 190 569 1202 574
rect 616 499 684 507
rect 616 494 621 499
rect 190 443 621 494
rect 679 494 684 499
rect 1132 494 1202 507
rect 679 443 1202 494
rect 190 434 1202 443
<< labels >>
flabel metal2 1086 277 1162 305 0 FreeSans 160 0 0 0 q
port 2 nsew
flabel metal1 1086 377 1162 405 0 FreeSans 160 0 0 0 qn
port 4 nsew
flabel metal3 190 434 1200 494 0 FreeSans 160 0 0 0 s
port 6 nsew
flabel metal3 190 569 1200 629 0 FreeSans 160 0 0 0 r
port 7 nsew
flabel locali 208 744 1144 778 0 FreeSans 160 0 0 0 VDD
port 8 nsew
flabel locali 230 210 1122 244 0 FreeSans 160 0 0 0 VSS
port 9 nsew
flabel metal1 190 377 229 405 0 FreeSans 160 0 0 0 q
port 10 nsew
flabel metal2 190 277 229 305 0 FreeSans 160 0 0 0 qn
port 11 nsew
<< end >>
