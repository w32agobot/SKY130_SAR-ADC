* SPICE3 file created from adc_array_cap_16.ext - technology: sky130A

.subckt adc_array_circuit ROW_N COL_N COLON_N SAMPLE SAMPLE_N CBOT VCOM VDRV VDD VSS
X0 VINT2 COLON_N VDRV VSS sky130_fd_pr__nfet_01v8 ad=2.478e+11p pd=2.86e+06u as=2.52e+11p ps=2.88e+06u w=420000u l=180000u
X1 VINT2 ROW_N VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.26e+11p ps=1.44e+06u w=420000u l=180000u
X2 VSS COL_N VINT2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=180000u
X3 CBOT SAMPLE_N VCOM VDD sky130_fd_pr__pfet_01v8 ad=4.5e+11p pd=2.8e+06u as=4.5e+11p ps=2.8e+06u w=900000u l=180000u
X4 VDRV SAMPLE CBOT VDD sky130_fd_pr__pfet_01v8 ad=1.305e+12p pd=8.3e+06u as=0p ps=0u w=900000u l=180000u
X5 VINT COL_N VDRV VDD sky130_fd_pr__pfet_01v8 ad=4.5e+11p pd=2.8e+06u as=0p ps=0u w=900000u l=180000u
X6 CBOT SAMPLE_N VDRV VSS sky130_fd_pr__nfet_01v8 ad=1.26e+11p pd=1.44e+06u as=0p ps=0u w=420000u l=180000u
X7 VCOM SAMPLE CBOT VSS sky130_fd_pr__nfet_01v8 ad=1.26e+11p pd=1.44e+06u as=0p ps=0u w=420000u l=180000u
X8 VDD ROW_N VINT VDD sky130_fd_pr__pfet_01v8 ad=4.5e+11p pd=2.8e+06u as=0p ps=0u w=900000u l=180000u
X9 VDRV COLON_N VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=900000u l=180000u
C0 VDRV SAMPLE_N 0.25fF
C1 COLON_N COL_N 1.23fF
C2 VDRV COL_N 0.98fF
C3 VDD SAMPLE_N 1.16fF
C4 COLON_N SAMPLE 0.69fF
C5 VDRV SAMPLE 0.24fF
C6 VDRV VCOM 0.26fF
C7 VDD ROW_N 0.27fF
C8 SAMPLE SAMPLE_N 0.21fF
C9 VDRV CBOT 0.23fF
C10 VCOM VSS 1.65fF
C11 COLON_N VSS 0.36fF
C12 COL_N VSS 0.34fF
C13 SAMPLE VSS 0.30fF
C14 ROW_N VSS 1.02fF
C15 SAMPLE_N VSS 0.36fF
C16 VDD VSS 2.65fF
C17 VDRV VSS 0.23fF
.ends

.subckt adc_array_cap_16 COL_N COLON_N CTOP ROW_N SAMPLE SAMPLE_N VCOM VDD CBOT VSS
Xadc_array_circuit_0 ROW_N COL_N COLON_N SAMPLE SAMPLE_N CBOT VCOM adc_array_circuit_0/VDRV
+ VDD VSS adc_array_circuit
C0 VDD CTOP 0.28fF
C1 COL_N CBOT 0.34fF
C2 VDD CBOT 0.91fF
C3 CBOT ROW_N 0.27fF
C4 COLON_N CBOT 0.35fF
C5 VCOM CBOT 0.47fF
C6 CBOT adc_array_circuit_0/VDRV 0.42fF
C7 CTOP CBOT 7.87fF
C8 CBOT SAMPLE 0.36fF
C9 CBOT SAMPLE_N 0.39fF
C10 CTOP VSS 0.91fF
C11 CBOT VSS 2.82fF
C12 VCOM VSS 1.65fF
C13 COLON_N VSS 0.36fF
C14 COL_N VSS 0.34fF
C15 SAMPLE VSS 0.30fF
C16 ROW_N VSS 1.02fF
C17 SAMPLE_N VSS 0.36fF
C18 VDD VSS 2.65fF
C19 adc_array_circuit_0/VDRV VSS 0.23fF
.ends

