VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_mm_sc_hd_dly5ns
  CLASS CORE ;
  FOREIGN sky130_mm_sc_hd_dly5ns ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.200 BY 2.720 ;
  SITE unithd ;
  PIN in
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.880000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.990 0.325 1.320 ;
    END
  END in
  PIN out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.366000 ;
    ANTENNADIFFAREA 0.361800 ;
    PORT
      LAYER li1 ;
        RECT 6.330 1.460 6.500 2.300 ;
        RECT 6.740 1.010 6.910 1.340 ;
        RECT 8.620 0.980 8.850 1.290 ;
        RECT 6.440 0.380 6.610 0.890 ;
      LAYER mcon ;
        RECT 6.330 1.540 6.500 1.820 ;
        RECT 6.740 1.090 6.910 1.260 ;
        RECT 8.650 1.100 8.820 1.270 ;
        RECT 6.440 0.720 6.610 0.890 ;
      LAYER met1 ;
        RECT 6.300 1.240 6.530 1.970 ;
        RECT 6.710 1.240 6.940 1.320 ;
        RECT 8.590 1.240 8.880 1.300 ;
        RECT 6.300 1.100 8.880 1.240 ;
        RECT 6.410 1.030 6.940 1.100 ;
        RECT 8.590 1.070 8.880 1.100 ;
        RECT 6.410 0.660 6.640 1.030 ;
    END
  END out
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.635 9.200 2.805 ;
        RECT 0.530 1.395 0.700 2.235 ;
        RECT 5.370 1.460 5.540 2.635 ;
        RECT 7.080 1.290 7.250 2.635 ;
        RECT 7.080 1.120 7.630 1.290 ;
        RECT 7.460 0.380 7.630 1.120 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 0.530 1.475 0.700 2.155 ;
      LAYER met1 ;
        RECT 0.000 2.480 9.200 2.960 ;
        RECT 0.500 1.415 0.730 2.480 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 7.930 1.180 8.100 2.300 ;
        RECT 7.930 1.010 8.450 1.180 ;
        RECT 0.530 0.455 0.700 0.915 ;
        RECT 5.480 0.085 5.650 0.840 ;
        RECT 8.280 0.085 8.450 1.010 ;
        RECT 0.000 -0.085 9.200 0.085 ;
      LAYER mcon ;
        RECT 0.530 0.535 0.700 0.835 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
      LAYER met1 ;
        RECT 0.500 0.240 0.730 0.910 ;
        RECT 4.800 0.240 5.320 0.680 ;
        RECT 0.000 -0.240 9.200 0.240 ;
      LAYER via ;
        RECT 4.900 0.290 5.220 0.640 ;
      LAYER met2 ;
        RECT 4.800 0.240 5.320 0.680 ;
      LAYER via2 ;
        RECT 4.900 0.300 5.220 0.670 ;
      LAYER met3 ;
        RECT 0.695 0.700 4.670 2.280 ;
        RECT 5.870 0.700 8.530 2.280 ;
        RECT 0.695 0.270 8.530 0.700 ;
    END
  END VGND
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.235 9.390 2.910 ;
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 -0.085 9.195 1.070 ;
    END
  END VNB
  OBS
      LAYER li1 ;
        RECT 4.820 1.180 4.990 2.235 ;
        RECT 5.850 1.460 6.020 2.300 ;
        RECT 7.420 1.460 7.620 2.300 ;
        RECT 8.410 1.460 8.610 2.300 ;
        RECT 5.410 1.180 5.770 1.290 ;
        RECT 4.820 1.010 5.770 1.180 ;
        RECT 4.820 0.365 4.990 1.010 ;
        RECT 5.960 0.380 6.130 0.840 ;
        RECT 6.980 0.380 7.150 0.840 ;
        RECT 7.940 0.380 8.110 0.840 ;
      LAYER mcon ;
        RECT 4.820 1.475 4.990 2.085 ;
        RECT 5.850 1.540 6.020 2.220 ;
        RECT 7.450 1.640 7.620 2.220 ;
        RECT 8.410 1.640 8.580 2.220 ;
        RECT 5.410 1.070 5.690 1.240 ;
        RECT 5.960 0.460 6.130 0.760 ;
        RECT 6.980 0.460 7.150 0.660 ;
        RECT 7.940 0.460 8.110 0.660 ;
      LAYER met1 ;
        RECT 4.790 1.290 5.020 2.195 ;
        RECT 5.820 2.110 8.610 2.280 ;
        RECT 5.820 1.480 6.050 2.110 ;
        RECT 7.420 1.580 7.650 2.110 ;
        RECT 8.380 1.580 8.610 2.110 ;
        RECT 4.790 1.010 5.770 1.290 ;
        RECT 5.930 0.520 6.160 0.820 ;
        RECT 6.950 0.520 7.180 0.720 ;
        RECT 7.910 0.520 8.140 0.720 ;
        RECT 5.930 0.380 8.140 0.520 ;
      LAYER via ;
        RECT 5.410 1.020 5.690 1.280 ;
      LAYER met2 ;
        RECT 5.040 0.840 5.770 1.430 ;
      LAYER via2 ;
        RECT 5.090 1.070 5.380 1.350 ;
      LAYER met3 ;
        RECT 5.030 1.000 5.440 1.600 ;
      LAYER via3 ;
        RECT 5.080 1.050 5.400 1.370 ;
      LAYER met4 ;
        RECT 5.030 1.340 5.440 1.430 ;
        RECT 4.110 0.970 6.470 1.340 ;
        RECT 5.030 0.840 5.440 0.970 ;
  END
END sky130_mm_sc_hd_dly5ns
END LIBRARY

