magic
tech sky130A
magscale 1 2
timestamp 1658918966
<< error_p >>
rect -161 -116 161 116
<< nwell >>
rect -161 -116 161 116
<< pmos >>
rect -63 -80 -33 80
rect 33 -80 63 80
<< pdiff >>
rect -125 68 -63 80
rect -125 -68 -113 68
rect -79 -68 -63 68
rect -125 -80 -63 -68
rect -33 68 33 80
rect -33 -68 -17 68
rect 17 -68 33 68
rect -33 -80 33 -68
rect 63 68 125 80
rect 63 -68 79 68
rect 113 -68 125 68
rect 63 -80 125 -68
<< pdiffc >>
rect -113 -68 -79 68
rect -17 -68 17 68
rect 79 -68 113 68
<< poly >>
rect -63 80 -33 106
rect 33 80 63 106
rect -63 -106 -33 -80
rect 33 -106 63 -80
<< locali >>
rect -113 68 -79 84
rect -113 -84 -79 -68
rect -17 68 17 84
rect -17 -84 17 -68
rect 79 68 113 84
rect 79 -84 113 -68
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.8 l 0.15 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
