* SPICE3 file created from adc_array_wafflecap_8(8)x563aF_25um2.ext - technology: sky130A

.subckt adc_array_wafflecap_8(8)x563aF_25um2 ctop cbot
C0 ctop cbot 4.51fF
C1 ctop VSUBS 0.69fF
C2 cbot VSUBS 2.01fF
.ends
