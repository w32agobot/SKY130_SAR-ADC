* SPICE3 file created from adc_array_fingercap_8(4)x343aF_topB_22um2.ext - technology: sky130A

C0 cbot floatingmetal 1.37fF
C1 VSS floatingmetal 0.50fF
C2 ctop cbot 1.37fF
C3 ctop VSS 0.52fF
C4 ctop floatingmetal 0.30fF
C5 cbot VSS 3.09fF
C6 floatingmetal VSUBS 0.46fF
C7 ctop VSUBS 0.51fF
C8 cbot VSUBS 0.43fF
C9 VSS VSUBS 1.80fF
