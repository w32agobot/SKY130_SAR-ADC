magic
tech sky130A
timestamp 1659097417
<< metal1 >>
rect 172 632 533 635
rect 172 606 225 632
rect 252 606 291 632
rect 318 606 424 632
rect 451 606 490 632
rect 517 606 533 632
rect 172 604 533 606
rect 169 29 533 32
rect 169 3 225 29
rect 252 3 291 29
rect 318 3 424 29
rect 451 3 490 29
rect 517 3 533 29
rect 169 2 533 3
rect 169 1 530 2
<< via1 >>
rect 225 606 252 632
rect 291 606 318 632
rect 424 606 451 632
rect 490 606 517 632
rect 225 3 252 29
rect 291 3 318 29
rect 424 3 451 29
rect 490 3 517 29
<< metal2 >>
rect 172 632 571 635
rect 172 606 225 632
rect 252 606 291 632
rect 318 606 424 632
rect 451 606 490 632
rect 517 606 571 632
rect 172 604 571 606
rect 172 592 343 604
rect 399 592 571 604
rect 172 524 328 592
rect 357 577 385 590
rect 343 574 399 577
rect 343 543 348 574
rect 394 543 399 574
rect 343 539 399 543
rect 172 471 343 524
rect 172 403 328 471
rect 357 456 385 539
rect 414 524 571 592
rect 399 471 571 524
rect 343 453 399 456
rect 343 422 348 453
rect 394 422 399 453
rect 343 418 399 422
rect 172 351 343 403
rect 172 283 328 351
rect 357 336 385 418
rect 414 403 571 471
rect 399 351 571 403
rect 343 333 399 336
rect 343 302 348 333
rect 394 302 399 333
rect 343 298 399 302
rect 172 231 343 283
rect 172 163 328 231
rect 357 216 385 298
rect 414 283 571 351
rect 399 231 571 283
rect 343 213 399 216
rect 343 182 348 213
rect 394 182 399 213
rect 343 178 399 182
rect 172 111 343 163
rect 172 44 328 111
rect 357 96 385 178
rect 414 163 571 231
rect 399 111 571 163
rect 343 93 399 96
rect 343 62 348 93
rect 394 62 399 93
rect 343 58 399 62
rect 357 53 385 58
rect 414 44 571 111
rect 172 32 343 44
rect 399 32 571 44
rect 172 29 571 32
rect 172 3 225 29
rect 252 3 291 29
rect 318 3 424 29
rect 451 3 490 29
rect 517 3 571 29
rect 172 1 571 3
<< via2 >>
rect 348 543 394 574
rect 348 422 394 453
rect 348 302 394 333
rect 348 182 394 213
rect 348 62 394 93
<< metal3 >>
rect 343 574 399 577
rect 343 573 348 574
rect 244 543 348 573
rect 394 573 399 574
rect 394 543 499 573
rect 343 539 399 543
rect 172 481 175 513
rect 207 512 210 513
rect 533 512 536 513
rect 207 482 328 512
rect 414 482 536 512
rect 207 481 210 482
rect 533 481 536 482
rect 568 481 571 513
rect 343 453 399 456
rect 343 452 348 453
rect 244 422 348 452
rect 394 452 399 453
rect 394 422 499 452
rect 343 418 399 422
rect 172 361 175 393
rect 207 392 210 393
rect 533 392 536 393
rect 207 362 328 392
rect 414 362 536 392
rect 207 361 210 362
rect 533 361 536 362
rect 568 361 571 393
rect 343 333 399 336
rect 343 332 348 333
rect 244 302 348 332
rect 394 332 399 333
rect 394 302 499 332
rect 343 298 399 302
rect 172 241 175 273
rect 207 272 210 273
rect 533 272 536 273
rect 207 242 328 272
rect 414 242 536 272
rect 207 241 210 242
rect 533 241 536 242
rect 568 241 571 273
rect 343 213 399 216
rect 343 212 348 213
rect 244 182 348 212
rect 394 212 399 213
rect 394 182 499 212
rect 343 178 399 182
rect 172 121 175 153
rect 207 152 210 153
rect 533 152 536 153
rect 207 122 328 152
rect 414 122 536 152
rect 207 121 210 122
rect 533 121 536 122
rect 568 121 571 153
rect 343 93 399 96
rect 343 92 348 93
rect 244 62 348 92
rect 394 92 399 93
rect 394 62 499 92
rect 343 58 399 62
<< via3 >>
rect 175 481 207 513
rect 536 481 568 513
rect 175 361 207 393
rect 536 361 568 393
rect 175 241 207 273
rect 536 241 568 273
rect 175 121 207 153
rect 536 121 568 153
<< metal4 >>
rect 172 603 571 635
rect 172 513 210 603
rect 172 481 175 513
rect 207 481 210 513
rect 172 393 210 481
rect 172 361 175 393
rect 207 361 210 393
rect 172 273 210 361
rect 172 241 175 273
rect 207 241 210 273
rect 172 153 210 241
rect 172 121 175 153
rect 207 121 210 153
rect 172 89 210 121
rect 169 58 210 89
rect 172 32 210 58
rect 533 513 571 603
rect 533 481 536 513
rect 568 481 571 513
rect 533 393 571 481
rect 533 361 536 393
rect 568 361 571 393
rect 533 273 571 361
rect 533 241 536 273
rect 568 241 571 273
rect 533 153 571 241
rect 533 121 536 153
rect 568 121 571 153
rect 533 32 571 121
rect 172 0 571 32
<< labels >>
rlabel metal2 357 53 385 53 1 cbot
rlabel metal4 169 58 169 89 7 ctop
rlabel metal1 169 1 169 32 3 VSS
<< end >>
