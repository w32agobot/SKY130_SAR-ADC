magic
tech sky130A
timestamp 1662367448
<< nwell >>
rect 1786 2998 1845 3202
rect 167 2759 349 2804
rect 144 2747 349 2759
rect 144 2618 172 2747
rect 227 2692 349 2747
rect 221 2673 349 2692
rect 227 2618 349 2673
rect 144 2605 349 2618
rect 1785 2426 1925 2628
<< poly >>
rect 1840 2954 1856 2968
rect 1840 2872 1855 2954
rect 1840 2863 1877 2872
rect 1840 2846 1855 2863
rect 1872 2846 1877 2863
rect 1840 2838 1877 2846
rect 1039 2460 1078 2465
rect 1039 2443 1047 2460
rect 1064 2443 1078 2460
rect 1039 2438 1078 2443
<< polycont >>
rect 1855 2846 1872 2863
rect 139 2585 156 2602
rect 1047 2443 1064 2460
<< locali >>
rect 291 3138 399 3141
rect 291 3120 297 3138
rect 314 3120 336 3138
rect 353 3120 372 3138
rect 389 3120 399 3138
rect 291 3117 399 3120
rect 291 2804 334 3117
rect 2271 2968 2338 2971
rect 2271 2950 2277 2968
rect 2295 2950 2314 2968
rect 2332 2950 2338 2968
rect 2271 2947 2338 2950
rect 175 2784 334 2804
rect 1851 2863 1875 2871
rect 1851 2846 1855 2863
rect 1872 2846 1875 2863
rect 1904 2846 2454 2872
rect 244 2692 266 2784
rect 244 2673 290 2692
rect 1851 2680 1875 2846
rect 1851 2662 1854 2680
rect 1872 2662 1875 2680
rect 131 2602 158 2610
rect 131 2585 139 2602
rect 156 2585 158 2602
rect 131 2577 158 2585
rect 248 2602 275 2610
rect 248 2585 256 2602
rect 273 2585 275 2602
rect 248 2577 275 2585
rect 1851 2504 1875 2662
rect 1892 2818 1916 2824
rect 1892 2800 1895 2818
rect 1913 2800 1916 2818
rect 1892 2650 1916 2800
rect 1985 2763 2028 2846
rect 2158 2673 2258 2676
rect 2158 2657 2196 2673
rect 2190 2655 2196 2657
rect 2214 2655 2234 2673
rect 2252 2655 2258 2673
rect 2190 2652 2258 2655
rect 1892 2632 1895 2650
rect 1913 2632 1916 2650
rect 1892 2626 1916 2632
rect 1851 2478 1980 2504
rect 1039 2460 1078 2465
rect 1039 2443 1047 2460
rect 1064 2443 1078 2460
rect 1802 2444 1970 2461
rect 1039 2438 1078 2443
<< viali >>
rect 297 3120 314 3138
rect 336 3120 353 3138
rect 372 3120 389 3138
rect 2277 2950 2295 2968
rect 2314 2950 2332 2968
rect 1854 2662 1872 2680
rect 139 2585 156 2602
rect 256 2585 273 2602
rect 1895 2800 1913 2818
rect 2196 2655 2214 2673
rect 2234 2655 2252 2673
rect 1895 2632 1913 2650
rect 1047 2443 1064 2460
rect 1086 2443 1103 2460
<< metal1 >>
rect -61 3168 -47 3283
rect 291 3138 399 3168
rect 291 3120 297 3138
rect 314 3120 336 3138
rect 353 3120 372 3138
rect 389 3120 399 3138
rect 291 3117 399 3120
rect 1781 3136 1842 3153
rect -61 2939 -54 2953
rect -61 2911 -54 2925
rect 1781 2824 1799 3136
rect 2328 2986 2538 3000
rect 2271 2968 2338 2971
rect 2271 2950 2277 2968
rect 2295 2950 2314 2968
rect 2332 2966 2338 2968
rect 2332 2952 2538 2966
rect 2332 2950 2338 2952
rect 2271 2947 2338 2950
rect 1781 2818 1916 2824
rect 1781 2805 1895 2818
rect 1892 2800 1895 2805
rect 1913 2800 1916 2818
rect 1892 2794 1916 2800
rect 1851 2680 1875 2686
rect 1851 2675 1854 2680
rect 1753 2662 1854 2675
rect 1872 2662 1875 2680
rect 1753 2656 1875 2662
rect 2190 2673 2258 2676
rect 1892 2650 1916 2656
rect 2190 2655 2196 2673
rect 2214 2655 2234 2673
rect 2252 2671 2258 2673
rect 2252 2657 2538 2671
rect 2252 2655 2258 2657
rect 2190 2652 2258 2655
rect 1892 2632 1895 2650
rect 1913 2643 1916 2650
rect 1913 2632 1941 2643
rect 1892 2624 1941 2632
rect 128 2602 159 2610
rect 128 2601 139 2602
rect -61 2587 139 2601
rect 128 2585 139 2587
rect 156 2585 159 2602
rect 128 2577 159 2585
rect 248 2602 276 2610
rect 248 2585 256 2602
rect 273 2593 276 2602
rect 273 2585 378 2593
rect 248 2577 378 2585
rect -61 2308 -50 2424
rect 114 2423 342 2476
rect 357 2465 378 2577
rect 357 2460 1111 2465
rect 357 2443 1047 2460
rect 1064 2443 1086 2460
rect 1103 2443 1111 2460
rect 357 2438 1111 2443
use NOR-Latch  NOR-Latch_0 ../NOR-Latch
timestamp 1661515501
transform 1 0 1845 0 1 2854
box -3 0 505 348
use NOR  NOR_0 ../NOR
timestamp 1661513809
transform 1 0 1929 0 -1 2656
box -4 -118 253 230
use adc_comp_circuit  adc_comp_circuit_0 ../adc_comp_circuit
timestamp 1662367448
transform 1 0 358 0 1 3087
box -419 -2565 2180 1987
use inverter  inverter_0 ../inverter
timestamp 1662366209
transform 1 0 144 0 1 2516
box -13 -65 104 291
use inverter  inverter_1
timestamp 1662366209
transform 1 0 261 0 1 2516
box -13 -65 104 291
<< labels >>
rlabel metal1 -61 2587 -61 2601 7 clk
port 1 w
rlabel metal1 2538 2657 2538 2671 3 comp_trig
port 11 e
rlabel metal1 2538 2986 2538 3000 3 latch_q
port 12 e
rlabel metal1 2538 2952 2538 2966 3 latch_qn
port 13 e
rlabel metal1 -61 2939 -61 2953 7 inp
port 15 w
rlabel metal1 -61 2911 -61 2925 7 inn
port 16 w
rlabel metal1 -61 3168 -61 3283 7 VDD
port 18 w
rlabel metal1 -61 2308 -61 2424 7 VSS
port 19 w
<< end >>
