magic
tech sky130A
magscale 1 2
timestamp 1663599054
<< nmos >>
rect -129 -50 -29 50
rect 29 -50 129 50
<< ndiff >>
rect -187 38 -129 50
rect -187 -38 -175 38
rect -141 -38 -129 38
rect -187 -50 -129 -38
rect -29 38 29 50
rect -29 -38 -17 38
rect 17 -38 29 38
rect -29 -50 29 -38
rect 129 38 187 50
rect 129 -38 141 38
rect 175 -38 187 38
rect 129 -50 187 -38
<< ndiffc >>
rect -175 -38 -141 38
rect -17 -38 17 38
rect 141 -38 175 38
<< poly >>
rect -129 50 -29 76
rect 29 50 129 76
rect -129 -76 -29 -50
rect 29 -76 129 -50
<< locali >>
rect -175 38 -141 54
rect -175 -54 -141 -38
rect -17 38 17 54
rect -17 -54 17 -38
rect 141 38 175 54
rect 141 -54 175 -38
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.5 l 0.5 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
