magic
tech sky130A
magscale 1 2
timestamp 1661178173
<< error_p >>
rect -1589 -1100 -1529 1100
rect -1509 -1100 -1449 1100
rect -70 -1100 -10 1100
rect 10 -1100 70 1100
rect 1449 -1100 1509 1100
rect 1529 -1100 1589 1100
<< metal3 >>
rect -3028 1072 -1529 1100
rect -3028 -1072 -1613 1072
rect -1549 -1072 -1529 1072
rect -3028 -1100 -1529 -1072
rect -1509 1072 -10 1100
rect -1509 -1072 -94 1072
rect -30 -1072 -10 1072
rect -1509 -1100 -10 -1072
rect 10 1072 1509 1100
rect 10 -1072 1425 1072
rect 1489 -1072 1509 1072
rect 10 -1100 1509 -1072
rect 1529 1072 3028 1100
rect 1529 -1072 2944 1072
rect 3008 -1072 3028 1072
rect 1529 -1100 3028 -1072
<< via3 >>
rect -1613 -1072 -1549 1072
rect -94 -1072 -30 1072
rect 1425 -1072 1489 1072
rect 2944 -1072 3008 1072
<< mimcap >>
rect -2928 960 -1728 1000
rect -2928 -960 -2888 960
rect -1768 -960 -1728 960
rect -2928 -1000 -1728 -960
rect -1409 960 -209 1000
rect -1409 -960 -1369 960
rect -249 -960 -209 960
rect -1409 -1000 -209 -960
rect 110 960 1310 1000
rect 110 -960 150 960
rect 1270 -960 1310 960
rect 110 -1000 1310 -960
rect 1629 960 2829 1000
rect 1629 -960 1669 960
rect 2789 -960 2829 960
rect 1629 -1000 2829 -960
<< mimcapcontact >>
rect -2888 -960 -1768 960
rect -1369 -960 -249 960
rect 150 -960 1270 960
rect 1669 -960 2789 960
<< metal4 >>
rect -1629 1072 -1533 1088
rect -2889 960 -1767 961
rect -2889 -960 -2888 960
rect -1768 -960 -1767 960
rect -2889 -961 -1767 -960
rect -1629 -1072 -1613 1072
rect -1549 -1072 -1533 1072
rect -110 1072 -14 1088
rect -1370 960 -248 961
rect -1370 -960 -1369 960
rect -249 -960 -248 960
rect -1370 -961 -248 -960
rect -1629 -1088 -1533 -1072
rect -110 -1072 -94 1072
rect -30 -1072 -14 1072
rect 1409 1072 1505 1088
rect 149 960 1271 961
rect 149 -960 150 960
rect 1270 -960 1271 960
rect 149 -961 1271 -960
rect -110 -1088 -14 -1072
rect 1409 -1072 1425 1072
rect 1489 -1072 1505 1072
rect 2928 1072 3024 1088
rect 1668 960 2790 961
rect 1668 -960 1669 960
rect 2789 -960 2790 960
rect 1668 -961 2790 -960
rect 1409 -1088 1505 -1072
rect 2928 -1072 2944 1072
rect 3008 -1072 3024 1072
rect 2928 -1088 3024 -1072
<< properties >>
string FIXED_BBOX 1529 -1100 2929 1100
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 6 l 10 val 126.08 carea 2.00 cperi 0.19 nx 4 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
