magic
tech sky130A
timestamp 1659880747
<< locali >>
rect -19 1934 0 1935
rect 175 1934 203 1935
rect 554 1934 582 1935
rect 933 1934 961 1935
rect 1312 1934 1340 1935
rect 1681 1934 1895 1935
rect 2070 1934 2098 1935
rect 2449 1934 2477 1935
rect 2828 1934 2856 1935
rect 3207 1934 3235 1935
rect 3576 1934 3790 1935
rect 3965 1934 3993 1935
rect 4344 1934 4372 1935
rect 4723 1934 4751 1935
rect 5102 1934 5130 1935
rect 5471 1934 5685 1935
rect 5860 1934 5888 1935
rect 6239 1934 6267 1935
rect 6618 1934 6646 1935
rect 6997 1934 7025 1935
rect 7366 1934 7580 1935
rect -19 1929 7599 1934
rect -19 1902 176 1929
rect 202 1902 555 1929
rect 581 1902 934 1929
rect 960 1902 1313 1929
rect 1339 1928 2071 1929
rect 1339 1902 1692 1928
rect -19 1901 1692 1902
rect 1718 1902 2071 1928
rect 2097 1902 2450 1929
rect 2476 1902 2829 1929
rect 2855 1902 3208 1929
rect 3234 1928 3966 1929
rect 3234 1902 3587 1928
rect 1718 1901 3587 1902
rect 3613 1902 3966 1928
rect 3992 1902 4345 1929
rect 4371 1902 4724 1929
rect 4750 1902 5103 1929
rect 5129 1928 5861 1929
rect 5129 1902 5482 1928
rect 3613 1901 5482 1902
rect 5508 1902 5861 1928
rect 5887 1902 6240 1929
rect 6266 1902 6619 1929
rect 6645 1902 6998 1929
rect 7024 1928 7599 1929
rect 7024 1902 7377 1928
rect 5508 1901 7377 1902
rect 7403 1901 7599 1928
rect -19 1896 7599 1901
rect 0 1895 209 1896
rect 166 1343 203 1895
rect 1684 1352 1721 1896
rect 1895 1895 2104 1896
rect 159 1336 203 1343
rect 554 1337 582 1341
rect 933 1337 961 1339
rect 159 1309 176 1336
rect 202 1309 203 1336
rect 159 1303 203 1309
rect 548 1335 1342 1337
rect 548 1308 555 1335
rect 581 1333 1342 1335
rect 581 1308 934 1333
rect 548 1306 934 1308
rect 960 1331 1342 1333
rect 960 1306 1313 1331
rect 548 1304 1313 1306
rect 1339 1304 1342 1331
rect 548 1303 1342 1304
rect 1681 1331 1723 1352
rect 2061 1343 2098 1895
rect 3579 1349 3616 1896
rect 3790 1895 3999 1896
rect 1681 1304 1692 1331
rect 1718 1304 1723 1331
rect 159 725 201 1303
rect 554 1302 582 1303
rect 554 726 582 729
rect 825 726 880 1303
rect 933 1300 961 1303
rect 1312 1298 1340 1303
rect 933 726 961 729
rect 1312 726 1340 729
rect 159 717 206 725
rect 159 690 176 717
rect 202 690 206 717
rect 550 723 1344 726
rect 550 696 555 723
rect 581 696 934 723
rect 960 696 1313 723
rect 1339 696 1344 723
rect 1681 724 1723 1304
rect 1681 697 1692 724
rect 1718 697 1723 724
rect 1681 696 1723 697
rect 2056 1336 2098 1343
rect 2449 1337 2477 1341
rect 2828 1337 2856 1339
rect 2056 1309 2071 1336
rect 2097 1309 2098 1336
rect 2056 725 2098 1309
rect 2443 1335 3237 1337
rect 2443 1308 2450 1335
rect 2476 1333 3237 1335
rect 2476 1308 2829 1333
rect 2443 1306 2829 1308
rect 2855 1331 3237 1333
rect 2855 1306 3208 1331
rect 2443 1304 3208 1306
rect 3234 1304 3237 1331
rect 2443 1303 3237 1304
rect 3574 1331 3616 1349
rect 3956 1342 3993 1895
rect 5474 1360 5511 1896
rect 5685 1895 5894 1896
rect 5851 1360 5888 1895
rect 7369 1366 7406 1896
rect 7580 1895 7599 1896
rect 3574 1304 3587 1331
rect 3613 1304 3616 1331
rect 2449 1302 2477 1303
rect 2449 726 2477 729
rect 2681 726 2736 1303
rect 2828 1300 2856 1303
rect 3207 1298 3235 1303
rect 2828 726 2856 729
rect 3207 726 3235 729
rect 3574 728 3616 1304
rect 3951 1336 3993 1342
rect 4344 1337 4372 1341
rect 4723 1337 4751 1339
rect 3951 1309 3966 1336
rect 3992 1309 3993 1336
rect 2056 717 2101 725
rect 550 692 1344 696
rect 554 690 582 692
rect 933 690 961 692
rect 1312 690 1340 692
rect 159 687 206 690
rect 168 523 206 687
rect 166 522 1372 523
rect 1684 522 1722 696
rect 2056 690 2071 717
rect 2097 690 2101 717
rect 2445 723 3239 726
rect 2445 696 2450 723
rect 2476 696 2829 723
rect 2855 696 3208 723
rect 3234 696 3239 723
rect 2445 692 3239 696
rect 3574 724 3617 728
rect 3574 697 3587 724
rect 3613 697 3617 724
rect 3574 693 3617 697
rect 2449 690 2477 692
rect 2056 687 2101 690
rect 166 511 1723 522
rect 2063 520 2101 687
rect 166 484 176 511
rect 202 484 555 511
rect 581 484 934 511
rect 960 484 1313 511
rect 1339 510 1723 511
rect 1339 484 1692 510
rect 166 483 1692 484
rect 1718 483 1723 510
rect 166 477 1723 483
rect 2062 513 2480 520
rect 2062 511 2450 513
rect 2062 484 2071 511
rect 2097 486 2450 511
rect 2476 486 2480 513
rect 2097 484 2480 486
rect 2062 479 2480 484
rect 2824 515 2857 692
rect 3207 690 3235 692
rect 2824 509 2858 515
rect 3579 512 3617 693
rect 3951 725 3993 1309
rect 4338 1335 5132 1337
rect 4338 1308 4345 1335
rect 4371 1333 5132 1335
rect 4371 1308 4724 1333
rect 4338 1306 4724 1308
rect 4750 1331 5132 1333
rect 4750 1306 5103 1331
rect 4338 1304 5103 1306
rect 5129 1304 5132 1331
rect 4338 1303 5132 1304
rect 5471 1331 5513 1360
rect 5471 1304 5482 1331
rect 5508 1304 5513 1331
rect 4344 1302 4372 1303
rect 4344 726 4372 729
rect 4577 726 4632 1303
rect 4723 1300 4751 1303
rect 5102 1298 5130 1303
rect 4723 726 4751 729
rect 5102 726 5130 729
rect 3951 717 3996 725
rect 3951 690 3966 717
rect 3992 690 3996 717
rect 4340 723 5134 726
rect 4340 696 4345 723
rect 4371 696 4724 723
rect 4750 696 5103 723
rect 5129 696 5134 723
rect 5471 724 5513 1304
rect 5471 704 5482 724
rect 4340 692 5134 696
rect 5474 697 5482 704
rect 5508 704 5513 724
rect 5851 1336 5893 1360
rect 6239 1337 6267 1341
rect 6618 1337 6646 1339
rect 5851 1309 5861 1336
rect 5887 1309 5893 1336
rect 5851 717 5893 1309
rect 6233 1335 7027 1337
rect 6233 1308 6240 1335
rect 6266 1333 7027 1335
rect 6266 1308 6619 1333
rect 6233 1306 6619 1308
rect 6645 1331 7027 1333
rect 6645 1306 6998 1331
rect 6233 1304 6998 1306
rect 7024 1304 7027 1331
rect 6233 1303 7027 1304
rect 7365 1331 7407 1366
rect 7365 1304 7377 1331
rect 7403 1304 7407 1331
rect 6239 1302 6267 1303
rect 6239 726 6267 729
rect 6480 726 6535 1303
rect 6618 1300 6646 1303
rect 6997 1298 7025 1303
rect 6618 728 6646 729
rect 6612 726 6648 728
rect 6997 726 7025 729
rect 5851 704 5861 717
rect 5508 697 5512 704
rect 4344 690 4372 692
rect 3951 686 3996 690
rect 3958 514 3996 686
rect 2824 482 2829 509
rect 2855 482 2858 509
rect 2063 478 2101 479
rect 166 473 1372 477
rect 2824 476 2858 482
rect 3202 510 3620 512
rect 3202 505 3587 510
rect 3202 478 3208 505
rect 3234 483 3587 505
rect 3613 483 3620 510
rect 3234 478 3620 483
rect 2824 475 2857 476
rect 3202 475 3620 478
rect 3956 511 4374 514
rect 3956 484 3966 511
rect 3992 506 4374 511
rect 3992 484 4345 506
rect 3956 479 4345 484
rect 4371 479 4374 506
rect 3956 477 4374 479
rect 3205 472 3237 475
rect 4342 473 4374 477
rect 4720 506 4753 692
rect 5102 690 5130 692
rect 5474 513 5512 697
rect 5853 690 5861 704
rect 5887 704 5893 717
rect 6235 723 7029 726
rect 5887 690 5891 704
rect 6235 696 6240 723
rect 6266 696 6619 723
rect 6645 696 6998 723
rect 7024 696 7029 723
rect 7365 724 7407 1304
rect 7365 710 7377 724
rect 6235 692 7029 696
rect 7369 697 7377 710
rect 7403 697 7407 724
rect 6239 690 6267 692
rect 5853 517 5891 690
rect 4720 479 4724 506
rect 4750 479 4753 506
rect 4720 471 4753 479
rect 5098 510 5512 513
rect 5098 507 5482 510
rect 5098 480 5103 507
rect 5129 483 5482 507
rect 5508 483 5512 510
rect 5129 481 5512 483
rect 5851 511 6270 517
rect 5851 484 5861 511
rect 5887 510 6270 511
rect 5887 484 6240 510
rect 5851 483 6240 484
rect 6266 483 6270 510
rect 5129 480 5511 481
rect 5851 480 6270 483
rect 6612 513 6648 692
rect 6997 690 7025 692
rect 6612 486 6619 513
rect 6645 486 6648 513
rect 5098 475 5511 480
rect 5853 478 5891 480
rect 6237 477 6269 480
rect 6612 479 6648 486
rect 6995 515 7027 516
rect 7369 515 7407 697
rect 6995 510 7407 515
rect 6995 483 6998 510
rect 7024 483 7377 510
rect 7403 483 7407 510
rect 6995 477 7407 483
rect 5100 474 5132 475
<< viali >>
rect 176 1902 202 1929
rect 555 1902 581 1929
rect 934 1902 960 1929
rect 1313 1902 1339 1929
rect 1692 1901 1718 1928
rect 2071 1902 2097 1929
rect 2450 1902 2476 1929
rect 2829 1902 2855 1929
rect 3208 1902 3234 1929
rect 3587 1901 3613 1928
rect 3966 1902 3992 1929
rect 4345 1902 4371 1929
rect 4724 1902 4750 1929
rect 5103 1902 5129 1929
rect 5482 1901 5508 1928
rect 5861 1902 5887 1929
rect 6240 1902 6266 1929
rect 6619 1902 6645 1929
rect 6998 1902 7024 1929
rect 7377 1901 7403 1928
rect 176 1309 202 1336
rect 555 1308 581 1335
rect 934 1306 960 1333
rect 1313 1304 1339 1331
rect 1692 1304 1718 1331
rect 176 690 202 717
rect 555 696 581 723
rect 934 696 960 723
rect 1313 696 1339 723
rect 1692 697 1718 724
rect 2071 1309 2097 1336
rect 2450 1308 2476 1335
rect 2829 1306 2855 1333
rect 3208 1304 3234 1331
rect 3587 1304 3613 1331
rect 3966 1309 3992 1336
rect 2071 690 2097 717
rect 2450 696 2476 723
rect 2829 696 2855 723
rect 3208 696 3234 723
rect 3587 697 3613 724
rect 176 484 202 511
rect 555 484 581 511
rect 934 484 960 511
rect 1313 484 1339 511
rect 1692 483 1718 510
rect 2071 484 2097 511
rect 2450 486 2476 513
rect 4345 1308 4371 1335
rect 4724 1306 4750 1333
rect 5103 1304 5129 1331
rect 5482 1304 5508 1331
rect 3966 690 3992 717
rect 4345 696 4371 723
rect 4724 696 4750 723
rect 5103 696 5129 723
rect 5482 697 5508 724
rect 5861 1309 5887 1336
rect 6240 1308 6266 1335
rect 6619 1306 6645 1333
rect 6998 1304 7024 1331
rect 7377 1304 7403 1331
rect 2829 482 2855 509
rect 3208 478 3234 505
rect 3587 483 3613 510
rect 3966 484 3992 511
rect 4345 479 4371 506
rect 5861 690 5887 717
rect 6240 696 6266 723
rect 6619 696 6645 723
rect 6998 696 7024 723
rect 7377 697 7403 724
rect 4724 479 4750 506
rect 5103 480 5129 507
rect 5482 483 5508 510
rect 5861 484 5887 511
rect 6240 483 6266 510
rect 6619 486 6645 513
rect 6998 483 7024 510
rect 7377 483 7403 510
<< metal1 >>
rect 0 2425 360 2428
rect 0 2399 34 2425
rect 61 2399 109 2425
rect 136 2399 242 2425
rect 269 2399 317 2425
rect 344 2399 360 2425
rect 0 2397 360 2399
rect 379 2425 739 2428
rect 379 2399 413 2425
rect 440 2399 488 2425
rect 515 2399 621 2425
rect 648 2399 696 2425
rect 723 2399 739 2425
rect 379 2397 739 2399
rect 758 2425 1118 2428
rect 758 2399 792 2425
rect 819 2399 867 2425
rect 894 2399 1000 2425
rect 1027 2399 1075 2425
rect 1102 2399 1118 2425
rect 758 2397 1118 2399
rect 1137 2425 1497 2428
rect 1137 2399 1171 2425
rect 1198 2399 1246 2425
rect 1273 2399 1379 2425
rect 1406 2399 1454 2425
rect 1481 2399 1497 2425
rect 1137 2397 1497 2399
rect 1516 2425 1876 2428
rect 1516 2399 1550 2425
rect 1577 2399 1625 2425
rect 1652 2399 1758 2425
rect 1785 2399 1833 2425
rect 1860 2399 1876 2425
rect 1516 2397 1876 2399
rect 1895 2425 2255 2428
rect 1895 2399 1929 2425
rect 1956 2399 2004 2425
rect 2031 2399 2137 2425
rect 2164 2399 2212 2425
rect 2239 2399 2255 2425
rect 1895 2397 2255 2399
rect 2274 2425 2634 2428
rect 2274 2399 2308 2425
rect 2335 2399 2383 2425
rect 2410 2399 2516 2425
rect 2543 2399 2591 2425
rect 2618 2399 2634 2425
rect 2274 2397 2634 2399
rect 2653 2425 3013 2428
rect 2653 2399 2687 2425
rect 2714 2399 2762 2425
rect 2789 2399 2895 2425
rect 2922 2399 2970 2425
rect 2997 2399 3013 2425
rect 2653 2397 3013 2399
rect 3032 2425 3392 2428
rect 3032 2399 3066 2425
rect 3093 2399 3141 2425
rect 3168 2399 3274 2425
rect 3301 2399 3349 2425
rect 3376 2399 3392 2425
rect 3032 2397 3392 2399
rect 3411 2425 3771 2428
rect 3411 2399 3445 2425
rect 3472 2399 3520 2425
rect 3547 2399 3653 2425
rect 3680 2399 3728 2425
rect 3755 2399 3771 2425
rect 3411 2397 3771 2399
rect 3790 2425 4150 2428
rect 3790 2399 3824 2425
rect 3851 2399 3899 2425
rect 3926 2399 4032 2425
rect 4059 2399 4107 2425
rect 4134 2399 4150 2425
rect 3790 2397 4150 2399
rect 4169 2425 4529 2428
rect 4169 2399 4203 2425
rect 4230 2399 4278 2425
rect 4305 2399 4411 2425
rect 4438 2399 4486 2425
rect 4513 2399 4529 2425
rect 4169 2397 4529 2399
rect 4548 2425 4908 2428
rect 4548 2399 4582 2425
rect 4609 2399 4657 2425
rect 4684 2399 4790 2425
rect 4817 2399 4865 2425
rect 4892 2399 4908 2425
rect 4548 2397 4908 2399
rect 4927 2425 5287 2428
rect 4927 2399 4961 2425
rect 4988 2399 5036 2425
rect 5063 2399 5169 2425
rect 5196 2399 5244 2425
rect 5271 2399 5287 2425
rect 4927 2397 5287 2399
rect 5306 2425 5666 2428
rect 5306 2399 5340 2425
rect 5367 2399 5415 2425
rect 5442 2399 5548 2425
rect 5575 2399 5623 2425
rect 5650 2399 5666 2425
rect 5306 2397 5666 2399
rect 5685 2425 6045 2428
rect 5685 2399 5719 2425
rect 5746 2399 5794 2425
rect 5821 2399 5927 2425
rect 5954 2399 6002 2425
rect 6029 2399 6045 2425
rect 6080 2425 6424 2428
rect 6080 2412 6109 2425
rect 6136 2412 6184 2425
rect 6211 2412 6317 2425
rect 6344 2412 6392 2425
rect 5685 2397 6045 2399
rect 6064 2399 6098 2412
rect 6136 2399 6173 2412
rect 6211 2399 6306 2412
rect 6344 2399 6381 2412
rect 6419 2399 6424 2425
rect 6461 2425 6803 2428
rect 6461 2412 6488 2425
rect 6515 2412 6563 2425
rect 6590 2412 6696 2425
rect 6723 2412 6771 2425
rect 6064 2397 6424 2399
rect 6443 2399 6477 2412
rect 6515 2399 6552 2412
rect 6590 2399 6685 2412
rect 6723 2399 6760 2412
rect 6798 2399 6803 2425
rect 6840 2425 7182 2428
rect 6840 2412 6867 2425
rect 6894 2412 6942 2425
rect 6969 2412 7075 2425
rect 7102 2412 7150 2425
rect 6443 2397 6803 2399
rect 6822 2399 6856 2412
rect 6894 2399 6931 2412
rect 6969 2399 7064 2412
rect 7102 2399 7139 2412
rect 7177 2399 7182 2425
rect 6822 2397 7182 2399
rect 7201 2425 7561 2428
rect 7201 2399 7235 2425
rect 7262 2399 7310 2425
rect 7337 2399 7443 2425
rect 7470 2399 7518 2425
rect 7545 2399 7561 2425
rect 7201 2397 7561 2399
rect 173 1929 205 1935
rect 173 1902 176 1929
rect 202 1902 205 1929
rect 173 1896 205 1902
rect 552 1929 584 1935
rect 552 1902 555 1929
rect 581 1902 584 1929
rect 552 1896 584 1902
rect 931 1929 963 1935
rect 931 1902 934 1929
rect 960 1902 963 1929
rect 931 1896 963 1902
rect 1310 1929 1342 1935
rect 1310 1902 1313 1929
rect 1339 1902 1342 1929
rect 1310 1896 1342 1902
rect 1689 1928 1721 1934
rect 1689 1901 1692 1928
rect 1718 1901 1721 1928
rect 1689 1895 1721 1901
rect 2068 1929 2100 1935
rect 2068 1902 2071 1929
rect 2097 1902 2100 1929
rect 2068 1896 2100 1902
rect 2447 1929 2479 1935
rect 2447 1902 2450 1929
rect 2476 1902 2479 1929
rect 2447 1896 2479 1902
rect 2826 1929 2858 1935
rect 2826 1902 2829 1929
rect 2855 1902 2858 1929
rect 2826 1896 2858 1902
rect 3205 1929 3237 1935
rect 3205 1902 3208 1929
rect 3234 1902 3237 1929
rect 3205 1896 3237 1902
rect 3584 1928 3616 1934
rect 3584 1901 3587 1928
rect 3613 1901 3616 1928
rect 3584 1895 3616 1901
rect 3963 1929 3995 1935
rect 3963 1902 3966 1929
rect 3992 1902 3995 1929
rect 3963 1896 3995 1902
rect 4342 1929 4374 1935
rect 4342 1902 4345 1929
rect 4371 1902 4374 1929
rect 4342 1896 4374 1902
rect 4721 1929 4753 1935
rect 4721 1902 4724 1929
rect 4750 1902 4753 1929
rect 4721 1896 4753 1902
rect 5100 1929 5132 1935
rect 5100 1902 5103 1929
rect 5129 1902 5132 1929
rect 5100 1896 5132 1902
rect 5479 1928 5511 1934
rect 5479 1901 5482 1928
rect 5508 1901 5511 1928
rect 5479 1895 5511 1901
rect 5858 1929 5890 1935
rect 5858 1902 5861 1929
rect 5887 1902 5890 1929
rect 5858 1896 5890 1902
rect 6237 1929 6269 1935
rect 6237 1902 6240 1929
rect 6266 1902 6269 1929
rect 6237 1896 6269 1902
rect 6616 1929 6648 1935
rect 6616 1902 6619 1929
rect 6645 1902 6648 1929
rect 6616 1896 6648 1902
rect 6995 1929 7027 1935
rect 6995 1902 6998 1929
rect 7024 1902 7027 1929
rect 6995 1896 7027 1902
rect 7374 1928 7406 1934
rect 7374 1901 7377 1928
rect 7403 1901 7406 1928
rect 7374 1895 7406 1901
rect 0 1822 360 1825
rect 0 1796 34 1822
rect 61 1796 109 1822
rect 136 1796 242 1822
rect 269 1796 317 1822
rect 344 1796 360 1822
rect 0 1794 360 1796
rect 379 1822 739 1825
rect 379 1796 413 1822
rect 440 1796 488 1822
rect 515 1796 621 1822
rect 648 1796 696 1822
rect 723 1796 739 1822
rect 379 1794 739 1796
rect 758 1822 1118 1825
rect 758 1796 792 1822
rect 819 1796 867 1822
rect 894 1796 1000 1822
rect 1027 1796 1075 1822
rect 1102 1796 1118 1822
rect 758 1794 1118 1796
rect 1137 1822 1497 1825
rect 1137 1796 1171 1822
rect 1198 1796 1246 1822
rect 1273 1796 1379 1822
rect 1406 1796 1454 1822
rect 1481 1796 1497 1822
rect 1137 1794 1497 1796
rect 1516 1822 1876 1825
rect 1516 1796 1550 1822
rect 1577 1796 1625 1822
rect 1652 1796 1758 1822
rect 1785 1796 1833 1822
rect 1860 1796 1876 1822
rect 1516 1794 1876 1796
rect 1895 1822 2255 1825
rect 1895 1796 1929 1822
rect 1956 1796 2004 1822
rect 2031 1796 2137 1822
rect 2164 1796 2212 1822
rect 2239 1796 2255 1822
rect 1895 1794 2255 1796
rect 2274 1822 2634 1825
rect 2274 1796 2308 1822
rect 2335 1796 2383 1822
rect 2410 1796 2516 1822
rect 2543 1796 2591 1822
rect 2618 1796 2634 1822
rect 2274 1794 2634 1796
rect 2653 1822 3013 1825
rect 2653 1796 2687 1822
rect 2714 1796 2762 1822
rect 2789 1796 2895 1822
rect 2922 1796 2970 1822
rect 2997 1796 3013 1822
rect 2653 1794 3013 1796
rect 3032 1822 3392 1825
rect 3032 1796 3066 1822
rect 3093 1796 3141 1822
rect 3168 1796 3274 1822
rect 3301 1796 3349 1822
rect 3376 1796 3392 1822
rect 3032 1794 3392 1796
rect 3411 1822 3771 1825
rect 3411 1796 3445 1822
rect 3472 1796 3520 1822
rect 3547 1796 3653 1822
rect 3680 1796 3728 1822
rect 3755 1796 3771 1822
rect 3411 1794 3771 1796
rect 3790 1822 4150 1825
rect 3790 1796 3824 1822
rect 3851 1796 3899 1822
rect 3926 1796 4032 1822
rect 4059 1796 4107 1822
rect 4134 1796 4150 1822
rect 3790 1794 4150 1796
rect 4169 1822 4529 1825
rect 4169 1796 4203 1822
rect 4230 1796 4278 1822
rect 4305 1796 4411 1822
rect 4438 1796 4486 1822
rect 4513 1796 4529 1822
rect 4169 1794 4529 1796
rect 4548 1822 4908 1825
rect 4548 1796 4582 1822
rect 4609 1796 4657 1822
rect 4684 1796 4790 1822
rect 4817 1796 4865 1822
rect 4892 1796 4908 1822
rect 4548 1794 4908 1796
rect 4927 1822 5287 1825
rect 4927 1796 4961 1822
rect 4988 1796 5036 1822
rect 5063 1796 5169 1822
rect 5196 1796 5244 1822
rect 5271 1796 5287 1822
rect 4927 1794 5287 1796
rect 5306 1822 5666 1825
rect 5306 1796 5340 1822
rect 5367 1796 5415 1822
rect 5442 1796 5548 1822
rect 5575 1796 5623 1822
rect 5650 1796 5666 1822
rect 5306 1794 5666 1796
rect 5685 1822 6045 1825
rect 5685 1796 5719 1822
rect 5746 1796 5794 1822
rect 5821 1796 5927 1822
rect 5954 1796 6002 1822
rect 6029 1796 6045 1822
rect 5685 1794 6045 1796
rect 6064 1822 6424 1825
rect 6064 1796 6098 1822
rect 6125 1796 6173 1822
rect 6200 1796 6306 1822
rect 6333 1796 6381 1822
rect 6408 1796 6424 1822
rect 6064 1794 6424 1796
rect 6443 1822 6803 1825
rect 6443 1796 6477 1822
rect 6504 1796 6552 1822
rect 6579 1796 6685 1822
rect 6712 1796 6760 1822
rect 6787 1796 6803 1822
rect 6443 1794 6803 1796
rect 6822 1822 7182 1825
rect 6822 1796 6856 1822
rect 6883 1796 6931 1822
rect 6958 1796 7064 1822
rect 7091 1796 7139 1822
rect 7166 1796 7182 1822
rect 6822 1794 7182 1796
rect 7201 1822 7561 1825
rect 7201 1796 7235 1822
rect 7262 1796 7310 1822
rect 7337 1796 7443 1822
rect 7470 1796 7518 1822
rect 7545 1796 7561 1822
rect 7201 1794 7561 1796
rect 173 1336 205 1342
rect 173 1309 176 1336
rect 202 1309 205 1336
rect 173 1303 205 1309
rect 552 1335 584 1341
rect 552 1308 555 1335
rect 581 1308 584 1335
rect 552 1302 584 1308
rect 931 1333 963 1339
rect 931 1306 934 1333
rect 960 1306 963 1333
rect 931 1300 963 1306
rect 1310 1331 1342 1337
rect 1310 1304 1313 1331
rect 1339 1304 1342 1331
rect 1310 1298 1342 1304
rect 1689 1331 1721 1337
rect 1689 1304 1692 1331
rect 1718 1304 1721 1331
rect 1689 1298 1721 1304
rect 2068 1336 2100 1342
rect 2068 1309 2071 1336
rect 2097 1309 2100 1336
rect 2068 1303 2100 1309
rect 2447 1335 2479 1341
rect 2447 1308 2450 1335
rect 2476 1308 2479 1335
rect 2447 1302 2479 1308
rect 2826 1333 2858 1339
rect 2826 1306 2829 1333
rect 2855 1306 2858 1333
rect 2826 1300 2858 1306
rect 3205 1331 3237 1337
rect 3205 1304 3208 1331
rect 3234 1304 3237 1331
rect 3205 1298 3237 1304
rect 3584 1331 3616 1337
rect 3584 1304 3587 1331
rect 3613 1304 3616 1331
rect 3584 1298 3616 1304
rect 3963 1336 3995 1342
rect 3963 1309 3966 1336
rect 3992 1309 3995 1336
rect 3963 1303 3995 1309
rect 4342 1335 4374 1341
rect 4342 1308 4345 1335
rect 4371 1308 4374 1335
rect 4342 1302 4374 1308
rect 4721 1333 4753 1339
rect 4721 1306 4724 1333
rect 4750 1306 4753 1333
rect 4721 1300 4753 1306
rect 5100 1331 5132 1337
rect 5100 1304 5103 1331
rect 5129 1304 5132 1331
rect 5100 1298 5132 1304
rect 5479 1331 5511 1337
rect 5479 1304 5482 1331
rect 5508 1304 5511 1331
rect 5479 1298 5511 1304
rect 5858 1336 5890 1342
rect 5858 1309 5861 1336
rect 5887 1309 5890 1336
rect 5858 1303 5890 1309
rect 6237 1335 6269 1341
rect 6237 1308 6240 1335
rect 6266 1308 6269 1335
rect 6237 1302 6269 1308
rect 6480 1222 6535 1336
rect 6616 1333 6648 1339
rect 6616 1306 6619 1333
rect 6645 1306 6648 1333
rect 6616 1300 6648 1306
rect 6995 1331 7027 1337
rect 6995 1304 6998 1331
rect 7024 1304 7027 1331
rect 6995 1298 7027 1304
rect 7374 1331 7406 1337
rect 7374 1304 7377 1331
rect 7403 1304 7406 1331
rect 7374 1298 7406 1304
rect 0 1219 360 1222
rect 0 1193 34 1219
rect 61 1193 109 1219
rect 136 1193 242 1219
rect 269 1193 317 1219
rect 344 1193 360 1219
rect 0 1191 360 1193
rect 379 1219 739 1222
rect 379 1193 413 1219
rect 440 1193 488 1219
rect 515 1193 621 1219
rect 648 1193 696 1219
rect 723 1193 739 1219
rect 379 1191 739 1193
rect 758 1219 1118 1222
rect 758 1193 792 1219
rect 819 1193 867 1219
rect 894 1193 1000 1219
rect 1027 1193 1075 1219
rect 1102 1193 1118 1219
rect 758 1191 1118 1193
rect 1137 1219 1497 1222
rect 1137 1193 1171 1219
rect 1198 1193 1246 1219
rect 1273 1193 1379 1219
rect 1406 1193 1454 1219
rect 1481 1193 1497 1219
rect 1137 1191 1497 1193
rect 1516 1219 1876 1222
rect 1516 1193 1550 1219
rect 1577 1193 1625 1219
rect 1652 1193 1758 1219
rect 1785 1193 1833 1219
rect 1860 1193 1876 1219
rect 1516 1191 1876 1193
rect 1895 1219 2255 1222
rect 1895 1193 1929 1219
rect 1956 1193 2004 1219
rect 2031 1193 2137 1219
rect 2164 1193 2212 1219
rect 2239 1193 2255 1219
rect 1895 1191 2255 1193
rect 2274 1219 2634 1222
rect 2274 1193 2308 1219
rect 2335 1193 2383 1219
rect 2410 1193 2516 1219
rect 2543 1193 2591 1219
rect 2618 1193 2634 1219
rect 2274 1191 2634 1193
rect 2653 1219 3013 1222
rect 2653 1193 2687 1219
rect 2714 1193 2762 1219
rect 2789 1193 2895 1219
rect 2922 1193 2970 1219
rect 2997 1193 3013 1219
rect 2653 1191 3013 1193
rect 3032 1219 3392 1222
rect 3032 1193 3066 1219
rect 3093 1193 3141 1219
rect 3168 1193 3274 1219
rect 3301 1193 3349 1219
rect 3376 1193 3392 1219
rect 3032 1191 3392 1193
rect 3411 1219 3771 1222
rect 3411 1193 3445 1219
rect 3472 1193 3520 1219
rect 3547 1193 3653 1219
rect 3680 1193 3728 1219
rect 3755 1193 3771 1219
rect 3411 1191 3771 1193
rect 3790 1219 4150 1222
rect 3790 1193 3824 1219
rect 3851 1193 3899 1219
rect 3926 1193 4032 1219
rect 4059 1193 4107 1219
rect 4134 1193 4150 1219
rect 3790 1191 4150 1193
rect 4169 1219 4529 1222
rect 4169 1193 4203 1219
rect 4230 1193 4278 1219
rect 4305 1193 4411 1219
rect 4438 1193 4486 1219
rect 4513 1193 4529 1219
rect 4169 1191 4529 1193
rect 4548 1219 4908 1222
rect 4548 1193 4582 1219
rect 4609 1193 4657 1219
rect 4684 1193 4790 1219
rect 4817 1193 4865 1219
rect 4892 1193 4908 1219
rect 4548 1191 4908 1193
rect 4927 1219 5287 1222
rect 4927 1193 4961 1219
rect 4988 1193 5036 1219
rect 5063 1193 5169 1219
rect 5196 1193 5244 1219
rect 5271 1193 5287 1219
rect 4927 1191 5287 1193
rect 5306 1219 5666 1222
rect 5306 1193 5340 1219
rect 5367 1193 5415 1219
rect 5442 1193 5548 1219
rect 5575 1193 5623 1219
rect 5650 1193 5666 1219
rect 5306 1191 5666 1193
rect 5685 1219 6045 1222
rect 5685 1193 5719 1219
rect 5746 1193 5794 1219
rect 5821 1193 5927 1219
rect 5954 1193 6002 1219
rect 6029 1193 6045 1219
rect 5685 1191 6045 1193
rect 6064 1219 6424 1222
rect 6064 1193 6098 1219
rect 6125 1193 6173 1219
rect 6200 1193 6306 1219
rect 6333 1193 6381 1219
rect 6408 1193 6424 1219
rect 6064 1191 6424 1193
rect 6443 1219 6803 1222
rect 6443 1193 6477 1219
rect 6504 1193 6552 1219
rect 6579 1193 6685 1219
rect 6712 1193 6760 1219
rect 6787 1193 6803 1219
rect 6443 1191 6803 1193
rect 6822 1219 7182 1222
rect 6822 1193 6856 1219
rect 6883 1193 6931 1219
rect 6958 1193 7064 1219
rect 7091 1193 7139 1219
rect 7166 1193 7182 1219
rect 6822 1191 7182 1193
rect 7201 1219 7561 1222
rect 7201 1193 7235 1219
rect 7262 1193 7310 1219
rect 7337 1193 7443 1219
rect 7470 1193 7518 1219
rect 7545 1193 7561 1219
rect 7201 1191 7561 1193
rect 552 723 584 729
rect 173 717 205 723
rect 173 690 176 717
rect 202 690 205 717
rect 552 696 555 723
rect 581 696 584 723
rect 552 690 584 696
rect 931 723 963 729
rect 931 696 934 723
rect 960 696 963 723
rect 931 690 963 696
rect 1310 723 1342 729
rect 1310 696 1313 723
rect 1339 696 1342 723
rect 1310 690 1342 696
rect 1689 724 1721 730
rect 1689 697 1692 724
rect 1718 697 1721 724
rect 2447 723 2479 729
rect 1689 691 1721 697
rect 2068 717 2100 723
rect 2068 690 2071 717
rect 2097 690 2100 717
rect 2447 696 2450 723
rect 2476 696 2479 723
rect 2447 690 2479 696
rect 2826 723 2858 729
rect 2826 696 2829 723
rect 2855 696 2858 723
rect 2826 690 2858 696
rect 3205 723 3237 729
rect 3205 696 3208 723
rect 3234 696 3237 723
rect 3205 690 3237 696
rect 3584 724 3616 730
rect 3584 697 3587 724
rect 3613 697 3616 724
rect 4342 723 4374 729
rect 3584 691 3616 697
rect 3963 717 3995 723
rect 3963 690 3966 717
rect 3992 690 3995 717
rect 4342 696 4345 723
rect 4371 696 4374 723
rect 4342 690 4374 696
rect 4721 723 4753 729
rect 4721 696 4724 723
rect 4750 696 4753 723
rect 4721 690 4753 696
rect 5100 723 5132 729
rect 5100 696 5103 723
rect 5129 696 5132 723
rect 5100 690 5132 696
rect 5479 724 5511 730
rect 5479 697 5482 724
rect 5508 697 5511 724
rect 6237 723 6269 729
rect 5479 691 5511 697
rect 5858 717 5890 723
rect 5858 690 5861 717
rect 5887 690 5890 717
rect 6237 696 6240 723
rect 6266 696 6269 723
rect 6480 699 6535 1191
rect 6616 723 6648 729
rect 6237 690 6269 696
rect 6616 696 6619 723
rect 6645 696 6648 723
rect 6616 690 6648 696
rect 6995 723 7027 729
rect 6995 696 6998 723
rect 7024 696 7027 723
rect 6995 690 7027 696
rect 7374 724 7406 730
rect 7374 697 7377 724
rect 7403 697 7406 724
rect 7374 691 7406 697
rect 173 684 205 690
rect 2068 684 2100 690
rect 3963 684 3995 690
rect 5858 684 5890 690
rect 0 616 360 619
rect 0 590 34 616
rect 61 590 109 616
rect 136 590 242 616
rect 269 590 317 616
rect 344 590 360 616
rect 0 588 360 590
rect 379 616 739 619
rect 379 590 413 616
rect 440 590 488 616
rect 515 590 621 616
rect 648 590 696 616
rect 723 590 739 616
rect 379 588 739 590
rect 758 616 1118 619
rect 758 590 792 616
rect 819 590 867 616
rect 894 590 1000 616
rect 1027 590 1075 616
rect 1102 590 1118 616
rect 758 588 1118 590
rect 1137 616 1497 619
rect 1137 590 1171 616
rect 1198 590 1246 616
rect 1273 590 1379 616
rect 1406 590 1454 616
rect 1481 590 1497 616
rect 1137 588 1497 590
rect 1516 616 1876 619
rect 1516 590 1550 616
rect 1577 590 1625 616
rect 1652 590 1758 616
rect 1785 590 1833 616
rect 1860 590 1876 616
rect 1516 588 1876 590
rect 1895 616 2255 619
rect 1895 590 1929 616
rect 1956 590 2004 616
rect 2031 590 2137 616
rect 2164 590 2212 616
rect 2239 590 2255 616
rect 1895 588 2255 590
rect 2274 616 2634 619
rect 2274 590 2308 616
rect 2335 590 2383 616
rect 2410 590 2516 616
rect 2543 590 2591 616
rect 2618 590 2634 616
rect 2274 588 2634 590
rect 2653 616 3013 619
rect 2653 590 2687 616
rect 2714 590 2762 616
rect 2789 590 2895 616
rect 2922 590 2970 616
rect 2997 590 3013 616
rect 2653 588 3013 590
rect 3032 616 3392 619
rect 3032 590 3066 616
rect 3093 590 3141 616
rect 3168 590 3274 616
rect 3301 590 3349 616
rect 3376 590 3392 616
rect 3032 588 3392 590
rect 3411 616 3771 619
rect 3411 590 3445 616
rect 3472 590 3520 616
rect 3547 590 3653 616
rect 3680 590 3728 616
rect 3755 590 3771 616
rect 3411 588 3771 590
rect 3790 616 4150 619
rect 3790 590 3824 616
rect 3851 590 3899 616
rect 3926 590 4032 616
rect 4059 590 4107 616
rect 4134 590 4150 616
rect 3790 588 4150 590
rect 4169 616 4529 619
rect 4169 590 4203 616
rect 4230 590 4278 616
rect 4305 590 4411 616
rect 4438 590 4486 616
rect 4513 590 4529 616
rect 4169 588 4529 590
rect 4548 616 4908 619
rect 4548 590 4582 616
rect 4609 590 4657 616
rect 4684 590 4790 616
rect 4817 590 4865 616
rect 4892 590 4908 616
rect 4548 588 4908 590
rect 4927 616 5287 619
rect 4927 590 4961 616
rect 4988 590 5036 616
rect 5063 590 5169 616
rect 5196 590 5244 616
rect 5271 590 5287 616
rect 4927 588 5287 590
rect 5306 616 5666 619
rect 5306 590 5340 616
rect 5367 590 5415 616
rect 5442 590 5548 616
rect 5575 590 5623 616
rect 5650 590 5666 616
rect 5306 588 5666 590
rect 5685 616 6045 619
rect 5685 590 5719 616
rect 5746 590 5794 616
rect 5821 590 5927 616
rect 5954 590 6002 616
rect 6029 590 6045 616
rect 5685 588 6045 590
rect 6064 616 6424 619
rect 6064 590 6098 616
rect 6125 590 6173 616
rect 6200 590 6306 616
rect 6333 590 6381 616
rect 6408 590 6424 616
rect 6064 588 6424 590
rect 6443 616 6803 619
rect 6443 590 6477 616
rect 6504 590 6552 616
rect 6579 590 6685 616
rect 6712 590 6760 616
rect 6787 590 6803 616
rect 6443 588 6803 590
rect 6822 616 7182 619
rect 6822 590 6856 616
rect 6883 590 6931 616
rect 6958 590 7064 616
rect 7091 590 7139 616
rect 7166 590 7182 616
rect 6822 588 7182 590
rect 7201 616 7561 619
rect 7201 590 7235 616
rect 7262 590 7310 616
rect 7337 590 7443 616
rect 7470 590 7518 616
rect 7545 590 7561 616
rect 7201 588 7561 590
rect 173 511 205 517
rect 173 484 176 511
rect 202 484 205 511
rect 173 478 205 484
rect 552 511 584 517
rect 552 484 555 511
rect 581 484 584 511
rect 552 478 584 484
rect 931 511 963 517
rect 931 484 934 511
rect 960 484 963 511
rect 931 478 963 484
rect 1310 511 1342 517
rect 1310 484 1313 511
rect 1339 484 1342 511
rect 1310 478 1342 484
rect 1689 510 1721 516
rect 1689 483 1692 510
rect 1718 483 1721 510
rect 1689 477 1721 483
rect 2068 511 2100 517
rect 2068 484 2071 511
rect 2097 484 2100 511
rect 2068 478 2100 484
rect 2447 513 2479 519
rect 2447 486 2450 513
rect 2476 486 2479 513
rect 2447 480 2479 486
rect 2826 509 2858 515
rect 2826 482 2829 509
rect 2855 482 2858 509
rect 2826 476 2858 482
rect 3205 505 3237 511
rect 3205 478 3208 505
rect 3234 478 3237 505
rect 3205 472 3237 478
rect 3584 510 3616 516
rect 3584 483 3587 510
rect 3613 483 3616 510
rect 3584 477 3616 483
rect 3963 511 3995 517
rect 3963 484 3966 511
rect 3992 484 3995 511
rect 3963 478 3995 484
rect 4342 506 4374 512
rect 4342 479 4345 506
rect 4371 479 4374 506
rect 4342 473 4374 479
rect 4721 506 4753 512
rect 4721 479 4724 506
rect 4750 479 4753 506
rect 4721 473 4753 479
rect 5100 507 5132 513
rect 5100 480 5103 507
rect 5129 480 5132 507
rect 5100 474 5132 480
rect 5479 510 5511 516
rect 5479 483 5482 510
rect 5508 483 5511 510
rect 5479 477 5511 483
rect 5858 511 5890 517
rect 5858 484 5861 511
rect 5887 484 5890 511
rect 5858 478 5890 484
rect 6237 510 6269 516
rect 6237 483 6240 510
rect 6266 483 6269 510
rect 6237 477 6269 483
rect 6616 513 6648 519
rect 6616 486 6619 513
rect 6645 486 6648 513
rect 6616 480 6648 486
rect 6995 510 7027 516
rect 6995 483 6998 510
rect 7024 483 7027 510
rect 6995 477 7027 483
rect 7374 510 7406 516
rect 7374 483 7377 510
rect 7403 483 7406 510
rect 7374 477 7406 483
rect 0 13 360 16
rect 0 -13 34 13
rect 61 -13 109 13
rect 136 -13 242 13
rect 269 -13 317 13
rect 344 -13 360 13
rect 0 -15 360 -13
rect 379 13 739 16
rect 379 -13 413 13
rect 440 -13 488 13
rect 515 -13 621 13
rect 648 -13 696 13
rect 723 -13 739 13
rect 379 -15 739 -13
rect 758 13 1118 16
rect 758 -13 792 13
rect 819 -13 867 13
rect 894 -13 1000 13
rect 1027 -13 1075 13
rect 1102 -13 1118 13
rect 758 -15 1118 -13
rect 1137 13 1497 16
rect 1137 -13 1171 13
rect 1198 -13 1246 13
rect 1273 -13 1379 13
rect 1406 -13 1454 13
rect 1481 -13 1497 13
rect 1137 -15 1497 -13
rect 1516 13 1876 16
rect 1516 -13 1550 13
rect 1577 -13 1625 13
rect 1652 -13 1758 13
rect 1785 -13 1833 13
rect 1860 -13 1876 13
rect 1516 -15 1876 -13
rect 1895 13 2255 16
rect 1895 -13 1929 13
rect 1956 -13 2004 13
rect 2031 -13 2137 13
rect 2164 -13 2212 13
rect 2239 -13 2255 13
rect 1895 -15 2255 -13
rect 2274 13 2634 16
rect 2274 -13 2308 13
rect 2335 -13 2383 13
rect 2410 -13 2516 13
rect 2543 -13 2591 13
rect 2618 -13 2634 13
rect 2274 -15 2634 -13
rect 2653 13 3013 16
rect 2653 -13 2687 13
rect 2714 -13 2762 13
rect 2789 -13 2895 13
rect 2922 -13 2970 13
rect 2997 -13 3013 13
rect 2653 -15 3013 -13
rect 3032 13 3392 16
rect 3032 -13 3066 13
rect 3093 -13 3141 13
rect 3168 -13 3274 13
rect 3301 -13 3349 13
rect 3376 -13 3392 13
rect 3032 -15 3392 -13
rect 3411 13 3771 16
rect 3411 -13 3445 13
rect 3472 -13 3520 13
rect 3547 -13 3653 13
rect 3680 -13 3728 13
rect 3755 -13 3771 13
rect 3411 -15 3771 -13
rect 3790 13 4150 16
rect 3790 -13 3824 13
rect 3851 -13 3899 13
rect 3926 -13 4032 13
rect 4059 -13 4107 13
rect 4134 -13 4150 13
rect 3790 -15 4150 -13
rect 4169 13 4529 16
rect 4169 -13 4203 13
rect 4230 -13 4278 13
rect 4305 -13 4411 13
rect 4438 -13 4486 13
rect 4513 -13 4529 13
rect 4169 -15 4529 -13
rect 4548 13 4908 16
rect 4548 -13 4582 13
rect 4609 -13 4657 13
rect 4684 -13 4790 13
rect 4817 -13 4865 13
rect 4892 -13 4908 13
rect 4548 -15 4908 -13
rect 4927 13 5287 16
rect 4927 -13 4961 13
rect 4988 -13 5036 13
rect 5063 -13 5169 13
rect 5196 -13 5244 13
rect 5271 -13 5287 13
rect 4927 -15 5287 -13
rect 5306 13 5666 16
rect 5306 -13 5340 13
rect 5367 -13 5415 13
rect 5442 -13 5548 13
rect 5575 -13 5623 13
rect 5650 -13 5666 13
rect 5306 -15 5666 -13
rect 5685 13 6045 16
rect 5685 -13 5719 13
rect 5746 -13 5794 13
rect 5821 -13 5927 13
rect 5954 -13 6002 13
rect 6029 -13 6045 13
rect 5685 -15 6045 -13
rect 6064 13 6424 16
rect 6064 -13 6098 13
rect 6125 -13 6173 13
rect 6200 -13 6306 13
rect 6333 -13 6381 13
rect 6408 -13 6424 13
rect 6064 -15 6424 -13
rect 6443 13 6803 16
rect 6443 -13 6477 13
rect 6504 -13 6552 13
rect 6579 -13 6685 13
rect 6712 -13 6760 13
rect 6787 -13 6803 13
rect 6443 -15 6803 -13
rect 6822 13 7182 16
rect 6822 -13 6856 13
rect 6883 -13 6931 13
rect 6958 -13 7064 13
rect 7091 -13 7139 13
rect 7166 -13 7182 13
rect 6822 -15 7182 -13
rect 7201 13 7561 16
rect 7201 -13 7235 13
rect 7262 -13 7310 13
rect 7337 -13 7443 13
rect 7470 -13 7518 13
rect 7545 -13 7561 13
rect 7201 -15 7561 -13
<< via1 >>
rect 34 2399 61 2425
rect 109 2399 136 2425
rect 242 2399 269 2425
rect 317 2399 344 2425
rect 413 2399 440 2425
rect 488 2399 515 2425
rect 621 2399 648 2425
rect 696 2399 723 2425
rect 792 2399 819 2425
rect 867 2399 894 2425
rect 1000 2399 1027 2425
rect 1075 2399 1102 2425
rect 1171 2399 1198 2425
rect 1246 2399 1273 2425
rect 1379 2399 1406 2425
rect 1454 2399 1481 2425
rect 1550 2399 1577 2425
rect 1625 2399 1652 2425
rect 1758 2399 1785 2425
rect 1833 2399 1860 2425
rect 1929 2399 1956 2425
rect 2004 2399 2031 2425
rect 2137 2399 2164 2425
rect 2212 2399 2239 2425
rect 2308 2399 2335 2425
rect 2383 2399 2410 2425
rect 2516 2399 2543 2425
rect 2591 2399 2618 2425
rect 2687 2399 2714 2425
rect 2762 2399 2789 2425
rect 2895 2399 2922 2425
rect 2970 2399 2997 2425
rect 3066 2399 3093 2425
rect 3141 2399 3168 2425
rect 3274 2399 3301 2425
rect 3349 2399 3376 2425
rect 3445 2399 3472 2425
rect 3520 2399 3547 2425
rect 3653 2399 3680 2425
rect 3728 2399 3755 2425
rect 3824 2399 3851 2425
rect 3899 2399 3926 2425
rect 4032 2399 4059 2425
rect 4107 2399 4134 2425
rect 4203 2399 4230 2425
rect 4278 2399 4305 2425
rect 4411 2399 4438 2425
rect 4486 2399 4513 2425
rect 4582 2399 4609 2425
rect 4657 2399 4684 2425
rect 4790 2399 4817 2425
rect 4865 2399 4892 2425
rect 4961 2399 4988 2425
rect 5036 2399 5063 2425
rect 5169 2399 5196 2425
rect 5244 2399 5271 2425
rect 5340 2399 5367 2425
rect 5415 2399 5442 2425
rect 5548 2399 5575 2425
rect 5623 2399 5650 2425
rect 5719 2399 5746 2425
rect 5794 2399 5821 2425
rect 5927 2399 5954 2425
rect 6002 2399 6029 2425
rect 6109 2412 6136 2425
rect 6184 2412 6211 2425
rect 6317 2412 6344 2425
rect 6392 2412 6419 2425
rect 6098 2399 6136 2412
rect 6173 2399 6211 2412
rect 6306 2399 6344 2412
rect 6381 2399 6419 2412
rect 6488 2412 6515 2425
rect 6563 2412 6590 2425
rect 6696 2412 6723 2425
rect 6771 2412 6798 2425
rect 6477 2399 6515 2412
rect 6552 2399 6590 2412
rect 6685 2399 6723 2412
rect 6760 2399 6798 2412
rect 6867 2412 6894 2425
rect 6942 2412 6969 2425
rect 7075 2412 7102 2425
rect 7150 2412 7177 2425
rect 6856 2399 6894 2412
rect 6931 2399 6969 2412
rect 7064 2399 7102 2412
rect 7139 2399 7177 2412
rect 7235 2399 7262 2425
rect 7310 2399 7337 2425
rect 7443 2399 7470 2425
rect 7518 2399 7545 2425
rect 176 1902 202 1929
rect 555 1902 581 1929
rect 934 1902 960 1929
rect 1313 1902 1339 1929
rect 1692 1901 1718 1928
rect 2071 1902 2097 1929
rect 2450 1902 2476 1929
rect 2829 1902 2855 1929
rect 3208 1902 3234 1929
rect 3587 1901 3613 1928
rect 3966 1902 3992 1929
rect 4345 1902 4371 1929
rect 4724 1902 4750 1929
rect 5103 1902 5129 1929
rect 5482 1901 5508 1928
rect 5861 1902 5887 1929
rect 6240 1902 6266 1929
rect 6619 1902 6645 1929
rect 6998 1902 7024 1929
rect 7377 1901 7403 1928
rect 34 1796 61 1822
rect 109 1796 136 1822
rect 242 1796 269 1822
rect 317 1796 344 1822
rect 413 1796 440 1822
rect 488 1796 515 1822
rect 621 1796 648 1822
rect 696 1796 723 1822
rect 792 1796 819 1822
rect 867 1796 894 1822
rect 1000 1796 1027 1822
rect 1075 1796 1102 1822
rect 1171 1796 1198 1822
rect 1246 1796 1273 1822
rect 1379 1796 1406 1822
rect 1454 1796 1481 1822
rect 1550 1796 1577 1822
rect 1625 1796 1652 1822
rect 1758 1796 1785 1822
rect 1833 1796 1860 1822
rect 1929 1796 1956 1822
rect 2004 1796 2031 1822
rect 2137 1796 2164 1822
rect 2212 1796 2239 1822
rect 2308 1796 2335 1822
rect 2383 1796 2410 1822
rect 2516 1796 2543 1822
rect 2591 1796 2618 1822
rect 2687 1796 2714 1822
rect 2762 1796 2789 1822
rect 2895 1796 2922 1822
rect 2970 1796 2997 1822
rect 3066 1796 3093 1822
rect 3141 1796 3168 1822
rect 3274 1796 3301 1822
rect 3349 1796 3376 1822
rect 3445 1796 3472 1822
rect 3520 1796 3547 1822
rect 3653 1796 3680 1822
rect 3728 1796 3755 1822
rect 3824 1796 3851 1822
rect 3899 1796 3926 1822
rect 4032 1796 4059 1822
rect 4107 1796 4134 1822
rect 4203 1796 4230 1822
rect 4278 1796 4305 1822
rect 4411 1796 4438 1822
rect 4486 1796 4513 1822
rect 4582 1796 4609 1822
rect 4657 1796 4684 1822
rect 4790 1796 4817 1822
rect 4865 1796 4892 1822
rect 4961 1796 4988 1822
rect 5036 1796 5063 1822
rect 5169 1796 5196 1822
rect 5244 1796 5271 1822
rect 5340 1796 5367 1822
rect 5415 1796 5442 1822
rect 5548 1796 5575 1822
rect 5623 1796 5650 1822
rect 5719 1796 5746 1822
rect 5794 1796 5821 1822
rect 5927 1796 5954 1822
rect 6002 1796 6029 1822
rect 6098 1796 6125 1822
rect 6173 1796 6200 1822
rect 6306 1796 6333 1822
rect 6381 1796 6408 1822
rect 6477 1796 6504 1822
rect 6552 1796 6579 1822
rect 6685 1796 6712 1822
rect 6760 1796 6787 1822
rect 6856 1796 6883 1822
rect 6931 1796 6958 1822
rect 7064 1796 7091 1822
rect 7139 1796 7166 1822
rect 7235 1796 7262 1822
rect 7310 1796 7337 1822
rect 7443 1796 7470 1822
rect 7518 1796 7545 1822
rect 176 1309 202 1336
rect 555 1308 581 1335
rect 934 1306 960 1333
rect 1313 1304 1339 1331
rect 1692 1304 1718 1331
rect 2071 1309 2097 1336
rect 2450 1308 2476 1335
rect 2829 1306 2855 1333
rect 3208 1304 3234 1331
rect 3587 1304 3613 1331
rect 3966 1309 3992 1336
rect 4345 1308 4371 1335
rect 4724 1306 4750 1333
rect 5103 1304 5129 1331
rect 5482 1304 5508 1331
rect 5861 1309 5887 1336
rect 6240 1308 6266 1335
rect 6619 1306 6645 1333
rect 6998 1304 7024 1331
rect 7377 1304 7403 1331
rect 34 1193 61 1219
rect 109 1193 136 1219
rect 242 1193 269 1219
rect 317 1193 344 1219
rect 413 1193 440 1219
rect 488 1193 515 1219
rect 621 1193 648 1219
rect 696 1193 723 1219
rect 792 1193 819 1219
rect 867 1193 894 1219
rect 1000 1193 1027 1219
rect 1075 1193 1102 1219
rect 1171 1193 1198 1219
rect 1246 1193 1273 1219
rect 1379 1193 1406 1219
rect 1454 1193 1481 1219
rect 1550 1193 1577 1219
rect 1625 1193 1652 1219
rect 1758 1193 1785 1219
rect 1833 1193 1860 1219
rect 1929 1193 1956 1219
rect 2004 1193 2031 1219
rect 2137 1193 2164 1219
rect 2212 1193 2239 1219
rect 2308 1193 2335 1219
rect 2383 1193 2410 1219
rect 2516 1193 2543 1219
rect 2591 1193 2618 1219
rect 2687 1193 2714 1219
rect 2762 1193 2789 1219
rect 2895 1193 2922 1219
rect 2970 1193 2997 1219
rect 3066 1193 3093 1219
rect 3141 1193 3168 1219
rect 3274 1193 3301 1219
rect 3349 1193 3376 1219
rect 3445 1193 3472 1219
rect 3520 1193 3547 1219
rect 3653 1193 3680 1219
rect 3728 1193 3755 1219
rect 3824 1193 3851 1219
rect 3899 1193 3926 1219
rect 4032 1193 4059 1219
rect 4107 1193 4134 1219
rect 4203 1193 4230 1219
rect 4278 1193 4305 1219
rect 4411 1193 4438 1219
rect 4486 1193 4513 1219
rect 4582 1193 4609 1219
rect 4657 1193 4684 1219
rect 4790 1193 4817 1219
rect 4865 1193 4892 1219
rect 4961 1193 4988 1219
rect 5036 1193 5063 1219
rect 5169 1193 5196 1219
rect 5244 1193 5271 1219
rect 5340 1193 5367 1219
rect 5415 1193 5442 1219
rect 5548 1193 5575 1219
rect 5623 1193 5650 1219
rect 5719 1193 5746 1219
rect 5794 1193 5821 1219
rect 5927 1193 5954 1219
rect 6002 1193 6029 1219
rect 6098 1193 6125 1219
rect 6173 1193 6200 1219
rect 6306 1193 6333 1219
rect 6381 1193 6408 1219
rect 6477 1193 6504 1219
rect 6552 1193 6579 1219
rect 6685 1193 6712 1219
rect 6760 1193 6787 1219
rect 6856 1193 6883 1219
rect 6931 1193 6958 1219
rect 7064 1193 7091 1219
rect 7139 1193 7166 1219
rect 7235 1193 7262 1219
rect 7310 1193 7337 1219
rect 7443 1193 7470 1219
rect 7518 1193 7545 1219
rect 176 690 202 717
rect 555 696 581 723
rect 934 696 960 723
rect 1313 696 1339 723
rect 1692 697 1718 724
rect 2071 690 2097 717
rect 2450 696 2476 723
rect 2829 696 2855 723
rect 3208 696 3234 723
rect 3587 697 3613 724
rect 3966 690 3992 717
rect 4345 696 4371 723
rect 4724 696 4750 723
rect 5103 696 5129 723
rect 5482 697 5508 724
rect 5861 690 5887 717
rect 6240 696 6266 723
rect 6619 696 6645 723
rect 6998 696 7024 723
rect 7377 697 7403 724
rect 34 590 61 616
rect 109 590 136 616
rect 242 590 269 616
rect 317 590 344 616
rect 413 590 440 616
rect 488 590 515 616
rect 621 590 648 616
rect 696 590 723 616
rect 792 590 819 616
rect 867 590 894 616
rect 1000 590 1027 616
rect 1075 590 1102 616
rect 1171 590 1198 616
rect 1246 590 1273 616
rect 1379 590 1406 616
rect 1454 590 1481 616
rect 1550 590 1577 616
rect 1625 590 1652 616
rect 1758 590 1785 616
rect 1833 590 1860 616
rect 1929 590 1956 616
rect 2004 590 2031 616
rect 2137 590 2164 616
rect 2212 590 2239 616
rect 2308 590 2335 616
rect 2383 590 2410 616
rect 2516 590 2543 616
rect 2591 590 2618 616
rect 2687 590 2714 616
rect 2762 590 2789 616
rect 2895 590 2922 616
rect 2970 590 2997 616
rect 3066 590 3093 616
rect 3141 590 3168 616
rect 3274 590 3301 616
rect 3349 590 3376 616
rect 3445 590 3472 616
rect 3520 590 3547 616
rect 3653 590 3680 616
rect 3728 590 3755 616
rect 3824 590 3851 616
rect 3899 590 3926 616
rect 4032 590 4059 616
rect 4107 590 4134 616
rect 4203 590 4230 616
rect 4278 590 4305 616
rect 4411 590 4438 616
rect 4486 590 4513 616
rect 4582 590 4609 616
rect 4657 590 4684 616
rect 4790 590 4817 616
rect 4865 590 4892 616
rect 4961 590 4988 616
rect 5036 590 5063 616
rect 5169 590 5196 616
rect 5244 590 5271 616
rect 5340 590 5367 616
rect 5415 590 5442 616
rect 5548 590 5575 616
rect 5623 590 5650 616
rect 5719 590 5746 616
rect 5794 590 5821 616
rect 5927 590 5954 616
rect 6002 590 6029 616
rect 6098 590 6125 616
rect 6173 590 6200 616
rect 6306 590 6333 616
rect 6381 590 6408 616
rect 6477 590 6504 616
rect 6552 590 6579 616
rect 6685 590 6712 616
rect 6760 590 6787 616
rect 6856 590 6883 616
rect 6931 590 6958 616
rect 7064 590 7091 616
rect 7139 590 7166 616
rect 7235 590 7262 616
rect 7310 590 7337 616
rect 7443 590 7470 616
rect 7518 590 7545 616
rect 176 484 202 511
rect 555 484 581 511
rect 934 484 960 511
rect 1313 484 1339 511
rect 1692 483 1718 510
rect 2071 484 2097 511
rect 2450 486 2476 513
rect 2829 482 2855 509
rect 3208 478 3234 505
rect 3587 483 3613 510
rect 3966 484 3992 511
rect 4345 479 4371 506
rect 4724 479 4750 506
rect 5103 480 5129 507
rect 5482 483 5508 510
rect 5861 484 5887 511
rect 6240 483 6266 510
rect 6619 486 6645 513
rect 6998 483 7024 510
rect 7377 483 7403 510
rect 34 -13 61 13
rect 109 -13 136 13
rect 242 -13 269 13
rect 317 -13 344 13
rect 413 -13 440 13
rect 488 -13 515 13
rect 621 -13 648 13
rect 696 -13 723 13
rect 792 -13 819 13
rect 867 -13 894 13
rect 1000 -13 1027 13
rect 1075 -13 1102 13
rect 1171 -13 1198 13
rect 1246 -13 1273 13
rect 1379 -13 1406 13
rect 1454 -13 1481 13
rect 1550 -13 1577 13
rect 1625 -13 1652 13
rect 1758 -13 1785 13
rect 1833 -13 1860 13
rect 1929 -13 1956 13
rect 2004 -13 2031 13
rect 2137 -13 2164 13
rect 2212 -13 2239 13
rect 2308 -13 2335 13
rect 2383 -13 2410 13
rect 2516 -13 2543 13
rect 2591 -13 2618 13
rect 2687 -13 2714 13
rect 2762 -13 2789 13
rect 2895 -13 2922 13
rect 2970 -13 2997 13
rect 3066 -13 3093 13
rect 3141 -13 3168 13
rect 3274 -13 3301 13
rect 3349 -13 3376 13
rect 3445 -13 3472 13
rect 3520 -13 3547 13
rect 3653 -13 3680 13
rect 3728 -13 3755 13
rect 3824 -13 3851 13
rect 3899 -13 3926 13
rect 4032 -13 4059 13
rect 4107 -13 4134 13
rect 4203 -13 4230 13
rect 4278 -13 4305 13
rect 4411 -13 4438 13
rect 4486 -13 4513 13
rect 4582 -13 4609 13
rect 4657 -13 4684 13
rect 4790 -13 4817 13
rect 4865 -13 4892 13
rect 4961 -13 4988 13
rect 5036 -13 5063 13
rect 5169 -13 5196 13
rect 5244 -13 5271 13
rect 5340 -13 5367 13
rect 5415 -13 5442 13
rect 5548 -13 5575 13
rect 5623 -13 5650 13
rect 5719 -13 5746 13
rect 5794 -13 5821 13
rect 5927 -13 5954 13
rect 6002 -13 6029 13
rect 6098 -13 6125 13
rect 6173 -13 6200 13
rect 6306 -13 6333 13
rect 6381 -13 6408 13
rect 6477 -13 6504 13
rect 6552 -13 6579 13
rect 6685 -13 6712 13
rect 6760 -13 6787 13
rect 6856 -13 6883 13
rect 6931 -13 6958 13
rect 7064 -13 7091 13
rect 7139 -13 7166 13
rect 7235 -13 7262 13
rect 7310 -13 7337 13
rect 7443 -13 7470 13
rect 7518 -13 7545 13
<< metal2 >>
rect -19 2425 7599 2428
rect -19 2399 34 2425
rect 61 2399 109 2425
rect 136 2399 242 2425
rect 269 2399 317 2425
rect 344 2399 413 2425
rect 440 2399 488 2425
rect 515 2399 621 2425
rect 648 2399 696 2425
rect 723 2399 792 2425
rect 819 2399 867 2425
rect 894 2399 1000 2425
rect 1027 2399 1075 2425
rect 1102 2399 1171 2425
rect 1198 2399 1246 2425
rect 1273 2399 1379 2425
rect 1406 2399 1454 2425
rect 1481 2399 1550 2425
rect 1577 2399 1625 2425
rect 1652 2399 1758 2425
rect 1785 2399 1833 2425
rect 1860 2399 1929 2425
rect 1956 2399 2004 2425
rect 2031 2399 2137 2425
rect 2164 2399 2212 2425
rect 2239 2399 2308 2425
rect 2335 2399 2383 2425
rect 2410 2399 2516 2425
rect 2543 2399 2591 2425
rect 2618 2399 2687 2425
rect 2714 2399 2762 2425
rect 2789 2399 2895 2425
rect 2922 2399 2970 2425
rect 2997 2399 3066 2425
rect 3093 2399 3141 2425
rect 3168 2399 3274 2425
rect 3301 2399 3349 2425
rect 3376 2399 3445 2425
rect 3472 2399 3520 2425
rect 3547 2399 3653 2425
rect 3680 2399 3728 2425
rect 3755 2399 3824 2425
rect 3851 2399 3899 2425
rect 3926 2399 4032 2425
rect 4059 2399 4107 2425
rect 4134 2399 4203 2425
rect 4230 2399 4278 2425
rect 4305 2399 4411 2425
rect 4438 2399 4486 2425
rect 4513 2399 4582 2425
rect 4609 2399 4657 2425
rect 4684 2399 4790 2425
rect 4817 2399 4865 2425
rect 4892 2399 4961 2425
rect 4988 2399 5036 2425
rect 5063 2399 5169 2425
rect 5196 2399 5244 2425
rect 5271 2399 5340 2425
rect 5367 2399 5415 2425
rect 5442 2399 5548 2425
rect 5575 2399 5623 2425
rect 5650 2399 5719 2425
rect 5746 2399 5794 2425
rect 5821 2399 5927 2425
rect 5954 2399 6002 2425
rect 6029 2412 6109 2425
rect 6136 2412 6184 2425
rect 6211 2412 6317 2425
rect 6344 2412 6392 2425
rect 6419 2412 6488 2425
rect 6515 2412 6563 2425
rect 6590 2412 6696 2425
rect 6723 2412 6771 2425
rect 6798 2412 6867 2425
rect 6894 2412 6942 2425
rect 6969 2412 7075 2425
rect 7102 2412 7150 2425
rect 6029 2399 6098 2412
rect 6136 2399 6173 2412
rect 6211 2399 6306 2412
rect 6344 2399 6381 2412
rect 6419 2399 6477 2412
rect 6515 2399 6552 2412
rect 6590 2399 6685 2412
rect 6723 2399 6760 2412
rect 6798 2399 6856 2412
rect 6894 2399 6931 2412
rect 6969 2399 7064 2412
rect 7102 2399 7139 2412
rect 7177 2399 7235 2425
rect 7262 2399 7310 2425
rect 7337 2399 7443 2425
rect 7470 2399 7518 2425
rect 7545 2399 7599 2425
rect -19 2396 7599 2399
rect -19 2385 161 2396
rect 217 2385 540 2396
rect 596 2385 919 2396
rect 975 2385 1298 2396
rect 1354 2385 1677 2396
rect 1733 2385 2056 2396
rect 2112 2385 2435 2396
rect 2491 2385 2814 2396
rect 2870 2385 3193 2396
rect 3249 2385 3572 2396
rect 3628 2385 3951 2396
rect 4007 2385 4330 2396
rect 4386 2385 4709 2396
rect 4765 2385 5088 2396
rect 5144 2385 5467 2396
rect 5523 2385 5846 2396
rect 5902 2385 6225 2396
rect 6281 2385 6604 2396
rect 6660 2385 6983 2396
rect 7039 2385 7362 2396
rect 7418 2385 7599 2396
rect -19 2317 146 2385
rect 175 2370 203 2382
rect 161 2367 217 2370
rect 161 2336 166 2367
rect 212 2336 217 2367
rect 161 2332 217 2336
rect -19 2264 161 2317
rect -19 2196 146 2264
rect 175 2249 203 2332
rect 232 2317 525 2385
rect 554 2370 582 2382
rect 540 2367 596 2370
rect 540 2336 545 2367
rect 591 2336 596 2367
rect 540 2332 596 2336
rect 217 2264 540 2317
rect 161 2246 217 2249
rect 161 2215 166 2246
rect 212 2215 217 2246
rect 161 2211 217 2215
rect -19 2144 161 2196
rect -19 2076 146 2144
rect 175 2129 203 2211
rect 232 2196 525 2264
rect 554 2249 582 2332
rect 611 2317 904 2385
rect 933 2370 961 2382
rect 919 2367 975 2370
rect 919 2336 924 2367
rect 970 2336 975 2367
rect 919 2332 975 2336
rect 596 2264 919 2317
rect 540 2246 596 2249
rect 540 2215 545 2246
rect 591 2215 596 2246
rect 540 2211 596 2215
rect 217 2144 540 2196
rect 161 2126 217 2129
rect 161 2095 166 2126
rect 212 2095 217 2126
rect 161 2091 217 2095
rect -19 2024 161 2076
rect -19 1956 146 2024
rect 175 2009 203 2091
rect 232 2076 525 2144
rect 554 2129 582 2211
rect 611 2196 904 2264
rect 933 2249 961 2332
rect 990 2317 1283 2385
rect 1312 2370 1340 2382
rect 1298 2367 1354 2370
rect 1298 2336 1303 2367
rect 1349 2336 1354 2367
rect 1298 2332 1354 2336
rect 975 2264 1298 2317
rect 919 2246 975 2249
rect 919 2215 924 2246
rect 970 2215 975 2246
rect 919 2211 975 2215
rect 596 2144 919 2196
rect 540 2126 596 2129
rect 540 2095 545 2126
rect 591 2095 596 2126
rect 540 2091 596 2095
rect 217 2024 540 2076
rect 161 2006 217 2009
rect 161 1975 166 2006
rect 212 1975 217 2006
rect 161 1971 217 1975
rect -19 1904 161 1956
rect 175 1929 203 1971
rect 232 1956 525 2024
rect 554 2009 582 2091
rect 611 2076 904 2144
rect 933 2129 961 2211
rect 990 2196 1283 2264
rect 1312 2249 1340 2332
rect 1369 2317 1662 2385
rect 1691 2370 1719 2382
rect 1677 2367 1733 2370
rect 1677 2336 1682 2367
rect 1728 2336 1733 2367
rect 1677 2332 1733 2336
rect 1354 2264 1677 2317
rect 1298 2246 1354 2249
rect 1298 2215 1303 2246
rect 1349 2215 1354 2246
rect 1298 2211 1354 2215
rect 975 2144 1298 2196
rect 919 2126 975 2129
rect 919 2095 924 2126
rect 970 2095 975 2126
rect 919 2091 975 2095
rect 596 2024 919 2076
rect 540 2006 596 2009
rect 540 1975 545 2006
rect 591 1975 596 2006
rect 540 1971 596 1975
rect -19 1837 146 1904
rect 175 1902 176 1929
rect 202 1902 203 1929
rect 217 1904 540 1956
rect 554 1929 582 1971
rect 611 1956 904 2024
rect 933 2009 961 2091
rect 990 2076 1283 2144
rect 1312 2129 1340 2211
rect 1369 2196 1662 2264
rect 1691 2249 1719 2332
rect 1748 2317 2041 2385
rect 2070 2370 2098 2382
rect 2056 2367 2112 2370
rect 2056 2336 2061 2367
rect 2107 2336 2112 2367
rect 2056 2332 2112 2336
rect 1733 2264 2056 2317
rect 1677 2246 1733 2249
rect 1677 2215 1682 2246
rect 1728 2215 1733 2246
rect 1677 2211 1733 2215
rect 1354 2144 1677 2196
rect 1298 2126 1354 2129
rect 1298 2095 1303 2126
rect 1349 2095 1354 2126
rect 1298 2091 1354 2095
rect 975 2024 1298 2076
rect 919 2006 975 2009
rect 919 1975 924 2006
rect 970 1975 975 2006
rect 919 1971 975 1975
rect 175 1889 203 1902
rect 161 1886 217 1889
rect 161 1855 166 1886
rect 212 1855 217 1886
rect 161 1851 217 1855
rect 175 1839 203 1851
rect 232 1837 525 1904
rect 554 1902 555 1929
rect 581 1902 582 1929
rect 596 1904 919 1956
rect 933 1929 961 1971
rect 990 1956 1283 2024
rect 1312 2009 1340 2091
rect 1369 2076 1662 2144
rect 1691 2129 1719 2211
rect 1748 2196 2041 2264
rect 2070 2249 2098 2332
rect 2127 2317 2420 2385
rect 2449 2370 2477 2382
rect 2435 2367 2491 2370
rect 2435 2336 2440 2367
rect 2486 2336 2491 2367
rect 2435 2332 2491 2336
rect 2112 2264 2435 2317
rect 2056 2246 2112 2249
rect 2056 2215 2061 2246
rect 2107 2215 2112 2246
rect 2056 2211 2112 2215
rect 1733 2144 2056 2196
rect 1677 2126 1733 2129
rect 1677 2095 1682 2126
rect 1728 2095 1733 2126
rect 1677 2091 1733 2095
rect 1354 2024 1677 2076
rect 1298 2006 1354 2009
rect 1298 1975 1303 2006
rect 1349 1975 1354 2006
rect 1298 1971 1354 1975
rect 554 1889 582 1902
rect 540 1886 596 1889
rect 540 1855 545 1886
rect 591 1855 596 1886
rect 540 1851 596 1855
rect 554 1839 582 1851
rect 611 1837 904 1904
rect 933 1902 934 1929
rect 960 1902 961 1929
rect 975 1904 1298 1956
rect 1312 1929 1340 1971
rect 1369 1956 1662 2024
rect 1691 2009 1719 2091
rect 1748 2076 2041 2144
rect 2070 2129 2098 2211
rect 2127 2196 2420 2264
rect 2449 2249 2477 2332
rect 2506 2317 2799 2385
rect 2828 2370 2856 2382
rect 2814 2367 2870 2370
rect 2814 2336 2819 2367
rect 2865 2336 2870 2367
rect 2814 2332 2870 2336
rect 2491 2264 2814 2317
rect 2435 2246 2491 2249
rect 2435 2215 2440 2246
rect 2486 2215 2491 2246
rect 2435 2211 2491 2215
rect 2112 2144 2435 2196
rect 2056 2126 2112 2129
rect 2056 2095 2061 2126
rect 2107 2095 2112 2126
rect 2056 2091 2112 2095
rect 1733 2024 2056 2076
rect 1677 2006 1733 2009
rect 1677 1975 1682 2006
rect 1728 1975 1733 2006
rect 1677 1971 1733 1975
rect 933 1889 961 1902
rect 919 1886 975 1889
rect 919 1855 924 1886
rect 970 1855 975 1886
rect 919 1851 975 1855
rect 933 1839 961 1851
rect 990 1837 1283 1904
rect 1312 1902 1313 1929
rect 1339 1902 1340 1929
rect 1354 1904 1677 1956
rect 1691 1928 1719 1971
rect 1748 1956 2041 2024
rect 2070 2009 2098 2091
rect 2127 2076 2420 2144
rect 2449 2129 2477 2211
rect 2506 2196 2799 2264
rect 2828 2249 2856 2332
rect 2885 2317 3178 2385
rect 3207 2370 3235 2382
rect 3193 2367 3249 2370
rect 3193 2336 3198 2367
rect 3244 2336 3249 2367
rect 3193 2332 3249 2336
rect 2870 2264 3193 2317
rect 2814 2246 2870 2249
rect 2814 2215 2819 2246
rect 2865 2215 2870 2246
rect 2814 2211 2870 2215
rect 2491 2144 2814 2196
rect 2435 2126 2491 2129
rect 2435 2095 2440 2126
rect 2486 2095 2491 2126
rect 2435 2091 2491 2095
rect 2112 2024 2435 2076
rect 2056 2006 2112 2009
rect 2056 1975 2061 2006
rect 2107 1975 2112 2006
rect 2056 1971 2112 1975
rect 1312 1889 1340 1902
rect 1298 1886 1354 1889
rect 1298 1855 1303 1886
rect 1349 1855 1354 1886
rect 1298 1851 1354 1855
rect 1312 1839 1340 1851
rect 1369 1837 1662 1904
rect 1691 1901 1692 1928
rect 1718 1901 1719 1928
rect 1733 1904 2056 1956
rect 2070 1929 2098 1971
rect 2127 1956 2420 2024
rect 2449 2009 2477 2091
rect 2506 2076 2799 2144
rect 2828 2129 2856 2211
rect 2885 2196 3178 2264
rect 3207 2249 3235 2332
rect 3264 2317 3557 2385
rect 3586 2370 3614 2382
rect 3572 2367 3628 2370
rect 3572 2336 3577 2367
rect 3623 2336 3628 2367
rect 3572 2332 3628 2336
rect 3249 2264 3572 2317
rect 3193 2246 3249 2249
rect 3193 2215 3198 2246
rect 3244 2215 3249 2246
rect 3193 2211 3249 2215
rect 2870 2144 3193 2196
rect 2814 2126 2870 2129
rect 2814 2095 2819 2126
rect 2865 2095 2870 2126
rect 2814 2091 2870 2095
rect 2491 2024 2814 2076
rect 2435 2006 2491 2009
rect 2435 1975 2440 2006
rect 2486 1975 2491 2006
rect 2435 1971 2491 1975
rect 1691 1889 1719 1901
rect 1677 1886 1733 1889
rect 1677 1855 1682 1886
rect 1728 1855 1733 1886
rect 1677 1851 1733 1855
rect 1691 1839 1719 1851
rect 1748 1837 2041 1904
rect 2070 1902 2071 1929
rect 2097 1902 2098 1929
rect 2112 1904 2435 1956
rect 2449 1929 2477 1971
rect 2506 1956 2799 2024
rect 2828 2009 2856 2091
rect 2885 2076 3178 2144
rect 3207 2129 3235 2211
rect 3264 2196 3557 2264
rect 3586 2249 3614 2332
rect 3643 2317 3936 2385
rect 3965 2370 3993 2382
rect 3951 2367 4007 2370
rect 3951 2336 3956 2367
rect 4002 2336 4007 2367
rect 3951 2332 4007 2336
rect 3628 2264 3951 2317
rect 3572 2246 3628 2249
rect 3572 2215 3577 2246
rect 3623 2215 3628 2246
rect 3572 2211 3628 2215
rect 3249 2144 3572 2196
rect 3193 2126 3249 2129
rect 3193 2095 3198 2126
rect 3244 2095 3249 2126
rect 3193 2091 3249 2095
rect 2870 2024 3193 2076
rect 2814 2006 2870 2009
rect 2814 1975 2819 2006
rect 2865 1975 2870 2006
rect 2814 1971 2870 1975
rect 2070 1889 2098 1902
rect 2056 1886 2112 1889
rect 2056 1855 2061 1886
rect 2107 1855 2112 1886
rect 2056 1851 2112 1855
rect 2070 1839 2098 1851
rect 2127 1837 2420 1904
rect 2449 1902 2450 1929
rect 2476 1902 2477 1929
rect 2491 1904 2814 1956
rect 2828 1929 2856 1971
rect 2885 1956 3178 2024
rect 3207 2009 3235 2091
rect 3264 2076 3557 2144
rect 3586 2129 3614 2211
rect 3643 2196 3936 2264
rect 3965 2249 3993 2332
rect 4022 2317 4315 2385
rect 4344 2370 4372 2382
rect 4330 2367 4386 2370
rect 4330 2336 4335 2367
rect 4381 2336 4386 2367
rect 4330 2332 4386 2336
rect 4007 2264 4330 2317
rect 3951 2246 4007 2249
rect 3951 2215 3956 2246
rect 4002 2215 4007 2246
rect 3951 2211 4007 2215
rect 3628 2144 3951 2196
rect 3572 2126 3628 2129
rect 3572 2095 3577 2126
rect 3623 2095 3628 2126
rect 3572 2091 3628 2095
rect 3249 2024 3572 2076
rect 3193 2006 3249 2009
rect 3193 1975 3198 2006
rect 3244 1975 3249 2006
rect 3193 1971 3249 1975
rect 2449 1889 2477 1902
rect 2435 1886 2491 1889
rect 2435 1855 2440 1886
rect 2486 1855 2491 1886
rect 2435 1851 2491 1855
rect 2449 1839 2477 1851
rect 2506 1837 2799 1904
rect 2828 1902 2829 1929
rect 2855 1902 2856 1929
rect 2870 1904 3193 1956
rect 3207 1929 3235 1971
rect 3264 1956 3557 2024
rect 3586 2009 3614 2091
rect 3643 2076 3936 2144
rect 3965 2129 3993 2211
rect 4022 2196 4315 2264
rect 4344 2249 4372 2332
rect 4401 2317 4694 2385
rect 4723 2370 4751 2382
rect 4709 2367 4765 2370
rect 4709 2336 4714 2367
rect 4760 2336 4765 2367
rect 4709 2332 4765 2336
rect 4386 2264 4709 2317
rect 4330 2246 4386 2249
rect 4330 2215 4335 2246
rect 4381 2215 4386 2246
rect 4330 2211 4386 2215
rect 4007 2144 4330 2196
rect 3951 2126 4007 2129
rect 3951 2095 3956 2126
rect 4002 2095 4007 2126
rect 3951 2091 4007 2095
rect 3628 2024 3951 2076
rect 3572 2006 3628 2009
rect 3572 1975 3577 2006
rect 3623 1975 3628 2006
rect 3572 1971 3628 1975
rect 2828 1889 2856 1902
rect 2814 1886 2870 1889
rect 2814 1855 2819 1886
rect 2865 1855 2870 1886
rect 2814 1851 2870 1855
rect 2828 1839 2856 1851
rect 2885 1837 3178 1904
rect 3207 1902 3208 1929
rect 3234 1902 3235 1929
rect 3249 1904 3572 1956
rect 3586 1928 3614 1971
rect 3643 1956 3936 2024
rect 3965 2009 3993 2091
rect 4022 2076 4315 2144
rect 4344 2129 4372 2211
rect 4401 2196 4694 2264
rect 4723 2249 4751 2332
rect 4780 2317 5073 2385
rect 5102 2370 5130 2382
rect 5088 2367 5144 2370
rect 5088 2336 5093 2367
rect 5139 2336 5144 2367
rect 5088 2332 5144 2336
rect 4765 2264 5088 2317
rect 4709 2246 4765 2249
rect 4709 2215 4714 2246
rect 4760 2215 4765 2246
rect 4709 2211 4765 2215
rect 4386 2144 4709 2196
rect 4330 2126 4386 2129
rect 4330 2095 4335 2126
rect 4381 2095 4386 2126
rect 4330 2091 4386 2095
rect 4007 2024 4330 2076
rect 3951 2006 4007 2009
rect 3951 1975 3956 2006
rect 4002 1975 4007 2006
rect 3951 1971 4007 1975
rect 3207 1889 3235 1902
rect 3193 1886 3249 1889
rect 3193 1855 3198 1886
rect 3244 1855 3249 1886
rect 3193 1851 3249 1855
rect 3207 1839 3235 1851
rect 3264 1837 3557 1904
rect 3586 1901 3587 1928
rect 3613 1901 3614 1928
rect 3628 1904 3951 1956
rect 3965 1929 3993 1971
rect 4022 1956 4315 2024
rect 4344 2009 4372 2091
rect 4401 2076 4694 2144
rect 4723 2129 4751 2211
rect 4780 2196 5073 2264
rect 5102 2249 5130 2332
rect 5159 2317 5452 2385
rect 5481 2370 5509 2382
rect 5467 2367 5523 2370
rect 5467 2336 5472 2367
rect 5518 2336 5523 2367
rect 5467 2332 5523 2336
rect 5144 2264 5467 2317
rect 5088 2246 5144 2249
rect 5088 2215 5093 2246
rect 5139 2215 5144 2246
rect 5088 2211 5144 2215
rect 4765 2144 5088 2196
rect 4709 2126 4765 2129
rect 4709 2095 4714 2126
rect 4760 2095 4765 2126
rect 4709 2091 4765 2095
rect 4386 2024 4709 2076
rect 4330 2006 4386 2009
rect 4330 1975 4335 2006
rect 4381 1975 4386 2006
rect 4330 1971 4386 1975
rect 3586 1889 3614 1901
rect 3572 1886 3628 1889
rect 3572 1855 3577 1886
rect 3623 1855 3628 1886
rect 3572 1851 3628 1855
rect 3586 1839 3614 1851
rect 3643 1837 3936 1904
rect 3965 1902 3966 1929
rect 3992 1902 3993 1929
rect 4007 1904 4330 1956
rect 4344 1929 4372 1971
rect 4401 1956 4694 2024
rect 4723 2009 4751 2091
rect 4780 2076 5073 2144
rect 5102 2129 5130 2211
rect 5159 2196 5452 2264
rect 5481 2249 5509 2332
rect 5538 2317 5831 2385
rect 5860 2370 5888 2382
rect 5846 2367 5902 2370
rect 5846 2336 5851 2367
rect 5897 2336 5902 2367
rect 5846 2332 5902 2336
rect 5523 2264 5846 2317
rect 5467 2246 5523 2249
rect 5467 2215 5472 2246
rect 5518 2215 5523 2246
rect 5467 2211 5523 2215
rect 5144 2144 5467 2196
rect 5088 2126 5144 2129
rect 5088 2095 5093 2126
rect 5139 2095 5144 2126
rect 5088 2091 5144 2095
rect 4765 2024 5088 2076
rect 4709 2006 4765 2009
rect 4709 1975 4714 2006
rect 4760 1975 4765 2006
rect 4709 1971 4765 1975
rect 3965 1889 3993 1902
rect 3951 1886 4007 1889
rect 3951 1855 3956 1886
rect 4002 1855 4007 1886
rect 3951 1851 4007 1855
rect 3965 1839 3993 1851
rect 4022 1837 4315 1904
rect 4344 1902 4345 1929
rect 4371 1902 4372 1929
rect 4386 1904 4709 1956
rect 4723 1929 4751 1971
rect 4780 1956 5073 2024
rect 5102 2009 5130 2091
rect 5159 2076 5452 2144
rect 5481 2129 5509 2211
rect 5538 2196 5831 2264
rect 5860 2249 5888 2332
rect 5917 2317 6210 2385
rect 6239 2370 6267 2382
rect 6225 2367 6281 2370
rect 6225 2336 6230 2367
rect 6276 2336 6281 2367
rect 6225 2332 6281 2336
rect 5902 2264 6225 2317
rect 5846 2246 5902 2249
rect 5846 2215 5851 2246
rect 5897 2215 5902 2246
rect 5846 2211 5902 2215
rect 5523 2144 5846 2196
rect 5467 2126 5523 2129
rect 5467 2095 5472 2126
rect 5518 2095 5523 2126
rect 5467 2091 5523 2095
rect 5144 2024 5467 2076
rect 5088 2006 5144 2009
rect 5088 1975 5093 2006
rect 5139 1975 5144 2006
rect 5088 1971 5144 1975
rect 4344 1889 4372 1902
rect 4330 1886 4386 1889
rect 4330 1855 4335 1886
rect 4381 1855 4386 1886
rect 4330 1851 4386 1855
rect 4344 1839 4372 1851
rect 4401 1837 4694 1904
rect 4723 1902 4724 1929
rect 4750 1902 4751 1929
rect 4765 1904 5088 1956
rect 5102 1929 5130 1971
rect 5159 1956 5452 2024
rect 5481 2009 5509 2091
rect 5538 2076 5831 2144
rect 5860 2129 5888 2211
rect 5917 2196 6210 2264
rect 6239 2249 6267 2332
rect 6296 2317 6589 2385
rect 6618 2370 6646 2382
rect 6604 2367 6660 2370
rect 6604 2336 6609 2367
rect 6655 2336 6660 2367
rect 6604 2332 6660 2336
rect 6281 2264 6604 2317
rect 6225 2246 6281 2249
rect 6225 2215 6230 2246
rect 6276 2215 6281 2246
rect 6225 2211 6281 2215
rect 5902 2144 6225 2196
rect 5846 2126 5902 2129
rect 5846 2095 5851 2126
rect 5897 2095 5902 2126
rect 5846 2091 5902 2095
rect 5523 2024 5846 2076
rect 5467 2006 5523 2009
rect 5467 1975 5472 2006
rect 5518 1975 5523 2006
rect 5467 1971 5523 1975
rect 4723 1889 4751 1902
rect 4709 1886 4765 1889
rect 4709 1855 4714 1886
rect 4760 1855 4765 1886
rect 4709 1851 4765 1855
rect 4723 1839 4751 1851
rect 4780 1837 5073 1904
rect 5102 1902 5103 1929
rect 5129 1902 5130 1929
rect 5144 1904 5467 1956
rect 5481 1928 5509 1971
rect 5538 1956 5831 2024
rect 5860 2009 5888 2091
rect 5917 2076 6210 2144
rect 6239 2129 6267 2211
rect 6296 2196 6589 2264
rect 6618 2249 6646 2332
rect 6675 2317 6968 2385
rect 6997 2370 7025 2382
rect 6983 2367 7039 2370
rect 6983 2336 6988 2367
rect 7034 2336 7039 2367
rect 6983 2332 7039 2336
rect 6660 2264 6983 2317
rect 6604 2246 6660 2249
rect 6604 2215 6609 2246
rect 6655 2215 6660 2246
rect 6604 2211 6660 2215
rect 6281 2144 6604 2196
rect 6225 2126 6281 2129
rect 6225 2095 6230 2126
rect 6276 2095 6281 2126
rect 6225 2091 6281 2095
rect 5902 2024 6225 2076
rect 5846 2006 5902 2009
rect 5846 1975 5851 2006
rect 5897 1975 5902 2006
rect 5846 1971 5902 1975
rect 5102 1889 5130 1902
rect 5088 1886 5144 1889
rect 5088 1855 5093 1886
rect 5139 1855 5144 1886
rect 5088 1851 5144 1855
rect 5102 1839 5130 1851
rect 5159 1837 5452 1904
rect 5481 1901 5482 1928
rect 5508 1901 5509 1928
rect 5523 1904 5846 1956
rect 5860 1929 5888 1971
rect 5917 1956 6210 2024
rect 6239 2009 6267 2091
rect 6296 2076 6589 2144
rect 6618 2129 6646 2211
rect 6675 2196 6968 2264
rect 6997 2249 7025 2332
rect 7054 2317 7347 2385
rect 7376 2370 7404 2382
rect 7362 2367 7418 2370
rect 7362 2336 7367 2367
rect 7413 2336 7418 2367
rect 7362 2332 7418 2336
rect 7039 2264 7362 2317
rect 6983 2246 7039 2249
rect 6983 2215 6988 2246
rect 7034 2215 7039 2246
rect 6983 2211 7039 2215
rect 6660 2144 6983 2196
rect 6604 2126 6660 2129
rect 6604 2095 6609 2126
rect 6655 2095 6660 2126
rect 6604 2091 6660 2095
rect 6281 2024 6604 2076
rect 6225 2006 6281 2009
rect 6225 1975 6230 2006
rect 6276 1975 6281 2006
rect 6225 1971 6281 1975
rect 5481 1889 5509 1901
rect 5467 1886 5523 1889
rect 5467 1855 5472 1886
rect 5518 1855 5523 1886
rect 5467 1851 5523 1855
rect 5481 1839 5509 1851
rect 5538 1837 5831 1904
rect 5860 1902 5861 1929
rect 5887 1902 5888 1929
rect 5902 1904 6225 1956
rect 6239 1929 6267 1971
rect 6296 1956 6589 2024
rect 6618 2009 6646 2091
rect 6675 2076 6968 2144
rect 6997 2129 7025 2211
rect 7054 2196 7347 2264
rect 7376 2249 7404 2332
rect 7433 2317 7599 2385
rect 7418 2264 7599 2317
rect 7362 2246 7418 2249
rect 7362 2215 7367 2246
rect 7413 2215 7418 2246
rect 7362 2211 7418 2215
rect 7039 2144 7362 2196
rect 6983 2126 7039 2129
rect 6983 2095 6988 2126
rect 7034 2095 7039 2126
rect 6983 2091 7039 2095
rect 6660 2024 6983 2076
rect 6604 2006 6660 2009
rect 6604 1975 6609 2006
rect 6655 1975 6660 2006
rect 6604 1971 6660 1975
rect 5860 1889 5888 1902
rect 5846 1886 5902 1889
rect 5846 1855 5851 1886
rect 5897 1855 5902 1886
rect 5846 1851 5902 1855
rect 5860 1839 5888 1851
rect 5917 1837 6210 1904
rect 6239 1902 6240 1929
rect 6266 1902 6267 1929
rect 6281 1904 6604 1956
rect 6618 1929 6646 1971
rect 6675 1956 6968 2024
rect 6997 2009 7025 2091
rect 7054 2076 7347 2144
rect 7376 2129 7404 2211
rect 7433 2196 7599 2264
rect 7418 2144 7599 2196
rect 7362 2126 7418 2129
rect 7362 2095 7367 2126
rect 7413 2095 7418 2126
rect 7362 2091 7418 2095
rect 7039 2024 7362 2076
rect 6983 2006 7039 2009
rect 6983 1975 6988 2006
rect 7034 1975 7039 2006
rect 6983 1971 7039 1975
rect 6239 1889 6267 1902
rect 6225 1886 6281 1889
rect 6225 1855 6230 1886
rect 6276 1855 6281 1886
rect 6225 1851 6281 1855
rect 6239 1839 6267 1851
rect 6296 1837 6589 1904
rect 6618 1902 6619 1929
rect 6645 1902 6646 1929
rect 6660 1904 6983 1956
rect 6997 1929 7025 1971
rect 7054 1956 7347 2024
rect 7376 2009 7404 2091
rect 7433 2076 7599 2144
rect 7418 2024 7599 2076
rect 7362 2006 7418 2009
rect 7362 1975 7367 2006
rect 7413 1975 7418 2006
rect 7362 1971 7418 1975
rect 6618 1889 6646 1902
rect 6604 1886 6660 1889
rect 6604 1855 6609 1886
rect 6655 1855 6660 1886
rect 6604 1851 6660 1855
rect 6618 1839 6646 1851
rect 6675 1837 6968 1904
rect 6997 1902 6998 1929
rect 7024 1902 7025 1929
rect 7039 1904 7362 1956
rect 7376 1928 7404 1971
rect 7433 1956 7599 2024
rect 6997 1889 7025 1902
rect 6983 1886 7039 1889
rect 6983 1855 6988 1886
rect 7034 1855 7039 1886
rect 6983 1851 7039 1855
rect 6997 1839 7025 1851
rect 7054 1837 7347 1904
rect 7376 1901 7377 1928
rect 7403 1901 7404 1928
rect 7418 1904 7599 1956
rect 7376 1889 7404 1901
rect 7362 1886 7418 1889
rect 7362 1855 7367 1886
rect 7413 1855 7418 1886
rect 7362 1851 7418 1855
rect 7376 1839 7404 1851
rect 7433 1837 7599 1904
rect -19 1825 161 1837
rect 217 1825 540 1837
rect 596 1825 919 1837
rect 975 1825 1298 1837
rect 1354 1825 1677 1837
rect 1733 1825 2056 1837
rect 2112 1825 2435 1837
rect 2491 1825 2814 1837
rect 2870 1825 3193 1837
rect 3249 1825 3572 1837
rect 3628 1825 3951 1837
rect 4007 1825 4330 1837
rect 4386 1825 4709 1837
rect 4765 1825 5088 1837
rect 5144 1825 5467 1837
rect 5523 1825 5846 1837
rect 5902 1825 6225 1837
rect 6281 1825 6604 1837
rect 6660 1825 6983 1837
rect 7039 1825 7362 1837
rect 7418 1825 7599 1837
rect -19 1822 7599 1825
rect -19 1796 34 1822
rect 61 1796 109 1822
rect 136 1796 242 1822
rect 269 1796 317 1822
rect 344 1796 413 1822
rect 440 1796 488 1822
rect 515 1796 621 1822
rect 648 1796 696 1822
rect 723 1796 792 1822
rect 819 1796 867 1822
rect 894 1796 1000 1822
rect 1027 1796 1075 1822
rect 1102 1796 1171 1822
rect 1198 1796 1246 1822
rect 1273 1796 1379 1822
rect 1406 1796 1454 1822
rect 1481 1796 1550 1822
rect 1577 1796 1625 1822
rect 1652 1796 1758 1822
rect 1785 1796 1833 1822
rect 1860 1796 1929 1822
rect 1956 1796 2004 1822
rect 2031 1796 2137 1822
rect 2164 1796 2212 1822
rect 2239 1796 2308 1822
rect 2335 1796 2383 1822
rect 2410 1796 2516 1822
rect 2543 1796 2591 1822
rect 2618 1796 2687 1822
rect 2714 1796 2762 1822
rect 2789 1796 2895 1822
rect 2922 1796 2970 1822
rect 2997 1796 3066 1822
rect 3093 1796 3141 1822
rect 3168 1796 3274 1822
rect 3301 1796 3349 1822
rect 3376 1796 3445 1822
rect 3472 1796 3520 1822
rect 3547 1796 3653 1822
rect 3680 1796 3728 1822
rect 3755 1796 3824 1822
rect 3851 1796 3899 1822
rect 3926 1796 4032 1822
rect 4059 1796 4107 1822
rect 4134 1796 4203 1822
rect 4230 1796 4278 1822
rect 4305 1796 4411 1822
rect 4438 1796 4486 1822
rect 4513 1796 4582 1822
rect 4609 1796 4657 1822
rect 4684 1796 4790 1822
rect 4817 1796 4865 1822
rect 4892 1796 4961 1822
rect 4988 1796 5036 1822
rect 5063 1796 5169 1822
rect 5196 1796 5244 1822
rect 5271 1796 5340 1822
rect 5367 1796 5415 1822
rect 5442 1796 5548 1822
rect 5575 1796 5623 1822
rect 5650 1796 5719 1822
rect 5746 1796 5794 1822
rect 5821 1796 5927 1822
rect 5954 1796 6002 1822
rect 6029 1796 6098 1822
rect 6125 1796 6173 1822
rect 6200 1796 6306 1822
rect 6333 1796 6381 1822
rect 6408 1796 6477 1822
rect 6504 1796 6552 1822
rect 6579 1796 6685 1822
rect 6712 1796 6760 1822
rect 6787 1796 6856 1822
rect 6883 1796 6931 1822
rect 6958 1796 7064 1822
rect 7091 1796 7139 1822
rect 7166 1796 7235 1822
rect 7262 1796 7310 1822
rect 7337 1796 7443 1822
rect 7470 1796 7518 1822
rect 7545 1796 7599 1822
rect -19 1793 7599 1796
rect -19 1782 161 1793
rect 217 1782 540 1793
rect 596 1782 919 1793
rect 975 1782 1298 1793
rect 1354 1782 1677 1793
rect 1733 1782 2056 1793
rect 2112 1782 2435 1793
rect 2491 1782 2814 1793
rect 2870 1782 3193 1793
rect 3249 1782 3572 1793
rect 3628 1782 3951 1793
rect 4007 1782 4330 1793
rect 4386 1782 4709 1793
rect 4765 1782 5088 1793
rect 5144 1782 5467 1793
rect 5523 1782 5846 1793
rect 5902 1782 6225 1793
rect 6281 1782 6604 1793
rect 6660 1782 6983 1793
rect 7039 1782 7362 1793
rect 7418 1782 7599 1793
rect -19 1714 146 1782
rect 175 1767 203 1779
rect 161 1764 217 1767
rect 161 1733 166 1764
rect 212 1733 217 1764
rect 161 1729 217 1733
rect -19 1661 161 1714
rect -19 1593 146 1661
rect 175 1646 203 1729
rect 232 1714 525 1782
rect 554 1767 582 1779
rect 540 1764 596 1767
rect 540 1733 545 1764
rect 591 1733 596 1764
rect 540 1729 596 1733
rect 217 1661 540 1714
rect 161 1643 217 1646
rect 161 1612 166 1643
rect 212 1612 217 1643
rect 161 1608 217 1612
rect -19 1541 161 1593
rect -19 1473 146 1541
rect 175 1526 203 1608
rect 232 1593 525 1661
rect 554 1646 582 1729
rect 611 1714 904 1782
rect 933 1767 961 1779
rect 919 1764 975 1767
rect 919 1733 924 1764
rect 970 1733 975 1764
rect 919 1729 975 1733
rect 596 1661 919 1714
rect 540 1643 596 1646
rect 540 1612 545 1643
rect 591 1612 596 1643
rect 540 1608 596 1612
rect 217 1541 540 1593
rect 161 1523 217 1526
rect 161 1492 166 1523
rect 212 1492 217 1523
rect 161 1488 217 1492
rect -19 1421 161 1473
rect -19 1353 146 1421
rect 175 1406 203 1488
rect 232 1473 525 1541
rect 554 1526 582 1608
rect 611 1593 904 1661
rect 933 1646 961 1729
rect 990 1714 1283 1782
rect 1312 1767 1340 1779
rect 1298 1764 1354 1767
rect 1298 1733 1303 1764
rect 1349 1733 1354 1764
rect 1298 1729 1354 1733
rect 975 1661 1298 1714
rect 919 1643 975 1646
rect 919 1612 924 1643
rect 970 1612 975 1643
rect 919 1608 975 1612
rect 596 1541 919 1593
rect 540 1523 596 1526
rect 540 1492 545 1523
rect 591 1492 596 1523
rect 540 1488 596 1492
rect 217 1421 540 1473
rect 161 1403 217 1406
rect 161 1372 166 1403
rect 212 1372 217 1403
rect 161 1368 217 1372
rect -19 1301 161 1353
rect 175 1336 203 1368
rect 232 1353 525 1421
rect 554 1406 582 1488
rect 611 1473 904 1541
rect 933 1526 961 1608
rect 990 1593 1283 1661
rect 1312 1646 1340 1729
rect 1369 1714 1662 1782
rect 1691 1767 1719 1779
rect 1677 1764 1733 1767
rect 1677 1733 1682 1764
rect 1728 1733 1733 1764
rect 1677 1729 1733 1733
rect 1354 1661 1677 1714
rect 1298 1643 1354 1646
rect 1298 1612 1303 1643
rect 1349 1612 1354 1643
rect 1298 1608 1354 1612
rect 975 1541 1298 1593
rect 919 1523 975 1526
rect 919 1492 924 1523
rect 970 1492 975 1523
rect 919 1488 975 1492
rect 596 1421 919 1473
rect 540 1403 596 1406
rect 540 1372 545 1403
rect 591 1372 596 1403
rect 540 1368 596 1372
rect 175 1309 176 1336
rect 202 1309 203 1336
rect -19 1234 146 1301
rect 175 1286 203 1309
rect 217 1301 540 1353
rect 554 1335 582 1368
rect 611 1353 904 1421
rect 933 1406 961 1488
rect 990 1473 1283 1541
rect 1312 1526 1340 1608
rect 1369 1593 1662 1661
rect 1691 1646 1719 1729
rect 1748 1714 2041 1782
rect 2070 1767 2098 1779
rect 2056 1764 2112 1767
rect 2056 1733 2061 1764
rect 2107 1733 2112 1764
rect 2056 1729 2112 1733
rect 1733 1661 2056 1714
rect 1677 1643 1733 1646
rect 1677 1612 1682 1643
rect 1728 1612 1733 1643
rect 1677 1608 1733 1612
rect 1354 1541 1677 1593
rect 1298 1523 1354 1526
rect 1298 1492 1303 1523
rect 1349 1492 1354 1523
rect 1298 1488 1354 1492
rect 975 1421 1298 1473
rect 919 1403 975 1406
rect 919 1372 924 1403
rect 970 1372 975 1403
rect 919 1368 975 1372
rect 554 1308 555 1335
rect 581 1308 582 1335
rect 161 1283 217 1286
rect 161 1252 166 1283
rect 212 1252 217 1283
rect 161 1248 217 1252
rect 175 1236 203 1248
rect 232 1234 525 1301
rect 554 1286 582 1308
rect 596 1301 919 1353
rect 933 1333 961 1368
rect 990 1353 1283 1421
rect 1312 1406 1340 1488
rect 1369 1473 1662 1541
rect 1691 1526 1719 1608
rect 1748 1593 2041 1661
rect 2070 1646 2098 1729
rect 2127 1714 2420 1782
rect 2449 1767 2477 1779
rect 2435 1764 2491 1767
rect 2435 1733 2440 1764
rect 2486 1733 2491 1764
rect 2435 1729 2491 1733
rect 2112 1661 2435 1714
rect 2056 1643 2112 1646
rect 2056 1612 2061 1643
rect 2107 1612 2112 1643
rect 2056 1608 2112 1612
rect 1733 1541 2056 1593
rect 1677 1523 1733 1526
rect 1677 1492 1682 1523
rect 1728 1492 1733 1523
rect 1677 1488 1733 1492
rect 1354 1421 1677 1473
rect 1298 1403 1354 1406
rect 1298 1372 1303 1403
rect 1349 1372 1354 1403
rect 1298 1368 1354 1372
rect 933 1306 934 1333
rect 960 1306 961 1333
rect 540 1283 596 1286
rect 540 1252 545 1283
rect 591 1252 596 1283
rect 540 1248 596 1252
rect 554 1236 582 1248
rect 611 1234 904 1301
rect 933 1286 961 1306
rect 975 1301 1298 1353
rect 1312 1331 1340 1368
rect 1369 1353 1662 1421
rect 1691 1406 1719 1488
rect 1748 1473 2041 1541
rect 2070 1526 2098 1608
rect 2127 1593 2420 1661
rect 2449 1646 2477 1729
rect 2506 1714 2799 1782
rect 2828 1767 2856 1779
rect 2814 1764 2870 1767
rect 2814 1733 2819 1764
rect 2865 1733 2870 1764
rect 2814 1729 2870 1733
rect 2491 1661 2814 1714
rect 2435 1643 2491 1646
rect 2435 1612 2440 1643
rect 2486 1612 2491 1643
rect 2435 1608 2491 1612
rect 2112 1541 2435 1593
rect 2056 1523 2112 1526
rect 2056 1492 2061 1523
rect 2107 1492 2112 1523
rect 2056 1488 2112 1492
rect 1733 1421 2056 1473
rect 1677 1403 1733 1406
rect 1677 1372 1682 1403
rect 1728 1372 1733 1403
rect 1677 1368 1733 1372
rect 1312 1304 1313 1331
rect 1339 1304 1340 1331
rect 919 1283 975 1286
rect 919 1252 924 1283
rect 970 1252 975 1283
rect 919 1248 975 1252
rect 933 1236 961 1248
rect 990 1234 1283 1301
rect 1312 1286 1340 1304
rect 1354 1301 1677 1353
rect 1691 1331 1719 1368
rect 1748 1353 2041 1421
rect 2070 1406 2098 1488
rect 2127 1473 2420 1541
rect 2449 1526 2477 1608
rect 2506 1593 2799 1661
rect 2828 1646 2856 1729
rect 2885 1714 3178 1782
rect 3207 1767 3235 1779
rect 3193 1764 3249 1767
rect 3193 1733 3198 1764
rect 3244 1733 3249 1764
rect 3193 1729 3249 1733
rect 2870 1661 3193 1714
rect 2814 1643 2870 1646
rect 2814 1612 2819 1643
rect 2865 1612 2870 1643
rect 2814 1608 2870 1612
rect 2491 1541 2814 1593
rect 2435 1523 2491 1526
rect 2435 1492 2440 1523
rect 2486 1492 2491 1523
rect 2435 1488 2491 1492
rect 2112 1421 2435 1473
rect 2056 1403 2112 1406
rect 2056 1372 2061 1403
rect 2107 1372 2112 1403
rect 2056 1368 2112 1372
rect 1691 1304 1692 1331
rect 1718 1304 1719 1331
rect 1298 1283 1354 1286
rect 1298 1252 1303 1283
rect 1349 1252 1354 1283
rect 1298 1248 1354 1252
rect 1312 1236 1340 1248
rect 1369 1234 1662 1301
rect 1691 1286 1719 1304
rect 1733 1301 2056 1353
rect 2070 1336 2098 1368
rect 2127 1353 2420 1421
rect 2449 1406 2477 1488
rect 2506 1473 2799 1541
rect 2828 1526 2856 1608
rect 2885 1593 3178 1661
rect 3207 1646 3235 1729
rect 3264 1714 3557 1782
rect 3586 1767 3614 1779
rect 3572 1764 3628 1767
rect 3572 1733 3577 1764
rect 3623 1733 3628 1764
rect 3572 1729 3628 1733
rect 3249 1661 3572 1714
rect 3193 1643 3249 1646
rect 3193 1612 3198 1643
rect 3244 1612 3249 1643
rect 3193 1608 3249 1612
rect 2870 1541 3193 1593
rect 2814 1523 2870 1526
rect 2814 1492 2819 1523
rect 2865 1492 2870 1523
rect 2814 1488 2870 1492
rect 2491 1421 2814 1473
rect 2435 1403 2491 1406
rect 2435 1372 2440 1403
rect 2486 1372 2491 1403
rect 2435 1368 2491 1372
rect 2070 1309 2071 1336
rect 2097 1309 2098 1336
rect 1677 1283 1733 1286
rect 1677 1252 1682 1283
rect 1728 1252 1733 1283
rect 1677 1248 1733 1252
rect 1691 1236 1719 1248
rect 1748 1234 2041 1301
rect 2070 1286 2098 1309
rect 2112 1301 2435 1353
rect 2449 1335 2477 1368
rect 2506 1353 2799 1421
rect 2828 1406 2856 1488
rect 2885 1473 3178 1541
rect 3207 1526 3235 1608
rect 3264 1593 3557 1661
rect 3586 1646 3614 1729
rect 3643 1714 3936 1782
rect 3965 1767 3993 1779
rect 3951 1764 4007 1767
rect 3951 1733 3956 1764
rect 4002 1733 4007 1764
rect 3951 1729 4007 1733
rect 3628 1661 3951 1714
rect 3572 1643 3628 1646
rect 3572 1612 3577 1643
rect 3623 1612 3628 1643
rect 3572 1608 3628 1612
rect 3249 1541 3572 1593
rect 3193 1523 3249 1526
rect 3193 1492 3198 1523
rect 3244 1492 3249 1523
rect 3193 1488 3249 1492
rect 2870 1421 3193 1473
rect 2814 1403 2870 1406
rect 2814 1372 2819 1403
rect 2865 1372 2870 1403
rect 2814 1368 2870 1372
rect 2449 1308 2450 1335
rect 2476 1308 2477 1335
rect 2056 1283 2112 1286
rect 2056 1252 2061 1283
rect 2107 1252 2112 1283
rect 2056 1248 2112 1252
rect 2070 1236 2098 1248
rect 2127 1234 2420 1301
rect 2449 1286 2477 1308
rect 2491 1301 2814 1353
rect 2828 1333 2856 1368
rect 2885 1353 3178 1421
rect 3207 1406 3235 1488
rect 3264 1473 3557 1541
rect 3586 1526 3614 1608
rect 3643 1593 3936 1661
rect 3965 1646 3993 1729
rect 4022 1714 4315 1782
rect 4344 1767 4372 1779
rect 4330 1764 4386 1767
rect 4330 1733 4335 1764
rect 4381 1733 4386 1764
rect 4330 1729 4386 1733
rect 4007 1661 4330 1714
rect 3951 1643 4007 1646
rect 3951 1612 3956 1643
rect 4002 1612 4007 1643
rect 3951 1608 4007 1612
rect 3628 1541 3951 1593
rect 3572 1523 3628 1526
rect 3572 1492 3577 1523
rect 3623 1492 3628 1523
rect 3572 1488 3628 1492
rect 3249 1421 3572 1473
rect 3193 1403 3249 1406
rect 3193 1372 3198 1403
rect 3244 1372 3249 1403
rect 3193 1368 3249 1372
rect 2828 1306 2829 1333
rect 2855 1306 2856 1333
rect 2435 1283 2491 1286
rect 2435 1252 2440 1283
rect 2486 1252 2491 1283
rect 2435 1248 2491 1252
rect 2449 1236 2477 1248
rect 2506 1234 2799 1301
rect 2828 1286 2856 1306
rect 2870 1301 3193 1353
rect 3207 1331 3235 1368
rect 3264 1353 3557 1421
rect 3586 1406 3614 1488
rect 3643 1473 3936 1541
rect 3965 1526 3993 1608
rect 4022 1593 4315 1661
rect 4344 1646 4372 1729
rect 4401 1714 4694 1782
rect 4723 1767 4751 1779
rect 4709 1764 4765 1767
rect 4709 1733 4714 1764
rect 4760 1733 4765 1764
rect 4709 1729 4765 1733
rect 4386 1661 4709 1714
rect 4330 1643 4386 1646
rect 4330 1612 4335 1643
rect 4381 1612 4386 1643
rect 4330 1608 4386 1612
rect 4007 1541 4330 1593
rect 3951 1523 4007 1526
rect 3951 1492 3956 1523
rect 4002 1492 4007 1523
rect 3951 1488 4007 1492
rect 3628 1421 3951 1473
rect 3572 1403 3628 1406
rect 3572 1372 3577 1403
rect 3623 1372 3628 1403
rect 3572 1368 3628 1372
rect 3207 1304 3208 1331
rect 3234 1304 3235 1331
rect 2814 1283 2870 1286
rect 2814 1252 2819 1283
rect 2865 1252 2870 1283
rect 2814 1248 2870 1252
rect 2828 1236 2856 1248
rect 2885 1234 3178 1301
rect 3207 1286 3235 1304
rect 3249 1301 3572 1353
rect 3586 1331 3614 1368
rect 3643 1353 3936 1421
rect 3965 1406 3993 1488
rect 4022 1473 4315 1541
rect 4344 1526 4372 1608
rect 4401 1593 4694 1661
rect 4723 1646 4751 1729
rect 4780 1714 5073 1782
rect 5102 1767 5130 1779
rect 5088 1764 5144 1767
rect 5088 1733 5093 1764
rect 5139 1733 5144 1764
rect 5088 1729 5144 1733
rect 4765 1661 5088 1714
rect 4709 1643 4765 1646
rect 4709 1612 4714 1643
rect 4760 1612 4765 1643
rect 4709 1608 4765 1612
rect 4386 1541 4709 1593
rect 4330 1523 4386 1526
rect 4330 1492 4335 1523
rect 4381 1492 4386 1523
rect 4330 1488 4386 1492
rect 4007 1421 4330 1473
rect 3951 1403 4007 1406
rect 3951 1372 3956 1403
rect 4002 1372 4007 1403
rect 3951 1368 4007 1372
rect 3586 1304 3587 1331
rect 3613 1304 3614 1331
rect 3193 1283 3249 1286
rect 3193 1252 3198 1283
rect 3244 1252 3249 1283
rect 3193 1248 3249 1252
rect 3207 1236 3235 1248
rect 3264 1234 3557 1301
rect 3586 1286 3614 1304
rect 3628 1301 3951 1353
rect 3965 1336 3993 1368
rect 4022 1353 4315 1421
rect 4344 1406 4372 1488
rect 4401 1473 4694 1541
rect 4723 1526 4751 1608
rect 4780 1593 5073 1661
rect 5102 1646 5130 1729
rect 5159 1714 5452 1782
rect 5481 1767 5509 1779
rect 5467 1764 5523 1767
rect 5467 1733 5472 1764
rect 5518 1733 5523 1764
rect 5467 1729 5523 1733
rect 5144 1661 5467 1714
rect 5088 1643 5144 1646
rect 5088 1612 5093 1643
rect 5139 1612 5144 1643
rect 5088 1608 5144 1612
rect 4765 1541 5088 1593
rect 4709 1523 4765 1526
rect 4709 1492 4714 1523
rect 4760 1492 4765 1523
rect 4709 1488 4765 1492
rect 4386 1421 4709 1473
rect 4330 1403 4386 1406
rect 4330 1372 4335 1403
rect 4381 1372 4386 1403
rect 4330 1368 4386 1372
rect 3965 1309 3966 1336
rect 3992 1309 3993 1336
rect 3572 1283 3628 1286
rect 3572 1252 3577 1283
rect 3623 1252 3628 1283
rect 3572 1248 3628 1252
rect 3586 1236 3614 1248
rect 3643 1234 3936 1301
rect 3965 1286 3993 1309
rect 4007 1301 4330 1353
rect 4344 1335 4372 1368
rect 4401 1353 4694 1421
rect 4723 1406 4751 1488
rect 4780 1473 5073 1541
rect 5102 1526 5130 1608
rect 5159 1593 5452 1661
rect 5481 1646 5509 1729
rect 5538 1714 5831 1782
rect 5860 1767 5888 1779
rect 5846 1764 5902 1767
rect 5846 1733 5851 1764
rect 5897 1733 5902 1764
rect 5846 1729 5902 1733
rect 5523 1661 5846 1714
rect 5467 1643 5523 1646
rect 5467 1612 5472 1643
rect 5518 1612 5523 1643
rect 5467 1608 5523 1612
rect 5144 1541 5467 1593
rect 5088 1523 5144 1526
rect 5088 1492 5093 1523
rect 5139 1492 5144 1523
rect 5088 1488 5144 1492
rect 4765 1421 5088 1473
rect 4709 1403 4765 1406
rect 4709 1372 4714 1403
rect 4760 1372 4765 1403
rect 4709 1368 4765 1372
rect 4344 1308 4345 1335
rect 4371 1308 4372 1335
rect 3951 1283 4007 1286
rect 3951 1252 3956 1283
rect 4002 1252 4007 1283
rect 3951 1248 4007 1252
rect 3965 1236 3993 1248
rect 4022 1234 4315 1301
rect 4344 1286 4372 1308
rect 4386 1301 4709 1353
rect 4723 1333 4751 1368
rect 4780 1353 5073 1421
rect 5102 1406 5130 1488
rect 5159 1473 5452 1541
rect 5481 1526 5509 1608
rect 5538 1593 5831 1661
rect 5860 1646 5888 1729
rect 5917 1714 6210 1782
rect 6239 1767 6267 1779
rect 6225 1764 6281 1767
rect 6225 1733 6230 1764
rect 6276 1733 6281 1764
rect 6225 1729 6281 1733
rect 5902 1661 6225 1714
rect 5846 1643 5902 1646
rect 5846 1612 5851 1643
rect 5897 1612 5902 1643
rect 5846 1608 5902 1612
rect 5523 1541 5846 1593
rect 5467 1523 5523 1526
rect 5467 1492 5472 1523
rect 5518 1492 5523 1523
rect 5467 1488 5523 1492
rect 5144 1421 5467 1473
rect 5088 1403 5144 1406
rect 5088 1372 5093 1403
rect 5139 1372 5144 1403
rect 5088 1368 5144 1372
rect 4723 1306 4724 1333
rect 4750 1306 4751 1333
rect 4330 1283 4386 1286
rect 4330 1252 4335 1283
rect 4381 1252 4386 1283
rect 4330 1248 4386 1252
rect 4344 1236 4372 1248
rect 4401 1234 4694 1301
rect 4723 1286 4751 1306
rect 4765 1301 5088 1353
rect 5102 1331 5130 1368
rect 5159 1353 5452 1421
rect 5481 1406 5509 1488
rect 5538 1473 5831 1541
rect 5860 1526 5888 1608
rect 5917 1593 6210 1661
rect 6239 1646 6267 1729
rect 6296 1714 6589 1782
rect 6618 1767 6646 1779
rect 6604 1764 6660 1767
rect 6604 1733 6609 1764
rect 6655 1733 6660 1764
rect 6604 1729 6660 1733
rect 6281 1661 6604 1714
rect 6225 1643 6281 1646
rect 6225 1612 6230 1643
rect 6276 1612 6281 1643
rect 6225 1608 6281 1612
rect 5902 1541 6225 1593
rect 5846 1523 5902 1526
rect 5846 1492 5851 1523
rect 5897 1492 5902 1523
rect 5846 1488 5902 1492
rect 5523 1421 5846 1473
rect 5467 1403 5523 1406
rect 5467 1372 5472 1403
rect 5518 1372 5523 1403
rect 5467 1368 5523 1372
rect 5102 1304 5103 1331
rect 5129 1304 5130 1331
rect 4709 1283 4765 1286
rect 4709 1252 4714 1283
rect 4760 1252 4765 1283
rect 4709 1248 4765 1252
rect 4723 1236 4751 1248
rect 4780 1234 5073 1301
rect 5102 1286 5130 1304
rect 5144 1301 5467 1353
rect 5481 1331 5509 1368
rect 5538 1353 5831 1421
rect 5860 1406 5888 1488
rect 5917 1473 6210 1541
rect 6239 1526 6267 1608
rect 6296 1593 6589 1661
rect 6618 1646 6646 1729
rect 6675 1714 6968 1782
rect 6997 1767 7025 1779
rect 6983 1764 7039 1767
rect 6983 1733 6988 1764
rect 7034 1733 7039 1764
rect 6983 1729 7039 1733
rect 6660 1661 6983 1714
rect 6604 1643 6660 1646
rect 6604 1612 6609 1643
rect 6655 1612 6660 1643
rect 6604 1608 6660 1612
rect 6281 1541 6604 1593
rect 6225 1523 6281 1526
rect 6225 1492 6230 1523
rect 6276 1492 6281 1523
rect 6225 1488 6281 1492
rect 5902 1421 6225 1473
rect 5846 1403 5902 1406
rect 5846 1372 5851 1403
rect 5897 1372 5902 1403
rect 5846 1368 5902 1372
rect 5481 1304 5482 1331
rect 5508 1304 5509 1331
rect 5088 1283 5144 1286
rect 5088 1252 5093 1283
rect 5139 1252 5144 1283
rect 5088 1248 5144 1252
rect 5102 1236 5130 1248
rect 5159 1234 5452 1301
rect 5481 1286 5509 1304
rect 5523 1301 5846 1353
rect 5860 1336 5888 1368
rect 5917 1353 6210 1421
rect 6239 1406 6267 1488
rect 6296 1473 6589 1541
rect 6618 1526 6646 1608
rect 6675 1593 6968 1661
rect 6997 1646 7025 1729
rect 7054 1714 7347 1782
rect 7376 1767 7404 1779
rect 7362 1764 7418 1767
rect 7362 1733 7367 1764
rect 7413 1733 7418 1764
rect 7362 1729 7418 1733
rect 7039 1661 7362 1714
rect 6983 1643 7039 1646
rect 6983 1612 6988 1643
rect 7034 1612 7039 1643
rect 6983 1608 7039 1612
rect 6660 1541 6983 1593
rect 6604 1523 6660 1526
rect 6604 1492 6609 1523
rect 6655 1492 6660 1523
rect 6604 1488 6660 1492
rect 6281 1421 6604 1473
rect 6225 1403 6281 1406
rect 6225 1372 6230 1403
rect 6276 1372 6281 1403
rect 6225 1368 6281 1372
rect 5860 1309 5861 1336
rect 5887 1309 5888 1336
rect 5467 1283 5523 1286
rect 5467 1252 5472 1283
rect 5518 1252 5523 1283
rect 5467 1248 5523 1252
rect 5481 1236 5509 1248
rect 5538 1234 5831 1301
rect 5860 1286 5888 1309
rect 5902 1301 6225 1353
rect 6239 1335 6267 1368
rect 6296 1353 6589 1421
rect 6618 1406 6646 1488
rect 6675 1473 6968 1541
rect 6997 1526 7025 1608
rect 7054 1593 7347 1661
rect 7376 1646 7404 1729
rect 7433 1714 7599 1782
rect 7418 1661 7599 1714
rect 7362 1643 7418 1646
rect 7362 1612 7367 1643
rect 7413 1612 7418 1643
rect 7362 1608 7418 1612
rect 7039 1541 7362 1593
rect 6983 1523 7039 1526
rect 6983 1492 6988 1523
rect 7034 1492 7039 1523
rect 6983 1488 7039 1492
rect 6660 1421 6983 1473
rect 6604 1403 6660 1406
rect 6604 1372 6609 1403
rect 6655 1372 6660 1403
rect 6604 1368 6660 1372
rect 6239 1308 6240 1335
rect 6266 1308 6267 1335
rect 5846 1283 5902 1286
rect 5846 1252 5851 1283
rect 5897 1252 5902 1283
rect 5846 1248 5902 1252
rect 5860 1236 5888 1248
rect 5917 1234 6210 1301
rect 6239 1286 6267 1308
rect 6281 1301 6604 1353
rect 6618 1333 6646 1368
rect 6675 1353 6968 1421
rect 6997 1406 7025 1488
rect 7054 1473 7347 1541
rect 7376 1526 7404 1608
rect 7433 1593 7599 1661
rect 7418 1541 7599 1593
rect 7362 1523 7418 1526
rect 7362 1492 7367 1523
rect 7413 1492 7418 1523
rect 7362 1488 7418 1492
rect 7039 1421 7362 1473
rect 6983 1403 7039 1406
rect 6983 1372 6988 1403
rect 7034 1372 7039 1403
rect 6983 1368 7039 1372
rect 6618 1306 6619 1333
rect 6645 1306 6646 1333
rect 6225 1283 6281 1286
rect 6225 1252 6230 1283
rect 6276 1252 6281 1283
rect 6225 1248 6281 1252
rect 6239 1236 6267 1248
rect 6296 1234 6589 1301
rect 6618 1286 6646 1306
rect 6660 1301 6983 1353
rect 6997 1331 7025 1368
rect 7054 1353 7347 1421
rect 7376 1406 7404 1488
rect 7433 1473 7599 1541
rect 7418 1421 7599 1473
rect 7362 1403 7418 1406
rect 7362 1372 7367 1403
rect 7413 1372 7418 1403
rect 7362 1368 7418 1372
rect 6997 1304 6998 1331
rect 7024 1304 7025 1331
rect 6604 1283 6660 1286
rect 6604 1252 6609 1283
rect 6655 1252 6660 1283
rect 6604 1248 6660 1252
rect 6618 1236 6646 1248
rect 6675 1234 6968 1301
rect 6997 1286 7025 1304
rect 7039 1301 7362 1353
rect 7376 1331 7404 1368
rect 7433 1353 7599 1421
rect 7376 1304 7377 1331
rect 7403 1304 7404 1331
rect 6983 1283 7039 1286
rect 6983 1252 6988 1283
rect 7034 1252 7039 1283
rect 6983 1248 7039 1252
rect 6997 1236 7025 1248
rect 7054 1234 7347 1301
rect 7376 1286 7404 1304
rect 7418 1301 7599 1353
rect 7362 1283 7418 1286
rect 7362 1252 7367 1283
rect 7413 1252 7418 1283
rect 7362 1248 7418 1252
rect 7376 1236 7404 1248
rect 7433 1234 7599 1301
rect -19 1222 161 1234
rect 217 1222 540 1234
rect 596 1222 919 1234
rect 975 1222 1298 1234
rect 1354 1222 1677 1234
rect 1733 1222 2056 1234
rect 2112 1222 2435 1234
rect 2491 1222 2814 1234
rect 2870 1222 3193 1234
rect 3249 1222 3572 1234
rect 3628 1222 3951 1234
rect 4007 1222 4330 1234
rect 4386 1222 4709 1234
rect 4765 1222 5088 1234
rect 5144 1222 5467 1234
rect 5523 1222 5846 1234
rect 5902 1222 6225 1234
rect 6281 1222 6604 1234
rect 6660 1222 6983 1234
rect 7039 1222 7362 1234
rect 7418 1222 7599 1234
rect -19 1219 7599 1222
rect -19 1193 34 1219
rect 61 1193 109 1219
rect 136 1193 242 1219
rect 269 1193 317 1219
rect 344 1193 413 1219
rect 440 1193 488 1219
rect 515 1193 621 1219
rect 648 1193 696 1219
rect 723 1193 792 1219
rect 819 1193 867 1219
rect 894 1193 1000 1219
rect 1027 1193 1075 1219
rect 1102 1193 1171 1219
rect 1198 1193 1246 1219
rect 1273 1193 1379 1219
rect 1406 1193 1454 1219
rect 1481 1193 1550 1219
rect 1577 1193 1625 1219
rect 1652 1193 1758 1219
rect 1785 1193 1833 1219
rect 1860 1193 1929 1219
rect 1956 1193 2004 1219
rect 2031 1193 2137 1219
rect 2164 1193 2212 1219
rect 2239 1193 2308 1219
rect 2335 1193 2383 1219
rect 2410 1193 2516 1219
rect 2543 1193 2591 1219
rect 2618 1193 2687 1219
rect 2714 1193 2762 1219
rect 2789 1193 2895 1219
rect 2922 1193 2970 1219
rect 2997 1193 3066 1219
rect 3093 1193 3141 1219
rect 3168 1193 3274 1219
rect 3301 1193 3349 1219
rect 3376 1193 3445 1219
rect 3472 1193 3520 1219
rect 3547 1193 3653 1219
rect 3680 1193 3728 1219
rect 3755 1193 3824 1219
rect 3851 1193 3899 1219
rect 3926 1193 4032 1219
rect 4059 1193 4107 1219
rect 4134 1193 4203 1219
rect 4230 1193 4278 1219
rect 4305 1193 4411 1219
rect 4438 1193 4486 1219
rect 4513 1193 4582 1219
rect 4609 1193 4657 1219
rect 4684 1193 4790 1219
rect 4817 1193 4865 1219
rect 4892 1193 4961 1219
rect 4988 1193 5036 1219
rect 5063 1193 5169 1219
rect 5196 1193 5244 1219
rect 5271 1193 5340 1219
rect 5367 1193 5415 1219
rect 5442 1193 5548 1219
rect 5575 1193 5623 1219
rect 5650 1193 5719 1219
rect 5746 1193 5794 1219
rect 5821 1193 5927 1219
rect 5954 1193 6002 1219
rect 6029 1193 6098 1219
rect 6125 1193 6173 1219
rect 6200 1193 6306 1219
rect 6333 1193 6381 1219
rect 6408 1193 6477 1219
rect 6504 1193 6552 1219
rect 6579 1193 6685 1219
rect 6712 1193 6760 1219
rect 6787 1193 6856 1219
rect 6883 1193 6931 1219
rect 6958 1193 7064 1219
rect 7091 1193 7139 1219
rect 7166 1193 7235 1219
rect 7262 1193 7310 1219
rect 7337 1193 7443 1219
rect 7470 1193 7518 1219
rect 7545 1193 7599 1219
rect -19 1190 7599 1193
rect -19 1179 161 1190
rect 217 1179 540 1190
rect 596 1179 919 1190
rect 975 1179 1298 1190
rect 1354 1179 1677 1190
rect 1733 1179 2056 1190
rect 2112 1179 2435 1190
rect 2491 1179 2814 1190
rect 2870 1179 3193 1190
rect 3249 1179 3572 1190
rect 3628 1179 3951 1190
rect 4007 1179 4330 1190
rect 4386 1179 4709 1190
rect 4765 1179 5088 1190
rect 5144 1179 5467 1190
rect 5523 1179 5846 1190
rect 5902 1179 6225 1190
rect 6281 1179 6604 1190
rect 6660 1179 6983 1190
rect 7039 1179 7362 1190
rect 7418 1179 7599 1190
rect -19 1111 146 1179
rect 175 1164 203 1176
rect 161 1161 217 1164
rect 161 1130 166 1161
rect 212 1130 217 1161
rect 161 1126 217 1130
rect -19 1058 161 1111
rect -19 990 146 1058
rect 175 1043 203 1126
rect 232 1111 525 1179
rect 554 1164 582 1176
rect 540 1161 596 1164
rect 540 1130 545 1161
rect 591 1130 596 1161
rect 540 1126 596 1130
rect 217 1058 540 1111
rect 161 1040 217 1043
rect 161 1009 166 1040
rect 212 1009 217 1040
rect 161 1005 217 1009
rect -19 938 161 990
rect -19 870 146 938
rect 175 923 203 1005
rect 232 990 525 1058
rect 554 1043 582 1126
rect 611 1111 904 1179
rect 933 1164 961 1176
rect 919 1161 975 1164
rect 919 1130 924 1161
rect 970 1130 975 1161
rect 919 1126 975 1130
rect 596 1058 919 1111
rect 540 1040 596 1043
rect 540 1009 545 1040
rect 591 1009 596 1040
rect 540 1005 596 1009
rect 217 938 540 990
rect 161 920 217 923
rect 161 889 166 920
rect 212 889 217 920
rect 161 885 217 889
rect -19 818 161 870
rect -19 750 146 818
rect 175 803 203 885
rect 232 870 525 938
rect 554 923 582 1005
rect 611 990 904 1058
rect 933 1043 961 1126
rect 990 1111 1283 1179
rect 1312 1164 1340 1176
rect 1298 1161 1354 1164
rect 1298 1130 1303 1161
rect 1349 1130 1354 1161
rect 1298 1126 1354 1130
rect 975 1058 1298 1111
rect 919 1040 975 1043
rect 919 1009 924 1040
rect 970 1009 975 1040
rect 919 1005 975 1009
rect 596 938 919 990
rect 540 920 596 923
rect 540 889 545 920
rect 591 889 596 920
rect 540 885 596 889
rect 217 818 540 870
rect 161 800 217 803
rect 161 769 166 800
rect 212 769 217 800
rect 161 765 217 769
rect -19 698 161 750
rect 175 717 203 765
rect 232 750 525 818
rect 554 803 582 885
rect 611 870 904 938
rect 933 923 961 1005
rect 990 990 1283 1058
rect 1312 1043 1340 1126
rect 1369 1111 1662 1179
rect 1691 1164 1719 1176
rect 1677 1161 1733 1164
rect 1677 1130 1682 1161
rect 1728 1130 1733 1161
rect 1677 1126 1733 1130
rect 1354 1058 1677 1111
rect 1298 1040 1354 1043
rect 1298 1009 1303 1040
rect 1349 1009 1354 1040
rect 1298 1005 1354 1009
rect 975 938 1298 990
rect 919 920 975 923
rect 919 889 924 920
rect 970 889 975 920
rect 919 885 975 889
rect 596 818 919 870
rect 540 800 596 803
rect 540 769 545 800
rect 591 769 596 800
rect 540 765 596 769
rect -19 631 146 698
rect 175 690 176 717
rect 202 690 203 717
rect 217 698 540 750
rect 554 723 582 765
rect 611 750 904 818
rect 933 803 961 885
rect 990 870 1283 938
rect 1312 923 1340 1005
rect 1369 990 1662 1058
rect 1691 1043 1719 1126
rect 1748 1111 2041 1179
rect 2070 1164 2098 1176
rect 2056 1161 2112 1164
rect 2056 1130 2061 1161
rect 2107 1130 2112 1161
rect 2056 1126 2112 1130
rect 1733 1058 2056 1111
rect 1677 1040 1733 1043
rect 1677 1009 1682 1040
rect 1728 1009 1733 1040
rect 1677 1005 1733 1009
rect 1354 938 1677 990
rect 1298 920 1354 923
rect 1298 889 1303 920
rect 1349 889 1354 920
rect 1298 885 1354 889
rect 975 818 1298 870
rect 919 800 975 803
rect 919 769 924 800
rect 970 769 975 800
rect 919 765 975 769
rect 175 683 203 690
rect 161 680 217 683
rect 161 649 166 680
rect 212 649 217 680
rect 161 645 217 649
rect 175 633 203 645
rect 232 631 525 698
rect 554 696 555 723
rect 581 696 582 723
rect 596 698 919 750
rect 933 723 961 765
rect 990 750 1283 818
rect 1312 803 1340 885
rect 1369 870 1662 938
rect 1691 923 1719 1005
rect 1748 990 2041 1058
rect 2070 1043 2098 1126
rect 2127 1111 2420 1179
rect 2449 1164 2477 1176
rect 2435 1161 2491 1164
rect 2435 1130 2440 1161
rect 2486 1130 2491 1161
rect 2435 1126 2491 1130
rect 2112 1058 2435 1111
rect 2056 1040 2112 1043
rect 2056 1009 2061 1040
rect 2107 1009 2112 1040
rect 2056 1005 2112 1009
rect 1733 938 2056 990
rect 1677 920 1733 923
rect 1677 889 1682 920
rect 1728 889 1733 920
rect 1677 885 1733 889
rect 1354 818 1677 870
rect 1298 800 1354 803
rect 1298 769 1303 800
rect 1349 769 1354 800
rect 1298 765 1354 769
rect 554 683 582 696
rect 540 680 596 683
rect 540 649 545 680
rect 591 649 596 680
rect 540 645 596 649
rect 554 633 582 645
rect 611 631 904 698
rect 933 696 934 723
rect 960 696 961 723
rect 975 698 1298 750
rect 1312 723 1340 765
rect 1369 750 1662 818
rect 1691 803 1719 885
rect 1748 870 2041 938
rect 2070 923 2098 1005
rect 2127 990 2420 1058
rect 2449 1043 2477 1126
rect 2506 1111 2799 1179
rect 2828 1164 2856 1176
rect 2814 1161 2870 1164
rect 2814 1130 2819 1161
rect 2865 1130 2870 1161
rect 2814 1126 2870 1130
rect 2491 1058 2814 1111
rect 2435 1040 2491 1043
rect 2435 1009 2440 1040
rect 2486 1009 2491 1040
rect 2435 1005 2491 1009
rect 2112 938 2435 990
rect 2056 920 2112 923
rect 2056 889 2061 920
rect 2107 889 2112 920
rect 2056 885 2112 889
rect 1733 818 2056 870
rect 1677 800 1733 803
rect 1677 769 1682 800
rect 1728 769 1733 800
rect 1677 765 1733 769
rect 933 683 961 696
rect 919 680 975 683
rect 919 649 924 680
rect 970 649 975 680
rect 919 645 975 649
rect 933 633 961 645
rect 990 631 1283 698
rect 1312 696 1313 723
rect 1339 696 1340 723
rect 1354 698 1677 750
rect 1691 724 1719 765
rect 1748 750 2041 818
rect 2070 803 2098 885
rect 2127 870 2420 938
rect 2449 923 2477 1005
rect 2506 990 2799 1058
rect 2828 1043 2856 1126
rect 2885 1111 3178 1179
rect 3207 1164 3235 1176
rect 3193 1161 3249 1164
rect 3193 1130 3198 1161
rect 3244 1130 3249 1161
rect 3193 1126 3249 1130
rect 2870 1058 3193 1111
rect 2814 1040 2870 1043
rect 2814 1009 2819 1040
rect 2865 1009 2870 1040
rect 2814 1005 2870 1009
rect 2491 938 2814 990
rect 2435 920 2491 923
rect 2435 889 2440 920
rect 2486 889 2491 920
rect 2435 885 2491 889
rect 2112 818 2435 870
rect 2056 800 2112 803
rect 2056 769 2061 800
rect 2107 769 2112 800
rect 2056 765 2112 769
rect 1312 683 1340 696
rect 1298 680 1354 683
rect 1298 649 1303 680
rect 1349 649 1354 680
rect 1298 645 1354 649
rect 1312 633 1340 645
rect 1369 631 1662 698
rect 1691 697 1692 724
rect 1718 697 1719 724
rect 1733 698 2056 750
rect 2070 717 2098 765
rect 2127 750 2420 818
rect 2449 803 2477 885
rect 2506 870 2799 938
rect 2828 923 2856 1005
rect 2885 990 3178 1058
rect 3207 1043 3235 1126
rect 3264 1111 3557 1179
rect 3586 1164 3614 1176
rect 3572 1161 3628 1164
rect 3572 1130 3577 1161
rect 3623 1130 3628 1161
rect 3572 1126 3628 1130
rect 3249 1058 3572 1111
rect 3193 1040 3249 1043
rect 3193 1009 3198 1040
rect 3244 1009 3249 1040
rect 3193 1005 3249 1009
rect 2870 938 3193 990
rect 2814 920 2870 923
rect 2814 889 2819 920
rect 2865 889 2870 920
rect 2814 885 2870 889
rect 2491 818 2814 870
rect 2435 800 2491 803
rect 2435 769 2440 800
rect 2486 769 2491 800
rect 2435 765 2491 769
rect 1691 683 1719 697
rect 1677 680 1733 683
rect 1677 649 1682 680
rect 1728 649 1733 680
rect 1677 645 1733 649
rect 1691 633 1719 645
rect 1748 631 2041 698
rect 2070 690 2071 717
rect 2097 690 2098 717
rect 2112 698 2435 750
rect 2449 723 2477 765
rect 2506 750 2799 818
rect 2828 803 2856 885
rect 2885 870 3178 938
rect 3207 923 3235 1005
rect 3264 990 3557 1058
rect 3586 1043 3614 1126
rect 3643 1111 3936 1179
rect 3965 1164 3993 1176
rect 3951 1161 4007 1164
rect 3951 1130 3956 1161
rect 4002 1130 4007 1161
rect 3951 1126 4007 1130
rect 3628 1058 3951 1111
rect 3572 1040 3628 1043
rect 3572 1009 3577 1040
rect 3623 1009 3628 1040
rect 3572 1005 3628 1009
rect 3249 938 3572 990
rect 3193 920 3249 923
rect 3193 889 3198 920
rect 3244 889 3249 920
rect 3193 885 3249 889
rect 2870 818 3193 870
rect 2814 800 2870 803
rect 2814 769 2819 800
rect 2865 769 2870 800
rect 2814 765 2870 769
rect 2070 683 2098 690
rect 2056 680 2112 683
rect 2056 649 2061 680
rect 2107 649 2112 680
rect 2056 645 2112 649
rect 2070 633 2098 645
rect 2127 631 2420 698
rect 2449 696 2450 723
rect 2476 696 2477 723
rect 2491 698 2814 750
rect 2828 723 2856 765
rect 2885 750 3178 818
rect 3207 803 3235 885
rect 3264 870 3557 938
rect 3586 923 3614 1005
rect 3643 990 3936 1058
rect 3965 1043 3993 1126
rect 4022 1111 4315 1179
rect 4344 1164 4372 1176
rect 4330 1161 4386 1164
rect 4330 1130 4335 1161
rect 4381 1130 4386 1161
rect 4330 1126 4386 1130
rect 4007 1058 4330 1111
rect 3951 1040 4007 1043
rect 3951 1009 3956 1040
rect 4002 1009 4007 1040
rect 3951 1005 4007 1009
rect 3628 938 3951 990
rect 3572 920 3628 923
rect 3572 889 3577 920
rect 3623 889 3628 920
rect 3572 885 3628 889
rect 3249 818 3572 870
rect 3193 800 3249 803
rect 3193 769 3198 800
rect 3244 769 3249 800
rect 3193 765 3249 769
rect 2449 683 2477 696
rect 2435 680 2491 683
rect 2435 649 2440 680
rect 2486 649 2491 680
rect 2435 645 2491 649
rect 2449 633 2477 645
rect 2506 631 2799 698
rect 2828 696 2829 723
rect 2855 696 2856 723
rect 2870 698 3193 750
rect 3207 723 3235 765
rect 3264 750 3557 818
rect 3586 803 3614 885
rect 3643 870 3936 938
rect 3965 923 3993 1005
rect 4022 990 4315 1058
rect 4344 1043 4372 1126
rect 4401 1111 4694 1179
rect 4723 1164 4751 1176
rect 4709 1161 4765 1164
rect 4709 1130 4714 1161
rect 4760 1130 4765 1161
rect 4709 1126 4765 1130
rect 4386 1058 4709 1111
rect 4330 1040 4386 1043
rect 4330 1009 4335 1040
rect 4381 1009 4386 1040
rect 4330 1005 4386 1009
rect 4007 938 4330 990
rect 3951 920 4007 923
rect 3951 889 3956 920
rect 4002 889 4007 920
rect 3951 885 4007 889
rect 3628 818 3951 870
rect 3572 800 3628 803
rect 3572 769 3577 800
rect 3623 769 3628 800
rect 3572 765 3628 769
rect 2828 683 2856 696
rect 2814 680 2870 683
rect 2814 649 2819 680
rect 2865 649 2870 680
rect 2814 645 2870 649
rect 2828 633 2856 645
rect 2885 631 3178 698
rect 3207 696 3208 723
rect 3234 696 3235 723
rect 3249 698 3572 750
rect 3586 724 3614 765
rect 3643 750 3936 818
rect 3965 803 3993 885
rect 4022 870 4315 938
rect 4344 923 4372 1005
rect 4401 990 4694 1058
rect 4723 1043 4751 1126
rect 4780 1111 5073 1179
rect 5102 1164 5130 1176
rect 5088 1161 5144 1164
rect 5088 1130 5093 1161
rect 5139 1130 5144 1161
rect 5088 1126 5144 1130
rect 4765 1058 5088 1111
rect 4709 1040 4765 1043
rect 4709 1009 4714 1040
rect 4760 1009 4765 1040
rect 4709 1005 4765 1009
rect 4386 938 4709 990
rect 4330 920 4386 923
rect 4330 889 4335 920
rect 4381 889 4386 920
rect 4330 885 4386 889
rect 4007 818 4330 870
rect 3951 800 4007 803
rect 3951 769 3956 800
rect 4002 769 4007 800
rect 3951 765 4007 769
rect 3207 683 3235 696
rect 3193 680 3249 683
rect 3193 649 3198 680
rect 3244 649 3249 680
rect 3193 645 3249 649
rect 3207 633 3235 645
rect 3264 631 3557 698
rect 3586 697 3587 724
rect 3613 697 3614 724
rect 3628 698 3951 750
rect 3965 717 3993 765
rect 4022 750 4315 818
rect 4344 803 4372 885
rect 4401 870 4694 938
rect 4723 923 4751 1005
rect 4780 990 5073 1058
rect 5102 1043 5130 1126
rect 5159 1111 5452 1179
rect 5481 1164 5509 1176
rect 5467 1161 5523 1164
rect 5467 1130 5472 1161
rect 5518 1130 5523 1161
rect 5467 1126 5523 1130
rect 5144 1058 5467 1111
rect 5088 1040 5144 1043
rect 5088 1009 5093 1040
rect 5139 1009 5144 1040
rect 5088 1005 5144 1009
rect 4765 938 5088 990
rect 4709 920 4765 923
rect 4709 889 4714 920
rect 4760 889 4765 920
rect 4709 885 4765 889
rect 4386 818 4709 870
rect 4330 800 4386 803
rect 4330 769 4335 800
rect 4381 769 4386 800
rect 4330 765 4386 769
rect 3586 683 3614 697
rect 3572 680 3628 683
rect 3572 649 3577 680
rect 3623 649 3628 680
rect 3572 645 3628 649
rect 3586 633 3614 645
rect 3643 631 3936 698
rect 3965 690 3966 717
rect 3992 690 3993 717
rect 4007 698 4330 750
rect 4344 723 4372 765
rect 4401 750 4694 818
rect 4723 803 4751 885
rect 4780 870 5073 938
rect 5102 923 5130 1005
rect 5159 990 5452 1058
rect 5481 1043 5509 1126
rect 5538 1111 5831 1179
rect 5860 1164 5888 1176
rect 5846 1161 5902 1164
rect 5846 1130 5851 1161
rect 5897 1130 5902 1161
rect 5846 1126 5902 1130
rect 5523 1058 5846 1111
rect 5467 1040 5523 1043
rect 5467 1009 5472 1040
rect 5518 1009 5523 1040
rect 5467 1005 5523 1009
rect 5144 938 5467 990
rect 5088 920 5144 923
rect 5088 889 5093 920
rect 5139 889 5144 920
rect 5088 885 5144 889
rect 4765 818 5088 870
rect 4709 800 4765 803
rect 4709 769 4714 800
rect 4760 769 4765 800
rect 4709 765 4765 769
rect 3965 683 3993 690
rect 3951 680 4007 683
rect 3951 649 3956 680
rect 4002 649 4007 680
rect 3951 645 4007 649
rect 3965 633 3993 645
rect 4022 631 4315 698
rect 4344 696 4345 723
rect 4371 696 4372 723
rect 4386 698 4709 750
rect 4723 723 4751 765
rect 4780 750 5073 818
rect 5102 803 5130 885
rect 5159 870 5452 938
rect 5481 923 5509 1005
rect 5538 990 5831 1058
rect 5860 1043 5888 1126
rect 5917 1111 6210 1179
rect 6239 1164 6267 1176
rect 6225 1161 6281 1164
rect 6225 1130 6230 1161
rect 6276 1130 6281 1161
rect 6225 1126 6281 1130
rect 5902 1058 6225 1111
rect 5846 1040 5902 1043
rect 5846 1009 5851 1040
rect 5897 1009 5902 1040
rect 5846 1005 5902 1009
rect 5523 938 5846 990
rect 5467 920 5523 923
rect 5467 889 5472 920
rect 5518 889 5523 920
rect 5467 885 5523 889
rect 5144 818 5467 870
rect 5088 800 5144 803
rect 5088 769 5093 800
rect 5139 769 5144 800
rect 5088 765 5144 769
rect 4344 683 4372 696
rect 4330 680 4386 683
rect 4330 649 4335 680
rect 4381 649 4386 680
rect 4330 645 4386 649
rect 4344 633 4372 645
rect 4401 631 4694 698
rect 4723 696 4724 723
rect 4750 696 4751 723
rect 4765 698 5088 750
rect 5102 723 5130 765
rect 5159 750 5452 818
rect 5481 803 5509 885
rect 5538 870 5831 938
rect 5860 923 5888 1005
rect 5917 990 6210 1058
rect 6239 1043 6267 1126
rect 6296 1111 6589 1179
rect 6618 1164 6646 1176
rect 6604 1161 6660 1164
rect 6604 1130 6609 1161
rect 6655 1130 6660 1161
rect 6604 1126 6660 1130
rect 6281 1058 6604 1111
rect 6225 1040 6281 1043
rect 6225 1009 6230 1040
rect 6276 1009 6281 1040
rect 6225 1005 6281 1009
rect 5902 938 6225 990
rect 5846 920 5902 923
rect 5846 889 5851 920
rect 5897 889 5902 920
rect 5846 885 5902 889
rect 5523 818 5846 870
rect 5467 800 5523 803
rect 5467 769 5472 800
rect 5518 769 5523 800
rect 5467 765 5523 769
rect 4723 683 4751 696
rect 4709 680 4765 683
rect 4709 649 4714 680
rect 4760 649 4765 680
rect 4709 645 4765 649
rect 4723 633 4751 645
rect 4780 631 5073 698
rect 5102 696 5103 723
rect 5129 696 5130 723
rect 5144 698 5467 750
rect 5481 724 5509 765
rect 5538 750 5831 818
rect 5860 803 5888 885
rect 5917 870 6210 938
rect 6239 923 6267 1005
rect 6296 990 6589 1058
rect 6618 1043 6646 1126
rect 6675 1111 6968 1179
rect 6997 1164 7025 1176
rect 6983 1161 7039 1164
rect 6983 1130 6988 1161
rect 7034 1130 7039 1161
rect 6983 1126 7039 1130
rect 6660 1058 6983 1111
rect 6604 1040 6660 1043
rect 6604 1009 6609 1040
rect 6655 1009 6660 1040
rect 6604 1005 6660 1009
rect 6281 938 6604 990
rect 6225 920 6281 923
rect 6225 889 6230 920
rect 6276 889 6281 920
rect 6225 885 6281 889
rect 5902 818 6225 870
rect 5846 800 5902 803
rect 5846 769 5851 800
rect 5897 769 5902 800
rect 5846 765 5902 769
rect 5102 683 5130 696
rect 5088 680 5144 683
rect 5088 649 5093 680
rect 5139 649 5144 680
rect 5088 645 5144 649
rect 5102 633 5130 645
rect 5159 631 5452 698
rect 5481 697 5482 724
rect 5508 697 5509 724
rect 5523 698 5846 750
rect 5860 717 5888 765
rect 5917 750 6210 818
rect 6239 803 6267 885
rect 6296 870 6589 938
rect 6618 923 6646 1005
rect 6675 990 6968 1058
rect 6997 1043 7025 1126
rect 7054 1111 7347 1179
rect 7376 1164 7404 1176
rect 7362 1161 7418 1164
rect 7362 1130 7367 1161
rect 7413 1130 7418 1161
rect 7362 1126 7418 1130
rect 7039 1058 7362 1111
rect 6983 1040 7039 1043
rect 6983 1009 6988 1040
rect 7034 1009 7039 1040
rect 6983 1005 7039 1009
rect 6660 938 6983 990
rect 6604 920 6660 923
rect 6604 889 6609 920
rect 6655 889 6660 920
rect 6604 885 6660 889
rect 6281 818 6604 870
rect 6225 800 6281 803
rect 6225 769 6230 800
rect 6276 769 6281 800
rect 6225 765 6281 769
rect 5481 683 5509 697
rect 5467 680 5523 683
rect 5467 649 5472 680
rect 5518 649 5523 680
rect 5467 645 5523 649
rect 5481 633 5509 645
rect 5538 631 5831 698
rect 5860 690 5861 717
rect 5887 690 5888 717
rect 5902 698 6225 750
rect 6239 723 6267 765
rect 6296 750 6589 818
rect 6618 803 6646 885
rect 6675 870 6968 938
rect 6997 923 7025 1005
rect 7054 990 7347 1058
rect 7376 1043 7404 1126
rect 7433 1111 7599 1179
rect 7418 1058 7599 1111
rect 7362 1040 7418 1043
rect 7362 1009 7367 1040
rect 7413 1009 7418 1040
rect 7362 1005 7418 1009
rect 7039 938 7362 990
rect 6983 920 7039 923
rect 6983 889 6988 920
rect 7034 889 7039 920
rect 6983 885 7039 889
rect 6660 818 6983 870
rect 6604 800 6660 803
rect 6604 769 6609 800
rect 6655 769 6660 800
rect 6604 765 6660 769
rect 5860 683 5888 690
rect 5846 680 5902 683
rect 5846 649 5851 680
rect 5897 649 5902 680
rect 5846 645 5902 649
rect 5860 633 5888 645
rect 5917 631 6210 698
rect 6239 696 6240 723
rect 6266 696 6267 723
rect 6281 698 6604 750
rect 6618 723 6646 765
rect 6675 750 6968 818
rect 6997 803 7025 885
rect 7054 870 7347 938
rect 7376 923 7404 1005
rect 7433 990 7599 1058
rect 7418 938 7599 990
rect 7362 920 7418 923
rect 7362 889 7367 920
rect 7413 889 7418 920
rect 7362 885 7418 889
rect 7039 818 7362 870
rect 6983 800 7039 803
rect 6983 769 6988 800
rect 7034 769 7039 800
rect 6983 765 7039 769
rect 6239 683 6267 696
rect 6225 680 6281 683
rect 6225 649 6230 680
rect 6276 649 6281 680
rect 6225 645 6281 649
rect 6239 633 6267 645
rect 6296 631 6589 698
rect 6618 696 6619 723
rect 6645 696 6646 723
rect 6660 698 6983 750
rect 6997 723 7025 765
rect 7054 750 7347 818
rect 7376 803 7404 885
rect 7433 870 7599 938
rect 7418 818 7599 870
rect 7362 800 7418 803
rect 7362 769 7367 800
rect 7413 769 7418 800
rect 7362 765 7418 769
rect 6618 683 6646 696
rect 6604 680 6660 683
rect 6604 649 6609 680
rect 6655 649 6660 680
rect 6604 645 6660 649
rect 6618 633 6646 645
rect 6675 631 6968 698
rect 6997 696 6998 723
rect 7024 696 7025 723
rect 7039 698 7362 750
rect 7376 724 7404 765
rect 7433 750 7599 818
rect 6997 683 7025 696
rect 6983 680 7039 683
rect 6983 649 6988 680
rect 7034 649 7039 680
rect 6983 645 7039 649
rect 6997 633 7025 645
rect 7054 631 7347 698
rect 7376 697 7377 724
rect 7403 697 7404 724
rect 7418 698 7599 750
rect 7376 683 7404 697
rect 7362 680 7418 683
rect 7362 649 7367 680
rect 7413 649 7418 680
rect 7362 645 7418 649
rect 7376 633 7404 645
rect 7433 631 7599 698
rect -19 619 161 631
rect 217 619 540 631
rect 596 619 919 631
rect 975 619 1298 631
rect 1354 619 1677 631
rect 1733 619 2056 631
rect 2112 619 2435 631
rect 2491 619 2814 631
rect 2870 619 3193 631
rect 3249 619 3572 631
rect 3628 619 3951 631
rect 4007 619 4330 631
rect 4386 619 4709 631
rect 4765 619 5088 631
rect 5144 619 5467 631
rect 5523 619 5846 631
rect 5902 619 6225 631
rect 6281 619 6604 631
rect 6660 619 6983 631
rect 7039 619 7362 631
rect 7418 619 7599 631
rect -19 616 7599 619
rect -19 590 34 616
rect 61 590 109 616
rect 136 590 242 616
rect 269 590 317 616
rect 344 590 413 616
rect 440 590 488 616
rect 515 590 621 616
rect 648 590 696 616
rect 723 590 792 616
rect 819 590 867 616
rect 894 590 1000 616
rect 1027 590 1075 616
rect 1102 590 1171 616
rect 1198 590 1246 616
rect 1273 590 1379 616
rect 1406 590 1454 616
rect 1481 590 1550 616
rect 1577 590 1625 616
rect 1652 590 1758 616
rect 1785 590 1833 616
rect 1860 590 1929 616
rect 1956 590 2004 616
rect 2031 590 2137 616
rect 2164 590 2212 616
rect 2239 590 2308 616
rect 2335 590 2383 616
rect 2410 590 2516 616
rect 2543 590 2591 616
rect 2618 590 2687 616
rect 2714 590 2762 616
rect 2789 590 2895 616
rect 2922 590 2970 616
rect 2997 590 3066 616
rect 3093 590 3141 616
rect 3168 590 3274 616
rect 3301 590 3349 616
rect 3376 590 3445 616
rect 3472 590 3520 616
rect 3547 590 3653 616
rect 3680 590 3728 616
rect 3755 590 3824 616
rect 3851 590 3899 616
rect 3926 590 4032 616
rect 4059 590 4107 616
rect 4134 590 4203 616
rect 4230 590 4278 616
rect 4305 590 4411 616
rect 4438 590 4486 616
rect 4513 590 4582 616
rect 4609 590 4657 616
rect 4684 590 4790 616
rect 4817 590 4865 616
rect 4892 590 4961 616
rect 4988 590 5036 616
rect 5063 590 5169 616
rect 5196 590 5244 616
rect 5271 590 5340 616
rect 5367 590 5415 616
rect 5442 590 5548 616
rect 5575 590 5623 616
rect 5650 590 5719 616
rect 5746 590 5794 616
rect 5821 590 5927 616
rect 5954 590 6002 616
rect 6029 590 6098 616
rect 6125 590 6173 616
rect 6200 590 6306 616
rect 6333 590 6381 616
rect 6408 590 6477 616
rect 6504 590 6552 616
rect 6579 590 6685 616
rect 6712 590 6760 616
rect 6787 590 6856 616
rect 6883 590 6931 616
rect 6958 590 7064 616
rect 7091 590 7139 616
rect 7166 590 7235 616
rect 7262 590 7310 616
rect 7337 590 7443 616
rect 7470 590 7518 616
rect 7545 590 7599 616
rect -19 587 7599 590
rect -19 576 161 587
rect 217 576 540 587
rect 596 576 919 587
rect 975 576 1298 587
rect 1354 576 1677 587
rect 1733 576 2056 587
rect 2112 576 2435 587
rect 2491 576 2814 587
rect 2870 576 3193 587
rect 3249 576 3572 587
rect 3628 576 3951 587
rect 4007 576 4330 587
rect 4386 576 4709 587
rect 4765 576 5088 587
rect 5144 576 5467 587
rect 5523 576 5846 587
rect 5902 576 6225 587
rect 6281 576 6604 587
rect 6660 576 6983 587
rect 7039 576 7362 587
rect 7418 576 7599 587
rect -19 508 146 576
rect 175 561 203 573
rect 161 558 217 561
rect 161 527 166 558
rect 212 527 217 558
rect 161 523 217 527
rect 175 511 203 523
rect -19 455 161 508
rect 175 484 176 511
rect 202 484 203 511
rect 232 508 525 576
rect 554 561 582 573
rect 540 558 596 561
rect 540 527 545 558
rect 591 527 596 558
rect 540 523 596 527
rect 554 511 582 523
rect -19 387 146 455
rect 175 440 203 484
rect 217 455 540 508
rect 554 484 555 511
rect 581 484 582 511
rect 611 508 904 576
rect 933 561 961 573
rect 919 558 975 561
rect 919 527 924 558
rect 970 527 975 558
rect 919 523 975 527
rect 933 511 961 523
rect 161 437 217 440
rect 161 406 166 437
rect 212 406 217 437
rect 161 402 217 406
rect -19 335 161 387
rect -19 267 146 335
rect 175 320 203 402
rect 232 387 525 455
rect 554 440 582 484
rect 596 455 919 508
rect 933 484 934 511
rect 960 484 961 511
rect 990 508 1283 576
rect 1312 561 1340 573
rect 1298 558 1354 561
rect 1298 527 1303 558
rect 1349 527 1354 558
rect 1298 523 1354 527
rect 1312 511 1340 523
rect 540 437 596 440
rect 540 406 545 437
rect 591 406 596 437
rect 540 402 596 406
rect 217 335 540 387
rect 161 317 217 320
rect 161 286 166 317
rect 212 286 217 317
rect 161 282 217 286
rect -19 215 161 267
rect -19 147 146 215
rect 175 200 203 282
rect 232 267 525 335
rect 554 320 582 402
rect 611 387 904 455
rect 933 440 961 484
rect 975 455 1298 508
rect 1312 484 1313 511
rect 1339 484 1340 511
rect 1369 508 1662 576
rect 1691 561 1719 573
rect 1677 558 1733 561
rect 1677 527 1682 558
rect 1728 527 1733 558
rect 1677 523 1733 527
rect 1691 510 1719 523
rect 919 437 975 440
rect 919 406 924 437
rect 970 406 975 437
rect 919 402 975 406
rect 596 335 919 387
rect 540 317 596 320
rect 540 286 545 317
rect 591 286 596 317
rect 540 282 596 286
rect 217 215 540 267
rect 161 197 217 200
rect 161 166 166 197
rect 212 166 217 197
rect 161 162 217 166
rect -19 95 161 147
rect -19 28 146 95
rect 175 80 203 162
rect 232 147 525 215
rect 554 200 582 282
rect 611 267 904 335
rect 933 320 961 402
rect 990 387 1283 455
rect 1312 440 1340 484
rect 1354 455 1677 508
rect 1691 483 1692 510
rect 1718 483 1719 510
rect 1748 508 2041 576
rect 2070 561 2098 573
rect 2056 558 2112 561
rect 2056 527 2061 558
rect 2107 527 2112 558
rect 2056 523 2112 527
rect 2070 511 2098 523
rect 1298 437 1354 440
rect 1298 406 1303 437
rect 1349 406 1354 437
rect 1298 402 1354 406
rect 975 335 1298 387
rect 919 317 975 320
rect 919 286 924 317
rect 970 286 975 317
rect 919 282 975 286
rect 596 215 919 267
rect 540 197 596 200
rect 540 166 545 197
rect 591 166 596 197
rect 540 162 596 166
rect 217 95 540 147
rect 161 77 217 80
rect 161 46 166 77
rect 212 46 217 77
rect 161 42 217 46
rect 175 30 203 42
rect 232 28 525 95
rect 554 80 582 162
rect 611 147 904 215
rect 933 200 961 282
rect 990 267 1283 335
rect 1312 320 1340 402
rect 1369 387 1662 455
rect 1691 440 1719 483
rect 1733 455 2056 508
rect 2070 484 2071 511
rect 2097 484 2098 511
rect 2127 508 2420 576
rect 2449 561 2477 573
rect 2435 558 2491 561
rect 2435 527 2440 558
rect 2486 527 2491 558
rect 2435 523 2491 527
rect 2449 513 2477 523
rect 1677 437 1733 440
rect 1677 406 1682 437
rect 1728 406 1733 437
rect 1677 402 1733 406
rect 1354 335 1677 387
rect 1298 317 1354 320
rect 1298 286 1303 317
rect 1349 286 1354 317
rect 1298 282 1354 286
rect 975 215 1298 267
rect 919 197 975 200
rect 919 166 924 197
rect 970 166 975 197
rect 919 162 975 166
rect 596 95 919 147
rect 540 77 596 80
rect 540 46 545 77
rect 591 46 596 77
rect 540 42 596 46
rect 554 30 582 42
rect 611 28 904 95
rect 933 80 961 162
rect 990 147 1283 215
rect 1312 200 1340 282
rect 1369 267 1662 335
rect 1691 320 1719 402
rect 1748 387 2041 455
rect 2070 440 2098 484
rect 2112 455 2435 508
rect 2449 486 2450 513
rect 2476 486 2477 513
rect 2506 508 2799 576
rect 2828 561 2856 573
rect 2814 558 2870 561
rect 2814 527 2819 558
rect 2865 527 2870 558
rect 2814 523 2870 527
rect 2828 509 2856 523
rect 2056 437 2112 440
rect 2056 406 2061 437
rect 2107 406 2112 437
rect 2056 402 2112 406
rect 1733 335 2056 387
rect 1677 317 1733 320
rect 1677 286 1682 317
rect 1728 286 1733 317
rect 1677 282 1733 286
rect 1354 215 1677 267
rect 1298 197 1354 200
rect 1298 166 1303 197
rect 1349 166 1354 197
rect 1298 162 1354 166
rect 975 95 1298 147
rect 919 77 975 80
rect 919 46 924 77
rect 970 46 975 77
rect 919 42 975 46
rect 933 30 961 42
rect 990 28 1283 95
rect 1312 80 1340 162
rect 1369 147 1662 215
rect 1691 200 1719 282
rect 1748 267 2041 335
rect 2070 320 2098 402
rect 2127 387 2420 455
rect 2449 440 2477 486
rect 2491 455 2814 508
rect 2828 482 2829 509
rect 2855 482 2856 509
rect 2885 508 3178 576
rect 3207 561 3235 573
rect 3193 558 3249 561
rect 3193 527 3198 558
rect 3244 527 3249 558
rect 3193 523 3249 527
rect 2435 437 2491 440
rect 2435 406 2440 437
rect 2486 406 2491 437
rect 2435 402 2491 406
rect 2112 335 2435 387
rect 2056 317 2112 320
rect 2056 286 2061 317
rect 2107 286 2112 317
rect 2056 282 2112 286
rect 1733 215 2056 267
rect 1677 197 1733 200
rect 1677 166 1682 197
rect 1728 166 1733 197
rect 1677 162 1733 166
rect 1354 95 1677 147
rect 1298 77 1354 80
rect 1298 46 1303 77
rect 1349 46 1354 77
rect 1298 42 1354 46
rect 1312 30 1340 42
rect 1369 28 1662 95
rect 1691 80 1719 162
rect 1748 147 2041 215
rect 2070 200 2098 282
rect 2127 267 2420 335
rect 2449 320 2477 402
rect 2506 387 2799 455
rect 2828 440 2856 482
rect 2870 455 3193 508
rect 3207 505 3235 523
rect 3264 508 3557 576
rect 3586 561 3614 573
rect 3572 558 3628 561
rect 3572 527 3577 558
rect 3623 527 3628 558
rect 3572 523 3628 527
rect 3586 510 3614 523
rect 3207 478 3208 505
rect 3234 478 3235 505
rect 2814 437 2870 440
rect 2814 406 2819 437
rect 2865 406 2870 437
rect 2814 402 2870 406
rect 2491 335 2814 387
rect 2435 317 2491 320
rect 2435 286 2440 317
rect 2486 286 2491 317
rect 2435 282 2491 286
rect 2112 215 2435 267
rect 2056 197 2112 200
rect 2056 166 2061 197
rect 2107 166 2112 197
rect 2056 162 2112 166
rect 1733 95 2056 147
rect 1677 77 1733 80
rect 1677 46 1682 77
rect 1728 46 1733 77
rect 1677 42 1733 46
rect 1691 30 1719 42
rect 1748 28 2041 95
rect 2070 80 2098 162
rect 2127 147 2420 215
rect 2449 200 2477 282
rect 2506 267 2799 335
rect 2828 320 2856 402
rect 2885 387 3178 455
rect 3207 440 3235 478
rect 3249 455 3572 508
rect 3586 483 3587 510
rect 3613 483 3614 510
rect 3643 508 3936 576
rect 3965 561 3993 573
rect 3951 558 4007 561
rect 3951 527 3956 558
rect 4002 527 4007 558
rect 3951 523 4007 527
rect 3965 511 3993 523
rect 3193 437 3249 440
rect 3193 406 3198 437
rect 3244 406 3249 437
rect 3193 402 3249 406
rect 2870 335 3193 387
rect 2814 317 2870 320
rect 2814 286 2819 317
rect 2865 286 2870 317
rect 2814 282 2870 286
rect 2491 215 2814 267
rect 2435 197 2491 200
rect 2435 166 2440 197
rect 2486 166 2491 197
rect 2435 162 2491 166
rect 2112 95 2435 147
rect 2056 77 2112 80
rect 2056 46 2061 77
rect 2107 46 2112 77
rect 2056 42 2112 46
rect 2070 30 2098 42
rect 2127 28 2420 95
rect 2449 80 2477 162
rect 2506 147 2799 215
rect 2828 200 2856 282
rect 2885 267 3178 335
rect 3207 320 3235 402
rect 3264 387 3557 455
rect 3586 440 3614 483
rect 3628 455 3951 508
rect 3965 484 3966 511
rect 3992 484 3993 511
rect 4022 508 4315 576
rect 4344 561 4372 573
rect 4330 558 4386 561
rect 4330 527 4335 558
rect 4381 527 4386 558
rect 4330 523 4386 527
rect 3572 437 3628 440
rect 3572 406 3577 437
rect 3623 406 3628 437
rect 3572 402 3628 406
rect 3249 335 3572 387
rect 3193 317 3249 320
rect 3193 286 3198 317
rect 3244 286 3249 317
rect 3193 282 3249 286
rect 2870 215 3193 267
rect 2814 197 2870 200
rect 2814 166 2819 197
rect 2865 166 2870 197
rect 2814 162 2870 166
rect 2491 95 2814 147
rect 2435 77 2491 80
rect 2435 46 2440 77
rect 2486 46 2491 77
rect 2435 42 2491 46
rect 2449 30 2477 42
rect 2506 28 2799 95
rect 2828 80 2856 162
rect 2885 147 3178 215
rect 3207 200 3235 282
rect 3264 267 3557 335
rect 3586 320 3614 402
rect 3643 387 3936 455
rect 3965 440 3993 484
rect 4007 455 4330 508
rect 4344 506 4372 523
rect 4401 508 4694 576
rect 4723 561 4751 573
rect 4709 558 4765 561
rect 4709 527 4714 558
rect 4760 527 4765 558
rect 4709 523 4765 527
rect 4344 479 4345 506
rect 4371 479 4372 506
rect 3951 437 4007 440
rect 3951 406 3956 437
rect 4002 406 4007 437
rect 3951 402 4007 406
rect 3628 335 3951 387
rect 3572 317 3628 320
rect 3572 286 3577 317
rect 3623 286 3628 317
rect 3572 282 3628 286
rect 3249 215 3572 267
rect 3193 197 3249 200
rect 3193 166 3198 197
rect 3244 166 3249 197
rect 3193 162 3249 166
rect 2870 95 3193 147
rect 2814 77 2870 80
rect 2814 46 2819 77
rect 2865 46 2870 77
rect 2814 42 2870 46
rect 2828 30 2856 42
rect 2885 28 3178 95
rect 3207 80 3235 162
rect 3264 147 3557 215
rect 3586 200 3614 282
rect 3643 267 3936 335
rect 3965 320 3993 402
rect 4022 387 4315 455
rect 4344 440 4372 479
rect 4386 455 4709 508
rect 4723 506 4751 523
rect 4780 508 5073 576
rect 5102 561 5130 573
rect 5088 558 5144 561
rect 5088 527 5093 558
rect 5139 527 5144 558
rect 5088 523 5144 527
rect 4723 479 4724 506
rect 4750 479 4751 506
rect 4330 437 4386 440
rect 4330 406 4335 437
rect 4381 406 4386 437
rect 4330 402 4386 406
rect 4007 335 4330 387
rect 3951 317 4007 320
rect 3951 286 3956 317
rect 4002 286 4007 317
rect 3951 282 4007 286
rect 3628 215 3951 267
rect 3572 197 3628 200
rect 3572 166 3577 197
rect 3623 166 3628 197
rect 3572 162 3628 166
rect 3249 95 3572 147
rect 3193 77 3249 80
rect 3193 46 3198 77
rect 3244 46 3249 77
rect 3193 42 3249 46
rect 3207 30 3235 42
rect 3264 28 3557 95
rect 3586 80 3614 162
rect 3643 147 3936 215
rect 3965 200 3993 282
rect 4022 267 4315 335
rect 4344 320 4372 402
rect 4401 387 4694 455
rect 4723 440 4751 479
rect 4765 455 5088 508
rect 5102 507 5130 523
rect 5159 508 5452 576
rect 5481 561 5509 573
rect 5467 558 5523 561
rect 5467 527 5472 558
rect 5518 527 5523 558
rect 5467 523 5523 527
rect 5481 510 5509 523
rect 5102 480 5103 507
rect 5129 480 5130 507
rect 4709 437 4765 440
rect 4709 406 4714 437
rect 4760 406 4765 437
rect 4709 402 4765 406
rect 4386 335 4709 387
rect 4330 317 4386 320
rect 4330 286 4335 317
rect 4381 286 4386 317
rect 4330 282 4386 286
rect 4007 215 4330 267
rect 3951 197 4007 200
rect 3951 166 3956 197
rect 4002 166 4007 197
rect 3951 162 4007 166
rect 3628 95 3951 147
rect 3572 77 3628 80
rect 3572 46 3577 77
rect 3623 46 3628 77
rect 3572 42 3628 46
rect 3586 30 3614 42
rect 3643 28 3936 95
rect 3965 80 3993 162
rect 4022 147 4315 215
rect 4344 200 4372 282
rect 4401 267 4694 335
rect 4723 320 4751 402
rect 4780 387 5073 455
rect 5102 440 5130 480
rect 5144 455 5467 508
rect 5481 483 5482 510
rect 5508 483 5509 510
rect 5538 508 5831 576
rect 5860 561 5888 573
rect 5846 558 5902 561
rect 5846 527 5851 558
rect 5897 527 5902 558
rect 5846 523 5902 527
rect 5860 511 5888 523
rect 5088 437 5144 440
rect 5088 406 5093 437
rect 5139 406 5144 437
rect 5088 402 5144 406
rect 4765 335 5088 387
rect 4709 317 4765 320
rect 4709 286 4714 317
rect 4760 286 4765 317
rect 4709 282 4765 286
rect 4386 215 4709 267
rect 4330 197 4386 200
rect 4330 166 4335 197
rect 4381 166 4386 197
rect 4330 162 4386 166
rect 4007 95 4330 147
rect 3951 77 4007 80
rect 3951 46 3956 77
rect 4002 46 4007 77
rect 3951 42 4007 46
rect 3965 30 3993 42
rect 4022 28 4315 95
rect 4344 80 4372 162
rect 4401 147 4694 215
rect 4723 200 4751 282
rect 4780 267 5073 335
rect 5102 320 5130 402
rect 5159 387 5452 455
rect 5481 440 5509 483
rect 5523 455 5846 508
rect 5860 484 5861 511
rect 5887 484 5888 511
rect 5917 508 6210 576
rect 6239 561 6267 573
rect 6225 558 6281 561
rect 6225 527 6230 558
rect 6276 527 6281 558
rect 6225 523 6281 527
rect 6239 510 6267 523
rect 5467 437 5523 440
rect 5467 406 5472 437
rect 5518 406 5523 437
rect 5467 402 5523 406
rect 5144 335 5467 387
rect 5088 317 5144 320
rect 5088 286 5093 317
rect 5139 286 5144 317
rect 5088 282 5144 286
rect 4765 215 5088 267
rect 4709 197 4765 200
rect 4709 166 4714 197
rect 4760 166 4765 197
rect 4709 162 4765 166
rect 4386 95 4709 147
rect 4330 77 4386 80
rect 4330 46 4335 77
rect 4381 46 4386 77
rect 4330 42 4386 46
rect 4344 30 4372 42
rect 4401 28 4694 95
rect 4723 80 4751 162
rect 4780 147 5073 215
rect 5102 200 5130 282
rect 5159 267 5452 335
rect 5481 320 5509 402
rect 5538 387 5831 455
rect 5860 440 5888 484
rect 5902 455 6225 508
rect 6239 483 6240 510
rect 6266 483 6267 510
rect 6296 508 6589 576
rect 6618 561 6646 573
rect 6604 558 6660 561
rect 6604 527 6609 558
rect 6655 527 6660 558
rect 6604 523 6660 527
rect 6618 513 6646 523
rect 5846 437 5902 440
rect 5846 406 5851 437
rect 5897 406 5902 437
rect 5846 402 5902 406
rect 5523 335 5846 387
rect 5467 317 5523 320
rect 5467 286 5472 317
rect 5518 286 5523 317
rect 5467 282 5523 286
rect 5144 215 5467 267
rect 5088 197 5144 200
rect 5088 166 5093 197
rect 5139 166 5144 197
rect 5088 162 5144 166
rect 4765 95 5088 147
rect 4709 77 4765 80
rect 4709 46 4714 77
rect 4760 46 4765 77
rect 4709 42 4765 46
rect 4723 30 4751 42
rect 4780 28 5073 95
rect 5102 80 5130 162
rect 5159 147 5452 215
rect 5481 200 5509 282
rect 5538 267 5831 335
rect 5860 320 5888 402
rect 5917 387 6210 455
rect 6239 440 6267 483
rect 6281 455 6604 508
rect 6618 486 6619 513
rect 6645 486 6646 513
rect 6675 508 6968 576
rect 6997 561 7025 573
rect 6983 558 7039 561
rect 6983 527 6988 558
rect 7034 527 7039 558
rect 6983 523 7039 527
rect 6997 510 7025 523
rect 6225 437 6281 440
rect 6225 406 6230 437
rect 6276 406 6281 437
rect 6225 402 6281 406
rect 5902 335 6225 387
rect 5846 317 5902 320
rect 5846 286 5851 317
rect 5897 286 5902 317
rect 5846 282 5902 286
rect 5523 215 5846 267
rect 5467 197 5523 200
rect 5467 166 5472 197
rect 5518 166 5523 197
rect 5467 162 5523 166
rect 5144 95 5467 147
rect 5088 77 5144 80
rect 5088 46 5093 77
rect 5139 46 5144 77
rect 5088 42 5144 46
rect 5102 30 5130 42
rect 5159 28 5452 95
rect 5481 80 5509 162
rect 5538 147 5831 215
rect 5860 200 5888 282
rect 5917 267 6210 335
rect 6239 320 6267 402
rect 6296 387 6589 455
rect 6618 440 6646 486
rect 6660 455 6983 508
rect 6997 483 6998 510
rect 7024 483 7025 510
rect 7054 508 7347 576
rect 7376 561 7404 573
rect 7362 558 7418 561
rect 7362 527 7367 558
rect 7413 527 7418 558
rect 7362 523 7418 527
rect 7376 510 7404 523
rect 6604 437 6660 440
rect 6604 406 6609 437
rect 6655 406 6660 437
rect 6604 402 6660 406
rect 6281 335 6604 387
rect 6225 317 6281 320
rect 6225 286 6230 317
rect 6276 286 6281 317
rect 6225 282 6281 286
rect 5902 215 6225 267
rect 5846 197 5902 200
rect 5846 166 5851 197
rect 5897 166 5902 197
rect 5846 162 5902 166
rect 5523 95 5846 147
rect 5467 77 5523 80
rect 5467 46 5472 77
rect 5518 46 5523 77
rect 5467 42 5523 46
rect 5481 30 5509 42
rect 5538 28 5831 95
rect 5860 80 5888 162
rect 5917 147 6210 215
rect 6239 200 6267 282
rect 6296 267 6589 335
rect 6618 320 6646 402
rect 6675 387 6968 455
rect 6997 440 7025 483
rect 7039 455 7362 508
rect 7376 483 7377 510
rect 7403 483 7404 510
rect 7433 508 7599 576
rect 6983 437 7039 440
rect 6983 406 6988 437
rect 7034 406 7039 437
rect 6983 402 7039 406
rect 6660 335 6983 387
rect 6604 317 6660 320
rect 6604 286 6609 317
rect 6655 286 6660 317
rect 6604 282 6660 286
rect 6281 215 6604 267
rect 6225 197 6281 200
rect 6225 166 6230 197
rect 6276 166 6281 197
rect 6225 162 6281 166
rect 5902 95 6225 147
rect 5846 77 5902 80
rect 5846 46 5851 77
rect 5897 46 5902 77
rect 5846 42 5902 46
rect 5860 30 5888 42
rect 5917 28 6210 95
rect 6239 80 6267 162
rect 6296 147 6589 215
rect 6618 200 6646 282
rect 6675 267 6968 335
rect 6997 320 7025 402
rect 7054 387 7347 455
rect 7376 440 7404 483
rect 7418 455 7599 508
rect 7362 437 7418 440
rect 7362 406 7367 437
rect 7413 406 7418 437
rect 7362 402 7418 406
rect 7039 335 7362 387
rect 6983 317 7039 320
rect 6983 286 6988 317
rect 7034 286 7039 317
rect 6983 282 7039 286
rect 6660 215 6983 267
rect 6604 197 6660 200
rect 6604 166 6609 197
rect 6655 166 6660 197
rect 6604 162 6660 166
rect 6281 95 6604 147
rect 6225 77 6281 80
rect 6225 46 6230 77
rect 6276 46 6281 77
rect 6225 42 6281 46
rect 6239 30 6267 42
rect 6296 28 6589 95
rect 6618 80 6646 162
rect 6675 147 6968 215
rect 6997 200 7025 282
rect 7054 267 7347 335
rect 7376 320 7404 402
rect 7433 387 7599 455
rect 7418 335 7599 387
rect 7362 317 7418 320
rect 7362 286 7367 317
rect 7413 286 7418 317
rect 7362 282 7418 286
rect 7039 215 7362 267
rect 6983 197 7039 200
rect 6983 166 6988 197
rect 7034 166 7039 197
rect 6983 162 7039 166
rect 6660 95 6983 147
rect 6604 77 6660 80
rect 6604 46 6609 77
rect 6655 46 6660 77
rect 6604 42 6660 46
rect 6618 30 6646 42
rect 6675 28 6968 95
rect 6997 80 7025 162
rect 7054 147 7347 215
rect 7376 200 7404 282
rect 7433 267 7599 335
rect 7418 215 7599 267
rect 7362 197 7418 200
rect 7362 166 7367 197
rect 7413 166 7418 197
rect 7362 162 7418 166
rect 7039 95 7362 147
rect 6983 77 7039 80
rect 6983 46 6988 77
rect 7034 46 7039 77
rect 6983 42 7039 46
rect 6997 30 7025 42
rect 7054 28 7347 95
rect 7376 80 7404 162
rect 7433 147 7599 215
rect 7418 95 7599 147
rect 7362 77 7418 80
rect 7362 46 7367 77
rect 7413 46 7418 77
rect 7362 42 7418 46
rect 7376 30 7404 42
rect 7433 28 7599 95
rect -19 16 161 28
rect 217 16 540 28
rect 596 16 919 28
rect 975 16 1298 28
rect 1354 16 1677 28
rect 1733 16 2056 28
rect 2112 16 2435 28
rect 2491 16 2814 28
rect 2870 16 3193 28
rect 3249 16 3572 28
rect 3628 16 3951 28
rect 4007 16 4330 28
rect 4386 16 4709 28
rect 4765 16 5088 28
rect 5144 16 5467 28
rect 5523 16 5846 28
rect 5902 16 6225 28
rect 6281 16 6604 28
rect 6660 16 6983 28
rect 7039 16 7362 28
rect 7418 16 7599 28
rect -19 13 7599 16
rect -19 -13 34 13
rect 61 -13 109 13
rect 136 -13 242 13
rect 269 -13 317 13
rect 344 -13 413 13
rect 440 -13 488 13
rect 515 -13 621 13
rect 648 -13 696 13
rect 723 -13 792 13
rect 819 -13 867 13
rect 894 -13 1000 13
rect 1027 -13 1075 13
rect 1102 -13 1171 13
rect 1198 -13 1246 13
rect 1273 -13 1379 13
rect 1406 -13 1454 13
rect 1481 -13 1550 13
rect 1577 -13 1625 13
rect 1652 -13 1758 13
rect 1785 -13 1833 13
rect 1860 -13 1929 13
rect 1956 -13 2004 13
rect 2031 -13 2137 13
rect 2164 -13 2212 13
rect 2239 -13 2308 13
rect 2335 -13 2383 13
rect 2410 -13 2516 13
rect 2543 -13 2591 13
rect 2618 -13 2687 13
rect 2714 -13 2762 13
rect 2789 -13 2895 13
rect 2922 -13 2970 13
rect 2997 -13 3066 13
rect 3093 -13 3141 13
rect 3168 -13 3274 13
rect 3301 -13 3349 13
rect 3376 -13 3445 13
rect 3472 -13 3520 13
rect 3547 -13 3653 13
rect 3680 -13 3728 13
rect 3755 -13 3824 13
rect 3851 -13 3899 13
rect 3926 -13 4032 13
rect 4059 -13 4107 13
rect 4134 -13 4203 13
rect 4230 -13 4278 13
rect 4305 -13 4411 13
rect 4438 -13 4486 13
rect 4513 -13 4582 13
rect 4609 -13 4657 13
rect 4684 -13 4790 13
rect 4817 -13 4865 13
rect 4892 -13 4961 13
rect 4988 -13 5036 13
rect 5063 -13 5169 13
rect 5196 -13 5244 13
rect 5271 -13 5340 13
rect 5367 -13 5415 13
rect 5442 -13 5548 13
rect 5575 -13 5623 13
rect 5650 -13 5719 13
rect 5746 -13 5794 13
rect 5821 -13 5927 13
rect 5954 -13 6002 13
rect 6029 -13 6098 13
rect 6125 -13 6173 13
rect 6200 -13 6306 13
rect 6333 -13 6381 13
rect 6408 -13 6477 13
rect 6504 -13 6552 13
rect 6579 -13 6685 13
rect 6712 -13 6760 13
rect 6787 -13 6856 13
rect 6883 -13 6931 13
rect 6958 -13 7064 13
rect 7091 -13 7139 13
rect 7166 -13 7235 13
rect 7262 -13 7310 13
rect 7337 -13 7443 13
rect 7470 -13 7518 13
rect 7545 -13 7599 13
rect -19 -16 7599 -13
<< via2 >>
rect 166 2336 212 2367
rect 545 2336 591 2367
rect 166 2215 212 2246
rect 924 2336 970 2367
rect 545 2215 591 2246
rect 166 2095 212 2126
rect 1303 2336 1349 2367
rect 924 2215 970 2246
rect 545 2095 591 2126
rect 166 1975 212 2006
rect 1682 2336 1728 2367
rect 1303 2215 1349 2246
rect 924 2095 970 2126
rect 545 1975 591 2006
rect 2061 2336 2107 2367
rect 1682 2215 1728 2246
rect 1303 2095 1349 2126
rect 924 1975 970 2006
rect 166 1855 212 1886
rect 2440 2336 2486 2367
rect 2061 2215 2107 2246
rect 1682 2095 1728 2126
rect 1303 1975 1349 2006
rect 545 1855 591 1886
rect 2819 2336 2865 2367
rect 2440 2215 2486 2246
rect 2061 2095 2107 2126
rect 1682 1975 1728 2006
rect 924 1855 970 1886
rect 3198 2336 3244 2367
rect 2819 2215 2865 2246
rect 2440 2095 2486 2126
rect 2061 1975 2107 2006
rect 1303 1855 1349 1886
rect 3577 2336 3623 2367
rect 3198 2215 3244 2246
rect 2819 2095 2865 2126
rect 2440 1975 2486 2006
rect 1682 1855 1728 1886
rect 3956 2336 4002 2367
rect 3577 2215 3623 2246
rect 3198 2095 3244 2126
rect 2819 1975 2865 2006
rect 2061 1855 2107 1886
rect 4335 2336 4381 2367
rect 3956 2215 4002 2246
rect 3577 2095 3623 2126
rect 3198 1975 3244 2006
rect 2440 1855 2486 1886
rect 4714 2336 4760 2367
rect 4335 2215 4381 2246
rect 3956 2095 4002 2126
rect 3577 1975 3623 2006
rect 2819 1855 2865 1886
rect 5093 2336 5139 2367
rect 4714 2215 4760 2246
rect 4335 2095 4381 2126
rect 3956 1975 4002 2006
rect 3198 1855 3244 1886
rect 5472 2336 5518 2367
rect 5093 2215 5139 2246
rect 4714 2095 4760 2126
rect 4335 1975 4381 2006
rect 3577 1855 3623 1886
rect 5851 2336 5897 2367
rect 5472 2215 5518 2246
rect 5093 2095 5139 2126
rect 4714 1975 4760 2006
rect 3956 1855 4002 1886
rect 6230 2336 6276 2367
rect 5851 2215 5897 2246
rect 5472 2095 5518 2126
rect 5093 1975 5139 2006
rect 4335 1855 4381 1886
rect 6609 2336 6655 2367
rect 6230 2215 6276 2246
rect 5851 2095 5897 2126
rect 5472 1975 5518 2006
rect 4714 1855 4760 1886
rect 6988 2336 7034 2367
rect 6609 2215 6655 2246
rect 6230 2095 6276 2126
rect 5851 1975 5897 2006
rect 5093 1855 5139 1886
rect 7367 2336 7413 2367
rect 6988 2215 7034 2246
rect 6609 2095 6655 2126
rect 6230 1975 6276 2006
rect 5472 1855 5518 1886
rect 7367 2215 7413 2246
rect 6988 2095 7034 2126
rect 6609 1975 6655 2006
rect 5851 1855 5897 1886
rect 7367 2095 7413 2126
rect 6988 1975 7034 2006
rect 6230 1855 6276 1886
rect 7367 1975 7413 2006
rect 6609 1855 6655 1886
rect 6988 1855 7034 1886
rect 7367 1855 7413 1886
rect 166 1733 212 1764
rect 545 1733 591 1764
rect 166 1612 212 1643
rect 924 1733 970 1764
rect 545 1612 591 1643
rect 166 1492 212 1523
rect 1303 1733 1349 1764
rect 924 1612 970 1643
rect 545 1492 591 1523
rect 166 1372 212 1403
rect 1682 1733 1728 1764
rect 1303 1612 1349 1643
rect 924 1492 970 1523
rect 545 1372 591 1403
rect 2061 1733 2107 1764
rect 1682 1612 1728 1643
rect 1303 1492 1349 1523
rect 924 1372 970 1403
rect 166 1252 212 1283
rect 2440 1733 2486 1764
rect 2061 1612 2107 1643
rect 1682 1492 1728 1523
rect 1303 1372 1349 1403
rect 545 1252 591 1283
rect 2819 1733 2865 1764
rect 2440 1612 2486 1643
rect 2061 1492 2107 1523
rect 1682 1372 1728 1403
rect 924 1252 970 1283
rect 3198 1733 3244 1764
rect 2819 1612 2865 1643
rect 2440 1492 2486 1523
rect 2061 1372 2107 1403
rect 1303 1252 1349 1283
rect 3577 1733 3623 1764
rect 3198 1612 3244 1643
rect 2819 1492 2865 1523
rect 2440 1372 2486 1403
rect 1682 1252 1728 1283
rect 3956 1733 4002 1764
rect 3577 1612 3623 1643
rect 3198 1492 3244 1523
rect 2819 1372 2865 1403
rect 2061 1252 2107 1283
rect 4335 1733 4381 1764
rect 3956 1612 4002 1643
rect 3577 1492 3623 1523
rect 3198 1372 3244 1403
rect 2440 1252 2486 1283
rect 4714 1733 4760 1764
rect 4335 1612 4381 1643
rect 3956 1492 4002 1523
rect 3577 1372 3623 1403
rect 2819 1252 2865 1283
rect 5093 1733 5139 1764
rect 4714 1612 4760 1643
rect 4335 1492 4381 1523
rect 3956 1372 4002 1403
rect 3198 1252 3244 1283
rect 5472 1733 5518 1764
rect 5093 1612 5139 1643
rect 4714 1492 4760 1523
rect 4335 1372 4381 1403
rect 3577 1252 3623 1283
rect 5851 1733 5897 1764
rect 5472 1612 5518 1643
rect 5093 1492 5139 1523
rect 4714 1372 4760 1403
rect 3956 1252 4002 1283
rect 6230 1733 6276 1764
rect 5851 1612 5897 1643
rect 5472 1492 5518 1523
rect 5093 1372 5139 1403
rect 4335 1252 4381 1283
rect 6609 1733 6655 1764
rect 6230 1612 6276 1643
rect 5851 1492 5897 1523
rect 5472 1372 5518 1403
rect 4714 1252 4760 1283
rect 6988 1733 7034 1764
rect 6609 1612 6655 1643
rect 6230 1492 6276 1523
rect 5851 1372 5897 1403
rect 5093 1252 5139 1283
rect 7367 1733 7413 1764
rect 6988 1612 7034 1643
rect 6609 1492 6655 1523
rect 6230 1372 6276 1403
rect 5472 1252 5518 1283
rect 7367 1612 7413 1643
rect 6988 1492 7034 1523
rect 6609 1372 6655 1403
rect 5851 1252 5897 1283
rect 7367 1492 7413 1523
rect 6988 1372 7034 1403
rect 6230 1252 6276 1283
rect 7367 1372 7413 1403
rect 6609 1252 6655 1283
rect 6988 1252 7034 1283
rect 7367 1252 7413 1283
rect 166 1130 212 1161
rect 545 1130 591 1161
rect 166 1009 212 1040
rect 924 1130 970 1161
rect 545 1009 591 1040
rect 166 889 212 920
rect 1303 1130 1349 1161
rect 924 1009 970 1040
rect 545 889 591 920
rect 166 769 212 800
rect 1682 1130 1728 1161
rect 1303 1009 1349 1040
rect 924 889 970 920
rect 545 769 591 800
rect 2061 1130 2107 1161
rect 1682 1009 1728 1040
rect 1303 889 1349 920
rect 924 769 970 800
rect 166 649 212 680
rect 2440 1130 2486 1161
rect 2061 1009 2107 1040
rect 1682 889 1728 920
rect 1303 769 1349 800
rect 545 649 591 680
rect 2819 1130 2865 1161
rect 2440 1009 2486 1040
rect 2061 889 2107 920
rect 1682 769 1728 800
rect 924 649 970 680
rect 3198 1130 3244 1161
rect 2819 1009 2865 1040
rect 2440 889 2486 920
rect 2061 769 2107 800
rect 1303 649 1349 680
rect 3577 1130 3623 1161
rect 3198 1009 3244 1040
rect 2819 889 2865 920
rect 2440 769 2486 800
rect 1682 649 1728 680
rect 3956 1130 4002 1161
rect 3577 1009 3623 1040
rect 3198 889 3244 920
rect 2819 769 2865 800
rect 2061 649 2107 680
rect 4335 1130 4381 1161
rect 3956 1009 4002 1040
rect 3577 889 3623 920
rect 3198 769 3244 800
rect 2440 649 2486 680
rect 4714 1130 4760 1161
rect 4335 1009 4381 1040
rect 3956 889 4002 920
rect 3577 769 3623 800
rect 2819 649 2865 680
rect 5093 1130 5139 1161
rect 4714 1009 4760 1040
rect 4335 889 4381 920
rect 3956 769 4002 800
rect 3198 649 3244 680
rect 5472 1130 5518 1161
rect 5093 1009 5139 1040
rect 4714 889 4760 920
rect 4335 769 4381 800
rect 3577 649 3623 680
rect 5851 1130 5897 1161
rect 5472 1009 5518 1040
rect 5093 889 5139 920
rect 4714 769 4760 800
rect 3956 649 4002 680
rect 6230 1130 6276 1161
rect 5851 1009 5897 1040
rect 5472 889 5518 920
rect 5093 769 5139 800
rect 4335 649 4381 680
rect 6609 1130 6655 1161
rect 6230 1009 6276 1040
rect 5851 889 5897 920
rect 5472 769 5518 800
rect 4714 649 4760 680
rect 6988 1130 7034 1161
rect 6609 1009 6655 1040
rect 6230 889 6276 920
rect 5851 769 5897 800
rect 5093 649 5139 680
rect 7367 1130 7413 1161
rect 6988 1009 7034 1040
rect 6609 889 6655 920
rect 6230 769 6276 800
rect 5472 649 5518 680
rect 7367 1009 7413 1040
rect 6988 889 7034 920
rect 6609 769 6655 800
rect 5851 649 5897 680
rect 7367 889 7413 920
rect 6988 769 7034 800
rect 6230 649 6276 680
rect 7367 769 7413 800
rect 6609 649 6655 680
rect 6988 649 7034 680
rect 7367 649 7413 680
rect 166 527 212 558
rect 545 527 591 558
rect 924 527 970 558
rect 166 406 212 437
rect 1303 527 1349 558
rect 545 406 591 437
rect 166 286 212 317
rect 1682 527 1728 558
rect 924 406 970 437
rect 545 286 591 317
rect 166 166 212 197
rect 2061 527 2107 558
rect 1303 406 1349 437
rect 924 286 970 317
rect 545 166 591 197
rect 166 46 212 77
rect 2440 527 2486 558
rect 1682 406 1728 437
rect 1303 286 1349 317
rect 924 166 970 197
rect 545 46 591 77
rect 2819 527 2865 558
rect 2061 406 2107 437
rect 1682 286 1728 317
rect 1303 166 1349 197
rect 924 46 970 77
rect 3198 527 3244 558
rect 2440 406 2486 437
rect 2061 286 2107 317
rect 1682 166 1728 197
rect 1303 46 1349 77
rect 3577 527 3623 558
rect 2819 406 2865 437
rect 2440 286 2486 317
rect 2061 166 2107 197
rect 1682 46 1728 77
rect 3956 527 4002 558
rect 3198 406 3244 437
rect 2819 286 2865 317
rect 2440 166 2486 197
rect 2061 46 2107 77
rect 4335 527 4381 558
rect 3577 406 3623 437
rect 3198 286 3244 317
rect 2819 166 2865 197
rect 2440 46 2486 77
rect 4714 527 4760 558
rect 3956 406 4002 437
rect 3577 286 3623 317
rect 3198 166 3244 197
rect 2819 46 2865 77
rect 5093 527 5139 558
rect 4335 406 4381 437
rect 3956 286 4002 317
rect 3577 166 3623 197
rect 3198 46 3244 77
rect 5472 527 5518 558
rect 4714 406 4760 437
rect 4335 286 4381 317
rect 3956 166 4002 197
rect 3577 46 3623 77
rect 5851 527 5897 558
rect 5093 406 5139 437
rect 4714 286 4760 317
rect 4335 166 4381 197
rect 3956 46 4002 77
rect 6230 527 6276 558
rect 5472 406 5518 437
rect 5093 286 5139 317
rect 4714 166 4760 197
rect 4335 46 4381 77
rect 6609 527 6655 558
rect 5851 406 5897 437
rect 5472 286 5518 317
rect 5093 166 5139 197
rect 4714 46 4760 77
rect 6988 527 7034 558
rect 6230 406 6276 437
rect 5851 286 5897 317
rect 5472 166 5518 197
rect 5093 46 5139 77
rect 7367 527 7413 558
rect 6609 406 6655 437
rect 6230 286 6276 317
rect 5851 166 5897 197
rect 5472 46 5518 77
rect 6988 406 7034 437
rect 6609 286 6655 317
rect 6230 166 6276 197
rect 5851 46 5897 77
rect 7367 406 7413 437
rect 6988 286 7034 317
rect 6609 166 6655 197
rect 6230 46 6276 77
rect 7367 286 7413 317
rect 6988 166 7034 197
rect 6609 46 6655 77
rect 7367 166 7413 197
rect 6988 46 7034 77
rect 7367 46 7413 77
<< metal3 >>
rect 161 2367 217 2370
rect 161 2366 166 2367
rect 53 2336 166 2366
rect 212 2366 217 2367
rect 540 2367 596 2370
rect 540 2366 545 2367
rect 212 2336 326 2366
rect 432 2336 545 2366
rect 591 2366 596 2367
rect 919 2367 975 2370
rect 919 2366 924 2367
rect 591 2336 705 2366
rect 811 2336 924 2366
rect 970 2366 975 2367
rect 1298 2367 1354 2370
rect 1298 2366 1303 2367
rect 970 2336 1084 2366
rect 1190 2336 1303 2366
rect 1349 2366 1354 2367
rect 1677 2367 1733 2370
rect 1677 2366 1682 2367
rect 1349 2336 1463 2366
rect 1569 2336 1682 2366
rect 1728 2366 1733 2367
rect 2056 2367 2112 2370
rect 2056 2366 2061 2367
rect 1728 2336 1842 2366
rect 1948 2336 2061 2366
rect 2107 2366 2112 2367
rect 2435 2367 2491 2370
rect 2435 2366 2440 2367
rect 2107 2336 2221 2366
rect 2327 2336 2440 2366
rect 2486 2366 2491 2367
rect 2814 2367 2870 2370
rect 2814 2366 2819 2367
rect 2486 2336 2600 2366
rect 2706 2336 2819 2366
rect 2865 2366 2870 2367
rect 3193 2367 3249 2370
rect 3193 2366 3198 2367
rect 2865 2336 2979 2366
rect 3085 2336 3198 2366
rect 3244 2366 3249 2367
rect 3572 2367 3628 2370
rect 3572 2366 3577 2367
rect 3244 2336 3358 2366
rect 3464 2336 3577 2366
rect 3623 2366 3628 2367
rect 3951 2367 4007 2370
rect 3951 2366 3956 2367
rect 3623 2336 3737 2366
rect 3843 2336 3956 2366
rect 4002 2366 4007 2367
rect 4330 2367 4386 2370
rect 4330 2366 4335 2367
rect 4002 2336 4116 2366
rect 4222 2336 4335 2366
rect 4381 2366 4386 2367
rect 4709 2367 4765 2370
rect 4709 2366 4714 2367
rect 4381 2336 4495 2366
rect 4601 2336 4714 2366
rect 4760 2366 4765 2367
rect 5088 2367 5144 2370
rect 5088 2366 5093 2367
rect 4760 2336 4874 2366
rect 4980 2336 5093 2366
rect 5139 2366 5144 2367
rect 5467 2367 5523 2370
rect 5467 2366 5472 2367
rect 5139 2336 5253 2366
rect 5359 2336 5472 2366
rect 5518 2366 5523 2367
rect 5846 2367 5902 2370
rect 5846 2366 5851 2367
rect 5518 2336 5632 2366
rect 5738 2336 5851 2366
rect 5897 2366 5902 2367
rect 6225 2367 6281 2370
rect 6225 2366 6230 2367
rect 5897 2336 6011 2366
rect 6117 2336 6230 2366
rect 6276 2366 6281 2367
rect 6604 2367 6660 2370
rect 6604 2366 6609 2367
rect 6276 2336 6390 2366
rect 6496 2336 6609 2366
rect 6655 2366 6660 2367
rect 6983 2367 7039 2370
rect 6983 2366 6988 2367
rect 6655 2336 6769 2366
rect 6875 2336 6988 2366
rect 7034 2366 7039 2367
rect 7362 2367 7418 2370
rect 7362 2366 7367 2367
rect 7034 2336 7148 2366
rect 7254 2336 7367 2366
rect 7413 2366 7418 2367
rect 7413 2336 7527 2366
rect 161 2332 217 2336
rect 540 2332 596 2336
rect 919 2332 975 2336
rect 1298 2332 1354 2336
rect 1677 2332 1733 2336
rect 2056 2332 2112 2336
rect 2435 2332 2491 2336
rect 2814 2332 2870 2336
rect 3193 2332 3249 2336
rect 3572 2332 3628 2336
rect 3951 2332 4007 2336
rect 4330 2332 4386 2336
rect 4709 2332 4765 2336
rect 5088 2332 5144 2336
rect 5467 2332 5523 2336
rect 5846 2332 5902 2336
rect 6225 2332 6281 2336
rect 6604 2332 6660 2336
rect 6983 2332 7039 2336
rect 7362 2332 7418 2336
rect -19 2274 -16 2306
rect 16 2305 19 2306
rect 360 2305 363 2306
rect 16 2275 146 2305
rect 232 2275 363 2305
rect 16 2274 19 2275
rect 360 2274 363 2275
rect 395 2305 398 2306
rect 739 2305 742 2306
rect 395 2275 525 2305
rect 611 2275 742 2305
rect 395 2274 398 2275
rect 739 2274 742 2275
rect 774 2305 777 2306
rect 1118 2305 1121 2306
rect 774 2275 904 2305
rect 990 2275 1121 2305
rect 774 2274 777 2275
rect 1118 2274 1121 2275
rect 1153 2305 1156 2306
rect 1497 2305 1500 2306
rect 1153 2275 1283 2305
rect 1369 2275 1500 2305
rect 1153 2274 1156 2275
rect 1497 2274 1500 2275
rect 1532 2305 1535 2306
rect 1876 2305 1879 2306
rect 1532 2275 1662 2305
rect 1748 2275 1879 2305
rect 1532 2274 1535 2275
rect 1876 2274 1879 2275
rect 1911 2305 1914 2306
rect 2255 2305 2258 2306
rect 1911 2275 2041 2305
rect 2127 2275 2258 2305
rect 1911 2274 1914 2275
rect 2255 2274 2258 2275
rect 2290 2305 2293 2306
rect 2634 2305 2637 2306
rect 2290 2275 2420 2305
rect 2506 2275 2637 2305
rect 2290 2274 2293 2275
rect 2634 2274 2637 2275
rect 2669 2305 2672 2306
rect 3013 2305 3016 2306
rect 2669 2275 2799 2305
rect 2885 2275 3016 2305
rect 2669 2274 2672 2275
rect 3013 2274 3016 2275
rect 3048 2305 3051 2306
rect 3392 2305 3395 2306
rect 3048 2275 3178 2305
rect 3264 2275 3395 2305
rect 3048 2274 3051 2275
rect 3392 2274 3395 2275
rect 3427 2305 3430 2306
rect 3771 2305 3774 2306
rect 3427 2275 3557 2305
rect 3643 2275 3774 2305
rect 3427 2274 3430 2275
rect 3771 2274 3774 2275
rect 3806 2305 3809 2306
rect 4150 2305 4153 2306
rect 3806 2275 3936 2305
rect 4022 2275 4153 2305
rect 3806 2274 3809 2275
rect 4150 2274 4153 2275
rect 4185 2305 4188 2306
rect 4529 2305 4532 2306
rect 4185 2275 4315 2305
rect 4401 2275 4532 2305
rect 4185 2274 4188 2275
rect 4529 2274 4532 2275
rect 4564 2305 4567 2306
rect 4908 2305 4911 2306
rect 4564 2275 4694 2305
rect 4780 2275 4911 2305
rect 4564 2274 4567 2275
rect 4908 2274 4911 2275
rect 4943 2305 4946 2306
rect 5287 2305 5290 2306
rect 4943 2275 5073 2305
rect 5159 2275 5290 2305
rect 4943 2274 4946 2275
rect 5287 2274 5290 2275
rect 5322 2305 5325 2306
rect 5666 2305 5669 2306
rect 5322 2275 5452 2305
rect 5538 2275 5669 2305
rect 5322 2274 5325 2275
rect 5666 2274 5669 2275
rect 5701 2305 5704 2306
rect 6045 2305 6048 2306
rect 5701 2275 5831 2305
rect 5917 2275 6048 2305
rect 5701 2274 5704 2275
rect 6045 2274 6048 2275
rect 6080 2305 6083 2306
rect 6424 2305 6427 2306
rect 6080 2275 6210 2305
rect 6296 2275 6427 2305
rect 6080 2274 6083 2275
rect 6424 2274 6427 2275
rect 6459 2305 6462 2306
rect 6803 2305 6806 2306
rect 6459 2275 6589 2305
rect 6675 2275 6806 2305
rect 6459 2274 6462 2275
rect 6803 2274 6806 2275
rect 6838 2305 6841 2306
rect 7182 2305 7185 2306
rect 6838 2275 6968 2305
rect 7054 2275 7185 2305
rect 6838 2274 6841 2275
rect 7182 2274 7185 2275
rect 7217 2305 7220 2306
rect 7561 2305 7564 2306
rect 7217 2275 7347 2305
rect 7433 2275 7564 2305
rect 7217 2274 7220 2275
rect 7561 2274 7564 2275
rect 7596 2274 7599 2306
rect 161 2246 217 2249
rect 161 2245 166 2246
rect 53 2215 166 2245
rect 212 2245 217 2246
rect 540 2246 596 2249
rect 540 2245 545 2246
rect 212 2215 326 2245
rect 432 2215 545 2245
rect 591 2245 596 2246
rect 919 2246 975 2249
rect 919 2245 924 2246
rect 591 2215 705 2245
rect 811 2215 924 2245
rect 970 2245 975 2246
rect 1298 2246 1354 2249
rect 1298 2245 1303 2246
rect 970 2215 1084 2245
rect 1190 2215 1303 2245
rect 1349 2245 1354 2246
rect 1677 2246 1733 2249
rect 1677 2245 1682 2246
rect 1349 2215 1463 2245
rect 1569 2215 1682 2245
rect 1728 2245 1733 2246
rect 2056 2246 2112 2249
rect 2056 2245 2061 2246
rect 1728 2215 1842 2245
rect 1948 2215 2061 2245
rect 2107 2245 2112 2246
rect 2435 2246 2491 2249
rect 2435 2245 2440 2246
rect 2107 2215 2221 2245
rect 2327 2215 2440 2245
rect 2486 2245 2491 2246
rect 2814 2246 2870 2249
rect 2814 2245 2819 2246
rect 2486 2215 2600 2245
rect 2706 2215 2819 2245
rect 2865 2245 2870 2246
rect 3193 2246 3249 2249
rect 3193 2245 3198 2246
rect 2865 2215 2979 2245
rect 3085 2215 3198 2245
rect 3244 2245 3249 2246
rect 3572 2246 3628 2249
rect 3572 2245 3577 2246
rect 3244 2215 3358 2245
rect 3464 2215 3577 2245
rect 3623 2245 3628 2246
rect 3951 2246 4007 2249
rect 3951 2245 3956 2246
rect 3623 2215 3737 2245
rect 3843 2215 3956 2245
rect 4002 2245 4007 2246
rect 4330 2246 4386 2249
rect 4330 2245 4335 2246
rect 4002 2215 4116 2245
rect 4222 2215 4335 2245
rect 4381 2245 4386 2246
rect 4709 2246 4765 2249
rect 4709 2245 4714 2246
rect 4381 2215 4495 2245
rect 4601 2215 4714 2245
rect 4760 2245 4765 2246
rect 5088 2246 5144 2249
rect 5088 2245 5093 2246
rect 4760 2215 4874 2245
rect 4980 2215 5093 2245
rect 5139 2245 5144 2246
rect 5467 2246 5523 2249
rect 5467 2245 5472 2246
rect 5139 2215 5253 2245
rect 5359 2215 5472 2245
rect 5518 2245 5523 2246
rect 5846 2246 5902 2249
rect 5846 2245 5851 2246
rect 5518 2215 5632 2245
rect 5738 2215 5851 2245
rect 5897 2245 5902 2246
rect 6225 2246 6281 2249
rect 6225 2245 6230 2246
rect 5897 2215 6011 2245
rect 6117 2215 6230 2245
rect 6276 2245 6281 2246
rect 6604 2246 6660 2249
rect 6604 2245 6609 2246
rect 6276 2215 6390 2245
rect 6496 2215 6609 2245
rect 6655 2245 6660 2246
rect 6983 2246 7039 2249
rect 6983 2245 6988 2246
rect 6655 2215 6769 2245
rect 6875 2215 6988 2245
rect 7034 2245 7039 2246
rect 7362 2246 7418 2249
rect 7362 2245 7367 2246
rect 7034 2215 7148 2245
rect 7254 2215 7367 2245
rect 7413 2245 7418 2246
rect 7413 2215 7527 2245
rect 161 2211 217 2215
rect 540 2211 596 2215
rect 919 2211 975 2215
rect 1298 2211 1354 2215
rect 1677 2211 1733 2215
rect 2056 2211 2112 2215
rect 2435 2211 2491 2215
rect 2814 2211 2870 2215
rect 3193 2211 3249 2215
rect 3572 2211 3628 2215
rect 3951 2211 4007 2215
rect 4330 2211 4386 2215
rect 4709 2211 4765 2215
rect 5088 2211 5144 2215
rect 5467 2211 5523 2215
rect 5846 2211 5902 2215
rect 6225 2211 6281 2215
rect 6604 2211 6660 2215
rect 6983 2211 7039 2215
rect 7362 2211 7418 2215
rect -19 2154 -16 2186
rect 16 2185 19 2186
rect 360 2185 363 2186
rect 16 2155 146 2185
rect 232 2155 363 2185
rect 16 2154 19 2155
rect 360 2154 363 2155
rect 395 2185 398 2186
rect 739 2185 742 2186
rect 395 2155 525 2185
rect 611 2155 742 2185
rect 395 2154 398 2155
rect 739 2154 742 2155
rect 774 2185 777 2186
rect 1118 2185 1121 2186
rect 774 2155 904 2185
rect 990 2155 1121 2185
rect 774 2154 777 2155
rect 1118 2154 1121 2155
rect 1153 2185 1156 2186
rect 1497 2185 1500 2186
rect 1153 2155 1283 2185
rect 1369 2155 1500 2185
rect 1153 2154 1156 2155
rect 1497 2154 1500 2155
rect 1532 2185 1535 2186
rect 1876 2185 1879 2186
rect 1532 2155 1662 2185
rect 1748 2155 1879 2185
rect 1532 2154 1535 2155
rect 1876 2154 1879 2155
rect 1911 2185 1914 2186
rect 2255 2185 2258 2186
rect 1911 2155 2041 2185
rect 2127 2155 2258 2185
rect 1911 2154 1914 2155
rect 2255 2154 2258 2155
rect 2290 2185 2293 2186
rect 2634 2185 2637 2186
rect 2290 2155 2420 2185
rect 2506 2155 2637 2185
rect 2290 2154 2293 2155
rect 2634 2154 2637 2155
rect 2669 2185 2672 2186
rect 3013 2185 3016 2186
rect 2669 2155 2799 2185
rect 2885 2155 3016 2185
rect 2669 2154 2672 2155
rect 3013 2154 3016 2155
rect 3048 2185 3051 2186
rect 3392 2185 3395 2186
rect 3048 2155 3178 2185
rect 3264 2155 3395 2185
rect 3048 2154 3051 2155
rect 3392 2154 3395 2155
rect 3427 2185 3430 2186
rect 3771 2185 3774 2186
rect 3427 2155 3557 2185
rect 3643 2155 3774 2185
rect 3427 2154 3430 2155
rect 3771 2154 3774 2155
rect 3806 2185 3809 2186
rect 4150 2185 4153 2186
rect 3806 2155 3936 2185
rect 4022 2155 4153 2185
rect 3806 2154 3809 2155
rect 4150 2154 4153 2155
rect 4185 2185 4188 2186
rect 4529 2185 4532 2186
rect 4185 2155 4315 2185
rect 4401 2155 4532 2185
rect 4185 2154 4188 2155
rect 4529 2154 4532 2155
rect 4564 2185 4567 2186
rect 4908 2185 4911 2186
rect 4564 2155 4694 2185
rect 4780 2155 4911 2185
rect 4564 2154 4567 2155
rect 4908 2154 4911 2155
rect 4943 2185 4946 2186
rect 5287 2185 5290 2186
rect 4943 2155 5073 2185
rect 5159 2155 5290 2185
rect 4943 2154 4946 2155
rect 5287 2154 5290 2155
rect 5322 2185 5325 2186
rect 5666 2185 5669 2186
rect 5322 2155 5452 2185
rect 5538 2155 5669 2185
rect 5322 2154 5325 2155
rect 5666 2154 5669 2155
rect 5701 2185 5704 2186
rect 6045 2185 6048 2186
rect 5701 2155 5831 2185
rect 5917 2155 6048 2185
rect 5701 2154 5704 2155
rect 6045 2154 6048 2155
rect 6080 2185 6083 2186
rect 6424 2185 6427 2186
rect 6080 2155 6210 2185
rect 6296 2155 6427 2185
rect 6080 2154 6083 2155
rect 6424 2154 6427 2155
rect 6459 2185 6462 2186
rect 6803 2185 6806 2186
rect 6459 2155 6589 2185
rect 6675 2155 6806 2185
rect 6459 2154 6462 2155
rect 6803 2154 6806 2155
rect 6838 2185 6841 2186
rect 7182 2185 7185 2186
rect 6838 2155 6968 2185
rect 7054 2155 7185 2185
rect 6838 2154 6841 2155
rect 7182 2154 7185 2155
rect 7217 2185 7220 2186
rect 7561 2185 7564 2186
rect 7217 2155 7347 2185
rect 7433 2155 7564 2185
rect 7217 2154 7220 2155
rect 7561 2154 7564 2155
rect 7596 2154 7599 2186
rect 161 2126 217 2129
rect 161 2125 166 2126
rect 53 2095 166 2125
rect 212 2125 217 2126
rect 540 2126 596 2129
rect 540 2125 545 2126
rect 212 2095 326 2125
rect 432 2095 545 2125
rect 591 2125 596 2126
rect 919 2126 975 2129
rect 919 2125 924 2126
rect 591 2095 705 2125
rect 811 2095 924 2125
rect 970 2125 975 2126
rect 1298 2126 1354 2129
rect 1298 2125 1303 2126
rect 970 2095 1084 2125
rect 1190 2095 1303 2125
rect 1349 2125 1354 2126
rect 1677 2126 1733 2129
rect 1677 2125 1682 2126
rect 1349 2095 1463 2125
rect 1569 2095 1682 2125
rect 1728 2125 1733 2126
rect 2056 2126 2112 2129
rect 2056 2125 2061 2126
rect 1728 2095 1842 2125
rect 1948 2095 2061 2125
rect 2107 2125 2112 2126
rect 2435 2126 2491 2129
rect 2435 2125 2440 2126
rect 2107 2095 2221 2125
rect 2327 2095 2440 2125
rect 2486 2125 2491 2126
rect 2814 2126 2870 2129
rect 2814 2125 2819 2126
rect 2486 2095 2600 2125
rect 2706 2095 2819 2125
rect 2865 2125 2870 2126
rect 3193 2126 3249 2129
rect 3193 2125 3198 2126
rect 2865 2095 2979 2125
rect 3085 2095 3198 2125
rect 3244 2125 3249 2126
rect 3572 2126 3628 2129
rect 3572 2125 3577 2126
rect 3244 2095 3358 2125
rect 3464 2095 3577 2125
rect 3623 2125 3628 2126
rect 3951 2126 4007 2129
rect 3951 2125 3956 2126
rect 3623 2095 3737 2125
rect 3843 2095 3956 2125
rect 4002 2125 4007 2126
rect 4330 2126 4386 2129
rect 4330 2125 4335 2126
rect 4002 2095 4116 2125
rect 4222 2095 4335 2125
rect 4381 2125 4386 2126
rect 4709 2126 4765 2129
rect 4709 2125 4714 2126
rect 4381 2095 4495 2125
rect 4601 2095 4714 2125
rect 4760 2125 4765 2126
rect 5088 2126 5144 2129
rect 5088 2125 5093 2126
rect 4760 2095 4874 2125
rect 4980 2095 5093 2125
rect 5139 2125 5144 2126
rect 5467 2126 5523 2129
rect 5467 2125 5472 2126
rect 5139 2095 5253 2125
rect 5359 2095 5472 2125
rect 5518 2125 5523 2126
rect 5846 2126 5902 2129
rect 5846 2125 5851 2126
rect 5518 2095 5632 2125
rect 5738 2095 5851 2125
rect 5897 2125 5902 2126
rect 6225 2126 6281 2129
rect 6225 2125 6230 2126
rect 5897 2095 6011 2125
rect 6117 2095 6230 2125
rect 6276 2125 6281 2126
rect 6604 2126 6660 2129
rect 6604 2125 6609 2126
rect 6276 2095 6390 2125
rect 6496 2095 6609 2125
rect 6655 2125 6660 2126
rect 6983 2126 7039 2129
rect 6983 2125 6988 2126
rect 6655 2095 6769 2125
rect 6875 2095 6988 2125
rect 7034 2125 7039 2126
rect 7362 2126 7418 2129
rect 7362 2125 7367 2126
rect 7034 2095 7148 2125
rect 7254 2095 7367 2125
rect 7413 2125 7418 2126
rect 7413 2095 7527 2125
rect 161 2091 217 2095
rect 540 2091 596 2095
rect 919 2091 975 2095
rect 1298 2091 1354 2095
rect 1677 2091 1733 2095
rect 2056 2091 2112 2095
rect 2435 2091 2491 2095
rect 2814 2091 2870 2095
rect 3193 2091 3249 2095
rect 3572 2091 3628 2095
rect 3951 2091 4007 2095
rect 4330 2091 4386 2095
rect 4709 2091 4765 2095
rect 5088 2091 5144 2095
rect 5467 2091 5523 2095
rect 5846 2091 5902 2095
rect 6225 2091 6281 2095
rect 6604 2091 6660 2095
rect 6983 2091 7039 2095
rect 7362 2091 7418 2095
rect -19 2034 -16 2066
rect 16 2065 19 2066
rect 360 2065 363 2066
rect 16 2035 146 2065
rect 232 2035 363 2065
rect 16 2034 19 2035
rect 360 2034 363 2035
rect 395 2065 398 2066
rect 739 2065 742 2066
rect 395 2035 525 2065
rect 611 2035 742 2065
rect 395 2034 398 2035
rect 739 2034 742 2035
rect 774 2065 777 2066
rect 1118 2065 1121 2066
rect 774 2035 904 2065
rect 990 2035 1121 2065
rect 774 2034 777 2035
rect 1118 2034 1121 2035
rect 1153 2065 1156 2066
rect 1497 2065 1500 2066
rect 1153 2035 1283 2065
rect 1369 2035 1500 2065
rect 1153 2034 1156 2035
rect 1497 2034 1500 2035
rect 1532 2065 1535 2066
rect 1876 2065 1879 2066
rect 1532 2035 1662 2065
rect 1748 2035 1879 2065
rect 1532 2034 1535 2035
rect 1876 2034 1879 2035
rect 1911 2065 1914 2066
rect 2255 2065 2258 2066
rect 1911 2035 2041 2065
rect 2127 2035 2258 2065
rect 1911 2034 1914 2035
rect 2255 2034 2258 2035
rect 2290 2065 2293 2066
rect 2634 2065 2637 2066
rect 2290 2035 2420 2065
rect 2506 2035 2637 2065
rect 2290 2034 2293 2035
rect 2634 2034 2637 2035
rect 2669 2065 2672 2066
rect 3013 2065 3016 2066
rect 2669 2035 2799 2065
rect 2885 2035 3016 2065
rect 2669 2034 2672 2035
rect 3013 2034 3016 2035
rect 3048 2065 3051 2066
rect 3392 2065 3395 2066
rect 3048 2035 3178 2065
rect 3264 2035 3395 2065
rect 3048 2034 3051 2035
rect 3392 2034 3395 2035
rect 3427 2065 3430 2066
rect 3771 2065 3774 2066
rect 3427 2035 3557 2065
rect 3643 2035 3774 2065
rect 3427 2034 3430 2035
rect 3771 2034 3774 2035
rect 3806 2065 3809 2066
rect 4150 2065 4153 2066
rect 3806 2035 3936 2065
rect 4022 2035 4153 2065
rect 3806 2034 3809 2035
rect 4150 2034 4153 2035
rect 4185 2065 4188 2066
rect 4529 2065 4532 2066
rect 4185 2035 4315 2065
rect 4401 2035 4532 2065
rect 4185 2034 4188 2035
rect 4529 2034 4532 2035
rect 4564 2065 4567 2066
rect 4908 2065 4911 2066
rect 4564 2035 4694 2065
rect 4780 2035 4911 2065
rect 4564 2034 4567 2035
rect 4908 2034 4911 2035
rect 4943 2065 4946 2066
rect 5287 2065 5290 2066
rect 4943 2035 5073 2065
rect 5159 2035 5290 2065
rect 4943 2034 4946 2035
rect 5287 2034 5290 2035
rect 5322 2065 5325 2066
rect 5666 2065 5669 2066
rect 5322 2035 5452 2065
rect 5538 2035 5669 2065
rect 5322 2034 5325 2035
rect 5666 2034 5669 2035
rect 5701 2065 5704 2066
rect 6045 2065 6048 2066
rect 5701 2035 5831 2065
rect 5917 2035 6048 2065
rect 5701 2034 5704 2035
rect 6045 2034 6048 2035
rect 6080 2065 6083 2066
rect 6424 2065 6427 2066
rect 6080 2035 6210 2065
rect 6296 2035 6427 2065
rect 6080 2034 6083 2035
rect 6424 2034 6427 2035
rect 6459 2065 6462 2066
rect 6803 2065 6806 2066
rect 6459 2035 6589 2065
rect 6675 2035 6806 2065
rect 6459 2034 6462 2035
rect 6803 2034 6806 2035
rect 6838 2065 6841 2066
rect 7182 2065 7185 2066
rect 6838 2035 6968 2065
rect 7054 2035 7185 2065
rect 6838 2034 6841 2035
rect 7182 2034 7185 2035
rect 7217 2065 7220 2066
rect 7561 2065 7564 2066
rect 7217 2035 7347 2065
rect 7433 2035 7564 2065
rect 7217 2034 7220 2035
rect 7561 2034 7564 2035
rect 7596 2034 7599 2066
rect 161 2006 217 2009
rect 161 2005 166 2006
rect 53 1975 166 2005
rect 212 2005 217 2006
rect 540 2006 596 2009
rect 540 2005 545 2006
rect 212 1975 326 2005
rect 432 1975 545 2005
rect 591 2005 596 2006
rect 919 2006 975 2009
rect 919 2005 924 2006
rect 591 1975 705 2005
rect 811 1975 924 2005
rect 970 2005 975 2006
rect 1298 2006 1354 2009
rect 1298 2005 1303 2006
rect 970 1975 1084 2005
rect 1190 1975 1303 2005
rect 1349 2005 1354 2006
rect 1677 2006 1733 2009
rect 1677 2005 1682 2006
rect 1349 1975 1463 2005
rect 1569 1975 1682 2005
rect 1728 2005 1733 2006
rect 2056 2006 2112 2009
rect 2056 2005 2061 2006
rect 1728 1975 1842 2005
rect 1948 1975 2061 2005
rect 2107 2005 2112 2006
rect 2435 2006 2491 2009
rect 2435 2005 2440 2006
rect 2107 1975 2221 2005
rect 2327 1975 2440 2005
rect 2486 2005 2491 2006
rect 2814 2006 2870 2009
rect 2814 2005 2819 2006
rect 2486 1975 2600 2005
rect 2706 1975 2819 2005
rect 2865 2005 2870 2006
rect 3193 2006 3249 2009
rect 3193 2005 3198 2006
rect 2865 1975 2979 2005
rect 3085 1975 3198 2005
rect 3244 2005 3249 2006
rect 3572 2006 3628 2009
rect 3572 2005 3577 2006
rect 3244 1975 3358 2005
rect 3464 1975 3577 2005
rect 3623 2005 3628 2006
rect 3951 2006 4007 2009
rect 3951 2005 3956 2006
rect 3623 1975 3737 2005
rect 3843 1975 3956 2005
rect 4002 2005 4007 2006
rect 4330 2006 4386 2009
rect 4330 2005 4335 2006
rect 4002 1975 4116 2005
rect 4222 1975 4335 2005
rect 4381 2005 4386 2006
rect 4709 2006 4765 2009
rect 4709 2005 4714 2006
rect 4381 1975 4495 2005
rect 4601 1975 4714 2005
rect 4760 2005 4765 2006
rect 5088 2006 5144 2009
rect 5088 2005 5093 2006
rect 4760 1975 4874 2005
rect 4980 1975 5093 2005
rect 5139 2005 5144 2006
rect 5467 2006 5523 2009
rect 5467 2005 5472 2006
rect 5139 1975 5253 2005
rect 5359 1975 5472 2005
rect 5518 2005 5523 2006
rect 5846 2006 5902 2009
rect 5846 2005 5851 2006
rect 5518 1975 5632 2005
rect 5738 1975 5851 2005
rect 5897 2005 5902 2006
rect 6225 2006 6281 2009
rect 6225 2005 6230 2006
rect 5897 1975 6011 2005
rect 6117 1975 6230 2005
rect 6276 2005 6281 2006
rect 6604 2006 6660 2009
rect 6604 2005 6609 2006
rect 6276 1975 6390 2005
rect 6496 1975 6609 2005
rect 6655 2005 6660 2006
rect 6983 2006 7039 2009
rect 6983 2005 6988 2006
rect 6655 1975 6769 2005
rect 6875 1975 6988 2005
rect 7034 2005 7039 2006
rect 7362 2006 7418 2009
rect 7362 2005 7367 2006
rect 7034 1975 7148 2005
rect 7254 1975 7367 2005
rect 7413 2005 7418 2006
rect 7413 1975 7527 2005
rect 161 1971 217 1975
rect 540 1971 596 1975
rect 919 1971 975 1975
rect 1298 1971 1354 1975
rect 1677 1971 1733 1975
rect 2056 1971 2112 1975
rect 2435 1971 2491 1975
rect 2814 1971 2870 1975
rect 3193 1971 3249 1975
rect 3572 1971 3628 1975
rect 3951 1971 4007 1975
rect 4330 1971 4386 1975
rect 4709 1971 4765 1975
rect 5088 1971 5144 1975
rect 5467 1971 5523 1975
rect 5846 1971 5902 1975
rect 6225 1971 6281 1975
rect 6604 1971 6660 1975
rect 6983 1971 7039 1975
rect 7362 1971 7418 1975
rect -19 1914 -16 1946
rect 16 1945 19 1946
rect 360 1945 363 1946
rect 16 1915 146 1945
rect 232 1915 363 1945
rect 16 1914 19 1915
rect 360 1914 363 1915
rect 395 1945 398 1946
rect 739 1945 742 1946
rect 395 1915 525 1945
rect 611 1915 742 1945
rect 395 1914 398 1915
rect 739 1914 742 1915
rect 774 1945 777 1946
rect 1118 1945 1121 1946
rect 774 1915 904 1945
rect 990 1915 1121 1945
rect 774 1914 777 1915
rect 1118 1914 1121 1915
rect 1153 1945 1156 1946
rect 1497 1945 1500 1946
rect 1153 1915 1283 1945
rect 1369 1915 1500 1945
rect 1153 1914 1156 1915
rect 1497 1914 1500 1915
rect 1532 1945 1535 1946
rect 1876 1945 1879 1946
rect 1532 1915 1662 1945
rect 1748 1915 1879 1945
rect 1532 1914 1535 1915
rect 1876 1914 1879 1915
rect 1911 1945 1914 1946
rect 2255 1945 2258 1946
rect 1911 1915 2041 1945
rect 2127 1915 2258 1945
rect 1911 1914 1914 1915
rect 2255 1914 2258 1915
rect 2290 1945 2293 1946
rect 2634 1945 2637 1946
rect 2290 1915 2420 1945
rect 2506 1915 2637 1945
rect 2290 1914 2293 1915
rect 2634 1914 2637 1915
rect 2669 1945 2672 1946
rect 3013 1945 3016 1946
rect 2669 1915 2799 1945
rect 2885 1915 3016 1945
rect 2669 1914 2672 1915
rect 3013 1914 3016 1915
rect 3048 1945 3051 1946
rect 3392 1945 3395 1946
rect 3048 1915 3178 1945
rect 3264 1915 3395 1945
rect 3048 1914 3051 1915
rect 3392 1914 3395 1915
rect 3427 1945 3430 1946
rect 3771 1945 3774 1946
rect 3427 1915 3557 1945
rect 3643 1915 3774 1945
rect 3427 1914 3430 1915
rect 3771 1914 3774 1915
rect 3806 1945 3809 1946
rect 4150 1945 4153 1946
rect 3806 1915 3936 1945
rect 4022 1915 4153 1945
rect 3806 1914 3809 1915
rect 4150 1914 4153 1915
rect 4185 1945 4188 1946
rect 4529 1945 4532 1946
rect 4185 1915 4315 1945
rect 4401 1915 4532 1945
rect 4185 1914 4188 1915
rect 4529 1914 4532 1915
rect 4564 1945 4567 1946
rect 4908 1945 4911 1946
rect 4564 1915 4694 1945
rect 4780 1915 4911 1945
rect 4564 1914 4567 1915
rect 4908 1914 4911 1915
rect 4943 1945 4946 1946
rect 5287 1945 5290 1946
rect 4943 1915 5073 1945
rect 5159 1915 5290 1945
rect 4943 1914 4946 1915
rect 5287 1914 5290 1915
rect 5322 1945 5325 1946
rect 5666 1945 5669 1946
rect 5322 1915 5452 1945
rect 5538 1915 5669 1945
rect 5322 1914 5325 1915
rect 5666 1914 5669 1915
rect 5701 1945 5704 1946
rect 6045 1945 6048 1946
rect 5701 1915 5831 1945
rect 5917 1915 6048 1945
rect 5701 1914 5704 1915
rect 6045 1914 6048 1915
rect 6080 1945 6083 1946
rect 6424 1945 6427 1946
rect 6080 1915 6210 1945
rect 6296 1915 6427 1945
rect 6080 1914 6083 1915
rect 6424 1914 6427 1915
rect 6459 1945 6462 1946
rect 6803 1945 6806 1946
rect 6459 1915 6589 1945
rect 6675 1915 6806 1945
rect 6459 1914 6462 1915
rect 6803 1914 6806 1915
rect 6838 1945 6841 1946
rect 7182 1945 7185 1946
rect 6838 1915 6968 1945
rect 7054 1915 7185 1945
rect 6838 1914 6841 1915
rect 7182 1914 7185 1915
rect 7217 1945 7220 1946
rect 7561 1945 7564 1946
rect 7217 1915 7347 1945
rect 7433 1915 7564 1945
rect 7217 1914 7220 1915
rect 7561 1914 7564 1915
rect 7596 1914 7599 1946
rect 161 1886 217 1889
rect 161 1885 166 1886
rect 53 1855 166 1885
rect 212 1885 217 1886
rect 540 1886 596 1889
rect 540 1885 545 1886
rect 212 1855 326 1885
rect 432 1855 545 1885
rect 591 1885 596 1886
rect 919 1886 975 1889
rect 919 1885 924 1886
rect 591 1855 705 1885
rect 811 1855 924 1885
rect 970 1885 975 1886
rect 1298 1886 1354 1889
rect 1298 1885 1303 1886
rect 970 1855 1084 1885
rect 1190 1855 1303 1885
rect 1349 1885 1354 1886
rect 1677 1886 1733 1889
rect 1677 1885 1682 1886
rect 1349 1855 1463 1885
rect 1569 1855 1682 1885
rect 1728 1885 1733 1886
rect 2056 1886 2112 1889
rect 2056 1885 2061 1886
rect 1728 1855 1842 1885
rect 1948 1855 2061 1885
rect 2107 1885 2112 1886
rect 2435 1886 2491 1889
rect 2435 1885 2440 1886
rect 2107 1855 2221 1885
rect 2327 1855 2440 1885
rect 2486 1885 2491 1886
rect 2814 1886 2870 1889
rect 2814 1885 2819 1886
rect 2486 1855 2600 1885
rect 2706 1855 2819 1885
rect 2865 1885 2870 1886
rect 3193 1886 3249 1889
rect 3193 1885 3198 1886
rect 2865 1855 2979 1885
rect 3085 1855 3198 1885
rect 3244 1885 3249 1886
rect 3572 1886 3628 1889
rect 3572 1885 3577 1886
rect 3244 1855 3358 1885
rect 3464 1855 3577 1885
rect 3623 1885 3628 1886
rect 3951 1886 4007 1889
rect 3951 1885 3956 1886
rect 3623 1855 3737 1885
rect 3843 1855 3956 1885
rect 4002 1885 4007 1886
rect 4330 1886 4386 1889
rect 4330 1885 4335 1886
rect 4002 1855 4116 1885
rect 4222 1855 4335 1885
rect 4381 1885 4386 1886
rect 4709 1886 4765 1889
rect 4709 1885 4714 1886
rect 4381 1855 4495 1885
rect 4601 1855 4714 1885
rect 4760 1885 4765 1886
rect 5088 1886 5144 1889
rect 5088 1885 5093 1886
rect 4760 1855 4874 1885
rect 4980 1855 5093 1885
rect 5139 1885 5144 1886
rect 5467 1886 5523 1889
rect 5467 1885 5472 1886
rect 5139 1855 5253 1885
rect 5359 1855 5472 1885
rect 5518 1885 5523 1886
rect 5846 1886 5902 1889
rect 5846 1885 5851 1886
rect 5518 1855 5632 1885
rect 5738 1855 5851 1885
rect 5897 1885 5902 1886
rect 6225 1886 6281 1889
rect 6225 1885 6230 1886
rect 5897 1855 6011 1885
rect 6117 1855 6230 1885
rect 6276 1885 6281 1886
rect 6604 1886 6660 1889
rect 6604 1885 6609 1886
rect 6276 1855 6390 1885
rect 6496 1855 6609 1885
rect 6655 1885 6660 1886
rect 6983 1886 7039 1889
rect 6983 1885 6988 1886
rect 6655 1855 6769 1885
rect 6875 1855 6988 1885
rect 7034 1885 7039 1886
rect 7362 1886 7418 1889
rect 7362 1885 7367 1886
rect 7034 1855 7148 1885
rect 7254 1855 7367 1885
rect 7413 1885 7418 1886
rect 7413 1855 7527 1885
rect 161 1851 217 1855
rect 540 1851 596 1855
rect 919 1851 975 1855
rect 1298 1851 1354 1855
rect 1677 1851 1733 1855
rect 2056 1851 2112 1855
rect 2435 1851 2491 1855
rect 2814 1851 2870 1855
rect 3193 1851 3249 1855
rect 3572 1851 3628 1855
rect 3951 1851 4007 1855
rect 4330 1851 4386 1855
rect 4709 1851 4765 1855
rect 5088 1851 5144 1855
rect 5467 1851 5523 1855
rect 5846 1851 5902 1855
rect 6225 1851 6281 1855
rect 6604 1851 6660 1855
rect 6983 1851 7039 1855
rect 7362 1851 7418 1855
rect 161 1764 217 1767
rect 161 1763 166 1764
rect 53 1733 166 1763
rect 212 1763 217 1764
rect 540 1764 596 1767
rect 540 1763 545 1764
rect 212 1733 326 1763
rect 432 1733 545 1763
rect 591 1763 596 1764
rect 919 1764 975 1767
rect 919 1763 924 1764
rect 591 1733 705 1763
rect 811 1733 924 1763
rect 970 1763 975 1764
rect 1298 1764 1354 1767
rect 1298 1763 1303 1764
rect 970 1733 1084 1763
rect 1190 1733 1303 1763
rect 1349 1763 1354 1764
rect 1677 1764 1733 1767
rect 1677 1763 1682 1764
rect 1349 1733 1463 1763
rect 1569 1733 1682 1763
rect 1728 1763 1733 1764
rect 2056 1764 2112 1767
rect 2056 1763 2061 1764
rect 1728 1733 1842 1763
rect 1948 1733 2061 1763
rect 2107 1763 2112 1764
rect 2435 1764 2491 1767
rect 2435 1763 2440 1764
rect 2107 1733 2221 1763
rect 2327 1733 2440 1763
rect 2486 1763 2491 1764
rect 2814 1764 2870 1767
rect 2814 1763 2819 1764
rect 2486 1733 2600 1763
rect 2706 1733 2819 1763
rect 2865 1763 2870 1764
rect 3193 1764 3249 1767
rect 3193 1763 3198 1764
rect 2865 1733 2979 1763
rect 3085 1733 3198 1763
rect 3244 1763 3249 1764
rect 3572 1764 3628 1767
rect 3572 1763 3577 1764
rect 3244 1733 3358 1763
rect 3464 1733 3577 1763
rect 3623 1763 3628 1764
rect 3951 1764 4007 1767
rect 3951 1763 3956 1764
rect 3623 1733 3737 1763
rect 3843 1733 3956 1763
rect 4002 1763 4007 1764
rect 4330 1764 4386 1767
rect 4330 1763 4335 1764
rect 4002 1733 4116 1763
rect 4222 1733 4335 1763
rect 4381 1763 4386 1764
rect 4709 1764 4765 1767
rect 4709 1763 4714 1764
rect 4381 1733 4495 1763
rect 4601 1733 4714 1763
rect 4760 1763 4765 1764
rect 5088 1764 5144 1767
rect 5088 1763 5093 1764
rect 4760 1733 4874 1763
rect 4980 1733 5093 1763
rect 5139 1763 5144 1764
rect 5467 1764 5523 1767
rect 5467 1763 5472 1764
rect 5139 1733 5253 1763
rect 5359 1733 5472 1763
rect 5518 1763 5523 1764
rect 5846 1764 5902 1767
rect 5846 1763 5851 1764
rect 5518 1733 5632 1763
rect 5738 1733 5851 1763
rect 5897 1763 5902 1764
rect 6225 1764 6281 1767
rect 6225 1763 6230 1764
rect 5897 1733 6011 1763
rect 6117 1733 6230 1763
rect 6276 1763 6281 1764
rect 6604 1764 6660 1767
rect 6604 1763 6609 1764
rect 6276 1733 6390 1763
rect 6496 1733 6609 1763
rect 6655 1763 6660 1764
rect 6983 1764 7039 1767
rect 6983 1763 6988 1764
rect 6655 1733 6769 1763
rect 6875 1733 6988 1763
rect 7034 1763 7039 1764
rect 7362 1764 7418 1767
rect 7362 1763 7367 1764
rect 7034 1733 7148 1763
rect 7254 1733 7367 1763
rect 7413 1763 7418 1764
rect 7413 1733 7527 1763
rect 161 1729 217 1733
rect 540 1729 596 1733
rect 919 1729 975 1733
rect 1298 1729 1354 1733
rect 1677 1729 1733 1733
rect 2056 1729 2112 1733
rect 2435 1729 2491 1733
rect 2814 1729 2870 1733
rect 3193 1729 3249 1733
rect 3572 1729 3628 1733
rect 3951 1729 4007 1733
rect 4330 1729 4386 1733
rect 4709 1729 4765 1733
rect 5088 1729 5144 1733
rect 5467 1729 5523 1733
rect 5846 1729 5902 1733
rect 6225 1729 6281 1733
rect 6604 1729 6660 1733
rect 6983 1729 7039 1733
rect 7362 1729 7418 1733
rect -19 1671 -16 1703
rect 16 1702 19 1703
rect 360 1702 363 1703
rect 16 1672 146 1702
rect 232 1672 363 1702
rect 16 1671 19 1672
rect 360 1671 363 1672
rect 395 1702 398 1703
rect 739 1702 742 1703
rect 395 1672 525 1702
rect 611 1672 742 1702
rect 395 1671 398 1672
rect 739 1671 742 1672
rect 774 1702 777 1703
rect 1118 1702 1121 1703
rect 774 1672 904 1702
rect 990 1672 1121 1702
rect 774 1671 777 1672
rect 1118 1671 1121 1672
rect 1153 1702 1156 1703
rect 1497 1702 1500 1703
rect 1153 1672 1283 1702
rect 1369 1672 1500 1702
rect 1153 1671 1156 1672
rect 1497 1671 1500 1672
rect 1532 1702 1535 1703
rect 1876 1702 1879 1703
rect 1532 1672 1662 1702
rect 1748 1672 1879 1702
rect 1532 1671 1535 1672
rect 1876 1671 1879 1672
rect 1911 1702 1914 1703
rect 2255 1702 2258 1703
rect 1911 1672 2041 1702
rect 2127 1672 2258 1702
rect 1911 1671 1914 1672
rect 2255 1671 2258 1672
rect 2290 1702 2293 1703
rect 2634 1702 2637 1703
rect 2290 1672 2420 1702
rect 2506 1672 2637 1702
rect 2290 1671 2293 1672
rect 2634 1671 2637 1672
rect 2669 1702 2672 1703
rect 3013 1702 3016 1703
rect 2669 1672 2799 1702
rect 2885 1672 3016 1702
rect 2669 1671 2672 1672
rect 3013 1671 3016 1672
rect 3048 1702 3051 1703
rect 3392 1702 3395 1703
rect 3048 1672 3178 1702
rect 3264 1672 3395 1702
rect 3048 1671 3051 1672
rect 3392 1671 3395 1672
rect 3427 1702 3430 1703
rect 3771 1702 3774 1703
rect 3427 1672 3557 1702
rect 3643 1672 3774 1702
rect 3427 1671 3430 1672
rect 3771 1671 3774 1672
rect 3806 1702 3809 1703
rect 4150 1702 4153 1703
rect 3806 1672 3936 1702
rect 4022 1672 4153 1702
rect 3806 1671 3809 1672
rect 4150 1671 4153 1672
rect 4185 1702 4188 1703
rect 4529 1702 4532 1703
rect 4185 1672 4315 1702
rect 4401 1672 4532 1702
rect 4185 1671 4188 1672
rect 4529 1671 4532 1672
rect 4564 1702 4567 1703
rect 4908 1702 4911 1703
rect 4564 1672 4694 1702
rect 4780 1672 4911 1702
rect 4564 1671 4567 1672
rect 4908 1671 4911 1672
rect 4943 1702 4946 1703
rect 5287 1702 5290 1703
rect 4943 1672 5073 1702
rect 5159 1672 5290 1702
rect 4943 1671 4946 1672
rect 5287 1671 5290 1672
rect 5322 1702 5325 1703
rect 5666 1702 5669 1703
rect 5322 1672 5452 1702
rect 5538 1672 5669 1702
rect 5322 1671 5325 1672
rect 5666 1671 5669 1672
rect 5701 1702 5704 1703
rect 6045 1702 6048 1703
rect 5701 1672 5831 1702
rect 5917 1672 6048 1702
rect 5701 1671 5704 1672
rect 6045 1671 6048 1672
rect 6080 1702 6083 1703
rect 6424 1702 6427 1703
rect 6080 1672 6210 1702
rect 6296 1672 6427 1702
rect 6080 1671 6083 1672
rect 6424 1671 6427 1672
rect 6459 1702 6462 1703
rect 6803 1702 6806 1703
rect 6459 1672 6589 1702
rect 6675 1672 6806 1702
rect 6459 1671 6462 1672
rect 6803 1671 6806 1672
rect 6838 1702 6841 1703
rect 7182 1702 7185 1703
rect 6838 1672 6968 1702
rect 7054 1672 7185 1702
rect 6838 1671 6841 1672
rect 7182 1671 7185 1672
rect 7217 1702 7220 1703
rect 7561 1702 7564 1703
rect 7217 1672 7347 1702
rect 7433 1672 7564 1702
rect 7217 1671 7220 1672
rect 7561 1671 7564 1672
rect 7596 1671 7599 1703
rect 161 1643 217 1646
rect 161 1642 166 1643
rect 53 1612 166 1642
rect 212 1642 217 1643
rect 540 1643 596 1646
rect 540 1642 545 1643
rect 212 1612 326 1642
rect 432 1612 545 1642
rect 591 1642 596 1643
rect 919 1643 975 1646
rect 919 1642 924 1643
rect 591 1612 705 1642
rect 811 1612 924 1642
rect 970 1642 975 1643
rect 1298 1643 1354 1646
rect 1298 1642 1303 1643
rect 970 1612 1084 1642
rect 1190 1612 1303 1642
rect 1349 1642 1354 1643
rect 1677 1643 1733 1646
rect 1677 1642 1682 1643
rect 1349 1612 1463 1642
rect 1569 1612 1682 1642
rect 1728 1642 1733 1643
rect 2056 1643 2112 1646
rect 2056 1642 2061 1643
rect 1728 1612 1842 1642
rect 1948 1612 2061 1642
rect 2107 1642 2112 1643
rect 2435 1643 2491 1646
rect 2435 1642 2440 1643
rect 2107 1612 2221 1642
rect 2327 1612 2440 1642
rect 2486 1642 2491 1643
rect 2814 1643 2870 1646
rect 2814 1642 2819 1643
rect 2486 1612 2600 1642
rect 2706 1612 2819 1642
rect 2865 1642 2870 1643
rect 3193 1643 3249 1646
rect 3193 1642 3198 1643
rect 2865 1612 2979 1642
rect 3085 1612 3198 1642
rect 3244 1642 3249 1643
rect 3572 1643 3628 1646
rect 3572 1642 3577 1643
rect 3244 1612 3358 1642
rect 3464 1612 3577 1642
rect 3623 1642 3628 1643
rect 3951 1643 4007 1646
rect 3951 1642 3956 1643
rect 3623 1612 3737 1642
rect 3843 1612 3956 1642
rect 4002 1642 4007 1643
rect 4330 1643 4386 1646
rect 4330 1642 4335 1643
rect 4002 1612 4116 1642
rect 4222 1612 4335 1642
rect 4381 1642 4386 1643
rect 4709 1643 4765 1646
rect 4709 1642 4714 1643
rect 4381 1612 4495 1642
rect 4601 1612 4714 1642
rect 4760 1642 4765 1643
rect 5088 1643 5144 1646
rect 5088 1642 5093 1643
rect 4760 1612 4874 1642
rect 4980 1612 5093 1642
rect 5139 1642 5144 1643
rect 5467 1643 5523 1646
rect 5467 1642 5472 1643
rect 5139 1612 5253 1642
rect 5359 1612 5472 1642
rect 5518 1642 5523 1643
rect 5846 1643 5902 1646
rect 5846 1642 5851 1643
rect 5518 1612 5632 1642
rect 5738 1612 5851 1642
rect 5897 1642 5902 1643
rect 6225 1643 6281 1646
rect 6225 1642 6230 1643
rect 5897 1612 6011 1642
rect 6117 1612 6230 1642
rect 6276 1642 6281 1643
rect 6604 1643 6660 1646
rect 6604 1642 6609 1643
rect 6276 1612 6390 1642
rect 6496 1612 6609 1642
rect 6655 1642 6660 1643
rect 6983 1643 7039 1646
rect 6983 1642 6988 1643
rect 6655 1612 6769 1642
rect 6875 1612 6988 1642
rect 7034 1642 7039 1643
rect 7362 1643 7418 1646
rect 7362 1642 7367 1643
rect 7034 1612 7148 1642
rect 7254 1612 7367 1642
rect 7413 1642 7418 1643
rect 7413 1612 7527 1642
rect 161 1608 217 1612
rect 540 1608 596 1612
rect 919 1608 975 1612
rect 1298 1608 1354 1612
rect 1677 1608 1733 1612
rect 2056 1608 2112 1612
rect 2435 1608 2491 1612
rect 2814 1608 2870 1612
rect 3193 1608 3249 1612
rect 3572 1608 3628 1612
rect 3951 1608 4007 1612
rect 4330 1608 4386 1612
rect 4709 1608 4765 1612
rect 5088 1608 5144 1612
rect 5467 1608 5523 1612
rect 5846 1608 5902 1612
rect 6225 1608 6281 1612
rect 6604 1608 6660 1612
rect 6983 1608 7039 1612
rect 7362 1608 7418 1612
rect -19 1551 -16 1583
rect 16 1582 19 1583
rect 360 1582 363 1583
rect 16 1552 146 1582
rect 232 1552 363 1582
rect 16 1551 19 1552
rect 360 1551 363 1552
rect 395 1582 398 1583
rect 739 1582 742 1583
rect 395 1552 525 1582
rect 611 1552 742 1582
rect 395 1551 398 1552
rect 739 1551 742 1552
rect 774 1582 777 1583
rect 1118 1582 1121 1583
rect 774 1552 904 1582
rect 990 1552 1121 1582
rect 774 1551 777 1552
rect 1118 1551 1121 1552
rect 1153 1582 1156 1583
rect 1497 1582 1500 1583
rect 1153 1552 1283 1582
rect 1369 1552 1500 1582
rect 1153 1551 1156 1552
rect 1497 1551 1500 1552
rect 1532 1582 1535 1583
rect 1876 1582 1879 1583
rect 1532 1552 1662 1582
rect 1748 1552 1879 1582
rect 1532 1551 1535 1552
rect 1876 1551 1879 1552
rect 1911 1582 1914 1583
rect 2255 1582 2258 1583
rect 1911 1552 2041 1582
rect 2127 1552 2258 1582
rect 1911 1551 1914 1552
rect 2255 1551 2258 1552
rect 2290 1582 2293 1583
rect 2634 1582 2637 1583
rect 2290 1552 2420 1582
rect 2506 1552 2637 1582
rect 2290 1551 2293 1552
rect 2634 1551 2637 1552
rect 2669 1582 2672 1583
rect 3013 1582 3016 1583
rect 2669 1552 2799 1582
rect 2885 1552 3016 1582
rect 2669 1551 2672 1552
rect 3013 1551 3016 1552
rect 3048 1582 3051 1583
rect 3392 1582 3395 1583
rect 3048 1552 3178 1582
rect 3264 1552 3395 1582
rect 3048 1551 3051 1552
rect 3392 1551 3395 1552
rect 3427 1582 3430 1583
rect 3771 1582 3774 1583
rect 3427 1552 3557 1582
rect 3643 1552 3774 1582
rect 3427 1551 3430 1552
rect 3771 1551 3774 1552
rect 3806 1582 3809 1583
rect 4150 1582 4153 1583
rect 3806 1552 3936 1582
rect 4022 1552 4153 1582
rect 3806 1551 3809 1552
rect 4150 1551 4153 1552
rect 4185 1582 4188 1583
rect 4529 1582 4532 1583
rect 4185 1552 4315 1582
rect 4401 1552 4532 1582
rect 4185 1551 4188 1552
rect 4529 1551 4532 1552
rect 4564 1582 4567 1583
rect 4908 1582 4911 1583
rect 4564 1552 4694 1582
rect 4780 1552 4911 1582
rect 4564 1551 4567 1552
rect 4908 1551 4911 1552
rect 4943 1582 4946 1583
rect 5287 1582 5290 1583
rect 4943 1552 5073 1582
rect 5159 1552 5290 1582
rect 4943 1551 4946 1552
rect 5287 1551 5290 1552
rect 5322 1582 5325 1583
rect 5666 1582 5669 1583
rect 5322 1552 5452 1582
rect 5538 1552 5669 1582
rect 5322 1551 5325 1552
rect 5666 1551 5669 1552
rect 5701 1582 5704 1583
rect 6045 1582 6048 1583
rect 5701 1552 5831 1582
rect 5917 1552 6048 1582
rect 5701 1551 5704 1552
rect 6045 1551 6048 1552
rect 6080 1582 6083 1583
rect 6424 1582 6427 1583
rect 6080 1552 6210 1582
rect 6296 1552 6427 1582
rect 6080 1551 6083 1552
rect 6424 1551 6427 1552
rect 6459 1582 6462 1583
rect 6803 1582 6806 1583
rect 6459 1552 6589 1582
rect 6675 1552 6806 1582
rect 6459 1551 6462 1552
rect 6803 1551 6806 1552
rect 6838 1582 6841 1583
rect 7182 1582 7185 1583
rect 6838 1552 6968 1582
rect 7054 1552 7185 1582
rect 6838 1551 6841 1552
rect 7182 1551 7185 1552
rect 7217 1582 7220 1583
rect 7561 1582 7564 1583
rect 7217 1552 7347 1582
rect 7433 1552 7564 1582
rect 7217 1551 7220 1552
rect 7561 1551 7564 1552
rect 7596 1551 7599 1583
rect 161 1523 217 1526
rect 161 1522 166 1523
rect 53 1492 166 1522
rect 212 1522 217 1523
rect 540 1523 596 1526
rect 540 1522 545 1523
rect 212 1492 326 1522
rect 432 1492 545 1522
rect 591 1522 596 1523
rect 919 1523 975 1526
rect 919 1522 924 1523
rect 591 1492 705 1522
rect 811 1492 924 1522
rect 970 1522 975 1523
rect 1298 1523 1354 1526
rect 1298 1522 1303 1523
rect 970 1492 1084 1522
rect 1190 1492 1303 1522
rect 1349 1522 1354 1523
rect 1677 1523 1733 1526
rect 1677 1522 1682 1523
rect 1349 1492 1463 1522
rect 1569 1492 1682 1522
rect 1728 1522 1733 1523
rect 2056 1523 2112 1526
rect 2056 1522 2061 1523
rect 1728 1492 1842 1522
rect 1948 1492 2061 1522
rect 2107 1522 2112 1523
rect 2435 1523 2491 1526
rect 2435 1522 2440 1523
rect 2107 1492 2221 1522
rect 2327 1492 2440 1522
rect 2486 1522 2491 1523
rect 2814 1523 2870 1526
rect 2814 1522 2819 1523
rect 2486 1492 2600 1522
rect 2706 1492 2819 1522
rect 2865 1522 2870 1523
rect 3193 1523 3249 1526
rect 3193 1522 3198 1523
rect 2865 1492 2979 1522
rect 3085 1492 3198 1522
rect 3244 1522 3249 1523
rect 3572 1523 3628 1526
rect 3572 1522 3577 1523
rect 3244 1492 3358 1522
rect 3464 1492 3577 1522
rect 3623 1522 3628 1523
rect 3951 1523 4007 1526
rect 3951 1522 3956 1523
rect 3623 1492 3737 1522
rect 3843 1492 3956 1522
rect 4002 1522 4007 1523
rect 4330 1523 4386 1526
rect 4330 1522 4335 1523
rect 4002 1492 4116 1522
rect 4222 1492 4335 1522
rect 4381 1522 4386 1523
rect 4709 1523 4765 1526
rect 4709 1522 4714 1523
rect 4381 1492 4495 1522
rect 4601 1492 4714 1522
rect 4760 1522 4765 1523
rect 5088 1523 5144 1526
rect 5088 1522 5093 1523
rect 4760 1492 4874 1522
rect 4980 1492 5093 1522
rect 5139 1522 5144 1523
rect 5467 1523 5523 1526
rect 5467 1522 5472 1523
rect 5139 1492 5253 1522
rect 5359 1492 5472 1522
rect 5518 1522 5523 1523
rect 5846 1523 5902 1526
rect 5846 1522 5851 1523
rect 5518 1492 5632 1522
rect 5738 1492 5851 1522
rect 5897 1522 5902 1523
rect 6225 1523 6281 1526
rect 6225 1522 6230 1523
rect 5897 1492 6011 1522
rect 6117 1492 6230 1522
rect 6276 1522 6281 1523
rect 6604 1523 6660 1526
rect 6604 1522 6609 1523
rect 6276 1492 6390 1522
rect 6496 1492 6609 1522
rect 6655 1522 6660 1523
rect 6983 1523 7039 1526
rect 6983 1522 6988 1523
rect 6655 1492 6769 1522
rect 6875 1492 6988 1522
rect 7034 1522 7039 1523
rect 7362 1523 7418 1526
rect 7362 1522 7367 1523
rect 7034 1492 7148 1522
rect 7254 1492 7367 1522
rect 7413 1522 7418 1523
rect 7413 1492 7527 1522
rect 161 1488 217 1492
rect 540 1488 596 1492
rect 919 1488 975 1492
rect 1298 1488 1354 1492
rect 1677 1488 1733 1492
rect 2056 1488 2112 1492
rect 2435 1488 2491 1492
rect 2814 1488 2870 1492
rect 3193 1488 3249 1492
rect 3572 1488 3628 1492
rect 3951 1488 4007 1492
rect 4330 1488 4386 1492
rect 4709 1488 4765 1492
rect 5088 1488 5144 1492
rect 5467 1488 5523 1492
rect 5846 1488 5902 1492
rect 6225 1488 6281 1492
rect 6604 1488 6660 1492
rect 6983 1488 7039 1492
rect 7362 1488 7418 1492
rect -19 1431 -16 1463
rect 16 1462 19 1463
rect 360 1462 363 1463
rect 16 1432 146 1462
rect 232 1432 363 1462
rect 16 1431 19 1432
rect 360 1431 363 1432
rect 395 1462 398 1463
rect 739 1462 742 1463
rect 395 1432 525 1462
rect 611 1432 742 1462
rect 395 1431 398 1432
rect 739 1431 742 1432
rect 774 1462 777 1463
rect 1118 1462 1121 1463
rect 774 1432 904 1462
rect 990 1432 1121 1462
rect 774 1431 777 1432
rect 1118 1431 1121 1432
rect 1153 1462 1156 1463
rect 1497 1462 1500 1463
rect 1153 1432 1283 1462
rect 1369 1432 1500 1462
rect 1153 1431 1156 1432
rect 1497 1431 1500 1432
rect 1532 1462 1535 1463
rect 1876 1462 1879 1463
rect 1532 1432 1662 1462
rect 1748 1432 1879 1462
rect 1532 1431 1535 1432
rect 1876 1431 1879 1432
rect 1911 1462 1914 1463
rect 2255 1462 2258 1463
rect 1911 1432 2041 1462
rect 2127 1432 2258 1462
rect 1911 1431 1914 1432
rect 2255 1431 2258 1432
rect 2290 1462 2293 1463
rect 2634 1462 2637 1463
rect 2290 1432 2420 1462
rect 2506 1432 2637 1462
rect 2290 1431 2293 1432
rect 2634 1431 2637 1432
rect 2669 1462 2672 1463
rect 3013 1462 3016 1463
rect 2669 1432 2799 1462
rect 2885 1432 3016 1462
rect 2669 1431 2672 1432
rect 3013 1431 3016 1432
rect 3048 1462 3051 1463
rect 3392 1462 3395 1463
rect 3048 1432 3178 1462
rect 3264 1432 3395 1462
rect 3048 1431 3051 1432
rect 3392 1431 3395 1432
rect 3427 1462 3430 1463
rect 3771 1462 3774 1463
rect 3427 1432 3557 1462
rect 3643 1432 3774 1462
rect 3427 1431 3430 1432
rect 3771 1431 3774 1432
rect 3806 1462 3809 1463
rect 4150 1462 4153 1463
rect 3806 1432 3936 1462
rect 4022 1432 4153 1462
rect 3806 1431 3809 1432
rect 4150 1431 4153 1432
rect 4185 1462 4188 1463
rect 4529 1462 4532 1463
rect 4185 1432 4315 1462
rect 4401 1432 4532 1462
rect 4185 1431 4188 1432
rect 4529 1431 4532 1432
rect 4564 1462 4567 1463
rect 4908 1462 4911 1463
rect 4564 1432 4694 1462
rect 4780 1432 4911 1462
rect 4564 1431 4567 1432
rect 4908 1431 4911 1432
rect 4943 1462 4946 1463
rect 5287 1462 5290 1463
rect 4943 1432 5073 1462
rect 5159 1432 5290 1462
rect 4943 1431 4946 1432
rect 5287 1431 5290 1432
rect 5322 1462 5325 1463
rect 5666 1462 5669 1463
rect 5322 1432 5452 1462
rect 5538 1432 5669 1462
rect 5322 1431 5325 1432
rect 5666 1431 5669 1432
rect 5701 1462 5704 1463
rect 6045 1462 6048 1463
rect 5701 1432 5831 1462
rect 5917 1432 6048 1462
rect 5701 1431 5704 1432
rect 6045 1431 6048 1432
rect 6080 1462 6083 1463
rect 6424 1462 6427 1463
rect 6080 1432 6210 1462
rect 6296 1432 6427 1462
rect 6080 1431 6083 1432
rect 6424 1431 6427 1432
rect 6459 1462 6462 1463
rect 6803 1462 6806 1463
rect 6459 1432 6589 1462
rect 6675 1432 6806 1462
rect 6459 1431 6462 1432
rect 6803 1431 6806 1432
rect 6838 1462 6841 1463
rect 7182 1462 7185 1463
rect 6838 1432 6968 1462
rect 7054 1432 7185 1462
rect 6838 1431 6841 1432
rect 7182 1431 7185 1432
rect 7217 1462 7220 1463
rect 7561 1462 7564 1463
rect 7217 1432 7347 1462
rect 7433 1432 7564 1462
rect 7217 1431 7220 1432
rect 7561 1431 7564 1432
rect 7596 1431 7599 1463
rect 161 1403 217 1406
rect 161 1402 166 1403
rect 53 1372 166 1402
rect 212 1402 217 1403
rect 540 1403 596 1406
rect 540 1402 545 1403
rect 212 1372 326 1402
rect 432 1372 545 1402
rect 591 1402 596 1403
rect 919 1403 975 1406
rect 919 1402 924 1403
rect 591 1372 705 1402
rect 811 1372 924 1402
rect 970 1402 975 1403
rect 1298 1403 1354 1406
rect 1298 1402 1303 1403
rect 970 1372 1084 1402
rect 1190 1372 1303 1402
rect 1349 1402 1354 1403
rect 1677 1403 1733 1406
rect 1677 1402 1682 1403
rect 1349 1372 1463 1402
rect 1569 1372 1682 1402
rect 1728 1402 1733 1403
rect 2056 1403 2112 1406
rect 2056 1402 2061 1403
rect 1728 1372 1842 1402
rect 1948 1372 2061 1402
rect 2107 1402 2112 1403
rect 2435 1403 2491 1406
rect 2435 1402 2440 1403
rect 2107 1372 2221 1402
rect 2327 1372 2440 1402
rect 2486 1402 2491 1403
rect 2814 1403 2870 1406
rect 2814 1402 2819 1403
rect 2486 1372 2600 1402
rect 2706 1372 2819 1402
rect 2865 1402 2870 1403
rect 3193 1403 3249 1406
rect 3193 1402 3198 1403
rect 2865 1372 2979 1402
rect 3085 1372 3198 1402
rect 3244 1402 3249 1403
rect 3572 1403 3628 1406
rect 3572 1402 3577 1403
rect 3244 1372 3358 1402
rect 3464 1372 3577 1402
rect 3623 1402 3628 1403
rect 3951 1403 4007 1406
rect 3951 1402 3956 1403
rect 3623 1372 3737 1402
rect 3843 1372 3956 1402
rect 4002 1402 4007 1403
rect 4330 1403 4386 1406
rect 4330 1402 4335 1403
rect 4002 1372 4116 1402
rect 4222 1372 4335 1402
rect 4381 1402 4386 1403
rect 4709 1403 4765 1406
rect 4709 1402 4714 1403
rect 4381 1372 4495 1402
rect 4601 1372 4714 1402
rect 4760 1402 4765 1403
rect 5088 1403 5144 1406
rect 5088 1402 5093 1403
rect 4760 1372 4874 1402
rect 4980 1372 5093 1402
rect 5139 1402 5144 1403
rect 5467 1403 5523 1406
rect 5467 1402 5472 1403
rect 5139 1372 5253 1402
rect 5359 1372 5472 1402
rect 5518 1402 5523 1403
rect 5846 1403 5902 1406
rect 5846 1402 5851 1403
rect 5518 1372 5632 1402
rect 5738 1372 5851 1402
rect 5897 1402 5902 1403
rect 6225 1403 6281 1406
rect 6225 1402 6230 1403
rect 5897 1372 6011 1402
rect 6117 1372 6230 1402
rect 6276 1402 6281 1403
rect 6604 1403 6660 1406
rect 6604 1402 6609 1403
rect 6276 1372 6390 1402
rect 6496 1372 6609 1402
rect 6655 1402 6660 1403
rect 6983 1403 7039 1406
rect 6983 1402 6988 1403
rect 6655 1372 6769 1402
rect 6875 1372 6988 1402
rect 7034 1402 7039 1403
rect 7362 1403 7418 1406
rect 7362 1402 7367 1403
rect 7034 1372 7148 1402
rect 7254 1372 7367 1402
rect 7413 1402 7418 1403
rect 7413 1372 7527 1402
rect 161 1368 217 1372
rect 540 1368 596 1372
rect 919 1368 975 1372
rect 1298 1368 1354 1372
rect 1677 1368 1733 1372
rect 2056 1368 2112 1372
rect 2435 1368 2491 1372
rect 2814 1368 2870 1372
rect 3193 1368 3249 1372
rect 3572 1368 3628 1372
rect 3951 1368 4007 1372
rect 4330 1368 4386 1372
rect 4709 1368 4765 1372
rect 5088 1368 5144 1372
rect 5467 1368 5523 1372
rect 5846 1368 5902 1372
rect 6225 1368 6281 1372
rect 6604 1368 6660 1372
rect 6983 1368 7039 1372
rect 7362 1368 7418 1372
rect -19 1311 -16 1343
rect 16 1342 19 1343
rect 360 1342 363 1343
rect 16 1312 146 1342
rect 232 1312 363 1342
rect 16 1311 19 1312
rect 360 1311 363 1312
rect 395 1342 398 1343
rect 739 1342 742 1343
rect 395 1312 525 1342
rect 611 1312 742 1342
rect 395 1311 398 1312
rect 739 1311 742 1312
rect 774 1342 777 1343
rect 1118 1342 1121 1343
rect 774 1312 904 1342
rect 990 1312 1121 1342
rect 774 1311 777 1312
rect 1118 1311 1121 1312
rect 1153 1342 1156 1343
rect 1497 1342 1500 1343
rect 1153 1312 1283 1342
rect 1369 1312 1500 1342
rect 1153 1311 1156 1312
rect 1497 1311 1500 1312
rect 1532 1342 1535 1343
rect 1876 1342 1879 1343
rect 1532 1312 1662 1342
rect 1748 1312 1879 1342
rect 1532 1311 1535 1312
rect 1876 1311 1879 1312
rect 1911 1342 1914 1343
rect 2255 1342 2258 1343
rect 1911 1312 2041 1342
rect 2127 1312 2258 1342
rect 1911 1311 1914 1312
rect 2255 1311 2258 1312
rect 2290 1342 2293 1343
rect 2634 1342 2637 1343
rect 2290 1312 2420 1342
rect 2506 1312 2637 1342
rect 2290 1311 2293 1312
rect 2634 1311 2637 1312
rect 2669 1342 2672 1343
rect 3013 1342 3016 1343
rect 2669 1312 2799 1342
rect 2885 1312 3016 1342
rect 2669 1311 2672 1312
rect 3013 1311 3016 1312
rect 3048 1342 3051 1343
rect 3392 1342 3395 1343
rect 3048 1312 3178 1342
rect 3264 1312 3395 1342
rect 3048 1311 3051 1312
rect 3392 1311 3395 1312
rect 3427 1342 3430 1343
rect 3771 1342 3774 1343
rect 3427 1312 3557 1342
rect 3643 1312 3774 1342
rect 3427 1311 3430 1312
rect 3771 1311 3774 1312
rect 3806 1342 3809 1343
rect 4150 1342 4153 1343
rect 3806 1312 3936 1342
rect 4022 1312 4153 1342
rect 3806 1311 3809 1312
rect 4150 1311 4153 1312
rect 4185 1342 4188 1343
rect 4529 1342 4532 1343
rect 4185 1312 4315 1342
rect 4401 1312 4532 1342
rect 4185 1311 4188 1312
rect 4529 1311 4532 1312
rect 4564 1342 4567 1343
rect 4908 1342 4911 1343
rect 4564 1312 4694 1342
rect 4780 1312 4911 1342
rect 4564 1311 4567 1312
rect 4908 1311 4911 1312
rect 4943 1342 4946 1343
rect 5287 1342 5290 1343
rect 4943 1312 5073 1342
rect 5159 1312 5290 1342
rect 4943 1311 4946 1312
rect 5287 1311 5290 1312
rect 5322 1342 5325 1343
rect 5666 1342 5669 1343
rect 5322 1312 5452 1342
rect 5538 1312 5669 1342
rect 5322 1311 5325 1312
rect 5666 1311 5669 1312
rect 5701 1342 5704 1343
rect 6045 1342 6048 1343
rect 5701 1312 5831 1342
rect 5917 1312 6048 1342
rect 5701 1311 5704 1312
rect 6045 1311 6048 1312
rect 6080 1342 6083 1343
rect 6424 1342 6427 1343
rect 6080 1312 6210 1342
rect 6296 1312 6427 1342
rect 6080 1311 6083 1312
rect 6424 1311 6427 1312
rect 6459 1342 6462 1343
rect 6803 1342 6806 1343
rect 6459 1312 6589 1342
rect 6675 1312 6806 1342
rect 6459 1311 6462 1312
rect 6803 1311 6806 1312
rect 6838 1342 6841 1343
rect 7182 1342 7185 1343
rect 6838 1312 6968 1342
rect 7054 1312 7185 1342
rect 6838 1311 6841 1312
rect 7182 1311 7185 1312
rect 7217 1342 7220 1343
rect 7561 1342 7564 1343
rect 7217 1312 7347 1342
rect 7433 1312 7564 1342
rect 7217 1311 7220 1312
rect 7561 1311 7564 1312
rect 7596 1311 7599 1343
rect 161 1283 217 1286
rect 161 1282 166 1283
rect 53 1252 166 1282
rect 212 1282 217 1283
rect 540 1283 596 1286
rect 540 1282 545 1283
rect 212 1252 326 1282
rect 432 1252 545 1282
rect 591 1282 596 1283
rect 919 1283 975 1286
rect 919 1282 924 1283
rect 591 1252 705 1282
rect 811 1252 924 1282
rect 970 1282 975 1283
rect 1298 1283 1354 1286
rect 1298 1282 1303 1283
rect 970 1252 1084 1282
rect 1190 1252 1303 1282
rect 1349 1282 1354 1283
rect 1677 1283 1733 1286
rect 1677 1282 1682 1283
rect 1349 1252 1463 1282
rect 1569 1252 1682 1282
rect 1728 1282 1733 1283
rect 2056 1283 2112 1286
rect 2056 1282 2061 1283
rect 1728 1252 1842 1282
rect 1948 1252 2061 1282
rect 2107 1282 2112 1283
rect 2435 1283 2491 1286
rect 2435 1282 2440 1283
rect 2107 1252 2221 1282
rect 2327 1252 2440 1282
rect 2486 1282 2491 1283
rect 2814 1283 2870 1286
rect 2814 1282 2819 1283
rect 2486 1252 2600 1282
rect 2706 1252 2819 1282
rect 2865 1282 2870 1283
rect 3193 1283 3249 1286
rect 3193 1282 3198 1283
rect 2865 1252 2979 1282
rect 3085 1252 3198 1282
rect 3244 1282 3249 1283
rect 3572 1283 3628 1286
rect 3572 1282 3577 1283
rect 3244 1252 3358 1282
rect 3464 1252 3577 1282
rect 3623 1282 3628 1283
rect 3951 1283 4007 1286
rect 3951 1282 3956 1283
rect 3623 1252 3737 1282
rect 3843 1252 3956 1282
rect 4002 1282 4007 1283
rect 4330 1283 4386 1286
rect 4330 1282 4335 1283
rect 4002 1252 4116 1282
rect 4222 1252 4335 1282
rect 4381 1282 4386 1283
rect 4709 1283 4765 1286
rect 4709 1282 4714 1283
rect 4381 1252 4495 1282
rect 4601 1252 4714 1282
rect 4760 1282 4765 1283
rect 5088 1283 5144 1286
rect 5088 1282 5093 1283
rect 4760 1252 4874 1282
rect 4980 1252 5093 1282
rect 5139 1282 5144 1283
rect 5467 1283 5523 1286
rect 5467 1282 5472 1283
rect 5139 1252 5253 1282
rect 5359 1252 5472 1282
rect 5518 1282 5523 1283
rect 5846 1283 5902 1286
rect 5846 1282 5851 1283
rect 5518 1252 5632 1282
rect 5738 1252 5851 1282
rect 5897 1282 5902 1283
rect 6225 1283 6281 1286
rect 6225 1282 6230 1283
rect 5897 1252 6011 1282
rect 6117 1252 6230 1282
rect 6276 1282 6281 1283
rect 6604 1283 6660 1286
rect 6604 1282 6609 1283
rect 6276 1252 6390 1282
rect 6496 1252 6609 1282
rect 6655 1282 6660 1283
rect 6983 1283 7039 1286
rect 6983 1282 6988 1283
rect 6655 1252 6769 1282
rect 6875 1252 6988 1282
rect 7034 1282 7039 1283
rect 7362 1283 7418 1286
rect 7362 1282 7367 1283
rect 7034 1252 7148 1282
rect 7254 1252 7367 1282
rect 7413 1282 7418 1283
rect 7413 1252 7527 1282
rect 161 1248 217 1252
rect 540 1248 596 1252
rect 919 1248 975 1252
rect 1298 1248 1354 1252
rect 1677 1248 1733 1252
rect 2056 1248 2112 1252
rect 2435 1248 2491 1252
rect 2814 1248 2870 1252
rect 3193 1248 3249 1252
rect 3572 1248 3628 1252
rect 3951 1248 4007 1252
rect 4330 1248 4386 1252
rect 4709 1248 4765 1252
rect 5088 1248 5144 1252
rect 5467 1248 5523 1252
rect 5846 1248 5902 1252
rect 6225 1248 6281 1252
rect 6604 1248 6660 1252
rect 6983 1248 7039 1252
rect 7362 1248 7418 1252
rect 161 1161 217 1164
rect 161 1160 166 1161
rect 53 1130 166 1160
rect 212 1160 217 1161
rect 540 1161 596 1164
rect 540 1160 545 1161
rect 212 1130 326 1160
rect 432 1130 545 1160
rect 591 1160 596 1161
rect 919 1161 975 1164
rect 919 1160 924 1161
rect 591 1130 705 1160
rect 811 1130 924 1160
rect 970 1160 975 1161
rect 1298 1161 1354 1164
rect 1298 1160 1303 1161
rect 970 1130 1084 1160
rect 1190 1130 1303 1160
rect 1349 1160 1354 1161
rect 1677 1161 1733 1164
rect 1677 1160 1682 1161
rect 1349 1130 1463 1160
rect 1569 1130 1682 1160
rect 1728 1160 1733 1161
rect 2056 1161 2112 1164
rect 2056 1160 2061 1161
rect 1728 1130 1842 1160
rect 1948 1130 2061 1160
rect 2107 1160 2112 1161
rect 2435 1161 2491 1164
rect 2435 1160 2440 1161
rect 2107 1130 2221 1160
rect 2327 1130 2440 1160
rect 2486 1160 2491 1161
rect 2814 1161 2870 1164
rect 2814 1160 2819 1161
rect 2486 1130 2600 1160
rect 2706 1130 2819 1160
rect 2865 1160 2870 1161
rect 3193 1161 3249 1164
rect 3193 1160 3198 1161
rect 2865 1130 2979 1160
rect 3085 1130 3198 1160
rect 3244 1160 3249 1161
rect 3572 1161 3628 1164
rect 3572 1160 3577 1161
rect 3244 1130 3358 1160
rect 3464 1130 3577 1160
rect 3623 1160 3628 1161
rect 3951 1161 4007 1164
rect 3951 1160 3956 1161
rect 3623 1130 3737 1160
rect 3843 1130 3956 1160
rect 4002 1160 4007 1161
rect 4330 1161 4386 1164
rect 4330 1160 4335 1161
rect 4002 1130 4116 1160
rect 4222 1130 4335 1160
rect 4381 1160 4386 1161
rect 4709 1161 4765 1164
rect 4709 1160 4714 1161
rect 4381 1130 4495 1160
rect 4601 1130 4714 1160
rect 4760 1160 4765 1161
rect 5088 1161 5144 1164
rect 5088 1160 5093 1161
rect 4760 1130 4874 1160
rect 4980 1130 5093 1160
rect 5139 1160 5144 1161
rect 5467 1161 5523 1164
rect 5467 1160 5472 1161
rect 5139 1130 5253 1160
rect 5359 1130 5472 1160
rect 5518 1160 5523 1161
rect 5846 1161 5902 1164
rect 5846 1160 5851 1161
rect 5518 1130 5632 1160
rect 5738 1130 5851 1160
rect 5897 1160 5902 1161
rect 6225 1161 6281 1164
rect 6225 1160 6230 1161
rect 5897 1130 6011 1160
rect 6117 1130 6230 1160
rect 6276 1160 6281 1161
rect 6604 1161 6660 1164
rect 6604 1160 6609 1161
rect 6276 1130 6390 1160
rect 6496 1130 6609 1160
rect 6655 1160 6660 1161
rect 6983 1161 7039 1164
rect 6983 1160 6988 1161
rect 6655 1130 6769 1160
rect 6875 1130 6988 1160
rect 7034 1160 7039 1161
rect 7362 1161 7418 1164
rect 7362 1160 7367 1161
rect 7034 1130 7148 1160
rect 7254 1130 7367 1160
rect 7413 1160 7418 1161
rect 7413 1130 7527 1160
rect 161 1126 217 1130
rect 540 1126 596 1130
rect 919 1126 975 1130
rect 1298 1126 1354 1130
rect 1677 1126 1733 1130
rect 2056 1126 2112 1130
rect 2435 1126 2491 1130
rect 2814 1126 2870 1130
rect 3193 1126 3249 1130
rect 3572 1126 3628 1130
rect 3951 1126 4007 1130
rect 4330 1126 4386 1130
rect 4709 1126 4765 1130
rect 5088 1126 5144 1130
rect 5467 1126 5523 1130
rect 5846 1126 5902 1130
rect 6225 1126 6281 1130
rect 6604 1126 6660 1130
rect 6983 1126 7039 1130
rect 7362 1126 7418 1130
rect -19 1068 -16 1100
rect 16 1099 19 1100
rect 360 1099 363 1100
rect 16 1069 146 1099
rect 232 1069 363 1099
rect 16 1068 19 1069
rect 360 1068 363 1069
rect 395 1099 398 1100
rect 739 1099 742 1100
rect 395 1069 525 1099
rect 611 1069 742 1099
rect 395 1068 398 1069
rect 739 1068 742 1069
rect 774 1099 777 1100
rect 1118 1099 1121 1100
rect 774 1069 904 1099
rect 990 1069 1121 1099
rect 774 1068 777 1069
rect 1118 1068 1121 1069
rect 1153 1099 1156 1100
rect 1497 1099 1500 1100
rect 1153 1069 1283 1099
rect 1369 1069 1500 1099
rect 1153 1068 1156 1069
rect 1497 1068 1500 1069
rect 1532 1099 1535 1100
rect 1876 1099 1879 1100
rect 1532 1069 1662 1099
rect 1748 1069 1879 1099
rect 1532 1068 1535 1069
rect 1876 1068 1879 1069
rect 1911 1099 1914 1100
rect 2255 1099 2258 1100
rect 1911 1069 2041 1099
rect 2127 1069 2258 1099
rect 1911 1068 1914 1069
rect 2255 1068 2258 1069
rect 2290 1099 2293 1100
rect 2634 1099 2637 1100
rect 2290 1069 2420 1099
rect 2506 1069 2637 1099
rect 2290 1068 2293 1069
rect 2634 1068 2637 1069
rect 2669 1099 2672 1100
rect 3013 1099 3016 1100
rect 2669 1069 2799 1099
rect 2885 1069 3016 1099
rect 2669 1068 2672 1069
rect 3013 1068 3016 1069
rect 3048 1099 3051 1100
rect 3392 1099 3395 1100
rect 3048 1069 3178 1099
rect 3264 1069 3395 1099
rect 3048 1068 3051 1069
rect 3392 1068 3395 1069
rect 3427 1099 3430 1100
rect 3771 1099 3774 1100
rect 3427 1069 3557 1099
rect 3643 1069 3774 1099
rect 3427 1068 3430 1069
rect 3771 1068 3774 1069
rect 3806 1099 3809 1100
rect 4150 1099 4153 1100
rect 3806 1069 3936 1099
rect 4022 1069 4153 1099
rect 3806 1068 3809 1069
rect 4150 1068 4153 1069
rect 4185 1099 4188 1100
rect 4529 1099 4532 1100
rect 4185 1069 4315 1099
rect 4401 1069 4532 1099
rect 4185 1068 4188 1069
rect 4529 1068 4532 1069
rect 4564 1099 4567 1100
rect 4908 1099 4911 1100
rect 4564 1069 4694 1099
rect 4780 1069 4911 1099
rect 4564 1068 4567 1069
rect 4908 1068 4911 1069
rect 4943 1099 4946 1100
rect 5287 1099 5290 1100
rect 4943 1069 5073 1099
rect 5159 1069 5290 1099
rect 4943 1068 4946 1069
rect 5287 1068 5290 1069
rect 5322 1099 5325 1100
rect 5666 1099 5669 1100
rect 5322 1069 5452 1099
rect 5538 1069 5669 1099
rect 5322 1068 5325 1069
rect 5666 1068 5669 1069
rect 5701 1099 5704 1100
rect 6045 1099 6048 1100
rect 5701 1069 5831 1099
rect 5917 1069 6048 1099
rect 5701 1068 5704 1069
rect 6045 1068 6048 1069
rect 6080 1099 6083 1100
rect 6424 1099 6427 1100
rect 6080 1069 6210 1099
rect 6296 1069 6427 1099
rect 6080 1068 6083 1069
rect 6424 1068 6427 1069
rect 6459 1099 6462 1100
rect 6803 1099 6806 1100
rect 6459 1069 6589 1099
rect 6675 1069 6806 1099
rect 6459 1068 6462 1069
rect 6803 1068 6806 1069
rect 6838 1099 6841 1100
rect 7182 1099 7185 1100
rect 6838 1069 6968 1099
rect 7054 1069 7185 1099
rect 6838 1068 6841 1069
rect 7182 1068 7185 1069
rect 7217 1099 7220 1100
rect 7561 1099 7564 1100
rect 7217 1069 7347 1099
rect 7433 1069 7564 1099
rect 7217 1068 7220 1069
rect 7561 1068 7564 1069
rect 7596 1068 7599 1100
rect 161 1040 217 1043
rect 161 1039 166 1040
rect 53 1009 166 1039
rect 212 1039 217 1040
rect 540 1040 596 1043
rect 540 1039 545 1040
rect 212 1009 326 1039
rect 432 1009 545 1039
rect 591 1039 596 1040
rect 919 1040 975 1043
rect 919 1039 924 1040
rect 591 1009 705 1039
rect 811 1009 924 1039
rect 970 1039 975 1040
rect 1298 1040 1354 1043
rect 1298 1039 1303 1040
rect 970 1009 1084 1039
rect 1190 1009 1303 1039
rect 1349 1039 1354 1040
rect 1677 1040 1733 1043
rect 1677 1039 1682 1040
rect 1349 1009 1463 1039
rect 1569 1009 1682 1039
rect 1728 1039 1733 1040
rect 2056 1040 2112 1043
rect 2056 1039 2061 1040
rect 1728 1009 1842 1039
rect 1948 1009 2061 1039
rect 2107 1039 2112 1040
rect 2435 1040 2491 1043
rect 2435 1039 2440 1040
rect 2107 1009 2221 1039
rect 2327 1009 2440 1039
rect 2486 1039 2491 1040
rect 2814 1040 2870 1043
rect 2814 1039 2819 1040
rect 2486 1009 2600 1039
rect 2706 1009 2819 1039
rect 2865 1039 2870 1040
rect 3193 1040 3249 1043
rect 3193 1039 3198 1040
rect 2865 1009 2979 1039
rect 3085 1009 3198 1039
rect 3244 1039 3249 1040
rect 3572 1040 3628 1043
rect 3572 1039 3577 1040
rect 3244 1009 3358 1039
rect 3464 1009 3577 1039
rect 3623 1039 3628 1040
rect 3951 1040 4007 1043
rect 3951 1039 3956 1040
rect 3623 1009 3737 1039
rect 3843 1009 3956 1039
rect 4002 1039 4007 1040
rect 4330 1040 4386 1043
rect 4330 1039 4335 1040
rect 4002 1009 4116 1039
rect 4222 1009 4335 1039
rect 4381 1039 4386 1040
rect 4709 1040 4765 1043
rect 4709 1039 4714 1040
rect 4381 1009 4495 1039
rect 4601 1009 4714 1039
rect 4760 1039 4765 1040
rect 5088 1040 5144 1043
rect 5088 1039 5093 1040
rect 4760 1009 4874 1039
rect 4980 1009 5093 1039
rect 5139 1039 5144 1040
rect 5467 1040 5523 1043
rect 5467 1039 5472 1040
rect 5139 1009 5253 1039
rect 5359 1009 5472 1039
rect 5518 1039 5523 1040
rect 5846 1040 5902 1043
rect 5846 1039 5851 1040
rect 5518 1009 5632 1039
rect 5738 1009 5851 1039
rect 5897 1039 5902 1040
rect 6225 1040 6281 1043
rect 6225 1039 6230 1040
rect 5897 1009 6011 1039
rect 6117 1009 6230 1039
rect 6276 1039 6281 1040
rect 6604 1040 6660 1043
rect 6604 1039 6609 1040
rect 6276 1009 6390 1039
rect 6496 1009 6609 1039
rect 6655 1039 6660 1040
rect 6983 1040 7039 1043
rect 6983 1039 6988 1040
rect 6655 1009 6769 1039
rect 6875 1009 6988 1039
rect 7034 1039 7039 1040
rect 7362 1040 7418 1043
rect 7362 1039 7367 1040
rect 7034 1009 7148 1039
rect 7254 1009 7367 1039
rect 7413 1039 7418 1040
rect 7413 1009 7527 1039
rect 161 1005 217 1009
rect 540 1005 596 1009
rect 919 1005 975 1009
rect 1298 1005 1354 1009
rect 1677 1005 1733 1009
rect 2056 1005 2112 1009
rect 2435 1005 2491 1009
rect 2814 1005 2870 1009
rect 3193 1005 3249 1009
rect 3572 1005 3628 1009
rect 3951 1005 4007 1009
rect 4330 1005 4386 1009
rect 4709 1005 4765 1009
rect 5088 1005 5144 1009
rect 5467 1005 5523 1009
rect 5846 1005 5902 1009
rect 6225 1005 6281 1009
rect 6604 1005 6660 1009
rect 6983 1005 7039 1009
rect 7362 1005 7418 1009
rect -19 948 -16 980
rect 16 979 19 980
rect 360 979 363 980
rect 16 949 146 979
rect 232 949 363 979
rect 16 948 19 949
rect 360 948 363 949
rect 395 979 398 980
rect 739 979 742 980
rect 395 949 525 979
rect 611 949 742 979
rect 395 948 398 949
rect 739 948 742 949
rect 774 979 777 980
rect 1118 979 1121 980
rect 774 949 904 979
rect 990 949 1121 979
rect 774 948 777 949
rect 1118 948 1121 949
rect 1153 979 1156 980
rect 1497 979 1500 980
rect 1153 949 1283 979
rect 1369 949 1500 979
rect 1153 948 1156 949
rect 1497 948 1500 949
rect 1532 979 1535 980
rect 1876 979 1879 980
rect 1532 949 1662 979
rect 1748 949 1879 979
rect 1532 948 1535 949
rect 1876 948 1879 949
rect 1911 979 1914 980
rect 2255 979 2258 980
rect 1911 949 2041 979
rect 2127 949 2258 979
rect 1911 948 1914 949
rect 2255 948 2258 949
rect 2290 979 2293 980
rect 2634 979 2637 980
rect 2290 949 2420 979
rect 2506 949 2637 979
rect 2290 948 2293 949
rect 2634 948 2637 949
rect 2669 979 2672 980
rect 3013 979 3016 980
rect 2669 949 2799 979
rect 2885 949 3016 979
rect 2669 948 2672 949
rect 3013 948 3016 949
rect 3048 979 3051 980
rect 3392 979 3395 980
rect 3048 949 3178 979
rect 3264 949 3395 979
rect 3048 948 3051 949
rect 3392 948 3395 949
rect 3427 979 3430 980
rect 3771 979 3774 980
rect 3427 949 3557 979
rect 3643 949 3774 979
rect 3427 948 3430 949
rect 3771 948 3774 949
rect 3806 979 3809 980
rect 4150 979 4153 980
rect 3806 949 3936 979
rect 4022 949 4153 979
rect 3806 948 3809 949
rect 4150 948 4153 949
rect 4185 979 4188 980
rect 4529 979 4532 980
rect 4185 949 4315 979
rect 4401 949 4532 979
rect 4185 948 4188 949
rect 4529 948 4532 949
rect 4564 979 4567 980
rect 4908 979 4911 980
rect 4564 949 4694 979
rect 4780 949 4911 979
rect 4564 948 4567 949
rect 4908 948 4911 949
rect 4943 979 4946 980
rect 5287 979 5290 980
rect 4943 949 5073 979
rect 5159 949 5290 979
rect 4943 948 4946 949
rect 5287 948 5290 949
rect 5322 979 5325 980
rect 5666 979 5669 980
rect 5322 949 5452 979
rect 5538 949 5669 979
rect 5322 948 5325 949
rect 5666 948 5669 949
rect 5701 979 5704 980
rect 6045 979 6048 980
rect 5701 949 5831 979
rect 5917 949 6048 979
rect 5701 948 5704 949
rect 6045 948 6048 949
rect 6080 979 6083 980
rect 6424 979 6427 980
rect 6080 949 6210 979
rect 6296 949 6427 979
rect 6080 948 6083 949
rect 6424 948 6427 949
rect 6459 979 6462 980
rect 6803 979 6806 980
rect 6459 949 6589 979
rect 6675 949 6806 979
rect 6459 948 6462 949
rect 6803 948 6806 949
rect 6838 979 6841 980
rect 7182 979 7185 980
rect 6838 949 6968 979
rect 7054 949 7185 979
rect 6838 948 6841 949
rect 7182 948 7185 949
rect 7217 979 7220 980
rect 7561 979 7564 980
rect 7217 949 7347 979
rect 7433 949 7564 979
rect 7217 948 7220 949
rect 7561 948 7564 949
rect 7596 948 7599 980
rect 161 920 217 923
rect 161 919 166 920
rect 53 889 166 919
rect 212 919 217 920
rect 540 920 596 923
rect 540 919 545 920
rect 212 889 326 919
rect 432 889 545 919
rect 591 919 596 920
rect 919 920 975 923
rect 919 919 924 920
rect 591 889 705 919
rect 811 889 924 919
rect 970 919 975 920
rect 1298 920 1354 923
rect 1298 919 1303 920
rect 970 889 1084 919
rect 1190 889 1303 919
rect 1349 919 1354 920
rect 1677 920 1733 923
rect 1677 919 1682 920
rect 1349 889 1463 919
rect 1569 889 1682 919
rect 1728 919 1733 920
rect 2056 920 2112 923
rect 2056 919 2061 920
rect 1728 889 1842 919
rect 1948 889 2061 919
rect 2107 919 2112 920
rect 2435 920 2491 923
rect 2435 919 2440 920
rect 2107 889 2221 919
rect 2327 889 2440 919
rect 2486 919 2491 920
rect 2814 920 2870 923
rect 2814 919 2819 920
rect 2486 889 2600 919
rect 2706 889 2819 919
rect 2865 919 2870 920
rect 3193 920 3249 923
rect 3193 919 3198 920
rect 2865 889 2979 919
rect 3085 889 3198 919
rect 3244 919 3249 920
rect 3572 920 3628 923
rect 3572 919 3577 920
rect 3244 889 3358 919
rect 3464 889 3577 919
rect 3623 919 3628 920
rect 3951 920 4007 923
rect 3951 919 3956 920
rect 3623 889 3737 919
rect 3843 889 3956 919
rect 4002 919 4007 920
rect 4330 920 4386 923
rect 4330 919 4335 920
rect 4002 889 4116 919
rect 4222 889 4335 919
rect 4381 919 4386 920
rect 4709 920 4765 923
rect 4709 919 4714 920
rect 4381 889 4495 919
rect 4601 889 4714 919
rect 4760 919 4765 920
rect 5088 920 5144 923
rect 5088 919 5093 920
rect 4760 889 4874 919
rect 4980 889 5093 919
rect 5139 919 5144 920
rect 5467 920 5523 923
rect 5467 919 5472 920
rect 5139 889 5253 919
rect 5359 889 5472 919
rect 5518 919 5523 920
rect 5846 920 5902 923
rect 5846 919 5851 920
rect 5518 889 5632 919
rect 5738 889 5851 919
rect 5897 919 5902 920
rect 6225 920 6281 923
rect 6225 919 6230 920
rect 5897 889 6011 919
rect 6117 889 6230 919
rect 6276 919 6281 920
rect 6604 920 6660 923
rect 6604 919 6609 920
rect 6276 889 6390 919
rect 6496 889 6609 919
rect 6655 919 6660 920
rect 6983 920 7039 923
rect 6983 919 6988 920
rect 6655 889 6769 919
rect 6875 889 6988 919
rect 7034 919 7039 920
rect 7362 920 7418 923
rect 7362 919 7367 920
rect 7034 889 7148 919
rect 7254 889 7367 919
rect 7413 919 7418 920
rect 7413 889 7527 919
rect 161 885 217 889
rect 540 885 596 889
rect 919 885 975 889
rect 1298 885 1354 889
rect 1677 885 1733 889
rect 2056 885 2112 889
rect 2435 885 2491 889
rect 2814 885 2870 889
rect 3193 885 3249 889
rect 3572 885 3628 889
rect 3951 885 4007 889
rect 4330 885 4386 889
rect 4709 885 4765 889
rect 5088 885 5144 889
rect 5467 885 5523 889
rect 5846 885 5902 889
rect 6225 885 6281 889
rect 6604 885 6660 889
rect 6983 885 7039 889
rect 7362 885 7418 889
rect -19 828 -16 860
rect 16 859 19 860
rect 360 859 363 860
rect 16 829 146 859
rect 232 829 363 859
rect 16 828 19 829
rect 360 828 363 829
rect 395 859 398 860
rect 739 859 742 860
rect 395 829 525 859
rect 611 829 742 859
rect 395 828 398 829
rect 739 828 742 829
rect 774 859 777 860
rect 1118 859 1121 860
rect 774 829 904 859
rect 990 829 1121 859
rect 774 828 777 829
rect 1118 828 1121 829
rect 1153 859 1156 860
rect 1497 859 1500 860
rect 1153 829 1283 859
rect 1369 829 1500 859
rect 1153 828 1156 829
rect 1497 828 1500 829
rect 1532 859 1535 860
rect 1876 859 1879 860
rect 1532 829 1662 859
rect 1748 829 1879 859
rect 1532 828 1535 829
rect 1876 828 1879 829
rect 1911 859 1914 860
rect 2255 859 2258 860
rect 1911 829 2041 859
rect 2127 829 2258 859
rect 1911 828 1914 829
rect 2255 828 2258 829
rect 2290 859 2293 860
rect 2634 859 2637 860
rect 2290 829 2420 859
rect 2506 829 2637 859
rect 2290 828 2293 829
rect 2634 828 2637 829
rect 2669 859 2672 860
rect 3013 859 3016 860
rect 2669 829 2799 859
rect 2885 829 3016 859
rect 2669 828 2672 829
rect 3013 828 3016 829
rect 3048 859 3051 860
rect 3392 859 3395 860
rect 3048 829 3178 859
rect 3264 829 3395 859
rect 3048 828 3051 829
rect 3392 828 3395 829
rect 3427 859 3430 860
rect 3771 859 3774 860
rect 3427 829 3557 859
rect 3643 829 3774 859
rect 3427 828 3430 829
rect 3771 828 3774 829
rect 3806 859 3809 860
rect 4150 859 4153 860
rect 3806 829 3936 859
rect 4022 829 4153 859
rect 3806 828 3809 829
rect 4150 828 4153 829
rect 4185 859 4188 860
rect 4529 859 4532 860
rect 4185 829 4315 859
rect 4401 829 4532 859
rect 4185 828 4188 829
rect 4529 828 4532 829
rect 4564 859 4567 860
rect 4908 859 4911 860
rect 4564 829 4694 859
rect 4780 829 4911 859
rect 4564 828 4567 829
rect 4908 828 4911 829
rect 4943 859 4946 860
rect 5287 859 5290 860
rect 4943 829 5073 859
rect 5159 829 5290 859
rect 4943 828 4946 829
rect 5287 828 5290 829
rect 5322 859 5325 860
rect 5666 859 5669 860
rect 5322 829 5452 859
rect 5538 829 5669 859
rect 5322 828 5325 829
rect 5666 828 5669 829
rect 5701 859 5704 860
rect 6045 859 6048 860
rect 5701 829 5831 859
rect 5917 829 6048 859
rect 5701 828 5704 829
rect 6045 828 6048 829
rect 6080 859 6083 860
rect 6424 859 6427 860
rect 6080 829 6210 859
rect 6296 829 6427 859
rect 6080 828 6083 829
rect 6424 828 6427 829
rect 6459 859 6462 860
rect 6803 859 6806 860
rect 6459 829 6589 859
rect 6675 829 6806 859
rect 6459 828 6462 829
rect 6803 828 6806 829
rect 6838 859 6841 860
rect 7182 859 7185 860
rect 6838 829 6968 859
rect 7054 829 7185 859
rect 6838 828 6841 829
rect 7182 828 7185 829
rect 7217 859 7220 860
rect 7561 859 7564 860
rect 7217 829 7347 859
rect 7433 829 7564 859
rect 7217 828 7220 829
rect 7561 828 7564 829
rect 7596 828 7599 860
rect 161 800 217 803
rect 161 799 166 800
rect 53 769 166 799
rect 212 799 217 800
rect 540 800 596 803
rect 540 799 545 800
rect 212 769 326 799
rect 432 769 545 799
rect 591 799 596 800
rect 919 800 975 803
rect 919 799 924 800
rect 591 769 705 799
rect 811 769 924 799
rect 970 799 975 800
rect 1298 800 1354 803
rect 1298 799 1303 800
rect 970 769 1084 799
rect 1190 769 1303 799
rect 1349 799 1354 800
rect 1677 800 1733 803
rect 1677 799 1682 800
rect 1349 769 1463 799
rect 1569 769 1682 799
rect 1728 799 1733 800
rect 2056 800 2112 803
rect 2056 799 2061 800
rect 1728 769 1842 799
rect 1948 769 2061 799
rect 2107 799 2112 800
rect 2435 800 2491 803
rect 2435 799 2440 800
rect 2107 769 2221 799
rect 2327 769 2440 799
rect 2486 799 2491 800
rect 2814 800 2870 803
rect 2814 799 2819 800
rect 2486 769 2600 799
rect 2706 769 2819 799
rect 2865 799 2870 800
rect 3193 800 3249 803
rect 3193 799 3198 800
rect 2865 769 2979 799
rect 3085 769 3198 799
rect 3244 799 3249 800
rect 3572 800 3628 803
rect 3572 799 3577 800
rect 3244 769 3358 799
rect 3464 769 3577 799
rect 3623 799 3628 800
rect 3951 800 4007 803
rect 3951 799 3956 800
rect 3623 769 3737 799
rect 3843 769 3956 799
rect 4002 799 4007 800
rect 4330 800 4386 803
rect 4330 799 4335 800
rect 4002 769 4116 799
rect 4222 769 4335 799
rect 4381 799 4386 800
rect 4709 800 4765 803
rect 4709 799 4714 800
rect 4381 769 4495 799
rect 4601 769 4714 799
rect 4760 799 4765 800
rect 5088 800 5144 803
rect 5088 799 5093 800
rect 4760 769 4874 799
rect 4980 769 5093 799
rect 5139 799 5144 800
rect 5467 800 5523 803
rect 5467 799 5472 800
rect 5139 769 5253 799
rect 5359 769 5472 799
rect 5518 799 5523 800
rect 5846 800 5902 803
rect 5846 799 5851 800
rect 5518 769 5632 799
rect 5738 769 5851 799
rect 5897 799 5902 800
rect 6225 800 6281 803
rect 6225 799 6230 800
rect 5897 769 6011 799
rect 6117 769 6230 799
rect 6276 799 6281 800
rect 6604 800 6660 803
rect 6604 799 6609 800
rect 6276 769 6390 799
rect 6496 769 6609 799
rect 6655 799 6660 800
rect 6983 800 7039 803
rect 6983 799 6988 800
rect 6655 769 6769 799
rect 6875 769 6988 799
rect 7034 799 7039 800
rect 7362 800 7418 803
rect 7362 799 7367 800
rect 7034 769 7148 799
rect 7254 769 7367 799
rect 7413 799 7418 800
rect 7413 769 7527 799
rect 161 765 217 769
rect 540 765 596 769
rect 919 765 975 769
rect 1298 765 1354 769
rect 1677 765 1733 769
rect 2056 765 2112 769
rect 2435 765 2491 769
rect 2814 765 2870 769
rect 3193 765 3249 769
rect 3572 765 3628 769
rect 3951 765 4007 769
rect 4330 765 4386 769
rect 4709 765 4765 769
rect 5088 765 5144 769
rect 5467 765 5523 769
rect 5846 765 5902 769
rect 6225 765 6281 769
rect 6604 765 6660 769
rect 6983 765 7039 769
rect 7362 765 7418 769
rect -19 708 -16 740
rect 16 739 19 740
rect 360 739 363 740
rect 16 709 146 739
rect 232 709 363 739
rect 16 708 19 709
rect 360 708 363 709
rect 395 739 398 740
rect 739 739 742 740
rect 395 709 525 739
rect 611 709 742 739
rect 395 708 398 709
rect 739 708 742 709
rect 774 739 777 740
rect 1118 739 1121 740
rect 774 709 904 739
rect 990 709 1121 739
rect 774 708 777 709
rect 1118 708 1121 709
rect 1153 739 1156 740
rect 1497 739 1500 740
rect 1153 709 1283 739
rect 1369 709 1500 739
rect 1153 708 1156 709
rect 1497 708 1500 709
rect 1532 739 1535 740
rect 1876 739 1879 740
rect 1532 709 1662 739
rect 1748 709 1879 739
rect 1532 708 1535 709
rect 1876 708 1879 709
rect 1911 739 1914 740
rect 2255 739 2258 740
rect 1911 709 2041 739
rect 2127 709 2258 739
rect 1911 708 1914 709
rect 2255 708 2258 709
rect 2290 739 2293 740
rect 2634 739 2637 740
rect 2290 709 2420 739
rect 2506 709 2637 739
rect 2290 708 2293 709
rect 2634 708 2637 709
rect 2669 739 2672 740
rect 3013 739 3016 740
rect 2669 709 2799 739
rect 2885 709 3016 739
rect 2669 708 2672 709
rect 3013 708 3016 709
rect 3048 739 3051 740
rect 3392 739 3395 740
rect 3048 709 3178 739
rect 3264 709 3395 739
rect 3048 708 3051 709
rect 3392 708 3395 709
rect 3427 739 3430 740
rect 3771 739 3774 740
rect 3427 709 3557 739
rect 3643 709 3774 739
rect 3427 708 3430 709
rect 3771 708 3774 709
rect 3806 739 3809 740
rect 4150 739 4153 740
rect 3806 709 3936 739
rect 4022 709 4153 739
rect 3806 708 3809 709
rect 4150 708 4153 709
rect 4185 739 4188 740
rect 4529 739 4532 740
rect 4185 709 4315 739
rect 4401 709 4532 739
rect 4185 708 4188 709
rect 4529 708 4532 709
rect 4564 739 4567 740
rect 4908 739 4911 740
rect 4564 709 4694 739
rect 4780 709 4911 739
rect 4564 708 4567 709
rect 4908 708 4911 709
rect 4943 739 4946 740
rect 5287 739 5290 740
rect 4943 709 5073 739
rect 5159 709 5290 739
rect 4943 708 4946 709
rect 5287 708 5290 709
rect 5322 739 5325 740
rect 5666 739 5669 740
rect 5322 709 5452 739
rect 5538 709 5669 739
rect 5322 708 5325 709
rect 5666 708 5669 709
rect 5701 739 5704 740
rect 6045 739 6048 740
rect 5701 709 5831 739
rect 5917 709 6048 739
rect 5701 708 5704 709
rect 6045 708 6048 709
rect 6080 739 6083 740
rect 6424 739 6427 740
rect 6080 709 6210 739
rect 6296 709 6427 739
rect 6080 708 6083 709
rect 6424 708 6427 709
rect 6459 739 6462 740
rect 6803 739 6806 740
rect 6459 709 6589 739
rect 6675 709 6806 739
rect 6459 708 6462 709
rect 6803 708 6806 709
rect 6838 739 6841 740
rect 7182 739 7185 740
rect 6838 709 6968 739
rect 7054 709 7185 739
rect 6838 708 6841 709
rect 7182 708 7185 709
rect 7217 739 7220 740
rect 7561 739 7564 740
rect 7217 709 7347 739
rect 7433 709 7564 739
rect 7217 708 7220 709
rect 7561 708 7564 709
rect 7596 708 7599 740
rect 161 680 217 683
rect 161 679 166 680
rect 53 649 166 679
rect 212 679 217 680
rect 540 680 596 683
rect 540 679 545 680
rect 212 649 326 679
rect 432 649 545 679
rect 591 679 596 680
rect 919 680 975 683
rect 919 679 924 680
rect 591 649 705 679
rect 811 649 924 679
rect 970 679 975 680
rect 1298 680 1354 683
rect 1298 679 1303 680
rect 970 649 1084 679
rect 1190 649 1303 679
rect 1349 679 1354 680
rect 1677 680 1733 683
rect 1677 679 1682 680
rect 1349 649 1463 679
rect 1569 649 1682 679
rect 1728 679 1733 680
rect 2056 680 2112 683
rect 2056 679 2061 680
rect 1728 649 1842 679
rect 1948 649 2061 679
rect 2107 679 2112 680
rect 2435 680 2491 683
rect 2435 679 2440 680
rect 2107 649 2221 679
rect 2327 649 2440 679
rect 2486 679 2491 680
rect 2814 680 2870 683
rect 2814 679 2819 680
rect 2486 649 2600 679
rect 2706 649 2819 679
rect 2865 679 2870 680
rect 3193 680 3249 683
rect 3193 679 3198 680
rect 2865 649 2979 679
rect 3085 649 3198 679
rect 3244 679 3249 680
rect 3572 680 3628 683
rect 3572 679 3577 680
rect 3244 649 3358 679
rect 3464 649 3577 679
rect 3623 679 3628 680
rect 3951 680 4007 683
rect 3951 679 3956 680
rect 3623 649 3737 679
rect 3843 649 3956 679
rect 4002 679 4007 680
rect 4330 680 4386 683
rect 4330 679 4335 680
rect 4002 649 4116 679
rect 4222 649 4335 679
rect 4381 679 4386 680
rect 4709 680 4765 683
rect 4709 679 4714 680
rect 4381 649 4495 679
rect 4601 649 4714 679
rect 4760 679 4765 680
rect 5088 680 5144 683
rect 5088 679 5093 680
rect 4760 649 4874 679
rect 4980 649 5093 679
rect 5139 679 5144 680
rect 5467 680 5523 683
rect 5467 679 5472 680
rect 5139 649 5253 679
rect 5359 649 5472 679
rect 5518 679 5523 680
rect 5846 680 5902 683
rect 5846 679 5851 680
rect 5518 649 5632 679
rect 5738 649 5851 679
rect 5897 679 5902 680
rect 6225 680 6281 683
rect 6225 679 6230 680
rect 5897 649 6011 679
rect 6117 649 6230 679
rect 6276 679 6281 680
rect 6604 680 6660 683
rect 6604 679 6609 680
rect 6276 649 6390 679
rect 6496 649 6609 679
rect 6655 679 6660 680
rect 6983 680 7039 683
rect 6983 679 6988 680
rect 6655 649 6769 679
rect 6875 649 6988 679
rect 7034 679 7039 680
rect 7362 680 7418 683
rect 7362 679 7367 680
rect 7034 649 7148 679
rect 7254 649 7367 679
rect 7413 679 7418 680
rect 7413 649 7527 679
rect 161 645 217 649
rect 540 645 596 649
rect 919 645 975 649
rect 1298 645 1354 649
rect 1677 645 1733 649
rect 2056 645 2112 649
rect 2435 645 2491 649
rect 2814 645 2870 649
rect 3193 645 3249 649
rect 3572 645 3628 649
rect 3951 645 4007 649
rect 4330 645 4386 649
rect 4709 645 4765 649
rect 5088 645 5144 649
rect 5467 645 5523 649
rect 5846 645 5902 649
rect 6225 645 6281 649
rect 6604 645 6660 649
rect 6983 645 7039 649
rect 7362 645 7418 649
rect 161 558 217 561
rect 161 557 166 558
rect 53 527 166 557
rect 212 557 217 558
rect 540 558 596 561
rect 540 557 545 558
rect 212 527 326 557
rect 432 527 545 557
rect 591 557 596 558
rect 919 558 975 561
rect 919 557 924 558
rect 591 527 705 557
rect 811 527 924 557
rect 970 557 975 558
rect 1298 558 1354 561
rect 1298 557 1303 558
rect 970 527 1084 557
rect 1190 527 1303 557
rect 1349 557 1354 558
rect 1677 558 1733 561
rect 1677 557 1682 558
rect 1349 527 1463 557
rect 1569 527 1682 557
rect 1728 557 1733 558
rect 2056 558 2112 561
rect 2056 557 2061 558
rect 1728 527 1842 557
rect 1948 527 2061 557
rect 2107 557 2112 558
rect 2435 558 2491 561
rect 2435 557 2440 558
rect 2107 527 2221 557
rect 2327 527 2440 557
rect 2486 557 2491 558
rect 2814 558 2870 561
rect 2814 557 2819 558
rect 2486 527 2600 557
rect 2706 527 2819 557
rect 2865 557 2870 558
rect 3193 558 3249 561
rect 3193 557 3198 558
rect 2865 527 2979 557
rect 3085 527 3198 557
rect 3244 557 3249 558
rect 3572 558 3628 561
rect 3572 557 3577 558
rect 3244 527 3358 557
rect 3464 527 3577 557
rect 3623 557 3628 558
rect 3951 558 4007 561
rect 3951 557 3956 558
rect 3623 527 3737 557
rect 3843 527 3956 557
rect 4002 557 4007 558
rect 4330 558 4386 561
rect 4330 557 4335 558
rect 4002 527 4116 557
rect 4222 527 4335 557
rect 4381 557 4386 558
rect 4709 558 4765 561
rect 4709 557 4714 558
rect 4381 527 4495 557
rect 4601 527 4714 557
rect 4760 557 4765 558
rect 5088 558 5144 561
rect 5088 557 5093 558
rect 4760 527 4874 557
rect 4980 527 5093 557
rect 5139 557 5144 558
rect 5467 558 5523 561
rect 5467 557 5472 558
rect 5139 527 5253 557
rect 5359 527 5472 557
rect 5518 557 5523 558
rect 5846 558 5902 561
rect 5846 557 5851 558
rect 5518 527 5632 557
rect 5738 527 5851 557
rect 5897 557 5902 558
rect 6225 558 6281 561
rect 6225 557 6230 558
rect 5897 527 6011 557
rect 6117 527 6230 557
rect 6276 557 6281 558
rect 6604 558 6660 561
rect 6604 557 6609 558
rect 6276 527 6390 557
rect 6496 527 6609 557
rect 6655 557 6660 558
rect 6983 558 7039 561
rect 6983 557 6988 558
rect 6655 527 6769 557
rect 6875 527 6988 557
rect 7034 557 7039 558
rect 7362 558 7418 561
rect 7362 557 7367 558
rect 7034 527 7148 557
rect 7254 527 7367 557
rect 7413 557 7418 558
rect 7413 527 7527 557
rect 161 523 217 527
rect 540 523 596 527
rect 919 523 975 527
rect 1298 523 1354 527
rect 1677 523 1733 527
rect 2056 523 2112 527
rect 2435 523 2491 527
rect 2814 523 2870 527
rect 3193 523 3249 527
rect 3572 523 3628 527
rect 3951 523 4007 527
rect 4330 523 4386 527
rect 4709 523 4765 527
rect 5088 523 5144 527
rect 5467 523 5523 527
rect 5846 523 5902 527
rect 6225 523 6281 527
rect 6604 523 6660 527
rect 6983 523 7039 527
rect 7362 523 7418 527
rect -19 465 -16 497
rect 16 496 19 497
rect 360 496 363 497
rect 16 466 146 496
rect 232 466 363 496
rect 16 465 19 466
rect 360 465 363 466
rect 395 496 398 497
rect 739 496 742 497
rect 395 466 525 496
rect 611 466 742 496
rect 395 465 398 466
rect 739 465 742 466
rect 774 496 777 497
rect 1118 496 1121 497
rect 774 466 904 496
rect 990 466 1121 496
rect 774 465 777 466
rect 1118 465 1121 466
rect 1153 496 1156 497
rect 1497 496 1500 497
rect 1153 466 1283 496
rect 1369 466 1500 496
rect 1153 465 1156 466
rect 1497 465 1500 466
rect 1532 496 1535 497
rect 1876 496 1879 497
rect 1532 466 1662 496
rect 1748 466 1879 496
rect 1532 465 1535 466
rect 1876 465 1879 466
rect 1911 496 1914 497
rect 2255 496 2258 497
rect 1911 466 2041 496
rect 2127 466 2258 496
rect 1911 465 1914 466
rect 2255 465 2258 466
rect 2290 496 2293 497
rect 2634 496 2637 497
rect 2290 466 2420 496
rect 2506 466 2637 496
rect 2290 465 2293 466
rect 2634 465 2637 466
rect 2669 496 2672 497
rect 3013 496 3016 497
rect 2669 466 2799 496
rect 2885 466 3016 496
rect 2669 465 2672 466
rect 3013 465 3016 466
rect 3048 496 3051 497
rect 3392 496 3395 497
rect 3048 466 3178 496
rect 3264 466 3395 496
rect 3048 465 3051 466
rect 3392 465 3395 466
rect 3427 496 3430 497
rect 3771 496 3774 497
rect 3427 466 3557 496
rect 3643 466 3774 496
rect 3427 465 3430 466
rect 3771 465 3774 466
rect 3806 496 3809 497
rect 4150 496 4153 497
rect 3806 466 3936 496
rect 4022 466 4153 496
rect 3806 465 3809 466
rect 4150 465 4153 466
rect 4185 496 4188 497
rect 4529 496 4532 497
rect 4185 466 4315 496
rect 4401 466 4532 496
rect 4185 465 4188 466
rect 4529 465 4532 466
rect 4564 496 4567 497
rect 4908 496 4911 497
rect 4564 466 4694 496
rect 4780 466 4911 496
rect 4564 465 4567 466
rect 4908 465 4911 466
rect 4943 496 4946 497
rect 5287 496 5290 497
rect 4943 466 5073 496
rect 5159 466 5290 496
rect 4943 465 4946 466
rect 5287 465 5290 466
rect 5322 496 5325 497
rect 5666 496 5669 497
rect 5322 466 5452 496
rect 5538 466 5669 496
rect 5322 465 5325 466
rect 5666 465 5669 466
rect 5701 496 5704 497
rect 6045 496 6048 497
rect 5701 466 5831 496
rect 5917 466 6048 496
rect 5701 465 5704 466
rect 6045 465 6048 466
rect 6080 496 6083 497
rect 6424 496 6427 497
rect 6080 466 6210 496
rect 6296 466 6427 496
rect 6080 465 6083 466
rect 6424 465 6427 466
rect 6459 496 6462 497
rect 6803 496 6806 497
rect 6459 466 6589 496
rect 6675 466 6806 496
rect 6459 465 6462 466
rect 6803 465 6806 466
rect 6838 496 6841 497
rect 7182 496 7185 497
rect 6838 466 6968 496
rect 7054 466 7185 496
rect 6838 465 6841 466
rect 7182 465 7185 466
rect 7217 496 7220 497
rect 7561 496 7564 497
rect 7217 466 7347 496
rect 7433 466 7564 496
rect 7217 465 7220 466
rect 7561 465 7564 466
rect 7596 465 7599 497
rect 161 437 217 440
rect 161 436 166 437
rect 53 406 166 436
rect 212 436 217 437
rect 540 437 596 440
rect 540 436 545 437
rect 212 406 326 436
rect 432 406 545 436
rect 591 436 596 437
rect 919 437 975 440
rect 919 436 924 437
rect 591 406 705 436
rect 811 406 924 436
rect 970 436 975 437
rect 1298 437 1354 440
rect 1298 436 1303 437
rect 970 406 1084 436
rect 1190 406 1303 436
rect 1349 436 1354 437
rect 1677 437 1733 440
rect 1677 436 1682 437
rect 1349 406 1463 436
rect 1569 406 1682 436
rect 1728 436 1733 437
rect 2056 437 2112 440
rect 2056 436 2061 437
rect 1728 406 1842 436
rect 1948 406 2061 436
rect 2107 436 2112 437
rect 2435 437 2491 440
rect 2435 436 2440 437
rect 2107 406 2221 436
rect 2327 406 2440 436
rect 2486 436 2491 437
rect 2814 437 2870 440
rect 2814 436 2819 437
rect 2486 406 2600 436
rect 2706 406 2819 436
rect 2865 436 2870 437
rect 3193 437 3249 440
rect 3193 436 3198 437
rect 2865 406 2979 436
rect 3085 406 3198 436
rect 3244 436 3249 437
rect 3572 437 3628 440
rect 3572 436 3577 437
rect 3244 406 3358 436
rect 3464 406 3577 436
rect 3623 436 3628 437
rect 3951 437 4007 440
rect 3951 436 3956 437
rect 3623 406 3737 436
rect 3843 406 3956 436
rect 4002 436 4007 437
rect 4330 437 4386 440
rect 4330 436 4335 437
rect 4002 406 4116 436
rect 4222 406 4335 436
rect 4381 436 4386 437
rect 4709 437 4765 440
rect 4709 436 4714 437
rect 4381 406 4495 436
rect 4601 406 4714 436
rect 4760 436 4765 437
rect 5088 437 5144 440
rect 5088 436 5093 437
rect 4760 406 4874 436
rect 4980 406 5093 436
rect 5139 436 5144 437
rect 5467 437 5523 440
rect 5467 436 5472 437
rect 5139 406 5253 436
rect 5359 406 5472 436
rect 5518 436 5523 437
rect 5846 437 5902 440
rect 5846 436 5851 437
rect 5518 406 5632 436
rect 5738 406 5851 436
rect 5897 436 5902 437
rect 6225 437 6281 440
rect 6225 436 6230 437
rect 5897 406 6011 436
rect 6117 406 6230 436
rect 6276 436 6281 437
rect 6604 437 6660 440
rect 6604 436 6609 437
rect 6276 406 6390 436
rect 6496 406 6609 436
rect 6655 436 6660 437
rect 6983 437 7039 440
rect 6983 436 6988 437
rect 6655 406 6769 436
rect 6875 406 6988 436
rect 7034 436 7039 437
rect 7362 437 7418 440
rect 7362 436 7367 437
rect 7034 406 7148 436
rect 7254 406 7367 436
rect 7413 436 7418 437
rect 7413 406 7527 436
rect 161 402 217 406
rect 540 402 596 406
rect 919 402 975 406
rect 1298 402 1354 406
rect 1677 402 1733 406
rect 2056 402 2112 406
rect 2435 402 2491 406
rect 2814 402 2870 406
rect 3193 402 3249 406
rect 3572 402 3628 406
rect 3951 402 4007 406
rect 4330 402 4386 406
rect 4709 402 4765 406
rect 5088 402 5144 406
rect 5467 402 5523 406
rect 5846 402 5902 406
rect 6225 402 6281 406
rect 6604 402 6660 406
rect 6983 402 7039 406
rect 7362 402 7418 406
rect -19 345 -16 377
rect 16 376 19 377
rect 360 376 363 377
rect 16 346 146 376
rect 232 346 363 376
rect 16 345 19 346
rect 360 345 363 346
rect 395 376 398 377
rect 739 376 742 377
rect 395 346 525 376
rect 611 346 742 376
rect 395 345 398 346
rect 739 345 742 346
rect 774 376 777 377
rect 1118 376 1121 377
rect 774 346 904 376
rect 990 346 1121 376
rect 774 345 777 346
rect 1118 345 1121 346
rect 1153 376 1156 377
rect 1497 376 1500 377
rect 1153 346 1283 376
rect 1369 346 1500 376
rect 1153 345 1156 346
rect 1497 345 1500 346
rect 1532 376 1535 377
rect 1876 376 1879 377
rect 1532 346 1662 376
rect 1748 346 1879 376
rect 1532 345 1535 346
rect 1876 345 1879 346
rect 1911 376 1914 377
rect 2255 376 2258 377
rect 1911 346 2041 376
rect 2127 346 2258 376
rect 1911 345 1914 346
rect 2255 345 2258 346
rect 2290 376 2293 377
rect 2634 376 2637 377
rect 2290 346 2420 376
rect 2506 346 2637 376
rect 2290 345 2293 346
rect 2634 345 2637 346
rect 2669 376 2672 377
rect 3013 376 3016 377
rect 2669 346 2799 376
rect 2885 346 3016 376
rect 2669 345 2672 346
rect 3013 345 3016 346
rect 3048 376 3051 377
rect 3392 376 3395 377
rect 3048 346 3178 376
rect 3264 346 3395 376
rect 3048 345 3051 346
rect 3392 345 3395 346
rect 3427 376 3430 377
rect 3771 376 3774 377
rect 3427 346 3557 376
rect 3643 346 3774 376
rect 3427 345 3430 346
rect 3771 345 3774 346
rect 3806 376 3809 377
rect 4150 376 4153 377
rect 3806 346 3936 376
rect 4022 346 4153 376
rect 3806 345 3809 346
rect 4150 345 4153 346
rect 4185 376 4188 377
rect 4529 376 4532 377
rect 4185 346 4315 376
rect 4401 346 4532 376
rect 4185 345 4188 346
rect 4529 345 4532 346
rect 4564 376 4567 377
rect 4908 376 4911 377
rect 4564 346 4694 376
rect 4780 346 4911 376
rect 4564 345 4567 346
rect 4908 345 4911 346
rect 4943 376 4946 377
rect 5287 376 5290 377
rect 4943 346 5073 376
rect 5159 346 5290 376
rect 4943 345 4946 346
rect 5287 345 5290 346
rect 5322 376 5325 377
rect 5666 376 5669 377
rect 5322 346 5452 376
rect 5538 346 5669 376
rect 5322 345 5325 346
rect 5666 345 5669 346
rect 5701 376 5704 377
rect 6045 376 6048 377
rect 5701 346 5831 376
rect 5917 346 6048 376
rect 5701 345 5704 346
rect 6045 345 6048 346
rect 6080 376 6083 377
rect 6424 376 6427 377
rect 6080 346 6210 376
rect 6296 346 6427 376
rect 6080 345 6083 346
rect 6424 345 6427 346
rect 6459 376 6462 377
rect 6803 376 6806 377
rect 6459 346 6589 376
rect 6675 346 6806 376
rect 6459 345 6462 346
rect 6803 345 6806 346
rect 6838 376 6841 377
rect 7182 376 7185 377
rect 6838 346 6968 376
rect 7054 346 7185 376
rect 6838 345 6841 346
rect 7182 345 7185 346
rect 7217 376 7220 377
rect 7561 376 7564 377
rect 7217 346 7347 376
rect 7433 346 7564 376
rect 7217 345 7220 346
rect 7561 345 7564 346
rect 7596 345 7599 377
rect 161 317 217 320
rect 161 316 166 317
rect 53 286 166 316
rect 212 316 217 317
rect 540 317 596 320
rect 540 316 545 317
rect 212 286 326 316
rect 432 286 545 316
rect 591 316 596 317
rect 919 317 975 320
rect 919 316 924 317
rect 591 286 705 316
rect 811 286 924 316
rect 970 316 975 317
rect 1298 317 1354 320
rect 1298 316 1303 317
rect 970 286 1084 316
rect 1190 286 1303 316
rect 1349 316 1354 317
rect 1677 317 1733 320
rect 1677 316 1682 317
rect 1349 286 1463 316
rect 1569 286 1682 316
rect 1728 316 1733 317
rect 2056 317 2112 320
rect 2056 316 2061 317
rect 1728 286 1842 316
rect 1948 286 2061 316
rect 2107 316 2112 317
rect 2435 317 2491 320
rect 2435 316 2440 317
rect 2107 286 2221 316
rect 2327 286 2440 316
rect 2486 316 2491 317
rect 2814 317 2870 320
rect 2814 316 2819 317
rect 2486 286 2600 316
rect 2706 286 2819 316
rect 2865 316 2870 317
rect 3193 317 3249 320
rect 3193 316 3198 317
rect 2865 286 2979 316
rect 3085 286 3198 316
rect 3244 316 3249 317
rect 3572 317 3628 320
rect 3572 316 3577 317
rect 3244 286 3358 316
rect 3464 286 3577 316
rect 3623 316 3628 317
rect 3951 317 4007 320
rect 3951 316 3956 317
rect 3623 286 3737 316
rect 3843 286 3956 316
rect 4002 316 4007 317
rect 4330 317 4386 320
rect 4330 316 4335 317
rect 4002 286 4116 316
rect 4222 286 4335 316
rect 4381 316 4386 317
rect 4709 317 4765 320
rect 4709 316 4714 317
rect 4381 286 4495 316
rect 4601 286 4714 316
rect 4760 316 4765 317
rect 5088 317 5144 320
rect 5088 316 5093 317
rect 4760 286 4874 316
rect 4980 286 5093 316
rect 5139 316 5144 317
rect 5467 317 5523 320
rect 5467 316 5472 317
rect 5139 286 5253 316
rect 5359 286 5472 316
rect 5518 316 5523 317
rect 5846 317 5902 320
rect 5846 316 5851 317
rect 5518 286 5632 316
rect 5738 286 5851 316
rect 5897 316 5902 317
rect 6225 317 6281 320
rect 6225 316 6230 317
rect 5897 286 6011 316
rect 6117 286 6230 316
rect 6276 316 6281 317
rect 6604 317 6660 320
rect 6604 316 6609 317
rect 6276 286 6390 316
rect 6496 286 6609 316
rect 6655 316 6660 317
rect 6983 317 7039 320
rect 6983 316 6988 317
rect 6655 286 6769 316
rect 6875 286 6988 316
rect 7034 316 7039 317
rect 7362 317 7418 320
rect 7362 316 7367 317
rect 7034 286 7148 316
rect 7254 286 7367 316
rect 7413 316 7418 317
rect 7413 286 7527 316
rect 161 282 217 286
rect 540 282 596 286
rect 919 282 975 286
rect 1298 282 1354 286
rect 1677 282 1733 286
rect 2056 282 2112 286
rect 2435 282 2491 286
rect 2814 282 2870 286
rect 3193 282 3249 286
rect 3572 282 3628 286
rect 3951 282 4007 286
rect 4330 282 4386 286
rect 4709 282 4765 286
rect 5088 282 5144 286
rect 5467 282 5523 286
rect 5846 282 5902 286
rect 6225 282 6281 286
rect 6604 282 6660 286
rect 6983 282 7039 286
rect 7362 282 7418 286
rect -19 225 -16 257
rect 16 256 19 257
rect 360 256 363 257
rect 16 226 146 256
rect 232 226 363 256
rect 16 225 19 226
rect 360 225 363 226
rect 395 256 398 257
rect 739 256 742 257
rect 395 226 525 256
rect 611 226 742 256
rect 395 225 398 226
rect 739 225 742 226
rect 774 256 777 257
rect 1118 256 1121 257
rect 774 226 904 256
rect 990 226 1121 256
rect 774 225 777 226
rect 1118 225 1121 226
rect 1153 256 1156 257
rect 1497 256 1500 257
rect 1153 226 1283 256
rect 1369 226 1500 256
rect 1153 225 1156 226
rect 1497 225 1500 226
rect 1532 256 1535 257
rect 1876 256 1879 257
rect 1532 226 1662 256
rect 1748 226 1879 256
rect 1532 225 1535 226
rect 1876 225 1879 226
rect 1911 256 1914 257
rect 2255 256 2258 257
rect 1911 226 2041 256
rect 2127 226 2258 256
rect 1911 225 1914 226
rect 2255 225 2258 226
rect 2290 256 2293 257
rect 2634 256 2637 257
rect 2290 226 2420 256
rect 2506 226 2637 256
rect 2290 225 2293 226
rect 2634 225 2637 226
rect 2669 256 2672 257
rect 3013 256 3016 257
rect 2669 226 2799 256
rect 2885 226 3016 256
rect 2669 225 2672 226
rect 3013 225 3016 226
rect 3048 256 3051 257
rect 3392 256 3395 257
rect 3048 226 3178 256
rect 3264 226 3395 256
rect 3048 225 3051 226
rect 3392 225 3395 226
rect 3427 256 3430 257
rect 3771 256 3774 257
rect 3427 226 3557 256
rect 3643 226 3774 256
rect 3427 225 3430 226
rect 3771 225 3774 226
rect 3806 256 3809 257
rect 4150 256 4153 257
rect 3806 226 3936 256
rect 4022 226 4153 256
rect 3806 225 3809 226
rect 4150 225 4153 226
rect 4185 256 4188 257
rect 4529 256 4532 257
rect 4185 226 4315 256
rect 4401 226 4532 256
rect 4185 225 4188 226
rect 4529 225 4532 226
rect 4564 256 4567 257
rect 4908 256 4911 257
rect 4564 226 4694 256
rect 4780 226 4911 256
rect 4564 225 4567 226
rect 4908 225 4911 226
rect 4943 256 4946 257
rect 5287 256 5290 257
rect 4943 226 5073 256
rect 5159 226 5290 256
rect 4943 225 4946 226
rect 5287 225 5290 226
rect 5322 256 5325 257
rect 5666 256 5669 257
rect 5322 226 5452 256
rect 5538 226 5669 256
rect 5322 225 5325 226
rect 5666 225 5669 226
rect 5701 256 5704 257
rect 6045 256 6048 257
rect 5701 226 5831 256
rect 5917 226 6048 256
rect 5701 225 5704 226
rect 6045 225 6048 226
rect 6080 256 6083 257
rect 6424 256 6427 257
rect 6080 226 6210 256
rect 6296 226 6427 256
rect 6080 225 6083 226
rect 6424 225 6427 226
rect 6459 256 6462 257
rect 6803 256 6806 257
rect 6459 226 6589 256
rect 6675 226 6806 256
rect 6459 225 6462 226
rect 6803 225 6806 226
rect 6838 256 6841 257
rect 7182 256 7185 257
rect 6838 226 6968 256
rect 7054 226 7185 256
rect 6838 225 6841 226
rect 7182 225 7185 226
rect 7217 256 7220 257
rect 7561 256 7564 257
rect 7217 226 7347 256
rect 7433 226 7564 256
rect 7217 225 7220 226
rect 7561 225 7564 226
rect 7596 225 7599 257
rect 161 197 217 200
rect 161 196 166 197
rect 53 166 166 196
rect 212 196 217 197
rect 540 197 596 200
rect 540 196 545 197
rect 212 166 326 196
rect 432 166 545 196
rect 591 196 596 197
rect 919 197 975 200
rect 919 196 924 197
rect 591 166 705 196
rect 811 166 924 196
rect 970 196 975 197
rect 1298 197 1354 200
rect 1298 196 1303 197
rect 970 166 1084 196
rect 1190 166 1303 196
rect 1349 196 1354 197
rect 1677 197 1733 200
rect 1677 196 1682 197
rect 1349 166 1463 196
rect 1569 166 1682 196
rect 1728 196 1733 197
rect 2056 197 2112 200
rect 2056 196 2061 197
rect 1728 166 1842 196
rect 1948 166 2061 196
rect 2107 196 2112 197
rect 2435 197 2491 200
rect 2435 196 2440 197
rect 2107 166 2221 196
rect 2327 166 2440 196
rect 2486 196 2491 197
rect 2814 197 2870 200
rect 2814 196 2819 197
rect 2486 166 2600 196
rect 2706 166 2819 196
rect 2865 196 2870 197
rect 3193 197 3249 200
rect 3193 196 3198 197
rect 2865 166 2979 196
rect 3085 166 3198 196
rect 3244 196 3249 197
rect 3572 197 3628 200
rect 3572 196 3577 197
rect 3244 166 3358 196
rect 3464 166 3577 196
rect 3623 196 3628 197
rect 3951 197 4007 200
rect 3951 196 3956 197
rect 3623 166 3737 196
rect 3843 166 3956 196
rect 4002 196 4007 197
rect 4330 197 4386 200
rect 4330 196 4335 197
rect 4002 166 4116 196
rect 4222 166 4335 196
rect 4381 196 4386 197
rect 4709 197 4765 200
rect 4709 196 4714 197
rect 4381 166 4495 196
rect 4601 166 4714 196
rect 4760 196 4765 197
rect 5088 197 5144 200
rect 5088 196 5093 197
rect 4760 166 4874 196
rect 4980 166 5093 196
rect 5139 196 5144 197
rect 5467 197 5523 200
rect 5467 196 5472 197
rect 5139 166 5253 196
rect 5359 166 5472 196
rect 5518 196 5523 197
rect 5846 197 5902 200
rect 5846 196 5851 197
rect 5518 166 5632 196
rect 5738 166 5851 196
rect 5897 196 5902 197
rect 6225 197 6281 200
rect 6225 196 6230 197
rect 5897 166 6011 196
rect 6117 166 6230 196
rect 6276 196 6281 197
rect 6604 197 6660 200
rect 6604 196 6609 197
rect 6276 166 6390 196
rect 6496 166 6609 196
rect 6655 196 6660 197
rect 6983 197 7039 200
rect 6983 196 6988 197
rect 6655 166 6769 196
rect 6875 166 6988 196
rect 7034 196 7039 197
rect 7362 197 7418 200
rect 7362 196 7367 197
rect 7034 166 7148 196
rect 7254 166 7367 196
rect 7413 196 7418 197
rect 7413 166 7527 196
rect 161 162 217 166
rect 540 162 596 166
rect 919 162 975 166
rect 1298 162 1354 166
rect 1677 162 1733 166
rect 2056 162 2112 166
rect 2435 162 2491 166
rect 2814 162 2870 166
rect 3193 162 3249 166
rect 3572 162 3628 166
rect 3951 162 4007 166
rect 4330 162 4386 166
rect 4709 162 4765 166
rect 5088 162 5144 166
rect 5467 162 5523 166
rect 5846 162 5902 166
rect 6225 162 6281 166
rect 6604 162 6660 166
rect 6983 162 7039 166
rect 7362 162 7418 166
rect -19 105 -16 137
rect 16 136 19 137
rect 360 136 363 137
rect 16 106 146 136
rect 232 106 363 136
rect 16 105 19 106
rect 360 105 363 106
rect 395 136 398 137
rect 739 136 742 137
rect 395 106 525 136
rect 611 106 742 136
rect 395 105 398 106
rect 739 105 742 106
rect 774 136 777 137
rect 1118 136 1121 137
rect 774 106 904 136
rect 990 106 1121 136
rect 774 105 777 106
rect 1118 105 1121 106
rect 1153 136 1156 137
rect 1497 136 1500 137
rect 1153 106 1283 136
rect 1369 106 1500 136
rect 1153 105 1156 106
rect 1497 105 1500 106
rect 1532 136 1535 137
rect 1876 136 1879 137
rect 1532 106 1662 136
rect 1748 106 1879 136
rect 1532 105 1535 106
rect 1876 105 1879 106
rect 1911 136 1914 137
rect 2255 136 2258 137
rect 1911 106 2041 136
rect 2127 106 2258 136
rect 1911 105 1914 106
rect 2255 105 2258 106
rect 2290 136 2293 137
rect 2634 136 2637 137
rect 2290 106 2420 136
rect 2506 106 2637 136
rect 2290 105 2293 106
rect 2634 105 2637 106
rect 2669 136 2672 137
rect 3013 136 3016 137
rect 2669 106 2799 136
rect 2885 106 3016 136
rect 2669 105 2672 106
rect 3013 105 3016 106
rect 3048 136 3051 137
rect 3392 136 3395 137
rect 3048 106 3178 136
rect 3264 106 3395 136
rect 3048 105 3051 106
rect 3392 105 3395 106
rect 3427 136 3430 137
rect 3771 136 3774 137
rect 3427 106 3557 136
rect 3643 106 3774 136
rect 3427 105 3430 106
rect 3771 105 3774 106
rect 3806 136 3809 137
rect 4150 136 4153 137
rect 3806 106 3936 136
rect 4022 106 4153 136
rect 3806 105 3809 106
rect 4150 105 4153 106
rect 4185 136 4188 137
rect 4529 136 4532 137
rect 4185 106 4315 136
rect 4401 106 4532 136
rect 4185 105 4188 106
rect 4529 105 4532 106
rect 4564 136 4567 137
rect 4908 136 4911 137
rect 4564 106 4694 136
rect 4780 106 4911 136
rect 4564 105 4567 106
rect 4908 105 4911 106
rect 4943 136 4946 137
rect 5287 136 5290 137
rect 4943 106 5073 136
rect 5159 106 5290 136
rect 4943 105 4946 106
rect 5287 105 5290 106
rect 5322 136 5325 137
rect 5666 136 5669 137
rect 5322 106 5452 136
rect 5538 106 5669 136
rect 5322 105 5325 106
rect 5666 105 5669 106
rect 5701 136 5704 137
rect 6045 136 6048 137
rect 5701 106 5831 136
rect 5917 106 6048 136
rect 5701 105 5704 106
rect 6045 105 6048 106
rect 6080 136 6083 137
rect 6424 136 6427 137
rect 6080 106 6210 136
rect 6296 106 6427 136
rect 6080 105 6083 106
rect 6424 105 6427 106
rect 6459 136 6462 137
rect 6803 136 6806 137
rect 6459 106 6589 136
rect 6675 106 6806 136
rect 6459 105 6462 106
rect 6803 105 6806 106
rect 6838 136 6841 137
rect 7182 136 7185 137
rect 6838 106 6968 136
rect 7054 106 7185 136
rect 6838 105 6841 106
rect 7182 105 7185 106
rect 7217 136 7220 137
rect 7561 136 7564 137
rect 7217 106 7347 136
rect 7433 106 7564 136
rect 7217 105 7220 106
rect 7561 105 7564 106
rect 7596 105 7599 137
rect 161 77 217 80
rect 161 76 166 77
rect 53 46 166 76
rect 212 76 217 77
rect 540 77 596 80
rect 540 76 545 77
rect 212 46 326 76
rect 432 46 545 76
rect 591 76 596 77
rect 919 77 975 80
rect 919 76 924 77
rect 591 46 705 76
rect 811 46 924 76
rect 970 76 975 77
rect 1298 77 1354 80
rect 1298 76 1303 77
rect 970 46 1084 76
rect 1190 46 1303 76
rect 1349 76 1354 77
rect 1677 77 1733 80
rect 1677 76 1682 77
rect 1349 46 1463 76
rect 1569 46 1682 76
rect 1728 76 1733 77
rect 2056 77 2112 80
rect 2056 76 2061 77
rect 1728 46 1842 76
rect 1948 46 2061 76
rect 2107 76 2112 77
rect 2435 77 2491 80
rect 2435 76 2440 77
rect 2107 46 2221 76
rect 2327 46 2440 76
rect 2486 76 2491 77
rect 2814 77 2870 80
rect 2814 76 2819 77
rect 2486 46 2600 76
rect 2706 46 2819 76
rect 2865 76 2870 77
rect 3193 77 3249 80
rect 3193 76 3198 77
rect 2865 46 2979 76
rect 3085 46 3198 76
rect 3244 76 3249 77
rect 3572 77 3628 80
rect 3572 76 3577 77
rect 3244 46 3358 76
rect 3464 46 3577 76
rect 3623 76 3628 77
rect 3951 77 4007 80
rect 3951 76 3956 77
rect 3623 46 3737 76
rect 3843 46 3956 76
rect 4002 76 4007 77
rect 4330 77 4386 80
rect 4330 76 4335 77
rect 4002 46 4116 76
rect 4222 46 4335 76
rect 4381 76 4386 77
rect 4709 77 4765 80
rect 4709 76 4714 77
rect 4381 46 4495 76
rect 4601 46 4714 76
rect 4760 76 4765 77
rect 5088 77 5144 80
rect 5088 76 5093 77
rect 4760 46 4874 76
rect 4980 46 5093 76
rect 5139 76 5144 77
rect 5467 77 5523 80
rect 5467 76 5472 77
rect 5139 46 5253 76
rect 5359 46 5472 76
rect 5518 76 5523 77
rect 5846 77 5902 80
rect 5846 76 5851 77
rect 5518 46 5632 76
rect 5738 46 5851 76
rect 5897 76 5902 77
rect 6225 77 6281 80
rect 6225 76 6230 77
rect 5897 46 6011 76
rect 6117 46 6230 76
rect 6276 76 6281 77
rect 6604 77 6660 80
rect 6604 76 6609 77
rect 6276 46 6390 76
rect 6496 46 6609 76
rect 6655 76 6660 77
rect 6983 77 7039 80
rect 6983 76 6988 77
rect 6655 46 6769 76
rect 6875 46 6988 76
rect 7034 76 7039 77
rect 7362 77 7418 80
rect 7362 76 7367 77
rect 7034 46 7148 76
rect 7254 46 7367 76
rect 7413 76 7418 77
rect 7413 46 7527 76
rect 161 42 217 46
rect 540 42 596 46
rect 919 42 975 46
rect 1298 42 1354 46
rect 1677 42 1733 46
rect 2056 42 2112 46
rect 2435 42 2491 46
rect 2814 42 2870 46
rect 3193 42 3249 46
rect 3572 42 3628 46
rect 3951 42 4007 46
rect 4330 42 4386 46
rect 4709 42 4765 46
rect 5088 42 5144 46
rect 5467 42 5523 46
rect 5846 42 5902 46
rect 6225 42 6281 46
rect 6604 42 6660 46
rect 6983 42 7039 46
rect 7362 42 7418 46
<< via3 >>
rect -16 2274 16 2306
rect 363 2274 395 2306
rect 742 2274 774 2306
rect 1121 2274 1153 2306
rect 1500 2274 1532 2306
rect 1879 2274 1911 2306
rect 2258 2274 2290 2306
rect 2637 2274 2669 2306
rect 3016 2274 3048 2306
rect 3395 2274 3427 2306
rect 3774 2274 3806 2306
rect 4153 2274 4185 2306
rect 4532 2274 4564 2306
rect 4911 2274 4943 2306
rect 5290 2274 5322 2306
rect 5669 2274 5701 2306
rect 6048 2274 6080 2306
rect 6427 2274 6459 2306
rect 6806 2274 6838 2306
rect 7185 2274 7217 2306
rect 7564 2274 7596 2306
rect -16 2154 16 2186
rect 363 2154 395 2186
rect 742 2154 774 2186
rect 1121 2154 1153 2186
rect 1500 2154 1532 2186
rect 1879 2154 1911 2186
rect 2258 2154 2290 2186
rect 2637 2154 2669 2186
rect 3016 2154 3048 2186
rect 3395 2154 3427 2186
rect 3774 2154 3806 2186
rect 4153 2154 4185 2186
rect 4532 2154 4564 2186
rect 4911 2154 4943 2186
rect 5290 2154 5322 2186
rect 5669 2154 5701 2186
rect 6048 2154 6080 2186
rect 6427 2154 6459 2186
rect 6806 2154 6838 2186
rect 7185 2154 7217 2186
rect 7564 2154 7596 2186
rect -16 2034 16 2066
rect 363 2034 395 2066
rect 742 2034 774 2066
rect 1121 2034 1153 2066
rect 1500 2034 1532 2066
rect 1879 2034 1911 2066
rect 2258 2034 2290 2066
rect 2637 2034 2669 2066
rect 3016 2034 3048 2066
rect 3395 2034 3427 2066
rect 3774 2034 3806 2066
rect 4153 2034 4185 2066
rect 4532 2034 4564 2066
rect 4911 2034 4943 2066
rect 5290 2034 5322 2066
rect 5669 2034 5701 2066
rect 6048 2034 6080 2066
rect 6427 2034 6459 2066
rect 6806 2034 6838 2066
rect 7185 2034 7217 2066
rect 7564 2034 7596 2066
rect -16 1914 16 1946
rect 363 1914 395 1946
rect 742 1914 774 1946
rect 1121 1914 1153 1946
rect 1500 1914 1532 1946
rect 1879 1914 1911 1946
rect 2258 1914 2290 1946
rect 2637 1914 2669 1946
rect 3016 1914 3048 1946
rect 3395 1914 3427 1946
rect 3774 1914 3806 1946
rect 4153 1914 4185 1946
rect 4532 1914 4564 1946
rect 4911 1914 4943 1946
rect 5290 1914 5322 1946
rect 5669 1914 5701 1946
rect 6048 1914 6080 1946
rect 6427 1914 6459 1946
rect 6806 1914 6838 1946
rect 7185 1914 7217 1946
rect 7564 1914 7596 1946
rect -16 1671 16 1703
rect 363 1671 395 1703
rect 742 1671 774 1703
rect 1121 1671 1153 1703
rect 1500 1671 1532 1703
rect 1879 1671 1911 1703
rect 2258 1671 2290 1703
rect 2637 1671 2669 1703
rect 3016 1671 3048 1703
rect 3395 1671 3427 1703
rect 3774 1671 3806 1703
rect 4153 1671 4185 1703
rect 4532 1671 4564 1703
rect 4911 1671 4943 1703
rect 5290 1671 5322 1703
rect 5669 1671 5701 1703
rect 6048 1671 6080 1703
rect 6427 1671 6459 1703
rect 6806 1671 6838 1703
rect 7185 1671 7217 1703
rect 7564 1671 7596 1703
rect -16 1551 16 1583
rect 363 1551 395 1583
rect 742 1551 774 1583
rect 1121 1551 1153 1583
rect 1500 1551 1532 1583
rect 1879 1551 1911 1583
rect 2258 1551 2290 1583
rect 2637 1551 2669 1583
rect 3016 1551 3048 1583
rect 3395 1551 3427 1583
rect 3774 1551 3806 1583
rect 4153 1551 4185 1583
rect 4532 1551 4564 1583
rect 4911 1551 4943 1583
rect 5290 1551 5322 1583
rect 5669 1551 5701 1583
rect 6048 1551 6080 1583
rect 6427 1551 6459 1583
rect 6806 1551 6838 1583
rect 7185 1551 7217 1583
rect 7564 1551 7596 1583
rect -16 1431 16 1463
rect 363 1431 395 1463
rect 742 1431 774 1463
rect 1121 1431 1153 1463
rect 1500 1431 1532 1463
rect 1879 1431 1911 1463
rect 2258 1431 2290 1463
rect 2637 1431 2669 1463
rect 3016 1431 3048 1463
rect 3395 1431 3427 1463
rect 3774 1431 3806 1463
rect 4153 1431 4185 1463
rect 4532 1431 4564 1463
rect 4911 1431 4943 1463
rect 5290 1431 5322 1463
rect 5669 1431 5701 1463
rect 6048 1431 6080 1463
rect 6427 1431 6459 1463
rect 6806 1431 6838 1463
rect 7185 1431 7217 1463
rect 7564 1431 7596 1463
rect -16 1311 16 1343
rect 363 1311 395 1343
rect 742 1311 774 1343
rect 1121 1311 1153 1343
rect 1500 1311 1532 1343
rect 1879 1311 1911 1343
rect 2258 1311 2290 1343
rect 2637 1311 2669 1343
rect 3016 1311 3048 1343
rect 3395 1311 3427 1343
rect 3774 1311 3806 1343
rect 4153 1311 4185 1343
rect 4532 1311 4564 1343
rect 4911 1311 4943 1343
rect 5290 1311 5322 1343
rect 5669 1311 5701 1343
rect 6048 1311 6080 1343
rect 6427 1311 6459 1343
rect 6806 1311 6838 1343
rect 7185 1311 7217 1343
rect 7564 1311 7596 1343
rect -16 1068 16 1100
rect 363 1068 395 1100
rect 742 1068 774 1100
rect 1121 1068 1153 1100
rect 1500 1068 1532 1100
rect 1879 1068 1911 1100
rect 2258 1068 2290 1100
rect 2637 1068 2669 1100
rect 3016 1068 3048 1100
rect 3395 1068 3427 1100
rect 3774 1068 3806 1100
rect 4153 1068 4185 1100
rect 4532 1068 4564 1100
rect 4911 1068 4943 1100
rect 5290 1068 5322 1100
rect 5669 1068 5701 1100
rect 6048 1068 6080 1100
rect 6427 1068 6459 1100
rect 6806 1068 6838 1100
rect 7185 1068 7217 1100
rect 7564 1068 7596 1100
rect -16 948 16 980
rect 363 948 395 980
rect 742 948 774 980
rect 1121 948 1153 980
rect 1500 948 1532 980
rect 1879 948 1911 980
rect 2258 948 2290 980
rect 2637 948 2669 980
rect 3016 948 3048 980
rect 3395 948 3427 980
rect 3774 948 3806 980
rect 4153 948 4185 980
rect 4532 948 4564 980
rect 4911 948 4943 980
rect 5290 948 5322 980
rect 5669 948 5701 980
rect 6048 948 6080 980
rect 6427 948 6459 980
rect 6806 948 6838 980
rect 7185 948 7217 980
rect 7564 948 7596 980
rect -16 828 16 860
rect 363 828 395 860
rect 742 828 774 860
rect 1121 828 1153 860
rect 1500 828 1532 860
rect 1879 828 1911 860
rect 2258 828 2290 860
rect 2637 828 2669 860
rect 3016 828 3048 860
rect 3395 828 3427 860
rect 3774 828 3806 860
rect 4153 828 4185 860
rect 4532 828 4564 860
rect 4911 828 4943 860
rect 5290 828 5322 860
rect 5669 828 5701 860
rect 6048 828 6080 860
rect 6427 828 6459 860
rect 6806 828 6838 860
rect 7185 828 7217 860
rect 7564 828 7596 860
rect -16 708 16 740
rect 363 708 395 740
rect 742 708 774 740
rect 1121 708 1153 740
rect 1500 708 1532 740
rect 1879 708 1911 740
rect 2258 708 2290 740
rect 2637 708 2669 740
rect 3016 708 3048 740
rect 3395 708 3427 740
rect 3774 708 3806 740
rect 4153 708 4185 740
rect 4532 708 4564 740
rect 4911 708 4943 740
rect 5290 708 5322 740
rect 5669 708 5701 740
rect 6048 708 6080 740
rect 6427 708 6459 740
rect 6806 708 6838 740
rect 7185 708 7217 740
rect 7564 708 7596 740
rect -16 465 16 497
rect 363 465 395 497
rect 742 465 774 497
rect 1121 465 1153 497
rect 1500 465 1532 497
rect 1879 465 1911 497
rect 2258 465 2290 497
rect 2637 465 2669 497
rect 3016 465 3048 497
rect 3395 465 3427 497
rect 3774 465 3806 497
rect 4153 465 4185 497
rect 4532 465 4564 497
rect 4911 465 4943 497
rect 5290 465 5322 497
rect 5669 465 5701 497
rect 6048 465 6080 497
rect 6427 465 6459 497
rect 6806 465 6838 497
rect 7185 465 7217 497
rect 7564 465 7596 497
rect -16 345 16 377
rect 363 345 395 377
rect 742 345 774 377
rect 1121 345 1153 377
rect 1500 345 1532 377
rect 1879 345 1911 377
rect 2258 345 2290 377
rect 2637 345 2669 377
rect 3016 345 3048 377
rect 3395 345 3427 377
rect 3774 345 3806 377
rect 4153 345 4185 377
rect 4532 345 4564 377
rect 4911 345 4943 377
rect 5290 345 5322 377
rect 5669 345 5701 377
rect 6048 345 6080 377
rect 6427 345 6459 377
rect 6806 345 6838 377
rect 7185 345 7217 377
rect 7564 345 7596 377
rect -16 225 16 257
rect 363 225 395 257
rect 742 225 774 257
rect 1121 225 1153 257
rect 1500 225 1532 257
rect 1879 225 1911 257
rect 2258 225 2290 257
rect 2637 225 2669 257
rect 3016 225 3048 257
rect 3395 225 3427 257
rect 3774 225 3806 257
rect 4153 225 4185 257
rect 4532 225 4564 257
rect 4911 225 4943 257
rect 5290 225 5322 257
rect 5669 225 5701 257
rect 6048 225 6080 257
rect 6427 225 6459 257
rect 6806 225 6838 257
rect 7185 225 7217 257
rect 7564 225 7596 257
rect -16 105 16 137
rect 363 105 395 137
rect 742 105 774 137
rect 1121 105 1153 137
rect 1500 105 1532 137
rect 1879 105 1911 137
rect 2258 105 2290 137
rect 2637 105 2669 137
rect 3016 105 3048 137
rect 3395 105 3427 137
rect 3774 105 3806 137
rect 4153 105 4185 137
rect 4532 105 4564 137
rect 4911 105 4943 137
rect 5290 105 5322 137
rect 5669 105 5701 137
rect 6048 105 6080 137
rect 6427 105 6459 137
rect 6806 105 6838 137
rect 7185 105 7217 137
rect 7564 105 7596 137
<< metal4 >>
rect -19 2396 7599 2428
rect -19 2306 19 2396
rect -19 2274 -16 2306
rect 16 2274 19 2306
rect -19 2186 19 2274
rect -19 2154 -16 2186
rect 16 2154 19 2186
rect -19 2066 19 2154
rect -19 2034 -16 2066
rect 16 2034 19 2066
rect -19 1946 19 2034
rect -19 1914 -16 1946
rect 16 1914 19 1946
rect -19 1825 19 1914
rect 360 2306 398 2396
rect 360 2274 363 2306
rect 395 2274 398 2306
rect 360 2186 398 2274
rect 360 2154 363 2186
rect 395 2154 398 2186
rect 360 2066 398 2154
rect 360 2034 363 2066
rect 395 2034 398 2066
rect 360 1946 398 2034
rect 360 1914 363 1946
rect 395 1914 398 1946
rect 360 1867 398 1914
rect 739 2306 777 2396
rect 739 2274 742 2306
rect 774 2274 777 2306
rect 739 2186 777 2274
rect 739 2154 742 2186
rect 774 2154 777 2186
rect 739 2066 777 2154
rect 739 2034 742 2066
rect 774 2034 777 2066
rect 739 1946 777 2034
rect 739 1914 742 1946
rect 774 1914 777 1946
rect 739 1867 777 1914
rect 1118 2306 1156 2396
rect 1118 2274 1121 2306
rect 1153 2274 1156 2306
rect 1118 2186 1156 2274
rect 1118 2154 1121 2186
rect 1153 2154 1156 2186
rect 1118 2066 1156 2154
rect 1118 2034 1121 2066
rect 1153 2034 1156 2066
rect 1118 1946 1156 2034
rect 1118 1914 1121 1946
rect 1153 1914 1156 1946
rect 1118 1867 1156 1914
rect 1497 2306 1535 2396
rect 1497 2274 1500 2306
rect 1532 2274 1535 2306
rect 1497 2186 1535 2274
rect 1497 2154 1500 2186
rect 1532 2154 1535 2186
rect 1497 2066 1535 2154
rect 1497 2034 1500 2066
rect 1532 2034 1535 2066
rect 1497 1946 1535 2034
rect 1497 1914 1500 1946
rect 1532 1914 1535 1946
rect 1497 1867 1535 1914
rect 1876 2306 1914 2396
rect 1876 2274 1879 2306
rect 1911 2274 1914 2306
rect 1876 2186 1914 2274
rect 1876 2154 1879 2186
rect 1911 2154 1914 2186
rect 1876 2066 1914 2154
rect 1876 2034 1879 2066
rect 1911 2034 1914 2066
rect 1876 1946 1914 2034
rect 1876 1914 1879 1946
rect 1911 1914 1914 1946
rect 1876 1825 1914 1914
rect 2255 2306 2293 2396
rect 2255 2274 2258 2306
rect 2290 2274 2293 2306
rect 2255 2186 2293 2274
rect 2255 2154 2258 2186
rect 2290 2154 2293 2186
rect 2255 2066 2293 2154
rect 2255 2034 2258 2066
rect 2290 2034 2293 2066
rect 2255 1946 2293 2034
rect 2255 1914 2258 1946
rect 2290 1914 2293 1946
rect 2255 1867 2293 1914
rect 2634 2306 2672 2396
rect 2634 2274 2637 2306
rect 2669 2274 2672 2306
rect 2634 2186 2672 2274
rect 2634 2154 2637 2186
rect 2669 2154 2672 2186
rect 2634 2066 2672 2154
rect 2634 2034 2637 2066
rect 2669 2034 2672 2066
rect 2634 1946 2672 2034
rect 2634 1914 2637 1946
rect 2669 1914 2672 1946
rect 2634 1867 2672 1914
rect 3013 2306 3051 2396
rect 3013 2274 3016 2306
rect 3048 2274 3051 2306
rect 3013 2186 3051 2274
rect 3013 2154 3016 2186
rect 3048 2154 3051 2186
rect 3013 2066 3051 2154
rect 3013 2034 3016 2066
rect 3048 2034 3051 2066
rect 3013 1946 3051 2034
rect 3013 1914 3016 1946
rect 3048 1914 3051 1946
rect 3013 1867 3051 1914
rect 3392 2306 3430 2396
rect 3392 2274 3395 2306
rect 3427 2274 3430 2306
rect 3392 2186 3430 2274
rect 3392 2154 3395 2186
rect 3427 2154 3430 2186
rect 3392 2066 3430 2154
rect 3392 2034 3395 2066
rect 3427 2034 3430 2066
rect 3392 1946 3430 2034
rect 3392 1914 3395 1946
rect 3427 1914 3430 1946
rect 3392 1867 3430 1914
rect 3771 2306 3809 2396
rect 3771 2274 3774 2306
rect 3806 2274 3809 2306
rect 3771 2186 3809 2274
rect 3771 2154 3774 2186
rect 3806 2154 3809 2186
rect 3771 2066 3809 2154
rect 3771 2034 3774 2066
rect 3806 2034 3809 2066
rect 3771 1946 3809 2034
rect 3771 1914 3774 1946
rect 3806 1914 3809 1946
rect 3771 1825 3809 1914
rect 4150 2306 4188 2396
rect 4150 2274 4153 2306
rect 4185 2274 4188 2306
rect 4150 2186 4188 2274
rect 4150 2154 4153 2186
rect 4185 2154 4188 2186
rect 4150 2066 4188 2154
rect 4150 2034 4153 2066
rect 4185 2034 4188 2066
rect 4150 1946 4188 2034
rect 4150 1914 4153 1946
rect 4185 1914 4188 1946
rect 4150 1867 4188 1914
rect 4529 2306 4567 2396
rect 4529 2274 4532 2306
rect 4564 2274 4567 2306
rect 4529 2186 4567 2274
rect 4529 2154 4532 2186
rect 4564 2154 4567 2186
rect 4529 2066 4567 2154
rect 4529 2034 4532 2066
rect 4564 2034 4567 2066
rect 4529 1946 4567 2034
rect 4529 1914 4532 1946
rect 4564 1914 4567 1946
rect 4529 1867 4567 1914
rect 4908 2306 4946 2396
rect 4908 2274 4911 2306
rect 4943 2274 4946 2306
rect 4908 2186 4946 2274
rect 4908 2154 4911 2186
rect 4943 2154 4946 2186
rect 4908 2066 4946 2154
rect 4908 2034 4911 2066
rect 4943 2034 4946 2066
rect 4908 1946 4946 2034
rect 4908 1914 4911 1946
rect 4943 1914 4946 1946
rect 4908 1867 4946 1914
rect 5287 2306 5325 2396
rect 5287 2274 5290 2306
rect 5322 2274 5325 2306
rect 5287 2186 5325 2274
rect 5287 2154 5290 2186
rect 5322 2154 5325 2186
rect 5287 2066 5325 2154
rect 5287 2034 5290 2066
rect 5322 2034 5325 2066
rect 5287 1946 5325 2034
rect 5287 1914 5290 1946
rect 5322 1914 5325 1946
rect 5287 1867 5325 1914
rect 5666 2306 5704 2396
rect 5666 2274 5669 2306
rect 5701 2274 5704 2306
rect 5666 2186 5704 2274
rect 5666 2154 5669 2186
rect 5701 2154 5704 2186
rect 5666 2066 5704 2154
rect 5666 2034 5669 2066
rect 5701 2034 5704 2066
rect 5666 1946 5704 2034
rect 5666 1914 5669 1946
rect 5701 1914 5704 1946
rect 5666 1825 5704 1914
rect 6045 2306 6083 2396
rect 6045 2274 6048 2306
rect 6080 2274 6083 2306
rect 6045 2186 6083 2274
rect 6045 2154 6048 2186
rect 6080 2154 6083 2186
rect 6045 2066 6083 2154
rect 6045 2034 6048 2066
rect 6080 2034 6083 2066
rect 6045 1946 6083 2034
rect 6045 1914 6048 1946
rect 6080 1914 6083 1946
rect 6045 1867 6083 1914
rect 6424 2306 6462 2396
rect 6424 2274 6427 2306
rect 6459 2274 6462 2306
rect 6424 2186 6462 2274
rect 6424 2154 6427 2186
rect 6459 2154 6462 2186
rect 6424 2066 6462 2154
rect 6424 2034 6427 2066
rect 6459 2034 6462 2066
rect 6424 1946 6462 2034
rect 6424 1914 6427 1946
rect 6459 1914 6462 1946
rect 6424 1867 6462 1914
rect 6803 2306 6841 2396
rect 6803 2274 6806 2306
rect 6838 2274 6841 2306
rect 6803 2186 6841 2274
rect 6803 2154 6806 2186
rect 6838 2154 6841 2186
rect 6803 2066 6841 2154
rect 6803 2034 6806 2066
rect 6838 2034 6841 2066
rect 6803 1946 6841 2034
rect 6803 1914 6806 1946
rect 6838 1914 6841 1946
rect 6803 1867 6841 1914
rect 7182 2306 7220 2396
rect 7182 2274 7185 2306
rect 7217 2274 7220 2306
rect 7182 2186 7220 2274
rect 7182 2154 7185 2186
rect 7217 2154 7220 2186
rect 7182 2066 7220 2154
rect 7182 2034 7185 2066
rect 7217 2034 7220 2066
rect 7182 1946 7220 2034
rect 7182 1914 7185 1946
rect 7217 1914 7220 1946
rect 7182 1867 7220 1914
rect 7561 2306 7599 2396
rect 7561 2274 7564 2306
rect 7596 2274 7599 2306
rect 7561 2186 7599 2274
rect 7561 2154 7564 2186
rect 7596 2154 7599 2186
rect 7561 2066 7599 2154
rect 7561 2034 7564 2066
rect 7596 2034 7599 2066
rect 7561 1946 7599 2034
rect 7561 1914 7564 1946
rect 7596 1914 7599 1946
rect 7561 1825 7599 1914
rect -19 1793 318 1825
rect 360 1793 1535 1825
rect 1577 1793 2213 1825
rect 2255 1793 3430 1825
rect 3472 1793 4108 1825
rect 4150 1793 5325 1825
rect 5367 1793 6003 1825
rect 6045 1793 7220 1825
rect 7262 1793 7599 1825
rect -19 1703 19 1793
rect -19 1671 -16 1703
rect 16 1671 19 1703
rect -19 1583 19 1671
rect -19 1551 -16 1583
rect 16 1551 19 1583
rect -19 1463 19 1551
rect -19 1431 -16 1463
rect 16 1431 19 1463
rect -19 1343 19 1431
rect -19 1311 -16 1343
rect 16 1311 19 1343
rect -19 1222 19 1311
rect 360 1703 398 1793
rect 360 1671 363 1703
rect 395 1671 398 1703
rect 360 1583 398 1671
rect 360 1551 363 1583
rect 395 1551 398 1583
rect 360 1463 398 1551
rect 360 1431 363 1463
rect 395 1431 398 1463
rect 360 1343 398 1431
rect 360 1311 363 1343
rect 395 1311 398 1343
rect 360 1222 398 1311
rect 739 1703 777 1793
rect 739 1671 742 1703
rect 774 1671 777 1703
rect 739 1583 777 1671
rect 739 1551 742 1583
rect 774 1551 777 1583
rect 739 1463 777 1551
rect 739 1431 742 1463
rect 774 1431 777 1463
rect 739 1343 777 1431
rect 739 1311 742 1343
rect 774 1311 777 1343
rect 739 1222 777 1311
rect 1118 1703 1156 1793
rect 1118 1671 1121 1703
rect 1153 1671 1156 1703
rect 1118 1583 1156 1671
rect 1118 1551 1121 1583
rect 1153 1551 1156 1583
rect 1118 1463 1156 1551
rect 1118 1431 1121 1463
rect 1153 1431 1156 1463
rect 1118 1343 1156 1431
rect 1118 1311 1121 1343
rect 1153 1311 1156 1343
rect 1118 1222 1156 1311
rect 1497 1703 1535 1793
rect 1497 1671 1500 1703
rect 1532 1671 1535 1703
rect 1497 1583 1535 1671
rect 1497 1551 1500 1583
rect 1532 1551 1535 1583
rect 1497 1463 1535 1551
rect 1497 1431 1500 1463
rect 1532 1431 1535 1463
rect 1497 1343 1535 1431
rect 1497 1311 1500 1343
rect 1532 1311 1535 1343
rect 1497 1222 1535 1311
rect 1876 1703 1914 1793
rect 1876 1671 1879 1703
rect 1911 1671 1914 1703
rect 1876 1583 1914 1671
rect 1876 1551 1879 1583
rect 1911 1551 1914 1583
rect 1876 1463 1914 1551
rect 1876 1431 1879 1463
rect 1911 1431 1914 1463
rect 1876 1343 1914 1431
rect 1876 1311 1879 1343
rect 1911 1311 1914 1343
rect 1876 1222 1914 1311
rect 2255 1703 2293 1793
rect 2255 1671 2258 1703
rect 2290 1671 2293 1703
rect 2255 1583 2293 1671
rect 2255 1551 2258 1583
rect 2290 1551 2293 1583
rect 2255 1463 2293 1551
rect 2255 1431 2258 1463
rect 2290 1431 2293 1463
rect 2255 1343 2293 1431
rect 2255 1311 2258 1343
rect 2290 1311 2293 1343
rect 2255 1222 2293 1311
rect 2634 1703 2672 1793
rect 2634 1671 2637 1703
rect 2669 1671 2672 1703
rect 2634 1583 2672 1671
rect 2634 1551 2637 1583
rect 2669 1551 2672 1583
rect 2634 1463 2672 1551
rect 2634 1431 2637 1463
rect 2669 1431 2672 1463
rect 2634 1343 2672 1431
rect 2634 1311 2637 1343
rect 2669 1311 2672 1343
rect 2634 1222 2672 1311
rect 3013 1703 3051 1793
rect 3013 1671 3016 1703
rect 3048 1671 3051 1703
rect 3013 1583 3051 1671
rect 3013 1551 3016 1583
rect 3048 1551 3051 1583
rect 3013 1463 3051 1551
rect 3013 1431 3016 1463
rect 3048 1431 3051 1463
rect 3013 1343 3051 1431
rect 3013 1311 3016 1343
rect 3048 1311 3051 1343
rect 3013 1222 3051 1311
rect 3392 1703 3430 1793
rect 3392 1671 3395 1703
rect 3427 1671 3430 1703
rect 3392 1583 3430 1671
rect 3392 1551 3395 1583
rect 3427 1551 3430 1583
rect 3392 1463 3430 1551
rect 3392 1431 3395 1463
rect 3427 1431 3430 1463
rect 3392 1343 3430 1431
rect 3392 1311 3395 1343
rect 3427 1311 3430 1343
rect 3392 1222 3430 1311
rect 3771 1703 3809 1793
rect 3771 1671 3774 1703
rect 3806 1671 3809 1703
rect 3771 1583 3809 1671
rect 3771 1551 3774 1583
rect 3806 1551 3809 1583
rect 3771 1463 3809 1551
rect 3771 1431 3774 1463
rect 3806 1431 3809 1463
rect 3771 1343 3809 1431
rect 3771 1311 3774 1343
rect 3806 1311 3809 1343
rect 3771 1222 3809 1311
rect 4150 1703 4188 1793
rect 4150 1671 4153 1703
rect 4185 1671 4188 1703
rect 4150 1583 4188 1671
rect 4150 1551 4153 1583
rect 4185 1551 4188 1583
rect 4150 1463 4188 1551
rect 4150 1431 4153 1463
rect 4185 1431 4188 1463
rect 4150 1343 4188 1431
rect 4150 1311 4153 1343
rect 4185 1311 4188 1343
rect 4150 1222 4188 1311
rect 4529 1703 4567 1793
rect 4529 1671 4532 1703
rect 4564 1671 4567 1703
rect 4529 1583 4567 1671
rect 4529 1551 4532 1583
rect 4564 1551 4567 1583
rect 4529 1463 4567 1551
rect 4529 1431 4532 1463
rect 4564 1431 4567 1463
rect 4529 1343 4567 1431
rect 4529 1311 4532 1343
rect 4564 1311 4567 1343
rect 4529 1222 4567 1311
rect 4908 1703 4946 1793
rect 4908 1671 4911 1703
rect 4943 1671 4946 1703
rect 4908 1583 4946 1671
rect 4908 1551 4911 1583
rect 4943 1551 4946 1583
rect 4908 1463 4946 1551
rect 4908 1431 4911 1463
rect 4943 1431 4946 1463
rect 4908 1343 4946 1431
rect 4908 1311 4911 1343
rect 4943 1311 4946 1343
rect 4908 1222 4946 1311
rect 5287 1703 5325 1793
rect 5287 1671 5290 1703
rect 5322 1671 5325 1703
rect 5287 1583 5325 1671
rect 5287 1551 5290 1583
rect 5322 1551 5325 1583
rect 5287 1463 5325 1551
rect 5287 1431 5290 1463
rect 5322 1431 5325 1463
rect 5287 1343 5325 1431
rect 5287 1311 5290 1343
rect 5322 1311 5325 1343
rect 5287 1222 5325 1311
rect 5666 1703 5704 1793
rect 5666 1671 5669 1703
rect 5701 1671 5704 1703
rect 5666 1583 5704 1671
rect 5666 1551 5669 1583
rect 5701 1551 5704 1583
rect 5666 1463 5704 1551
rect 5666 1431 5669 1463
rect 5701 1431 5704 1463
rect 5666 1343 5704 1431
rect 5666 1311 5669 1343
rect 5701 1311 5704 1343
rect 5666 1222 5704 1311
rect 6045 1703 6083 1793
rect 6045 1671 6048 1703
rect 6080 1671 6083 1703
rect 6045 1583 6083 1671
rect 6045 1551 6048 1583
rect 6080 1551 6083 1583
rect 6045 1463 6083 1551
rect 6045 1431 6048 1463
rect 6080 1431 6083 1463
rect 6045 1343 6083 1431
rect 6045 1311 6048 1343
rect 6080 1311 6083 1343
rect 6045 1222 6083 1311
rect 6424 1703 6462 1793
rect 6424 1671 6427 1703
rect 6459 1671 6462 1703
rect 6424 1583 6462 1671
rect 6424 1551 6427 1583
rect 6459 1551 6462 1583
rect 6424 1463 6462 1551
rect 6424 1431 6427 1463
rect 6459 1431 6462 1463
rect 6424 1343 6462 1431
rect 6424 1311 6427 1343
rect 6459 1311 6462 1343
rect 6424 1222 6462 1311
rect 6803 1703 6841 1793
rect 6803 1671 6806 1703
rect 6838 1671 6841 1703
rect 6803 1583 6841 1671
rect 6803 1551 6806 1583
rect 6838 1551 6841 1583
rect 6803 1463 6841 1551
rect 6803 1431 6806 1463
rect 6838 1431 6841 1463
rect 6803 1343 6841 1431
rect 6803 1311 6806 1343
rect 6838 1311 6841 1343
rect 6803 1222 6841 1311
rect 7182 1703 7220 1793
rect 7182 1671 7185 1703
rect 7217 1671 7220 1703
rect 7182 1583 7220 1671
rect 7182 1551 7185 1583
rect 7217 1551 7220 1583
rect 7182 1463 7220 1551
rect 7182 1431 7185 1463
rect 7217 1431 7220 1463
rect 7182 1343 7220 1431
rect 7182 1311 7185 1343
rect 7217 1311 7220 1343
rect 7182 1222 7220 1311
rect 7561 1703 7599 1793
rect 7561 1671 7564 1703
rect 7596 1671 7599 1703
rect 7561 1583 7599 1671
rect 7561 1551 7564 1583
rect 7596 1551 7599 1583
rect 7561 1463 7599 1551
rect 7561 1431 7564 1463
rect 7596 1431 7599 1463
rect 7561 1343 7599 1431
rect 7561 1311 7564 1343
rect 7596 1311 7599 1343
rect -19 1190 318 1222
rect 360 1190 1535 1222
rect 1577 1190 1834 1222
rect 1876 1190 2213 1222
rect 2255 1190 3430 1222
rect 3472 1190 3729 1222
rect 3771 1190 4108 1222
rect 4150 1190 5325 1222
rect 5367 1190 5624 1222
rect 5666 1190 6003 1222
rect 6045 1190 7220 1222
rect 7262 1190 7519 1222
rect -19 1100 19 1190
rect -19 1068 -16 1100
rect 16 1068 19 1100
rect -19 980 19 1068
rect -19 948 -16 980
rect 16 948 19 980
rect -19 860 19 948
rect -19 828 -16 860
rect 16 828 19 860
rect -19 740 19 828
rect -19 708 -16 740
rect 16 708 19 740
rect -19 619 19 708
rect 360 1100 398 1190
rect 360 1068 363 1100
rect 395 1068 398 1100
rect 360 980 398 1068
rect 360 948 363 980
rect 395 948 398 980
rect 360 860 398 948
rect 360 828 363 860
rect 395 828 398 860
rect 360 740 398 828
rect 360 708 363 740
rect 395 708 398 740
rect 360 619 398 708
rect 739 1100 777 1190
rect 739 1068 742 1100
rect 774 1068 777 1100
rect 739 980 777 1068
rect 739 948 742 980
rect 774 948 777 980
rect 739 860 777 948
rect 739 828 742 860
rect 774 828 777 860
rect 739 740 777 828
rect 739 708 742 740
rect 774 708 777 740
rect 739 619 777 708
rect 1118 1100 1156 1190
rect 1118 1068 1121 1100
rect 1153 1068 1156 1100
rect 1118 980 1156 1068
rect 1118 948 1121 980
rect 1153 948 1156 980
rect 1118 860 1156 948
rect 1118 828 1121 860
rect 1153 828 1156 860
rect 1118 740 1156 828
rect 1118 708 1121 740
rect 1153 708 1156 740
rect 1118 619 1156 708
rect 1497 1100 1535 1190
rect 1497 1068 1500 1100
rect 1532 1068 1535 1100
rect 1497 980 1535 1068
rect 1497 948 1500 980
rect 1532 948 1535 980
rect 1497 860 1535 948
rect 1497 828 1500 860
rect 1532 828 1535 860
rect 1497 740 1535 828
rect 1497 708 1500 740
rect 1532 708 1535 740
rect 1497 619 1535 708
rect 1876 1100 1914 1190
rect 1876 1068 1879 1100
rect 1911 1068 1914 1100
rect 1876 980 1914 1068
rect 1876 948 1879 980
rect 1911 948 1914 980
rect 1876 860 1914 948
rect 1876 828 1879 860
rect 1911 828 1914 860
rect 1876 740 1914 828
rect 1876 708 1879 740
rect 1911 708 1914 740
rect 1876 619 1914 708
rect 2255 1100 2293 1190
rect 2255 1068 2258 1100
rect 2290 1068 2293 1100
rect 2255 980 2293 1068
rect 2255 948 2258 980
rect 2290 948 2293 980
rect 2255 860 2293 948
rect 2255 828 2258 860
rect 2290 828 2293 860
rect 2255 740 2293 828
rect 2255 708 2258 740
rect 2290 708 2293 740
rect 2255 619 2293 708
rect 2634 1100 2672 1190
rect 2634 1068 2637 1100
rect 2669 1068 2672 1100
rect 2634 980 2672 1068
rect 2634 948 2637 980
rect 2669 948 2672 980
rect 2634 860 2672 948
rect 2634 828 2637 860
rect 2669 828 2672 860
rect 2634 740 2672 828
rect 2634 708 2637 740
rect 2669 708 2672 740
rect 2634 619 2672 708
rect 3013 1100 3051 1190
rect 3013 1068 3016 1100
rect 3048 1068 3051 1100
rect 3013 980 3051 1068
rect 3013 948 3016 980
rect 3048 948 3051 980
rect 3013 860 3051 948
rect 3013 828 3016 860
rect 3048 828 3051 860
rect 3013 740 3051 828
rect 3013 708 3016 740
rect 3048 708 3051 740
rect 3013 619 3051 708
rect 3392 1100 3430 1190
rect 3392 1068 3395 1100
rect 3427 1068 3430 1100
rect 3392 980 3430 1068
rect 3392 948 3395 980
rect 3427 948 3430 980
rect 3392 860 3430 948
rect 3392 828 3395 860
rect 3427 828 3430 860
rect 3392 740 3430 828
rect 3392 708 3395 740
rect 3427 708 3430 740
rect 3392 619 3430 708
rect 3771 1100 3809 1190
rect 3771 1068 3774 1100
rect 3806 1068 3809 1100
rect 3771 980 3809 1068
rect 3771 948 3774 980
rect 3806 948 3809 980
rect 3771 860 3809 948
rect 3771 828 3774 860
rect 3806 828 3809 860
rect 3771 740 3809 828
rect 3771 708 3774 740
rect 3806 708 3809 740
rect 3771 619 3809 708
rect 4150 1100 4188 1190
rect 4150 1068 4153 1100
rect 4185 1068 4188 1100
rect 4150 980 4188 1068
rect 4150 948 4153 980
rect 4185 948 4188 980
rect 4150 860 4188 948
rect 4150 828 4153 860
rect 4185 828 4188 860
rect 4150 740 4188 828
rect 4150 708 4153 740
rect 4185 708 4188 740
rect 4150 619 4188 708
rect 4529 1100 4567 1190
rect 4529 1068 4532 1100
rect 4564 1068 4567 1100
rect 4529 980 4567 1068
rect 4529 948 4532 980
rect 4564 948 4567 980
rect 4529 860 4567 948
rect 4529 828 4532 860
rect 4564 828 4567 860
rect 4529 740 4567 828
rect 4529 708 4532 740
rect 4564 708 4567 740
rect 4529 619 4567 708
rect 4908 1100 4946 1190
rect 4908 1068 4911 1100
rect 4943 1068 4946 1100
rect 4908 980 4946 1068
rect 4908 948 4911 980
rect 4943 948 4946 980
rect 4908 860 4946 948
rect 4908 828 4911 860
rect 4943 828 4946 860
rect 4908 740 4946 828
rect 4908 708 4911 740
rect 4943 708 4946 740
rect 4908 619 4946 708
rect 5287 1100 5325 1190
rect 5287 1068 5290 1100
rect 5322 1068 5325 1100
rect 5287 980 5325 1068
rect 5287 948 5290 980
rect 5322 948 5325 980
rect 5287 860 5325 948
rect 5287 828 5290 860
rect 5322 828 5325 860
rect 5287 740 5325 828
rect 5287 708 5290 740
rect 5322 708 5325 740
rect 5287 619 5325 708
rect 5666 1100 5704 1190
rect 5666 1068 5669 1100
rect 5701 1068 5704 1100
rect 5666 980 5704 1068
rect 5666 948 5669 980
rect 5701 948 5704 980
rect 5666 860 5704 948
rect 5666 828 5669 860
rect 5701 828 5704 860
rect 5666 740 5704 828
rect 5666 708 5669 740
rect 5701 708 5704 740
rect 5666 619 5704 708
rect 6045 1100 6083 1190
rect 6045 1068 6048 1100
rect 6080 1068 6083 1100
rect 6045 980 6083 1068
rect 6045 948 6048 980
rect 6080 948 6083 980
rect 6045 860 6083 948
rect 6045 828 6048 860
rect 6080 828 6083 860
rect 6045 740 6083 828
rect 6045 708 6048 740
rect 6080 708 6083 740
rect 6045 619 6083 708
rect 6424 1100 6462 1190
rect 6424 1068 6427 1100
rect 6459 1068 6462 1100
rect 6424 980 6462 1068
rect 6424 948 6427 980
rect 6459 948 6462 980
rect 6424 860 6462 948
rect 6424 828 6427 860
rect 6459 828 6462 860
rect 6424 740 6462 828
rect 6424 708 6427 740
rect 6459 708 6462 740
rect 6424 619 6462 708
rect 6803 1100 6841 1190
rect 6803 1068 6806 1100
rect 6838 1068 6841 1100
rect 6803 980 6841 1068
rect 6803 948 6806 980
rect 6838 948 6841 980
rect 6803 860 6841 948
rect 6803 828 6806 860
rect 6838 828 6841 860
rect 6803 740 6841 828
rect 6803 708 6806 740
rect 6838 708 6841 740
rect 6803 619 6841 708
rect 7182 1100 7220 1190
rect 7182 1068 7185 1100
rect 7217 1068 7220 1100
rect 7182 980 7220 1068
rect 7182 948 7185 980
rect 7217 948 7220 980
rect 7182 860 7220 948
rect 7182 828 7185 860
rect 7217 828 7220 860
rect 7182 740 7220 828
rect 7182 708 7185 740
rect 7217 708 7220 740
rect 7182 619 7220 708
rect 7561 1100 7599 1311
rect 7561 1068 7564 1100
rect 7596 1068 7599 1100
rect 7561 980 7599 1068
rect 7561 948 7564 980
rect 7596 948 7599 980
rect 7561 860 7599 948
rect 7561 828 7564 860
rect 7596 828 7599 860
rect 7561 740 7599 828
rect 7561 708 7564 740
rect 7596 708 7599 740
rect 7561 619 7599 708
rect -19 587 318 619
rect 360 587 1535 619
rect 1577 587 2213 619
rect 2255 587 3430 619
rect 3472 587 4108 619
rect 4150 587 5325 619
rect 5367 587 6003 619
rect 6045 587 7220 619
rect 7262 587 7599 619
rect -19 497 19 587
rect -19 465 -16 497
rect 16 465 19 497
rect -19 377 19 465
rect -19 345 -16 377
rect 16 345 19 377
rect -19 257 19 345
rect -19 225 -16 257
rect 16 225 19 257
rect -19 137 19 225
rect -19 105 -16 137
rect 16 105 19 137
rect -19 16 19 105
rect 360 497 398 545
rect 360 465 363 497
rect 395 465 398 497
rect 360 377 398 465
rect 360 345 363 377
rect 395 345 398 377
rect 360 257 398 345
rect 360 225 363 257
rect 395 225 398 257
rect 360 137 398 225
rect 360 105 363 137
rect 395 105 398 137
rect 360 16 398 105
rect 739 497 777 545
rect 739 465 742 497
rect 774 465 777 497
rect 739 377 777 465
rect 739 345 742 377
rect 774 345 777 377
rect 739 257 777 345
rect 739 225 742 257
rect 774 225 777 257
rect 739 137 777 225
rect 739 105 742 137
rect 774 105 777 137
rect 739 16 777 105
rect 1118 497 1156 545
rect 1118 465 1121 497
rect 1153 465 1156 497
rect 1118 377 1156 465
rect 1118 345 1121 377
rect 1153 345 1156 377
rect 1118 257 1156 345
rect 1118 225 1121 257
rect 1153 225 1156 257
rect 1118 137 1156 225
rect 1118 105 1121 137
rect 1153 105 1156 137
rect 1118 16 1156 105
rect 1497 497 1535 545
rect 1497 465 1500 497
rect 1532 465 1535 497
rect 1497 377 1535 465
rect 1497 345 1500 377
rect 1532 345 1535 377
rect 1497 257 1535 345
rect 1497 225 1500 257
rect 1532 225 1535 257
rect 1497 137 1535 225
rect 1497 105 1500 137
rect 1532 105 1535 137
rect 1497 16 1535 105
rect 1876 497 1914 587
rect 1876 465 1879 497
rect 1911 465 1914 497
rect 1876 377 1914 465
rect 1876 345 1879 377
rect 1911 345 1914 377
rect 1876 257 1914 345
rect 1876 225 1879 257
rect 1911 225 1914 257
rect 1876 137 1914 225
rect 1876 105 1879 137
rect 1911 105 1914 137
rect 1876 16 1914 105
rect 2255 497 2293 545
rect 2255 465 2258 497
rect 2290 465 2293 497
rect 2255 377 2293 465
rect 2255 345 2258 377
rect 2290 345 2293 377
rect 2255 257 2293 345
rect 2634 497 2672 587
rect 2634 465 2637 497
rect 2669 465 2672 497
rect 2634 377 2672 465
rect 2634 345 2637 377
rect 2669 345 2672 377
rect 2634 299 2672 345
rect 3013 497 3051 587
rect 3013 465 3016 497
rect 3048 465 3051 497
rect 3013 377 3051 465
rect 3013 345 3016 377
rect 3048 345 3051 377
rect 3013 300 3051 345
rect 3392 497 3430 545
rect 3392 465 3395 497
rect 3427 465 3430 497
rect 3392 377 3430 465
rect 3392 345 3395 377
rect 3427 345 3430 377
rect 2255 225 2258 257
rect 2290 225 2293 257
rect 2255 137 2293 225
rect 2255 105 2258 137
rect 2290 105 2293 137
rect 2255 16 2293 105
rect 2634 257 2672 259
rect 2634 225 2637 257
rect 2669 225 2672 257
rect 2634 137 2672 225
rect 2634 105 2637 137
rect 2669 105 2672 137
rect 2634 16 2672 105
rect 3013 257 3051 260
rect 3013 225 3016 257
rect 3048 225 3051 257
rect 3013 137 3051 225
rect 3013 105 3016 137
rect 3048 105 3051 137
rect 3013 16 3051 105
rect 3392 257 3430 345
rect 3392 225 3395 257
rect 3427 225 3430 257
rect 3392 137 3430 225
rect 3392 105 3395 137
rect 3427 105 3430 137
rect 3392 16 3430 105
rect 3771 497 3809 587
rect 3771 465 3774 497
rect 3806 465 3809 497
rect 3771 377 3809 465
rect 3771 345 3774 377
rect 3806 345 3809 377
rect 3771 257 3809 345
rect 3771 225 3774 257
rect 3806 225 3809 257
rect 3771 137 3809 225
rect 3771 105 3774 137
rect 3806 105 3809 137
rect 3771 16 3809 105
rect 4150 497 4188 545
rect 4150 465 4153 497
rect 4185 465 4188 497
rect 4150 377 4188 465
rect 4529 497 4567 587
rect 4529 465 4532 497
rect 4564 465 4567 497
rect 4529 422 4567 465
rect 4908 497 4946 587
rect 4908 465 4911 497
rect 4943 465 4946 497
rect 4908 422 4946 465
rect 5287 497 5325 545
rect 5287 465 5290 497
rect 5322 465 5325 497
rect 4150 345 4153 377
rect 4185 345 4188 377
rect 4150 257 4188 345
rect 4150 225 4153 257
rect 4185 225 4188 257
rect 4150 137 4188 225
rect 4150 105 4153 137
rect 4185 105 4188 137
rect 4150 16 4188 105
rect 4529 377 4567 380
rect 4529 345 4532 377
rect 4564 345 4567 377
rect 4529 257 4567 345
rect 4529 225 4532 257
rect 4564 225 4567 257
rect 4529 137 4567 225
rect 4529 105 4532 137
rect 4564 105 4567 137
rect 4529 16 4567 105
rect 4908 377 4946 380
rect 4908 345 4911 377
rect 4943 345 4946 377
rect 4908 257 4946 345
rect 4908 225 4911 257
rect 4943 225 4946 257
rect 4908 137 4946 225
rect 4908 105 4911 137
rect 4943 105 4946 137
rect 4908 16 4946 105
rect 5287 377 5325 465
rect 5287 345 5290 377
rect 5322 345 5325 377
rect 5287 257 5325 345
rect 5287 225 5290 257
rect 5322 225 5325 257
rect 5287 137 5325 225
rect 5287 105 5290 137
rect 5322 105 5325 137
rect 5287 16 5325 105
rect 5666 497 5704 587
rect 5666 465 5669 497
rect 5701 465 5704 497
rect 5666 377 5704 465
rect 5666 345 5669 377
rect 5701 345 5704 377
rect 5666 257 5704 345
rect 5666 225 5669 257
rect 5701 225 5704 257
rect 5666 137 5704 225
rect 5666 105 5669 137
rect 5701 105 5704 137
rect 5666 16 5704 105
rect 6045 497 6083 545
rect 6045 465 6048 497
rect 6080 465 6083 497
rect 6045 377 6083 465
rect 6424 497 6462 587
rect 6424 465 6427 497
rect 6459 465 6462 497
rect 6424 422 6462 465
rect 6803 497 6841 540
rect 6803 465 6806 497
rect 6838 465 6841 497
rect 6045 345 6048 377
rect 6080 345 6083 377
rect 6045 257 6083 345
rect 6045 225 6048 257
rect 6080 225 6083 257
rect 6045 137 6083 225
rect 6045 105 6048 137
rect 6080 105 6083 137
rect 6045 16 6083 105
rect 6424 377 6462 380
rect 6424 345 6427 377
rect 6459 345 6462 377
rect 6424 257 6462 345
rect 6424 225 6427 257
rect 6459 225 6462 257
rect 6424 137 6462 225
rect 6424 105 6427 137
rect 6459 105 6462 137
rect 6424 16 6462 105
rect 6803 377 6841 465
rect 6803 345 6806 377
rect 6838 345 6841 377
rect 6803 257 6841 345
rect 6803 225 6806 257
rect 6838 225 6841 257
rect 6803 137 6841 225
rect 6803 105 6806 137
rect 6838 105 6841 137
rect 6803 16 6841 105
rect 7182 497 7220 545
rect 7182 465 7185 497
rect 7217 465 7220 497
rect 7182 377 7220 465
rect 7182 345 7185 377
rect 7217 345 7220 377
rect 7182 257 7220 345
rect 7182 225 7185 257
rect 7217 225 7220 257
rect 7182 137 7220 225
rect 7182 105 7185 137
rect 7217 105 7220 137
rect 7182 16 7220 105
rect 7561 497 7599 587
rect 7561 465 7564 497
rect 7596 465 7599 497
rect 7561 377 7599 465
rect 7561 345 7564 377
rect 7596 345 7599 377
rect 7561 257 7599 345
rect 7561 225 7564 257
rect 7596 225 7599 257
rect 7561 137 7599 225
rect 7561 105 7564 137
rect 7596 105 7599 137
rect 7561 16 7599 105
rect -19 -16 7599 16
<< labels >>
rlabel metal4 -19 2335 -19 2350 7 dummy_top
rlabel metal2 -19 2314 -19 2329 7 shielding
rlabel metal4 360 757 360 772 7 top_8
rlabel metal3 432 772 432 787 7 bot_8
rlabel metal4 2255 751 2255 766 7 top_4
rlabel metal3 2327 776 2327 791 7 bot_4
rlabel metal4 4150 766 4150 781 7 top_2
rlabel metal3 4222 776 4222 791 7 bot_2
rlabel metal4 6045 767 6045 782 7 top_1
rlabel metal3 6117 780 6117 795 7 bot_1
rlabel metal2 175 2290 175 2313 7 dummy_bot
<< end >>
