* NGSPICE file created from adc_array_matrix_flat.ext - technology: sky130A

.subckt adc_array_matrix_flat vcm ctop sample sample_n sw sw_n col_n[0] col_n[1] col_n[2]
+ col_n[3] col_n[4] col_n[5] col_n[6] col_n[7] col_n[8] col_n[9] col_n[10] col_n[11]
+ col_n[12] col_n[13] col_n[14] col_n[15] col_n[16] col_n[17] col_n[18] col_n[19]
+ col_n[20] col_n[21] col_n[22] col_n[23] col_n[24] col_n[25] col_n[26] col_n[27]
+ col_n[28] col_n[29] col_n[30] col_n[31] en_n_bit[2] en_n_bit[1] en_n_bit[0] row_n[0]
+ row_n[1] row_n[2] row_n[3] row_n[4] row_n[5] row_n[6] row_n[7] row_n[8] row_n[9]
+ row_n[10] row_n[11] row_n[12] row_n[13] row_n[14] row_n[15] rowon_n[0] rowon_n[1]
+ rowon_n[2] rowon_n[3] rowon_n[4] rowon_n[5] rowon_n[6] rowon_n[7] rowon_n[8] rowon_n[9]
+ rowon_n[10] rowon_n[11] rowon_n[12] rowon_n[13] rowon_n[14] rowon_n[15] analog_in
+ en_C0_n VSS VDD
X0 adc_array_wafflecap_8_8_0[10|4]/adc_array_circuit_150n_0/vdrv row_n[11] adc_array_wafflecap_8_8_0[10|4]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1 adc_array_wafflecap_8_8_0[10|14]/adc_array_circuit_150n_0/vdrv row_n[11] adc_array_wafflecap_8_8_0[10|14]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2 adc_array_wafflecap_8_8_0[8|18]/adc_array_circuit_150n_0/vint1 col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=1.72952e+14p ps=1.48678e+09u w=800000u l=150000u
X3 vcm adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|21]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=7.7469e+13p pd=8.687e+08u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4 adc_array_wafflecap_8_Dummy_4[17]/adc_array_circuit_150n_0/vint2 col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=4.352e+14p ps=2.01194e+09u w=420000u l=150000u
X5 adc_array_wafflecap_8_8_0[11|16]/adc_array_circuit_150n_0/vint1 col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X6 VDD rowon_n[4] adc_array_wafflecap_8_8_0[3|17]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X7 adc_array_wafflecap_8_8_0[7|17]/adc_array_circuit_150n_0/vdrv row_n[8] adc_array_wafflecap_8_8_0[7|17]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8 VSS row_n[8] adc_array_wafflecap_8_8_0[7|24]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X9 adc_array_wafflecap_8_8_0[0|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X10 VSS row_n[2] adc_array_wafflecap_8_8_0[1|27]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X11 VSS row_n[6] adc_array_wafflecap_8_8_0[5|26]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X12 VSS row_n[14] adc_array_wafflecap_8_8_0[13|23]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X13 vcm adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|15]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X14 adc_array_wafflecap_8_8_0[7|6]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|6]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X15 adc_array_wafflecap_8_8_0[7|16]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|16]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X16 adc_array_wafflecap_8_8_0[14|29]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|29]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X17 adc_array_wafflecap_8_8_0[13|16]/adc_array_circuit_150n_0/vdrv row_n[14] adc_array_wafflecap_8_8_0[13|16]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X18 vcm adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|5]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X19 adc_array_wafflecap_8_8_0[11|27]/adc_array_circuit_150n_0/vint2 rowon_n[12] adc_array_wafflecap_8_8_0[11|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X20 VDD rowon_n[10] adc_array_wafflecap_8_8_0[9|23]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X21 vcm adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|26]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X22 vcm adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|4]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X23 adc_array_wafflecap_8_8_0[0|6]/adc_array_circuit_150n_0/vint2 col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X24 VDD VDD adc_array_wafflecap_8_Dummy_4[23]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X25 adc_array_wafflecap_8_8_0[13|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=1.4756e+14p ps=1.3209e+09u w=800000u l=150000u
X26 adc_array_wafflecap_8_8_0[13|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X27 adc_array_wafflecap_8_8_0[12|22]/adc_array_circuit_150n_0/vint2 col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X28 adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X29 adc_array_wafflecap_8_8_0[1|27]/adc_array_circuit_150n_0/vint1 col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X30 VSS row_n[11] adc_array_wafflecap_8_8_0[10|26]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X31 adc_array_wafflecap_8_8_0[3|8]/adc_array_circuit_150n_0/vdrv row_n[4] adc_array_wafflecap_8_8_0[3|8]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X32 adc_array_wafflecap_8_Dummy_1[3]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_1[3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X33 adc_array_wafflecap_8_8_0[2|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X34 adc_array_wafflecap_8_8_0[3|9]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|9]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X35 adc_array_wafflecap_8_8_0[3|18]/adc_array_circuit_150n_0/vint1 col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X36 VSS row_n[4] adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X37 vcm VSS adc_array_wafflecap_8_Dummy_4[18]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X38 adc_array_wafflecap_8_8_0[14|21]/adc_array_circuit_150n_0/vint1 col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X39 adc_array_wafflecap_8_8_0[7|13]/adc_array_circuit_150n_0/vint2 col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X40 adc_array_wafflecap_8_Dummy_8[4]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_8[4]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X41 adc_array_wafflecap_8_8_0[7|3]/adc_array_circuit_150n_0/vint2 col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X42 adc_array_wafflecap_8_8_0[2|22]/adc_array_circuit_150n_0/vint2 rowon_n[3] adc_array_wafflecap_8_8_0[2|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X43 adc_array_wafflecap_8_8_0[10|22]/adc_array_circuit_150n_0/vdrv row_n[11] adc_array_wafflecap_8_8_0[10|22]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X44 adc_array_wafflecap_8_8_0[8|26]/adc_array_circuit_150n_0/vint1 col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X45 adc_array_wafflecap_8_Dummy_1[2]/adc_array_circuit_150n_0/vint2 col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X46 adc_array_wafflecap_8_8_0[2|10]/adc_array_circuit_150n_0/vint2 col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X47 adc_array_wafflecap_8_8_0[14|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X48 adc_array_wafflecap_8_8_0[9|12]/adc_array_circuit_150n_0/vint1 col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X49 adc_array_wafflecap_8_8_0[8|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X50 adc_array_wafflecap_8_8_0[6|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X51 adc_array_wafflecap_8_8_0[2|0]/adc_array_circuit_150n_0/vdrv row_n[3] adc_array_wafflecap_8_8_0[2|0]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X52 adc_array_wafflecap_8_8_1[22]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[22]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X53 vcm adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|30]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X54 adc_array_wafflecap_8_8_0[13|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X55 vcm adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|21]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X56 adc_array_wafflecap_8_8_0[9|2]/adc_array_circuit_150n_0/vint1 col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X57 VDD rowon_n[6] adc_array_wafflecap_8_8_0[5|24]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X58 adc_array_wafflecap_8_8_0[2|1]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|1]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X59 adc_array_wafflecap_8_8_0[0|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X60 adc_array_wafflecap_8_8_0[5|12]/adc_array_circuit_150n_0/vdrv row_n[6] adc_array_wafflecap_8_8_0[5|12]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X61 adc_array_wafflecap_8_8_0[5|13]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|13]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X62 adc_array_wafflecap_8_8_0[1|14]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|14]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X63 VDD rowon_n[1] adc_array_wafflecap_8_8_0[0|22]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X64 adc_array_wafflecap_8_8_0[8|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X65 adc_array_wafflecap_8_8_0[0|10]/adc_array_circuit_150n_0/vdrv row_n[1] adc_array_wafflecap_8_8_0[0|10]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X66 adc_array_wafflecap_8_8_0[8|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X67 adc_array_wafflecap_8_8_0[6|21]/adc_array_circuit_150n_0/vint2 col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X68 vcm adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[18]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X69 adc_array_wafflecap_8_8_0[0|15]/adc_array_circuit_150n_0/vint2 col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X70 adc_array_wafflecap_8_8_0[14|0]/adc_array_circuit_150n_0/vdrv row_n[15] adc_array_wafflecap_8_8_0[14|0]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X71 adc_array_wafflecap_8_8_0[14|10]/adc_array_circuit_150n_0/vdrv row_n[15] adc_array_wafflecap_8_8_0[14|10]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X72 adc_array_wafflecap_8_8_0[12|21]/adc_array_circuit_150n_0/vint2 rowon_n[13] adc_array_wafflecap_8_8_0[12|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X73 adc_array_wafflecap_8_8_0[4|5]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|5]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X74 adc_array_wafflecap_8_8_0[0|26]/adc_array_circuit_150n_0/vint2 rowon_n[1] adc_array_wafflecap_8_8_0[0|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X75 adc_array_wafflecap_8_8_0[0|6]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|6]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X76 vcm adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|9]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X77 adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X78 adc_array_wafflecap_8_8_0[11|25]/adc_array_circuit_150n_0/vint2 rowon_n[12] adc_array_wafflecap_8_8_0[11|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X79 adc_array_wafflecap_8_8_0[9|28]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|28]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X80 VSS row_n[9] adc_array_wafflecap_8_8_0[8|22]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X81 VSS row_n[7] adc_array_wafflecap_8_8_0[6|6]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X82 VSS sample_n adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X83 adc_array_wafflecap_8_8_0[10|6]/adc_array_circuit_150n_0/vint2 rowon_n[11] adc_array_wafflecap_8_8_0[10|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X84 adc_array_wafflecap_8_8_0[10|16]/adc_array_circuit_150n_0/vint2 rowon_n[11] adc_array_wafflecap_8_8_0[10|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X85 adc_array_wafflecap_8_8_0[8|14]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|14]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X86 adc_array_wafflecap_8_8_1[1]/adc_array_circuit_150n_0/vdrv row_n[0] adc_array_wafflecap_8_8_1[1]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X87 vcm adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|13]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X88 adc_array_wafflecap_8_8_0[11|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X89 adc_array_wafflecap_8_8_0[8|4]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|4]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X90 adc_array_wafflecap_8_8_0[6|21]/adc_array_circuit_150n_0/vdrv row_n[7] adc_array_wafflecap_8_8_0[6|21]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X91 adc_array_wafflecap_8_8_0[3|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X92 VDD rowon_n[4] adc_array_wafflecap_8_8_0[3|28]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X93 adc_array_wafflecap_8_Dummy_1[6]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_1[6]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X94 vcm adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|3]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X95 adc_array_wafflecap_8_8_0[4|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X96 adc_array_wafflecap_8_8_0[3|17]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|17]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X97 VDD rowon_n[11] adc_array_wafflecap_8_8_0[10|21]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X98 VDD VSS adc_array_wafflecap_8_Dummy_3[1]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X99 VDD rowon_n[10] adc_array_wafflecap_8_8_0[9|2]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X100 VDD rowon_n[10] adc_array_wafflecap_8_8_0[9|12]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X101 VDD rowon_n[5] adc_array_wafflecap_8_8_0[4|10]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X102 VDD rowon_n[9] adc_array_wafflecap_8_8_0[8|16]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X103 VSS VSS adc_array_wafflecap_8_Dummy_2[4]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X104 adc_array_wafflecap_8_8_0[13|20]/adc_array_circuit_150n_0/vint2 col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X105 VDD rowon_n[9] adc_array_wafflecap_8_8_0[8|6]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X106 adc_array_wafflecap_8_8_0[6|6]/adc_array_circuit_150n_0/vint1 col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X107 adc_array_wafflecap_8_8_0[2|7]/adc_array_circuit_150n_0/vint1 col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X108 adc_array_wafflecap_8_8_0[2|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X109 VDD rowon_n[0] adc_array_wafflecap_8_8_1[7]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X110 adc_array_wafflecap_8_8_0[2|30]/adc_array_circuit_150n_0/vint2 rowon_n[3] adc_array_wafflecap_8_8_0[2|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X111 VSS row_n[13] adc_array_wafflecap_8_8_0[12|10]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X112 adc_array_wafflecap_8_8_1[12]/adc_array_circuit_150n_0/vint2 rowon_n[0] adc_array_wafflecap_8_8_1[12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X113 adc_array_wafflecap_8_8_0[1|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X114 VSS row_n[13] adc_array_wafflecap_8_8_0[12|0]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X115 adc_array_wafflecap_8_Dummy_4[20]/adc_array_circuit_150n_0/vint1 col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X116 adc_array_wafflecap_8_8_0[13|7]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|7]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X117 VSS row_n[12] adc_array_wafflecap_8_8_0[11|14]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X118 adc_array_wafflecap_8_8_0[9|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X119 adc_array_wafflecap_8_8_0[8|11]/adc_array_circuit_150n_0/vint2 col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X120 adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/vint1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X121 adc_array_wafflecap_8_8_0[11|29]/adc_array_circuit_150n_0/vdrv row_n[12] adc_array_wafflecap_8_8_0[11|29]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X122 VSS row_n[12] adc_array_wafflecap_8_8_0[11|4]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X123 adc_array_wafflecap_8_8_0[8|1]/adc_array_circuit_150n_0/vint2 col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X124 VDD rowon_n[3] adc_array_wafflecap_8_8_0[2|15]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X125 adc_array_wafflecap_8_8_1[28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_1[28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X126 adc_array_wafflecap_8_8_1[23]/adc_array_circuit_150n_0/vdrv row_n[0] adc_array_wafflecap_8_8_1[23]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X127 VDD rowon_n[1] adc_array_wafflecap_8_8_0[0|30]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X128 vcm adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|10]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X129 adc_array_wafflecap_8_8_0[10|10]/adc_array_circuit_150n_0/vint1 col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X130 adc_array_wafflecap_8_8_0[4|11]/adc_array_circuit_150n_0/vint1 col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X131 adc_array_wafflecap_8_8_0[4|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X132 adc_array_wafflecap_8_8_0[0|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X133 adc_array_wafflecap_8_8_0[10|0]/adc_array_circuit_150n_0/vint1 col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X134 adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X135 adc_array_wafflecap_8_8_1[8]/adc_array_circuit_150n_0/vint1 col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X136 adc_array_wafflecap_8_8_0[6|2]/adc_array_circuit_150n_0/vint2 rowon_n[7] adc_array_wafflecap_8_8_0[6|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X137 adc_array_wafflecap_8_8_1[27]/adc_array_circuit_150n_0/vint2 col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X138 adc_array_wafflecap_8_8_0[6|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X139 VSS row_n[6] adc_array_wafflecap_8_8_0[5|20]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X140 adc_array_wafflecap_8_8_0[8|22]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|22]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X141 adc_array_wafflecap_8_8_0[7|20]/adc_array_circuit_150n_0/vint2 rowon_n[8] adc_array_wafflecap_8_8_0[7|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X142 adc_array_wafflecap_8_8_0[5|18]/adc_array_circuit_150n_0/vint2 col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X143 VSS row_n[0] adc_array_wafflecap_8_8_1[13]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X144 adc_array_wafflecap_8_8_0[1|19]/adc_array_circuit_150n_0/vint2 col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X145 adc_array_wafflecap_8_8_0[2|30]/adc_array_circuit_150n_0/vdrv row_n[3] adc_array_wafflecap_8_8_0[2|30]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X146 vcm adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|2]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X147 adc_array_wafflecap_8_Dummy_4[9]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[9]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X148 adc_array_wafflecap_8_8_0[13|19]/adc_array_circuit_150n_0/vint2 rowon_n[14] adc_array_wafflecap_8_8_0[13|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X149 adc_array_wafflecap_8_8_0[12|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X150 vcm adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|8]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X151 adc_array_wafflecap_8_8_0[7|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X152 adc_array_wafflecap_8_8_0[7|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X153 adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X154 adc_array_wafflecap_8_8_1[4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X155 adc_array_wafflecap_8_8_0[12|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X156 adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/vint2 rowon_n[13] adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X157 vcm adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|12]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X158 VDD rowon_n[7] adc_array_wafflecap_8_8_0[6|2]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X159 adc_array_wafflecap_8_Dummy_4[26]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[26]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X160 adc_array_wafflecap_8_8_0[13|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X161 adc_array_wafflecap_8_8_0[11|14]/adc_array_circuit_150n_0/vint2 rowon_n[12] adc_array_wafflecap_8_8_0[11|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X162 vcm adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|2]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X163 adc_array_wafflecap_8_Dummy_8[5]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_8[5]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X164 adc_array_wafflecap_8_8_0[11|4]/adc_array_circuit_150n_0/vint2 rowon_n[12] adc_array_wafflecap_8_8_0[11|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X165 adc_array_wafflecap_8_Dummy_2[0]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X166 adc_array_wafflecap_8_8_0[14|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X167 adc_array_wafflecap_8_8_0[14|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X168 VSS row_n[4] adc_array_wafflecap_8_8_0[3|25]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X169 adc_array_wafflecap_8_8_0[1|19]/adc_array_circuit_150n_0/vdrv row_n[2] adc_array_wafflecap_8_8_0[1|19]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X170 adc_array_wafflecap_8_8_0[10|16]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|16]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X171 VSS row_n[7] adc_array_wafflecap_8_8_0[6|3]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X172 adc_array_wafflecap_8_8_0[10|6]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|6]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X173 VDD rowon_n[11] adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X174 adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/vint2 VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X175 adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/vint2 col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X176 VSS row_n[8] adc_array_wafflecap_8_8_0[7|9]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X177 adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/vdrv row_n[0] adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X178 vcm adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|23]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X179 vcm adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|24]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X180 adc_array_wafflecap_8_8_0[0|17]/adc_array_circuit_150n_0/vint2 rowon_n[1] adc_array_wafflecap_8_8_0[0|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X181 VSS row_n[14] adc_array_wafflecap_8_8_0[13|8]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X182 adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/vint1 col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X183 adc_array_wafflecap_8_8_0[6|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X184 adc_array_wafflecap_8_8_0[6|3]/adc_array_circuit_150n_0/vint1 col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X185 vcm adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|14]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X186 adc_array_wafflecap_8_Dummy_4[31]/adc_array_circuit_150n_0/vint1 col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X187 adc_array_wafflecap_8_8_0[13|18]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|18]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X188 adc_array_wafflecap_8_8_0[9|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X189 adc_array_wafflecap_8_8_0[0|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X190 VSS row_n[2] adc_array_wafflecap_8_8_0[1|29]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X191 adc_array_wafflecap_8_8_0[12|7]/adc_array_circuit_150n_0/vint2 col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X192 VDD VSS adc_array_wafflecap_8_Dummy_2[0]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X193 adc_array_wafflecap_8_8_0[11|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X194 vcm adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|6]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X195 adc_array_wafflecap_8_8_0[4|19]/adc_array_circuit_150n_0/vint2 rowon_n[5] adc_array_wafflecap_8_8_0[4|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X196 adc_array_wafflecap_8_8_0[14|6]/adc_array_circuit_150n_0/vint1 col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X197 adc_array_wafflecap_8_8_0[4|7]/adc_array_circuit_150n_0/vint2 col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X198 VSS row_n[1] adc_array_wafflecap_8_8_0[0|18]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X199 adc_array_wafflecap_8_8_0[0|8]/adc_array_circuit_150n_0/vint2 col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X200 vcm adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|28]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X201 VSS row_n[5] adc_array_wafflecap_8_8_0[4|17]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X202 vcm VSS adc_array_wafflecap_8_Dummy_3[3]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X203 vcm adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|27]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X204 vcm adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X205 adc_array_wafflecap_8_8_0[10|7]/adc_array_circuit_150n_0/vdrv row_n[11] adc_array_wafflecap_8_8_0[10|7]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X206 adc_array_wafflecap_8_8_0[8|18]/adc_array_circuit_150n_0/vint2 rowon_n[9] adc_array_wafflecap_8_8_0[8|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X207 adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/vint2 rowon_n[8] adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X208 VDD rowon_n[4] adc_array_wafflecap_8_8_0[3|22]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X209 adc_array_wafflecap_8_8_1[0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_1[0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X210 VDD sample_n adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X211 adc_array_wafflecap_8_8_0[1|29]/adc_array_circuit_150n_0/vint1 col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X212 adc_array_wafflecap_8_8_0[8|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X213 adc_array_wafflecap_8_8_0[7|9]/adc_array_circuit_150n_0/vint2 rowon_n[8] adc_array_wafflecap_8_8_0[7|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X214 adc_array_wafflecap_8_8_0[3|10]/adc_array_circuit_150n_0/vdrv row_n[4] adc_array_wafflecap_8_8_0[3|10]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X215 adc_array_wafflecap_8_8_0[3|11]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|11]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X216 adc_array_wafflecap_8_Dummy_1[5]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_1[5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X217 adc_array_wafflecap_8_8_0[13|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X218 adc_array_wafflecap_8_8_0[8|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X219 adc_array_wafflecap_8_Dummy_4[20]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[20]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X220 adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X221 vcm adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|19]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X222 adc_array_wafflecap_8_4_0/adc_array_circuit_150n_0/vdrv en_n_bit[2] adc_array_wafflecap_8_4_0/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X223 adc_array_wafflecap_8_8_0[9|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X224 adc_array_wafflecap_8_Dummy_2[1]/adc_array_circuit_150n_0/vint1 col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X225 adc_array_wafflecap_8_8_0[9|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X226 adc_array_wafflecap_8_Dummy_7/adc_array_circuit_150n_0/vint2 col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X227 adc_array_wafflecap_8_8_0[2|24]/adc_array_circuit_150n_0/vint2 rowon_n[3] adc_array_wafflecap_8_8_0[2|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X228 adc_array_wafflecap_8_Dummy_4[14]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X229 adc_array_wafflecap_8_Dummy_1[4]/adc_array_circuit_150n_0/vint2 col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X230 adc_array_wafflecap_8_8_0[2|12]/adc_array_circuit_150n_0/vint2 col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X231 adc_array_wafflecap_8_Dummy_4[4]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X232 adc_array_wafflecap_8_8_1[24]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[24]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X233 vcm adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X234 adc_array_wafflecap_8_Dummy_4[11]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X235 adc_array_wafflecap_8_8_0[14|25]/adc_array_circuit_150n_0/vint2 col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X236 VSS row_n[13] adc_array_wafflecap_8_8_0[12|29]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X237 adc_array_wafflecap_8_8_0[11|14]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|14]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X238 adc_array_wafflecap_8_8_0[9|26]/adc_array_circuit_150n_0/vint2 col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X239 adc_array_wafflecap_8_8_0[6|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X240 adc_array_wafflecap_8_8_0[2|2]/adc_array_circuit_150n_0/vdrv row_n[3] adc_array_wafflecap_8_8_0[2|2]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X241 adc_array_wafflecap_8_8_0[2|3]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|3]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X242 adc_array_wafflecap_8_Dummy_8[2]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_8[2]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X243 adc_array_wafflecap_8_Dummy_4[1]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X244 adc_array_wafflecap_8_8_0[11|4]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|4]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X245 adc_array_wafflecap_8_8_0[1|16]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|16]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X246 adc_array_wafflecap_8_8_0[8|30]/adc_array_circuit_150n_0/vint2 col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X247 adc_array_wafflecap_8_8_0[5|15]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|15]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X248 adc_array_wafflecap_8_8_0[14|12]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|12]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X249 VSS row_n[9] adc_array_wafflecap_8_8_0[8|7]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X250 adc_array_wafflecap_8_8_1[22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_1[22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X251 VDD rowon_n[1] adc_array_wafflecap_8_8_0[0|24]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X252 adc_array_wafflecap_8_8_0[14|2]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|2]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X253 VDD rowon_n[15] adc_array_wafflecap_8_8_0[14|28]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X254 adc_array_wafflecap_8_8_0[0|12]/adc_array_circuit_150n_0/vdrv row_n[1] adc_array_wafflecap_8_8_0[0|12]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X255 adc_array_wafflecap_8_8_0[12|25]/adc_array_circuit_150n_0/vdrv row_n[13] adc_array_wafflecap_8_8_0[12|25]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X256 adc_array_wafflecap_8_8_0[10|29]/adc_array_circuit_150n_0/vint1 col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X257 adc_array_wafflecap_8_8_0[6|23]/adc_array_circuit_150n_0/vint2 col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X258 VDD rowon_n[14] adc_array_wafflecap_8_8_0[13|0]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X259 VDD rowon_n[14] adc_array_wafflecap_8_8_0[13|10]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X260 adc_array_wafflecap_8_8_0[7|26]/adc_array_circuit_150n_0/vdrv row_n[8] adc_array_wafflecap_8_8_0[7|26]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X261 adc_array_wafflecap_8_8_0[5|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X262 VDD rowon_n[3] adc_array_wafflecap_8_8_0[2|8]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X263 adc_array_wafflecap_8_8_0[1|0]/adc_array_circuit_150n_0/vint2 rowon_n[2] adc_array_wafflecap_8_8_0[1|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X264 adc_array_wafflecap_8_8_0[11|15]/adc_array_circuit_150n_0/vint1 col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X265 vcm adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|24]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X266 adc_array_wafflecap_8_8_0[11|5]/adc_array_circuit_150n_0/vint1 col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X267 adc_array_wafflecap_8_8_0[10|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X268 adc_array_wafflecap_8_8_0[0|28]/adc_array_circuit_150n_0/vint2 rowon_n[1] adc_array_wafflecap_8_8_0[0|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X269 adc_array_wafflecap_8_8_0[12|18]/adc_array_circuit_150n_0/vint2 col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X270 adc_array_wafflecap_8_8_0[3|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X271 VDD rowon_n[4] adc_array_wafflecap_8_8_0[3|30]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X272 adc_array_wafflecap_8_8_0[2|24]/adc_array_circuit_150n_0/vdrv row_n[3] adc_array_wafflecap_8_8_0[2|24]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X273 adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X274 adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X275 adc_array_wafflecap_8_8_0[6|23]/adc_array_circuit_150n_0/vdrv row_n[7] adc_array_wafflecap_8_8_0[6|23]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X276 adc_array_wafflecap_8_Dummy_4[28]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[28]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X277 vcm adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|27]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X278 adc_array_wafflecap_8_8_0[4|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X279 VSS row_n[0] adc_array_wafflecap_8_8_1[6]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X280 VDD rowon_n[2] adc_array_wafflecap_8_8_0[1|0]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X281 VSS sample adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X282 VDD VSS adc_array_wafflecap_8_Dummy_3[3]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X283 adc_array_wafflecap_8_8_0[14|17]/adc_array_circuit_150n_0/vint1 col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X284 adc_array_wafflecap_8_8_0[14|24]/adc_array_circuit_150n_0/vint2 rowon_n[15] adc_array_wafflecap_8_8_0[14|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X285 vcm adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|7]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X286 adc_array_wafflecap_8_8_0[2|9]/adc_array_circuit_150n_0/vint1 col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X287 adc_array_wafflecap_8_Dummy_4[22]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X288 adc_array_wafflecap_8_8_0[10|18]/adc_array_circuit_150n_0/vdrv row_n[11] adc_array_wafflecap_8_8_0[10|18]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X289 VSS row_n[11] adc_array_wafflecap_8_8_0[10|25]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X290 adc_array_wafflecap_8_8_0[8|7]/adc_array_circuit_150n_0/vint2 rowon_n[9] adc_array_wafflecap_8_8_0[8|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X291 adc_array_wafflecap_8_8_0[8|29]/adc_array_circuit_150n_0/vint2 rowon_n[9] adc_array_wafflecap_8_8_0[8|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X292 adc_array_wafflecap_8_8_0[3|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X293 adc_array_wafflecap_8_8_0[2|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X294 VDD rowon_n[0] adc_array_wafflecap_8_8_1[9]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X295 VSS row_n[2] adc_array_wafflecap_8_8_0[1|1]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X296 adc_array_wafflecap_8_8_0[11|22]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|22]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X297 adc_array_wafflecap_8_8_0[4|4]/adc_array_circuit_150n_0/vint2 col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X298 vcm VSS adc_array_wafflecap_8_Dummy_4[17]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X299 adc_array_wafflecap_8_8_1[14]/adc_array_circuit_150n_0/vint2 rowon_n[0] adc_array_wafflecap_8_8_1[14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X300 adc_array_wafflecap_8_8_0[1|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X301 vcm VSS adc_array_wafflecap_8_Dummy_4[7]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X302 VDD rowon_n[13] adc_array_wafflecap_8_8_0[12|24]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X303 adc_array_wafflecap_8_8_0[10|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X304 adc_array_wafflecap_8_8_0[10|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X305 adc_array_wafflecap_8_8_0[8|25]/adc_array_circuit_150n_0/vint1 col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X306 adc_array_wafflecap_8_8_0[3|16]/adc_array_circuit_150n_0/vint2 col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X307 adc_array_wafflecap_8_8_0[8|7]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|7]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X308 adc_array_wafflecap_8_8_0[4|27]/adc_array_circuit_150n_0/vdrv row_n[5] adc_array_wafflecap_8_8_0[4|27]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X309 adc_array_wafflecap_8_8_0[4|28]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|28]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X310 adc_array_wafflecap_8_8_1[30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_1[30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X311 vcm VSS adc_array_wafflecap_8_Dummy_0[1]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X312 adc_array_wafflecap_8_8_0[0|29]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|29]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X313 adc_array_wafflecap_8_8_0[1|1]/adc_array_circuit_150n_0/vint1 col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X314 adc_array_wafflecap_8_Dummy_4[24]/adc_array_circuit_150n_0/vint2 col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X315 VSS row_n[14] adc_array_wafflecap_8_8_0[13|27]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X316 vcm adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|12]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X317 adc_array_wafflecap_8_8_0[6|19]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|19]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X318 adc_array_wafflecap_8_8_0[4|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X319 adc_array_wafflecap_8_8_0[0|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X320 VSS row_n[15] adc_array_wafflecap_8_8_0[14|13]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X321 VSS row_n[15] adc_array_wafflecap_8_8_0[14|3]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X322 adc_array_wafflecap_8_8_0[6|4]/adc_array_circuit_150n_0/vint2 rowon_n[7] adc_array_wafflecap_8_8_0[6|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X323 adc_array_wafflecap_8_8_1[10]/adc_array_circuit_150n_0/vint1 col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X324 adc_array_wafflecap_8_Dummy_4[11]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[11]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X325 VDD VDD adc_array_wafflecap_8_Dummy_4[27]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X326 adc_array_wafflecap_8_8_0[10|14]/adc_array_circuit_150n_0/vint2 col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X327 VSS row_n[9] adc_array_wafflecap_8_8_0[8|18]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X328 VSS row_n[6] adc_array_wafflecap_8_8_0[5|22]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X329 adc_array_wafflecap_8_8_1[29]/adc_array_circuit_150n_0/vint2 col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X330 VSS row_n[2] adc_array_wafflecap_8_8_0[1|23]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X331 adc_array_wafflecap_8_Dummy_4[1]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[1]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X332 VDD rowon_n[15] adc_array_wafflecap_8_8_0[14|17]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X333 adc_array_wafflecap_8_8_0[10|4]/adc_array_circuit_150n_0/vint2 col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X334 adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/vint2 rowon_n[6] adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X335 adc_array_wafflecap_8_8_0[13|23]/adc_array_circuit_150n_0/vdrv row_n[14] adc_array_wafflecap_8_8_0[13|23]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X336 adc_array_wafflecap_8_8_0[10|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X337 vcm adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|23]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X338 adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/vdrv row_n[3] adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X339 adc_array_wafflecap_8_8_0[12|13]/adc_array_circuit_150n_0/vint1 col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X340 adc_array_wafflecap_8_8_0[12|3]/adc_array_circuit_150n_0/vint1 col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X341 adc_array_wafflecap_8_8_0[7|17]/adc_array_circuit_150n_0/vint2 col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X342 adc_array_wafflecap_8_8_0[8|4]/adc_array_circuit_150n_0/vdrv row_n[9] adc_array_wafflecap_8_8_0[8|4]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X343 adc_array_wafflecap_8_8_0[8|14]/adc_array_circuit_150n_0/vdrv row_n[9] adc_array_wafflecap_8_8_0[8|14]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X344 VDD rowon_n[7] adc_array_wafflecap_8_8_0[6|4]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X345 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X346 adc_array_wafflecap_8_8_0[1|23]/adc_array_circuit_150n_0/vint1 col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X347 vcm adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|21]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X348 adc_array_wafflecap_8_8_0[13|16]/adc_array_circuit_150n_0/vint2 col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X349 VSS sample_n adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X350 adc_array_wafflecap_8_8_0[11|12]/adc_array_circuit_150n_0/vdrv row_n[12] adc_array_wafflecap_8_8_0[11|12]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X351 adc_array_wafflecap_8_8_0[9|16]/adc_array_circuit_150n_0/vint1 col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X352 adc_array_wafflecap_8_8_0[9|23]/adc_array_circuit_150n_0/vint2 rowon_n[10] adc_array_wafflecap_8_8_0[9|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X353 adc_array_wafflecap_8_8_0[8|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X354 VSS row_n[7] adc_array_wafflecap_8_8_0[6|5]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X355 adc_array_wafflecap_8_8_0[11|2]/adc_array_circuit_150n_0/vdrv row_n[12] adc_array_wafflecap_8_8_0[11|2]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X356 adc_array_wafflecap_8_Dummy_8[5]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_8[5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X357 adc_array_wafflecap_8_Dummy_4[23]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X358 adc_array_wafflecap_8_8_0[14|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X359 adc_array_wafflecap_8_8_0[14|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X360 VSS row_n[4] adc_array_wafflecap_8_8_0[3|26]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X361 VSS row_n[12] adc_array_wafflecap_8_8_0[11|23]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X362 vcm adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|15]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X363 adc_array_wafflecap_8_Dummy_4[33]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X364 adc_array_wafflecap_8_8_0[12|29]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|29]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X365 vcm adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|5]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X366 VDD rowon_n[8] adc_array_wafflecap_8_8_0[7|23]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X367 adc_array_wafflecap_8_8_0[6|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X368 vcm adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|25]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X369 vcm adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|26]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X370 adc_array_wafflecap_8_8_0[6|5]/adc_array_circuit_150n_0/vint1 col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X371 vcm adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|4]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X372 adc_array_wafflecap_8_Dummy_8[4]/adc_array_circuit_150n_0/vint2 col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X373 VSS row_n[15] adc_array_wafflecap_8_8_0[14|21]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X374 VDD rowon_n[14] adc_array_wafflecap_8_8_0[13|22]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X375 adc_array_wafflecap_8_8_0[11|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X376 vcm adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|16]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X377 adc_array_wafflecap_8_8_0[11|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X378 adc_array_wafflecap_8_8_0[10|22]/adc_array_circuit_150n_0/vint2 col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X379 adc_array_wafflecap_8_8_1[27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X380 VSS row_n[9] adc_array_wafflecap_8_8_0[8|26]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X381 adc_array_wafflecap_8_8_0[5|7]/adc_array_circuit_150n_0/vdrv row_n[6] adc_array_wafflecap_8_8_0[5|7]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X382 VDD rowon_n[6] adc_array_wafflecap_8_8_0[5|19]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X383 adc_array_wafflecap_8_8_0[0|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X384 adc_array_wafflecap_8_8_0[8|18]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|18]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X385 adc_array_wafflecap_8_8_0[5|8]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|8]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X386 adc_array_wafflecap_8_8_0[5|17]/adc_array_circuit_150n_0/vint1 col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X387 VSS row_n[2] adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X388 adc_array_wafflecap_8_8_0[1|9]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|9]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X389 vcm adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|17]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X390 VSS row_n[10] adc_array_wafflecap_8_8_0[9|2]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X391 VSS row_n[10] adc_array_wafflecap_8_8_0[9|12]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X392 adc_array_wafflecap_8_8_0[5|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X393 adc_array_wafflecap_8_8_0[12|21]/adc_array_circuit_150n_0/vint1 col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X394 VDD rowon_n[15] adc_array_wafflecap_8_8_0[14|15]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X395 adc_array_wafflecap_8_8_0[0|22]/adc_array_circuit_150n_0/vint2 rowon_n[1] adc_array_wafflecap_8_8_0[0|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X396 VDD rowon_n[15] adc_array_wafflecap_8_8_0[14|5]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X397 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.64e+07u l=1.6e+07u
X398 adc_array_wafflecap_8_8_0[8|22]/adc_array_circuit_150n_0/vdrv row_n[9] adc_array_wafflecap_8_8_0[8|22]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X399 adc_array_wafflecap_8_8_0[4|21]/adc_array_circuit_150n_0/vint2 rowon_n[5] adc_array_wafflecap_8_8_0[4|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X400 adc_array_wafflecap_8_8_0[0|10]/adc_array_circuit_150n_0/vint2 col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X401 adc_array_wafflecap_8_8_0[12|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X402 adc_array_wafflecap_8_8_0[7|12]/adc_array_circuit_150n_0/vint1 col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X403 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X404 vcm VSS adc_array_wafflecap_8_Dummy_3[5]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X405 adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/vint1 col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X406 adc_array_wafflecap_8_8_0[11|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X407 vcm adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|21]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X408 adc_array_wafflecap_8_8_0[7|2]/adc_array_circuit_150n_0/vint1 col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X409 adc_array_wafflecap_8_8_0[4|0]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|0]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X410 adc_array_wafflecap_8_8_0[3|12]/adc_array_circuit_150n_0/vdrv row_n[4] adc_array_wafflecap_8_8_0[3|12]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X411 VDD rowon_n[4] adc_array_wafflecap_8_8_0[3|24]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X412 adc_array_wafflecap_8_2_0/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_2_0/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X413 adc_array_wafflecap_8_8_0[0|1]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|1]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X414 adc_array_wafflecap_8_8_0[14|10]/adc_array_circuit_150n_0/vint2 col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X415 adc_array_wafflecap_8_8_0[3|13]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|13]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X416 adc_array_wafflecap_8_8_0[14|0]/adc_array_circuit_150n_0/vint2 col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X417 VDD VSS adc_array_wafflecap_8_Dummy_2[5]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X418 adc_array_wafflecap_8_Dummy_1[1]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_1[1]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X419 adc_array_wafflecap_8_8_1[1]/adc_array_circuit_150n_0/vint2 col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X420 adc_array_wafflecap_8_Dummy_1[6]/adc_array_circuit_150n_0/vint2 col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X421 adc_array_wafflecap_8_8_0[12|0]/adc_array_circuit_150n_0/vdrv row_n[13] adc_array_wafflecap_8_8_0[12|0]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X422 adc_array_wafflecap_8_8_0[12|10]/adc_array_circuit_150n_0/vdrv row_n[13] adc_array_wafflecap_8_8_0[12|10]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X423 adc_array_wafflecap_8_8_0[10|21]/adc_array_circuit_150n_0/vint2 rowon_n[11] adc_array_wafflecap_8_8_0[10|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X424 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.64e+07u l=1.6e+07u
X425 adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X426 adc_array_wafflecap_8_8_0[9|2]/adc_array_circuit_150n_0/vint2 rowon_n[10] adc_array_wafflecap_8_8_0[9|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X427 adc_array_wafflecap_8_8_0[9|12]/adc_array_circuit_150n_0/vint2 rowon_n[10] adc_array_wafflecap_8_8_0[9|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X428 adc_array_wafflecap_8_8_0[6|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X429 adc_array_wafflecap_8_8_0[2|5]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|5]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X430 adc_array_wafflecap_8_Dummy_8[4]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_8[4]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X431 adc_array_wafflecap_8_Dummy_3[1]/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_3[1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X432 adc_array_wafflecap_8_Dummy_4[13]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X433 vcm adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|9]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X434 adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X435 adc_array_wafflecap_8_Dummy_4[3]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X436 VSS sample_n adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X437 adc_array_wafflecap_8_8_0[8|6]/adc_array_circuit_150n_0/vint2 rowon_n[9] adc_array_wafflecap_8_8_0[8|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X438 adc_array_wafflecap_8_8_0[8|16]/adc_array_circuit_150n_0/vint2 rowon_n[9] adc_array_wafflecap_8_8_0[8|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X439 adc_array_wafflecap_8_8_1[7]/adc_array_circuit_150n_0/vint2 rowon_n[0] adc_array_wafflecap_8_8_1[7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X440 adc_array_wafflecap_8_8_0[1|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X441 vcm adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|3]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X442 vcm adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|13]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X443 adc_array_wafflecap_8_8_0[4|21]/adc_array_circuit_150n_0/vdrv row_n[5] adc_array_wafflecap_8_8_0[4|21]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X444 adc_array_wafflecap_8_8_1[24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_1[24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X445 vcm adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|29]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X446 adc_array_wafflecap_8_8_0[1|17]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|17]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X447 adc_array_wafflecap_8_8_0[2|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X448 VDD rowon_n[9] adc_array_wafflecap_8_8_0[8|21]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X449 adc_array_wafflecap_8_8_0[6|25]/adc_array_circuit_150n_0/vint2 col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X450 adc_array_wafflecap_8_8_0[5|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X451 VDD rowon_n[3] adc_array_wafflecap_8_8_0[2|10]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X452 VSS VDD adc_array_wafflecap_8_Dummy_4[20]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X453 VDD rowon_n[8] adc_array_wafflecap_8_8_0[7|2]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X454 VDD rowon_n[8] adc_array_wafflecap_8_8_0[7|12]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X455 VSS row_n[15] adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X456 adc_array_wafflecap_8_8_0[11|20]/adc_array_circuit_150n_0/vint2 col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X457 adc_array_wafflecap_8_8_0[4|6]/adc_array_circuit_150n_0/vint1 col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X458 adc_array_wafflecap_8_8_0[4|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X459 adc_array_wafflecap_8_8_1[23]/adc_array_circuit_150n_0/vint2 col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X460 adc_array_wafflecap_8_8_0[0|30]/adc_array_circuit_150n_0/vint2 rowon_n[1] adc_array_wafflecap_8_8_0[0|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X461 adc_array_wafflecap_8_8_0[0|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X462 VSS row_n[11] adc_array_wafflecap_8_8_0[10|10]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X463 adc_array_wafflecap_8_8_0[5|14]/adc_array_circuit_150n_0/vint2 col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X464 VSS row_n[11] adc_array_wafflecap_8_8_0[10|0]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X465 adc_array_wafflecap_8_8_0[6|25]/adc_array_circuit_150n_0/vdrv row_n[7] adc_array_wafflecap_8_8_0[6|25]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X466 adc_array_wafflecap_8_8_0[13|19]/adc_array_circuit_150n_0/vint1 col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X467 adc_array_wafflecap_8_8_0[11|7]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|7]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X468 adc_array_wafflecap_8_8_0[7|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X469 adc_array_wafflecap_8_8_0[6|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X470 adc_array_wafflecap_8_8_0[5|4]/adc_array_circuit_150n_0/vdrv row_n[6] adc_array_wafflecap_8_8_0[5|4]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X471 VDD VDD adc_array_wafflecap_8_Dummy_4[14]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X472 adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/vint1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X473 adc_array_wafflecap_8_8_0[9|29]/adc_array_circuit_150n_0/vdrv row_n[10] adc_array_wafflecap_8_8_0[9|29]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X474 VSS row_n[0] adc_array_wafflecap_8_8_1[8]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X475 VDD VDD adc_array_wafflecap_8_Dummy_4[4]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X476 VDD VSS adc_array_wafflecap_8_Dummy_3[5]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X477 adc_array_wafflecap_8_Dummy_7/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X478 adc_array_wafflecap_8_8_0[9|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X479 adc_array_wafflecap_8_8_0[8|10]/adc_array_circuit_150n_0/vint1 col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X480 adc_array_wafflecap_8_8_0[2|11]/adc_array_circuit_150n_0/vint1 col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X481 adc_array_wafflecap_8_8_0[2|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X482 adc_array_wafflecap_8_Dummy_1[4]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X483 adc_array_wafflecap_8_8_0[8|0]/adc_array_circuit_150n_0/vint1 col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X484 adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X485 adc_array_wafflecap_8_Dummy_4[9]/adc_array_circuit_150n_0/vint2 col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X486 VSS row_n[4] adc_array_wafflecap_8_8_0[3|20]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X487 adc_array_wafflecap_8_8_0[3|18]/adc_array_circuit_150n_0/vint2 col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X488 vcm VSS adc_array_wafflecap_8_Dummy_8[0]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X489 adc_array_wafflecap_8_8_0[13|8]/adc_array_circuit_150n_0/vdrv row_n[14] adc_array_wafflecap_8_8_0[13|8]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X490 adc_array_wafflecap_8_8_0[11|19]/adc_array_circuit_150n_0/vint2 rowon_n[12] adc_array_wafflecap_8_8_0[11|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X491 adc_array_wafflecap_8_8_0[10|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X492 vcm adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|8]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X493 adc_array_wafflecap_8_8_0[6|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X494 adc_array_wafflecap_8_8_0[4|30]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|30]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X495 adc_array_wafflecap_8_8_0[4|12]/adc_array_circuit_150n_0/vint2 rowon_n[5] adc_array_wafflecap_8_8_0[4|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X496 adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X497 adc_array_wafflecap_8_8_0[14|21]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|21]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X498 adc_array_wafflecap_8_8_0[10|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X499 adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/vint2 rowon_n[11] adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X500 VDD rowon_n[5] adc_array_wafflecap_8_8_0[4|2]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X501 adc_array_wafflecap_8_8_0[4|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X502 adc_array_wafflecap_8_8_1[26]/adc_array_circuit_150n_0/vdrv row_n[0] adc_array_wafflecap_8_8_1[26]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X503 adc_array_wafflecap_8_8_0[13|25]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|25]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X504 adc_array_wafflecap_8_8_0[11|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X505 adc_array_wafflecap_8_8_0[6|6]/adc_array_circuit_150n_0/vint2 rowon_n[7] adc_array_wafflecap_8_8_0[6|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X506 adc_array_wafflecap_8_8_0[4|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X507 adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/vint2 VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X508 adc_array_wafflecap_8_8_0[12|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X509 adc_array_wafflecap_8_8_0[12|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X510 vcm adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|9]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X511 VSS row_n[6] adc_array_wafflecap_8_8_0[5|24]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X512 VSS row_n[2] adc_array_wafflecap_8_8_0[1|25]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X513 VSS row_n[10] adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X514 VDD rowon_n[9] adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X515 VSS VDD adc_array_wafflecap_8_Dummy_4[31]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X516 VDD rowon_n[12] adc_array_wafflecap_8_8_0[11|30]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X517 adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/vint2 col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X518 VDD rowon_n[7] adc_array_wafflecap_8_8_0[6|6]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X519 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.64e+07u l=1.6e+07u
X520 VDD rowon_n[12] adc_array_wafflecap_8_8_0[11|8]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X521 VSS row_n[5] adc_array_wafflecap_8_8_0[4|13]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X522 vcm VSS adc_array_wafflecap_8_1_0/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X523 adc_array_wafflecap_8_Dummy_2[0]/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_2[0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X524 adc_array_wafflecap_8_8_0[1|25]/adc_array_circuit_150n_0/vint1 col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X525 vcm adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|23]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X526 adc_array_wafflecap_8_Dummy_4[18]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X527 VSS row_n[12] adc_array_wafflecap_8_8_0[11|8]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X528 adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/vint1 col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X529 vcm adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|1]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X530 adc_array_wafflecap_8_8_0[4|3]/adc_array_circuit_150n_0/vint1 col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X531 adc_array_wafflecap_8_8_0[13|30]/adc_array_circuit_150n_0/vint1 col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X532 adc_array_wafflecap_8_8_0[11|18]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|18]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X533 vcm adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|26]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X534 adc_array_wafflecap_8_8_0[7|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X535 VSS row_n[15] adc_array_wafflecap_8_8_0[14|6]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X536 adc_array_wafflecap_8_Dummy_1[0]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_1[0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X537 adc_array_wafflecap_8_8_0[10|7]/adc_array_circuit_150n_0/vint2 col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X538 adc_array_wafflecap_8_Dummy_4[20]/adc_array_circuit_150n_0/vint2 col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X539 adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X540 vcm adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|6]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X541 adc_array_wafflecap_8_8_0[2|19]/adc_array_circuit_150n_0/vint2 rowon_n[3] adc_array_wafflecap_8_8_0[2|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X542 adc_array_wafflecap_8_8_0[12|6]/adc_array_circuit_150n_0/vint1 col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X543 adc_array_wafflecap_8_8_0[7|29]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|29]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X544 adc_array_wafflecap_8_4_0/adc_array_circuit_150n_0/vint2 en_n_bit[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X545 VSS VSS adc_array_wafflecap_8_Dummy_2[1]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X546 adc_array_wafflecap_8_8_0[2|7]/adc_array_circuit_150n_0/vint2 col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X547 adc_array_wafflecap_8_Dummy_4[32]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[32]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X548 vcm adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|28]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X549 adc_array_wafflecap_8_8_1[19]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[19]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X550 vcm adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|27]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X551 VSS row_n[3] adc_array_wafflecap_8_8_0[2|17]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X552 vcm adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X553 adc_array_wafflecap_8_8_0[9|20]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|20]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X554 adc_array_wafflecap_8_8_0[8|7]/adc_array_circuit_150n_0/vdrv row_n[9] adc_array_wafflecap_8_8_0[8|7]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X555 adc_array_wafflecap_8_8_0[6|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X556 VDD rowon_n[6] adc_array_wafflecap_8_8_0[5|21]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X557 adc_array_wafflecap_8_Dummy_0[0]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_0[0]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X558 adc_array_wafflecap_8_8_1[29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X559 adc_array_wafflecap_8_8_0[1|11]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|11]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X560 adc_array_wafflecap_8_8_0[11|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X561 vcm adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|17]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X562 adc_array_wafflecap_8_8_0[5|10]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|10]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X563 adc_array_wafflecap_8_8_0[13|19]/adc_array_circuit_150n_0/vdrv row_n[14] adc_array_wafflecap_8_8_0[13|19]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X564 adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X565 vcm adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|19]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X566 VDD rowon_n[1] adc_array_wafflecap_8_8_0[0|19]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X567 adc_array_wafflecap_8_8_0[0|17]/adc_array_circuit_150n_0/vint1 col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X568 adc_array_wafflecap_8_8_0[0|7]/adc_array_circuit_150n_0/vdrv row_n[1] adc_array_wafflecap_8_8_0[0|7]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X569 adc_array_wafflecap_8_8_0[4|23]/adc_array_circuit_150n_0/vint2 rowon_n[5] adc_array_wafflecap_8_8_0[4|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X570 adc_array_wafflecap_8_8_0[0|24]/adc_array_circuit_150n_0/vint2 rowon_n[1] adc_array_wafflecap_8_8_0[0|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X571 adc_array_wafflecap_8_8_0[14|28]/adc_array_circuit_150n_0/vint2 rowon_n[15] adc_array_wafflecap_8_8_0[14|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X572 adc_array_wafflecap_8_8_0[13|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X573 VSS row_n[7] adc_array_wafflecap_8_8_0[6|28]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X574 adc_array_wafflecap_8_8_0[5|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X575 adc_array_wafflecap_8_8_0[0|12]/adc_array_circuit_150n_0/vint2 col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X576 adc_array_wafflecap_8_8_0[13|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X577 vcm VSS adc_array_wafflecap_8_Dummy_6/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X578 adc_array_wafflecap_8_8_0[13|10]/adc_array_circuit_150n_0/vint2 rowon_n[14] adc_array_wafflecap_8_8_0[13|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X579 adc_array_wafflecap_8_8_0[12|25]/adc_array_circuit_150n_0/vint2 col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X580 VSS row_n[11] adc_array_wafflecap_8_8_0[10|29]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X581 adc_array_wafflecap_8_8_0[7|26]/adc_array_circuit_150n_0/vint2 col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X582 adc_array_wafflecap_8_8_0[0|3]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|3]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X583 adc_array_wafflecap_8_8_0[13|0]/adc_array_circuit_150n_0/vint2 rowon_n[14] adc_array_wafflecap_8_8_0[13|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X584 adc_array_wafflecap_8_8_0[4|2]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|2]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X585 adc_array_wafflecap_8_8_0[3|15]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|15]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X586 adc_array_wafflecap_8_8_0[12|12]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|12]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X587 VDD en_n_bit[0] adc_array_wafflecap_8_1_0/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X588 adc_array_wafflecap_8_8_0[14|24]/adc_array_circuit_150n_0/vint1 col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X589 adc_array_wafflecap_8_8_0[12|2]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|2]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X590 VDD rowon_n[13] adc_array_wafflecap_8_8_0[12|28]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X591 adc_array_wafflecap_8_8_0[11|21]/adc_array_circuit_150n_0/vdrv row_n[12] adc_array_wafflecap_8_8_0[11|21]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X592 adc_array_wafflecap_8_8_0[6|28]/adc_array_circuit_150n_0/vint1 col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X593 adc_array_wafflecap_8_Dummy_1[3]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_1[3]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X594 adc_array_wafflecap_8_8_0[10|25]/adc_array_circuit_150n_0/vdrv row_n[11] adc_array_wafflecap_8_8_0[10|25]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X595 adc_array_wafflecap_8_8_0[8|29]/adc_array_circuit_150n_0/vint1 col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X596 adc_array_wafflecap_8_8_0[4|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X597 adc_array_wafflecap_8_8_0[14|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X598 adc_array_wafflecap_8_8_0[3|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X599 adc_array_wafflecap_8_Dummy_4[28]/adc_array_circuit_150n_0/vint2 col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X600 adc_array_wafflecap_8_8_0[9|15]/adc_array_circuit_150n_0/vint1 col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X601 vcm adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|24]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X602 adc_array_wafflecap_8_8_0[9|5]/adc_array_circuit_150n_0/vint1 col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X603 adc_array_wafflecap_8_8_0[8|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X604 adc_array_wafflecap_8_Dummy_3[3]/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_3[3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X605 VSS row_n[15] adc_array_wafflecap_8_8_0[14|17]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X606 adc_array_wafflecap_8_8_0[10|18]/adc_array_circuit_150n_0/vint2 col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X607 adc_array_wafflecap_8_8_1[9]/adc_array_circuit_150n_0/vint2 rowon_n[0] adc_array_wafflecap_8_8_1[9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X608 adc_array_wafflecap_8_8_0[1|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X609 vcm adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X610 adc_array_wafflecap_8_8_0[4|23]/adc_array_circuit_150n_0/vdrv row_n[5] adc_array_wafflecap_8_8_0[4|23]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X611 adc_array_wafflecap_8_8_0[4|24]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|24]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X612 adc_array_wafflecap_8_8_0[13|27]/adc_array_circuit_150n_0/vdrv row_n[14] adc_array_wafflecap_8_8_0[13|27]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X613 vcm adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|27]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X614 adc_array_wafflecap_8_8_0[2|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X615 VSS sample adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X616 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X617 adc_array_wafflecap_8_8_1[20]/adc_array_circuit_150n_0/vdrv row_n[0] adc_array_wafflecap_8_8_1[20]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X618 adc_array_wafflecap_8_8_0[14|3]/adc_array_circuit_150n_0/vdrv row_n[15] adc_array_wafflecap_8_8_0[14|3]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X619 adc_array_wafflecap_8_8_0[14|13]/adc_array_circuit_150n_0/vdrv row_n[15] adc_array_wafflecap_8_8_0[14|13]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X620 adc_array_wafflecap_8_8_0[12|17]/adc_array_circuit_150n_0/vint1 col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X621 adc_array_wafflecap_8_8_0[12|24]/adc_array_circuit_150n_0/vint2 rowon_n[13] adc_array_wafflecap_8_8_0[12|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X622 vcm adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|7]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X623 adc_array_wafflecap_8_8_0[13|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X624 adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X625 adc_array_wafflecap_8_8_0[8|18]/adc_array_circuit_150n_0/vdrv row_n[9] adc_array_wafflecap_8_8_0[8|18]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X626 VSS row_n[9] adc_array_wafflecap_8_8_0[8|25]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X627 adc_array_wafflecap_8_8_0[4|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X628 adc_array_wafflecap_8_8_0[0|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X629 adc_array_wafflecap_8_8_0[1|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X630 adc_array_wafflecap_8_8_0[2|4]/adc_array_circuit_150n_0/vint2 col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X631 vcm adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|16]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X632 adc_array_wafflecap_8_8_0[9|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X633 adc_array_wafflecap_8_8_1[5]/adc_array_circuit_150n_0/vint1 col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X634 vcm adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|6]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X635 VDD rowon_n[11] adc_array_wafflecap_8_8_0[10|24]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X636 adc_array_wafflecap_8_8_0[5|27]/adc_array_circuit_150n_0/vint2 rowon_n[6] adc_array_wafflecap_8_8_0[5|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X637 VSS row_n[0] adc_array_wafflecap_8_8_1[10]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X638 adc_array_wafflecap_8_8_0[1|16]/adc_array_circuit_150n_0/vint2 col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X639 adc_array_wafflecap_8_Dummy_4[27]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X640 adc_array_wafflecap_8_8_0[2|27]/adc_array_circuit_150n_0/vdrv row_n[3] adc_array_wafflecap_8_8_0[2|27]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X641 adc_array_wafflecap_8_8_0[2|28]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|28]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X642 adc_array_wafflecap_8_Dummy_3[4]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_3[4]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X643 adc_array_wafflecap_8_8_0[0|4]/adc_array_circuit_150n_0/vdrv row_n[1] adc_array_wafflecap_8_8_0[0|4]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X644 adc_array_wafflecap_8_8_0[14|17]/adc_array_circuit_150n_0/vint2 rowon_n[15] adc_array_wafflecap_8_8_0[14|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X645 adc_array_wafflecap_8_8_0[13|23]/adc_array_circuit_150n_0/vint2 col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X646 VSS row_n[12] adc_array_wafflecap_8_8_0[11|27]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X647 adc_array_wafflecap_8_8_1[1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X648 adc_array_wafflecap_8_8_0[2|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X649 adc_array_wafflecap_8_Dummy_1[6]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X650 VSS row_n[13] adc_array_wafflecap_8_8_0[12|13]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X651 VSS row_n[13] adc_array_wafflecap_8_8_0[12|3]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X652 VDD rowon_n[6] adc_array_wafflecap_8_8_0[5|12]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X653 adc_array_wafflecap_8_Dummy_4[23]/adc_array_circuit_150n_0/vint1 col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X654 adc_array_wafflecap_8_8_0[13|10]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|10]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X655 VDD rowon_n[14] adc_array_wafflecap_8_8_0[13|26]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X656 adc_array_wafflecap_8_8_0[9|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X657 adc_array_wafflecap_8_8_0[8|14]/adc_array_circuit_150n_0/vint2 col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X658 VSS row_n[4] adc_array_wafflecap_8_8_0[3|22]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X659 adc_array_wafflecap_8_8_0[1|16]/adc_array_circuit_150n_0/vdrv row_n[2] adc_array_wafflecap_8_8_0[1|16]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X660 adc_array_wafflecap_8_8_0[13|0]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|0]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X661 VDD rowon_n[13] adc_array_wafflecap_8_8_0[12|17]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X662 adc_array_wafflecap_8_8_0[8|4]/adc_array_circuit_150n_0/vint2 col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X663 VSS row_n[7] adc_array_wafflecap_8_8_0[6|0]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X664 adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/vint2 rowon_n[4] adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X665 adc_array_wafflecap_8_8_0[8|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X666 adc_array_wafflecap_8_8_0[10|13]/adc_array_circuit_150n_0/vint1 col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X667 VSS row_n[10] adc_array_wafflecap_8_8_0[9|16]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X668 adc_array_wafflecap_8_8_0[6|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X669 adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X670 adc_array_wafflecap_8_8_0[4|14]/adc_array_circuit_150n_0/vint2 rowon_n[5] adc_array_wafflecap_8_8_0[4|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X671 adc_array_wafflecap_8_8_0[10|3]/adc_array_circuit_150n_0/vint1 col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X672 VDD rowon_n[5] adc_array_wafflecap_8_8_0[4|4]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X673 vcm adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|20]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X674 vcm adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|21]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X675 vcm adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|20]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X676 adc_array_wafflecap_8_8_0[11|16]/adc_array_circuit_150n_0/vint2 col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X677 adc_array_wafflecap_8_8_0[6|0]/adc_array_circuit_150n_0/vint1 col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X678 adc_array_wafflecap_8_8_0[4|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X679 VSS sample_n adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X680 VDD rowon_n[0] adc_array_wafflecap_8_8_1[1]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X681 adc_array_wafflecap_8_8_0[9|12]/adc_array_circuit_150n_0/vdrv row_n[10] adc_array_wafflecap_8_8_0[9|12]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X682 adc_array_wafflecap_8_8_0[8|25]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|25]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X683 adc_array_wafflecap_8_8_0[7|16]/adc_array_circuit_150n_0/vint1 col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X684 adc_array_wafflecap_8_8_0[7|23]/adc_array_circuit_150n_0/vint2 rowon_n[8] adc_array_wafflecap_8_8_0[7|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X685 vcm adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|11]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X686 adc_array_wafflecap_8_8_0[5|13]/adc_array_circuit_150n_0/vint1 col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X687 adc_array_wafflecap_8_8_0[9|2]/adc_array_circuit_150n_0/vdrv row_n[10] adc_array_wafflecap_8_8_0[9|2]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X688 adc_array_wafflecap_8_Dummy_4[12]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[12]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X689 adc_array_wafflecap_8_8_0[7|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X690 adc_array_wafflecap_8_8_0[7|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X691 adc_array_wafflecap_8_Dummy_4[2]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[2]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X692 adc_array_wafflecap_8_8_0[14|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X693 adc_array_wafflecap_8_8_0[13|22]/adc_array_circuit_150n_0/vint2 rowon_n[14] adc_array_wafflecap_8_8_0[13|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X694 adc_array_wafflecap_8_8_0[12|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X695 adc_array_wafflecap_8_8_0[12|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X696 vcm adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|1]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X697 vcm adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|11]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X698 VSS row_n[2] adc_array_wafflecap_8_8_0[1|26]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X699 vcm adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|15]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X700 adc_array_wafflecap_8_8_0[4|29]/adc_array_circuit_150n_0/vint2 col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X701 adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X702 adc_array_wafflecap_8_8_0[10|29]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|29]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X703 vcm adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|5]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X704 VSS row_n[5] adc_array_wafflecap_8_8_0[4|15]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X705 vcm VSS adc_array_wafflecap_8_Dummy_3[1]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X706 vcm adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|25]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X707 vcm adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|3]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X708 adc_array_wafflecap_8_8_0[4|5]/adc_array_circuit_150n_0/vint1 col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X709 vcm adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|4]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X710 VSS row_n[13] adc_array_wafflecap_8_8_0[12|21]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X711 adc_array_wafflecap_8_8_0[14|5]/adc_array_circuit_150n_0/vint2 rowon_n[15] adc_array_wafflecap_8_8_0[14|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X712 adc_array_wafflecap_8_8_0[14|15]/adc_array_circuit_150n_0/vint2 rowon_n[15] adc_array_wafflecap_8_8_0[14|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X713 adc_array_wafflecap_8_8_0[8|22]/adc_array_circuit_150n_0/vint2 col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X714 adc_array_wafflecap_8_8_0[1|26]/adc_array_circuit_150n_0/vint1 col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X715 adc_array_wafflecap_8_8_0[3|7]/adc_array_circuit_150n_0/vdrv row_n[4] adc_array_wafflecap_8_8_0[3|7]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X716 VDD rowon_n[4] adc_array_wafflecap_8_8_0[3|19]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X717 adc_array_wafflecap_8_Dummy_1[2]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_1[2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X718 adc_array_wafflecap_8_8_1[2]/adc_array_circuit_150n_0/vint1 col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X719 adc_array_wafflecap_8_8_0[3|8]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|8]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X720 adc_array_wafflecap_8_8_0[3|17]/adc_array_circuit_150n_0/vint1 col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X721 VDD rowon_n[15] adc_array_wafflecap_8_8_0[14|20]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X722 vcm adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|17]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X723 VSS row_n[8] adc_array_wafflecap_8_8_0[7|2]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X724 VSS row_n[8] adc_array_wafflecap_8_8_0[7|12]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X725 adc_array_wafflecap_8_8_0[3|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X726 adc_array_wafflecap_8_8_0[10|21]/adc_array_circuit_150n_0/vint1 col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X727 VDD rowon_n[13] adc_array_wafflecap_8_8_0[12|15]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X728 adc_array_wafflecap_8_Dummy_2[5]/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_2[5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X729 VDD rowon_n[13] adc_array_wafflecap_8_8_0[12|5]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X730 adc_array_wafflecap_8_Dummy_1[1]/adc_array_circuit_150n_0/vint2 col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X731 adc_array_wafflecap_8_8_0[2|21]/adc_array_circuit_150n_0/vint2 rowon_n[3] adc_array_wafflecap_8_8_0[2|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X732 adc_array_wafflecap_8_8_0[10|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X733 adc_array_wafflecap_8_8_1[21]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[21]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X734 adc_array_wafflecap_8_8_0[6|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X735 VDD rowon_n[6] adc_array_wafflecap_8_8_0[5|23]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X736 adc_array_wafflecap_8_8_0[2|0]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|0]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X737 adc_array_wafflecap_8_1_1/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_1_1/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X738 adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X739 adc_array_wafflecap_8_8_0[12|10]/adc_array_circuit_150n_0/vint2 col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X740 adc_array_wafflecap_8_8_0[5|12]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|12]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X741 adc_array_wafflecap_8_8_0[1|13]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|13]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X742 adc_array_wafflecap_8_8_0[12|0]/adc_array_circuit_150n_0/vint2 col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X743 VDD sample adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X744 VDD rowon_n[1] adc_array_wafflecap_8_8_0[0|21]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X745 adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/vdrv row_n[15] adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X746 adc_array_wafflecap_8_8_1[19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_1[19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X747 vcm adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[17]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X748 adc_array_wafflecap_8_8_0[14|9]/adc_array_circuit_150n_0/vint1 col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X749 adc_array_wafflecap_8_8_0[11|6]/adc_array_circuit_150n_0/vdrv row_n[12] adc_array_wafflecap_8_8_0[11|6]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X750 adc_array_wafflecap_8_8_0[6|20]/adc_array_circuit_150n_0/vint2 col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X751 VSS row_n[7] adc_array_wafflecap_8_8_0[6|30]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X752 adc_array_wafflecap_8_8_0[5|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X753 adc_array_wafflecap_8_8_0[4|25]/adc_array_circuit_150n_0/vint2 rowon_n[5] adc_array_wafflecap_8_8_0[4|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X754 vcm adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X755 adc_array_wafflecap_8_8_0[14|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X756 adc_array_wafflecap_8_8_0[14|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X757 adc_array_wafflecap_8_8_0[10|0]/adc_array_circuit_150n_0/vdrv row_n[11] adc_array_wafflecap_8_8_0[10|0]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X758 adc_array_wafflecap_8_8_0[10|10]/adc_array_circuit_150n_0/vdrv row_n[11] adc_array_wafflecap_8_8_0[10|10]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X759 adc_array_wafflecap_8_8_0[9|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X760 adc_array_wafflecap_8_8_0[8|21]/adc_array_circuit_150n_0/vint2 rowon_n[9] adc_array_wafflecap_8_8_0[8|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X761 adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X762 adc_array_wafflecap_8_8_0[8|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X763 adc_array_wafflecap_8_8_0[7|2]/adc_array_circuit_150n_0/vint2 rowon_n[8] adc_array_wafflecap_8_8_0[7|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X764 adc_array_wafflecap_8_8_0[7|12]/adc_array_circuit_150n_0/vint2 rowon_n[8] adc_array_wafflecap_8_8_0[7|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X765 adc_array_wafflecap_8_8_0[0|5]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|5]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X766 adc_array_wafflecap_8_8_0[13|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X767 vcm adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|9]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X768 adc_array_wafflecap_8_8_0[8|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X769 adc_array_wafflecap_8_8_0[13|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X770 VSS sample_n adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X771 adc_array_wafflecap_8_8_0[5|9]/adc_array_circuit_150n_0/vint2 col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X772 adc_array_wafflecap_8_8_0[6|20]/adc_array_circuit_150n_0/vdrv row_n[7] adc_array_wafflecap_8_8_0[6|20]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X773 adc_array_wafflecap_8_8_0[2|21]/adc_array_circuit_150n_0/vdrv row_n[3] adc_array_wafflecap_8_8_0[2|21]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X774 adc_array_wafflecap_8_8_0[6|30]/adc_array_circuit_150n_0/vint1 col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X775 adc_array_wafflecap_8_8_0[4|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X776 vcm adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|29]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X777 adc_array_wafflecap_8_8_0[0|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X778 adc_array_wafflecap_8_8_0[3|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X779 VSS row_n[14] adc_array_wafflecap_8_8_0[13|19]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X780 adc_array_wafflecap_8_8_0[7|2]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|2]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X781 adc_array_wafflecap_8_8_0[7|12]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|12]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X782 adc_array_wafflecap_8_Dummy_4[14]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X783 VSS row_n[13] adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X784 adc_array_wafflecap_8_8_0[9|29]/adc_array_circuit_150n_0/vint2 col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X785 adc_array_wafflecap_8_Dummy_4[4]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X786 adc_array_wafflecap_8_8_0[2|6]/adc_array_circuit_150n_0/vint1 col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X787 adc_array_wafflecap_8_8_0[2|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X788 adc_array_wafflecap_8_4_0/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X789 adc_array_wafflecap_8_Dummy_3[5]/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_3[5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X790 adc_array_wafflecap_8_8_0[4|1]/adc_array_circuit_150n_0/vint2 col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X791 VDD VDD adc_array_wafflecap_8_Dummy_4[19]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X792 VSS row_n[9] adc_array_wafflecap_8_8_0[8|10]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X793 adc_array_wafflecap_8_8_0[3|14]/adc_array_circuit_150n_0/vint2 col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X794 adc_array_wafflecap_8_8_0[14|5]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|5]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X795 VDD rowon_n[15] adc_array_wafflecap_8_8_0[14|9]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X796 adc_array_wafflecap_8_8_0[14|15]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|15]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X797 VDD rowon_n[15] adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X798 adc_array_wafflecap_8_8_0[11|28]/adc_array_circuit_150n_0/vint1 col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X799 VSS row_n[9] adc_array_wafflecap_8_8_0[8|0]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X800 adc_array_wafflecap_8_8_0[4|25]/adc_array_circuit_150n_0/vdrv row_n[5] adc_array_wafflecap_8_8_0[4|25]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X801 adc_array_wafflecap_8_8_0[4|26]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|26]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X802 adc_array_wafflecap_8_8_0[3|4]/adc_array_circuit_150n_0/vdrv row_n[4] adc_array_wafflecap_8_8_0[3|4]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X803 VDD rowon_n[14] adc_array_wafflecap_8_8_0[13|13]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X804 adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/vint1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X805 adc_array_wafflecap_8_8_0[7|29]/adc_array_circuit_150n_0/vdrv row_n[8] adc_array_wafflecap_8_8_0[7|29]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X806 VDD rowon_n[14] adc_array_wafflecap_8_8_0[13|3]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X807 adc_array_wafflecap_8_8_1[22]/adc_array_circuit_150n_0/vdrv row_n[0] adc_array_wafflecap_8_8_1[22]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X808 adc_array_wafflecap_8_8_0[4|7]/adc_array_circuit_150n_0/vint2 rowon_n[5] adc_array_wafflecap_8_8_0[4|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X809 adc_array_wafflecap_8_8_0[0|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X810 adc_array_wafflecap_8_8_0[4|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X811 adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X812 adc_array_wafflecap_8_8_0[13|8]/adc_array_circuit_150n_0/vint2 col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X813 adc_array_wafflecap_8_8_0[8|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X814 adc_array_wafflecap_8_8_0[6|1]/adc_array_circuit_150n_0/vint2 rowon_n[7] adc_array_wafflecap_8_8_0[6|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X815 adc_array_wafflecap_8_8_1[26]/adc_array_circuit_150n_0/vint2 col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X816 adc_array_wafflecap_8_Dummy_4[31]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[31]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X817 vcm adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|30]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X818 VSS row_n[6] adc_array_wafflecap_8_8_0[5|19]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X819 VSS row_n[2] adc_array_wafflecap_8_8_0[1|20]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X820 adc_array_wafflecap_8_8_0[5|29]/adc_array_circuit_150n_0/vint2 rowon_n[6] adc_array_wafflecap_8_8_0[5|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X821 adc_array_wafflecap_8_8_0[1|18]/adc_array_circuit_150n_0/vint2 col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X822 adc_array_wafflecap_8_Dummy_4[8]/adc_array_circuit_150n_0/vint1 col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X823 vcm VSS adc_array_wafflecap_8_Dummy_4[30]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X824 adc_array_wafflecap_8_8_0[9|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X825 adc_array_wafflecap_8_8_0[5|17]/adc_array_circuit_150n_0/vint2 col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X826 adc_array_wafflecap_8_8_0[8|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X827 adc_array_wafflecap_8_8_0[2|30]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|30]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X828 adc_array_wafflecap_8_8_1[3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X829 adc_array_wafflecap_8_8_0[2|12]/adc_array_circuit_150n_0/vint2 rowon_n[3] adc_array_wafflecap_8_8_0[2|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X830 adc_array_wafflecap_8_Dummy_4[25]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X831 adc_array_wafflecap_8_8_0[12|21]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|21]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X832 adc_array_wafflecap_8_8_0[8|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X833 adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/vint2 rowon_n[9] adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X834 adc_array_wafflecap_8_8_0[2|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X835 adc_array_wafflecap_8_8_0[11|25]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|25]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X836 VDD rowon_n[7] adc_array_wafflecap_8_8_0[6|1]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X837 VDD rowon_n[3] adc_array_wafflecap_8_8_0[2|2]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X838 VDD rowon_n[6] adc_array_wafflecap_8_8_0[5|14]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X839 VSS row_n[5] adc_array_wafflecap_8_8_0[4|8]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X840 adc_array_wafflecap_8_8_0[1|20]/adc_array_circuit_150n_0/vint1 col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X841 adc_array_wafflecap_8_8_0[2|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X842 adc_array_wafflecap_8_8_0[10|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X843 adc_array_wafflecap_8_8_0[10|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X844 VSS row_n[4] adc_array_wafflecap_8_8_0[3|24]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X845 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X846 adc_array_wafflecap_8_8_0[1|18]/adc_array_circuit_150n_0/vdrv row_n[2] adc_array_wafflecap_8_8_0[1|18]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X847 VSS row_n[8] adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X848 VSS row_n[7] adc_array_wafflecap_8_8_0[6|2]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X849 VDD rowon_n[1] adc_array_wafflecap_8_8_0[0|12]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X850 adc_array_wafflecap_8_8_0[8|10]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|10]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X851 VSS row_n[14] adc_array_wafflecap_8_8_0[13|30]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X852 adc_array_wafflecap_8_8_0[8|0]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|0]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X853 adc_array_wafflecap_8_8_0[4|16]/adc_array_circuit_150n_0/vint2 rowon_n[5] adc_array_wafflecap_8_8_0[4|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X854 VDD rowon_n[10] adc_array_wafflecap_8_8_0[9|30]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X855 VDD rowon_n[5] adc_array_wafflecap_8_8_0[4|6]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X856 VDD rowon_n[10] adc_array_wafflecap_8_8_0[9|8]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X857 vcm adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|22]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X858 vcm adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|23]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X859 VSS row_n[3] adc_array_wafflecap_8_8_0[2|13]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X860 adc_array_wafflecap_8_Dummy_4[14]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[14]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X861 VDD VDD adc_array_wafflecap_8_Dummy_4[30]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X862 adc_array_wafflecap_8_8_0[13|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X863 adc_array_wafflecap_8_8_0[5|29]/adc_array_circuit_150n_0/vdrv row_n[6] adc_array_wafflecap_8_8_0[5|29]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X864 adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X865 vcm adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|1]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X866 adc_array_wafflecap_8_8_0[2|3]/adc_array_circuit_150n_0/vint1 col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X867 adc_array_wafflecap_8_Dummy_4[4]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[4]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X868 VDD VDD adc_array_wafflecap_8_Dummy_4[8]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X869 adc_array_wafflecap_8_8_0[6|2]/adc_array_circuit_150n_0/vint1 col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X870 vcm adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|13]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X871 VDD rowon_n[0] adc_array_wafflecap_8_8_1[3]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X872 vcm adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|26]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X873 adc_array_wafflecap_8_8_0[5|15]/adc_array_circuit_150n_0/vint1 col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X874 VSS row_n[13] adc_array_wafflecap_8_8_0[12|6]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X875 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.64e+07u l=1.6e+07u
X876 adc_array_wafflecap_8_8_0[0|13]/adc_array_circuit_150n_0/vint1 col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X877 adc_array_wafflecap_8_8_0[8|7]/adc_array_circuit_150n_0/vint2 col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X878 adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/vint2 col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X879 adc_array_wafflecap_8_8_0[14|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X880 adc_array_wafflecap_8_8_0[13|19]/adc_array_circuit_150n_0/vint2 col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X881 vcm adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|5]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X882 adc_array_wafflecap_8_8_0[4|18]/adc_array_circuit_150n_0/vint2 rowon_n[5] adc_array_wafflecap_8_8_0[4|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X883 adc_array_wafflecap_8_8_0[0|19]/adc_array_circuit_150n_0/vint2 rowon_n[1] adc_array_wafflecap_8_8_0[0|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X884 vcm adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|6]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X885 adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X886 adc_array_wafflecap_8_8_0[11|15]/adc_array_circuit_150n_0/vdrv row_n[12] adc_array_wafflecap_8_8_0[11|15]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X887 adc_array_wafflecap_8_8_0[10|6]/adc_array_circuit_150n_0/vint1 col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X888 adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X889 adc_array_wafflecap_8_8_0[0|7]/adc_array_circuit_150n_0/vint2 col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X890 adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X891 adc_array_wafflecap_8_8_0[11|5]/adc_array_circuit_150n_0/vdrv row_n[12] adc_array_wafflecap_8_8_0[11|5]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X892 vcm adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|28]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X893 VSS row_n[5] adc_array_wafflecap_8_8_0[4|16]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X894 vcm VSS adc_array_wafflecap_8_Dummy_3[2]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X895 VSS row_n[1] adc_array_wafflecap_8_8_0[0|17]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X896 VDD rowon_n[4] adc_array_wafflecap_8_8_0[3|21]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X897 adc_array_wafflecap_8_8_1[4]/adc_array_circuit_150n_0/vint1 col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X898 adc_array_wafflecap_8_Dummy_4[19]/adc_array_circuit_150n_0/vint1 col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X899 adc_array_wafflecap_8_8_0[9|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X900 adc_array_wafflecap_8_8_0[3|10]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|10]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X901 VDD VSS adc_array_wafflecap_8_Dummy_2[2]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X902 adc_array_wafflecap_8_Dummy_8[5]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_8[5]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X903 adc_array_wafflecap_8_Dummy_2[0]/adc_array_circuit_150n_0/vint1 col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X904 adc_array_wafflecap_8_1_0/adc_array_circuit_150n_0/vint2 en_n_bit[0] adc_array_wafflecap_8_1_0/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X905 adc_array_wafflecap_8_8_0[2|23]/adc_array_circuit_150n_0/vint2 rowon_n[3] adc_array_wafflecap_8_8_0[2|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X906 adc_array_wafflecap_8_8_0[14|17]/adc_array_circuit_150n_0/vdrv row_n[15] adc_array_wafflecap_8_8_0[14|17]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X907 VSS row_n[15] adc_array_wafflecap_8_8_0[14|24]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X908 adc_array_wafflecap_8_8_0[12|28]/adc_array_circuit_150n_0/vint2 rowon_n[13] adc_array_wafflecap_8_8_0[12|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X909 adc_array_wafflecap_8_8_0[11|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X910 adc_array_wafflecap_8_8_0[3|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X911 adc_array_wafflecap_8_Dummy_1[3]/adc_array_circuit_150n_0/vint2 col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X912 adc_array_wafflecap_8_8_0[11|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X913 adc_array_wafflecap_8_8_0[10|25]/adc_array_circuit_150n_0/vint2 col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X914 adc_array_wafflecap_8_8_0[11|10]/adc_array_circuit_150n_0/vint2 rowon_n[12] adc_array_wafflecap_8_8_0[11|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X915 VSS row_n[9] adc_array_wafflecap_8_8_0[8|29]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X916 VDD rowon_n[6] adc_array_wafflecap_8_8_0[5|25]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X917 adc_array_wafflecap_8_Dummy_8[1]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_8[1]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X918 adc_array_wafflecap_8_8_0[11|0]/adc_array_circuit_150n_0/vint2 rowon_n[12] adc_array_wafflecap_8_8_0[11|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X919 adc_array_wafflecap_8_8_0[2|2]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|2]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X920 adc_array_wafflecap_8_8_0[14|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X921 adc_array_wafflecap_8_8_0[14|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X922 VSS row_n[10] adc_array_wafflecap_8_8_0[9|5]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X923 VSS row_n[10] adc_array_wafflecap_8_8_0[9|15]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X924 adc_array_wafflecap_8_8_0[1|15]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|15]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X925 adc_array_wafflecap_8_8_0[12|24]/adc_array_circuit_150n_0/vint1 col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X926 adc_array_wafflecap_8_8_0[10|12]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|12]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X927 adc_array_wafflecap_8_8_0[9|21]/adc_array_circuit_150n_0/vdrv row_n[10] adc_array_wafflecap_8_8_0[9|21]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X928 adc_array_wafflecap_8_8_1[21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_1[21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X929 VDD rowon_n[1] adc_array_wafflecap_8_8_0[0|23]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X930 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.64e+07u l=1.6e+07u
X931 adc_array_wafflecap_8_8_0[10|2]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|2]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X932 VDD rowon_n[11] adc_array_wafflecap_8_8_0[10|28]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X933 adc_array_wafflecap_8_8_0[4|28]/adc_array_circuit_150n_0/vint1 col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X934 adc_array_wafflecap_8_8_0[8|25]/adc_array_circuit_150n_0/vdrv row_n[9] adc_array_wafflecap_8_8_0[8|25]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X935 adc_array_wafflecap_8_8_0[6|22]/adc_array_circuit_150n_0/vint2 col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X936 adc_array_wafflecap_8_8_0[2|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X937 adc_array_wafflecap_8_8_0[12|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X938 VSS row_n[7] adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X939 adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X940 adc_array_wafflecap_8_8_0[5|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X941 adc_array_wafflecap_8_8_0[1|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X942 adc_array_wafflecap_8_8_0[13|27]/adc_array_circuit_150n_0/vint2 col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X943 adc_array_wafflecap_8_8_0[7|15]/adc_array_circuit_150n_0/vint1 col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X944 vcm adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|24]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X945 adc_array_wafflecap_8_8_0[7|5]/adc_array_circuit_150n_0/vint1 col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X946 adc_array_wafflecap_8_8_1[20]/adc_array_circuit_150n_0/vint2 col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X947 adc_array_wafflecap_8_8_0[14|13]/adc_array_circuit_150n_0/vint2 col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X948 VSS row_n[13] adc_array_wafflecap_8_8_0[12|17]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X949 adc_array_wafflecap_8_8_0[14|3]/adc_array_circuit_150n_0/vint2 col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X950 adc_array_wafflecap_8_Dummy_4[27]/adc_array_circuit_150n_0/vint1 col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X951 adc_array_wafflecap_8_8_0[8|18]/adc_array_circuit_150n_0/vint2 col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X952 adc_array_wafflecap_8_8_0[5|11]/adc_array_circuit_150n_0/vint2 col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X953 adc_array_wafflecap_8_8_0[6|22]/adc_array_circuit_150n_0/vdrv row_n[7] adc_array_wafflecap_8_8_0[6|22]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X954 vcm adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X955 adc_array_wafflecap_8_8_0[2|23]/adc_array_circuit_150n_0/vdrv row_n[3] adc_array_wafflecap_8_8_0[2|23]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X956 adc_array_wafflecap_8_8_0[2|24]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|24]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X957 adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/vint1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X958 adc_array_wafflecap_8_8_0[5|1]/adc_array_circuit_150n_0/vdrv row_n[6] adc_array_wafflecap_8_8_0[5|1]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X959 adc_array_wafflecap_8_8_0[4|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X960 VSS row_n[0] adc_array_wafflecap_8_8_1[5]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X961 adc_array_wafflecap_8_8_0[0|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X962 adc_array_wafflecap_8_8_0[12|3]/adc_array_circuit_150n_0/vdrv row_n[13] adc_array_wafflecap_8_8_0[12|3]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X963 adc_array_wafflecap_8_8_0[12|13]/adc_array_circuit_150n_0/vdrv row_n[13] adc_array_wafflecap_8_8_0[12|13]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X964 adc_array_wafflecap_8_8_0[10|17]/adc_array_circuit_150n_0/vint1 col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X965 adc_array_wafflecap_8_8_0[10|24]/adc_array_circuit_150n_0/vint2 rowon_n[11] adc_array_wafflecap_8_8_0[10|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X966 adc_array_wafflecap_8_8_0[9|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X967 adc_array_wafflecap_8_8_0[9|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X968 adc_array_wafflecap_8_Dummy_4[16]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X969 adc_array_wafflecap_8_8_0[11|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X970 adc_array_wafflecap_8_8_0[2|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X971 adc_array_wafflecap_8_Dummy_1[1]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X972 adc_array_wafflecap_8_Dummy_4[6]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X973 adc_array_wafflecap_8_8_0[4|3]/adc_array_circuit_150n_0/vint2 col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X974 adc_array_wafflecap_8_8_0[0|4]/adc_array_circuit_150n_0/vint2 col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X975 vcm adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|16]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X976 VDD rowon_n[6] adc_array_wafflecap_8_8_0[5|7]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X977 vcm adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|6]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X978 VDD rowon_n[9] adc_array_wafflecap_8_8_0[8|24]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X979 adc_array_wafflecap_8_8_0[3|27]/adc_array_circuit_150n_0/vint2 rowon_n[4] adc_array_wafflecap_8_8_0[3|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X980 VSS VDD adc_array_wafflecap_8_Dummy_4[23]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X981 adc_array_wafflecap_8_8_1[24]/adc_array_circuit_150n_0/vdrv row_n[0] adc_array_wafflecap_8_8_1[24]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X982 adc_array_wafflecap_8_8_0[13|26]/adc_array_circuit_150n_0/vint2 rowon_n[14] adc_array_wafflecap_8_8_0[13|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X983 adc_array_wafflecap_8_Dummy_8[2]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_8[2]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X984 adc_array_wafflecap_8_8_0[0|28]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|28]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X985 adc_array_wafflecap_8_8_0[12|17]/adc_array_circuit_150n_0/vint2 rowon_n[13] adc_array_wafflecap_8_8_0[12|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X986 adc_array_wafflecap_8_8_0[11|23]/adc_array_circuit_150n_0/vint2 col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X987 adc_array_wafflecap_8_8_0[6|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X988 adc_array_wafflecap_8_8_0[4|27]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|27]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X989 adc_array_wafflecap_8_8_0[4|9]/adc_array_circuit_150n_0/vint2 rowon_n[5] adc_array_wafflecap_8_8_0[4|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X990 adc_array_wafflecap_8_Dummy_4[33]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[33]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X991 adc_array_wafflecap_8_8_0[0|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X992 adc_array_wafflecap_8_Dummy_4[10]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X993 VSS row_n[11] adc_array_wafflecap_8_8_0[10|13]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X994 adc_array_wafflecap_8_8_0[6|18]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|18]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X995 adc_array_wafflecap_8_Dummy_4[0]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X996 VSS row_n[11] adc_array_wafflecap_8_8_0[10|3]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X997 adc_array_wafflecap_8_8_0[6|3]/adc_array_circuit_150n_0/vint2 rowon_n[7] adc_array_wafflecap_8_8_0[6|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X998 VDD rowon_n[4] adc_array_wafflecap_8_8_0[3|12]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X999 adc_array_wafflecap_8_8_0[13|22]/adc_array_circuit_150n_0/vint1 col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1000 adc_array_wafflecap_8_8_0[11|10]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|10]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1001 adc_array_wafflecap_8_8_0[7|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1002 VSS row_n[2] adc_array_wafflecap_8_8_0[1|22]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1003 VDD VDD adc_array_wafflecap_8_Dummy_4[17]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1004 adc_array_wafflecap_8_8_0[11|0]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|0]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1005 VDD rowon_n[11] adc_array_wafflecap_8_8_0[10|17]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1006 adc_array_wafflecap_8_8_0[5|8]/adc_array_circuit_150n_0/vint1 col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1007 VSS row_n[6] adc_array_wafflecap_8_8_0[5|21]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1008 adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/vint2 rowon_n[6] adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1009 adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/vint2 rowon_n[2] adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1010 VDD VDD adc_array_wafflecap_8_Dummy_4[7]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1011 adc_array_wafflecap_8_8_0[9|12]/adc_array_circuit_150n_0/vint2 col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1012 adc_array_wafflecap_8_8_1[1]/adc_array_circuit_150n_0/vint2 rowon_n[0] adc_array_wafflecap_8_8_1[1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1013 adc_array_wafflecap_8_8_0[9|2]/adc_array_circuit_150n_0/vint2 col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1014 adc_array_wafflecap_8_8_0[8|13]/adc_array_circuit_150n_0/vint1 col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1015 VSS row_n[8] adc_array_wafflecap_8_8_0[7|16]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1016 adc_array_wafflecap_8_8_1[5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1017 adc_array_wafflecap_8_8_0[2|14]/adc_array_circuit_150n_0/vint2 rowon_n[3] adc_array_wafflecap_8_8_0[2|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1018 adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1019 adc_array_wafflecap_8_8_0[8|3]/adc_array_circuit_150n_0/vint1 col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1020 adc_array_wafflecap_8_Dummy_4[2]/adc_array_circuit_150n_0/vint2 col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1021 adc_array_wafflecap_8_Dummy_4[12]/adc_array_circuit_150n_0/vint2 col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1022 VDD rowon_n[7] adc_array_wafflecap_8_8_0[6|3]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1023 VSS row_n[5] adc_array_wafflecap_8_8_0[4|10]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1024 VDD rowon_n[3] adc_array_wafflecap_8_8_0[2|4]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1025 vcm VSS adc_array_wafflecap_8_Dummy_2[4]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1026 adc_array_wafflecap_8_8_0[11|11]/adc_array_circuit_150n_0/vint1 col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1027 adc_array_wafflecap_8_8_0[7|21]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|21]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1028 VDD rowon_n[6] adc_array_wafflecap_8_8_0[5|16]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1029 adc_array_wafflecap_8_8_0[1|22]/adc_array_circuit_150n_0/vint1 col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1030 vcm adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|20]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1031 vcm adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|20]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1032 adc_array_wafflecap_8_8_0[11|1]/adc_array_circuit_150n_0/vint1 col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1033 adc_array_wafflecap_8_8_0[4|0]/adc_array_circuit_150n_0/vint1 col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1034 VDD rowon_n[2] adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1035 VSS sample_n adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1036 adc_array_wafflecap_8_8_0[2|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1037 adc_array_wafflecap_8_8_0[7|12]/adc_array_circuit_150n_0/vdrv row_n[8] adc_array_wafflecap_8_8_0[7|12]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1038 adc_array_wafflecap_8_8_0[3|13]/adc_array_circuit_150n_0/vint1 col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1039 adc_array_wafflecap_8_8_0[7|2]/adc_array_circuit_150n_0/vdrv row_n[8] adc_array_wafflecap_8_8_0[7|2]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1040 VSS row_n[7] adc_array_wafflecap_8_8_0[6|4]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1041 VDD rowon_n[1] adc_array_wafflecap_8_8_0[0|14]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1042 adc_array_wafflecap_8_8_0[13|11]/adc_array_circuit_150n_0/vdrv row_n[14] adc_array_wafflecap_8_8_0[13|11]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1043 adc_array_wafflecap_8_8_0[10|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1044 adc_array_wafflecap_8_8_0[14|24]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|24]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1045 adc_array_wafflecap_8_8_0[13|1]/adc_array_circuit_150n_0/vdrv row_n[14] adc_array_wafflecap_8_8_0[13|1]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1046 adc_array_wafflecap_8_8_0[12|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1047 adc_array_wafflecap_8_8_0[11|22]/adc_array_circuit_150n_0/vint2 rowon_n[12] adc_array_wafflecap_8_8_0[11|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1048 adc_array_wafflecap_8_8_0[10|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1049 vcm adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|1]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1050 vcm adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|11]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1051 VSS row_n[0] adc_array_wafflecap_8_8_1[2]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1052 adc_array_wafflecap_8_8_0[2|29]/adc_array_circuit_150n_0/vint2 col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1053 adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1054 VSS row_n[3] adc_array_wafflecap_8_8_0[2|15]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1055 adc_array_wafflecap_8_8_0[14|20]/adc_array_circuit_150n_0/vint2 rowon_n[15] adc_array_wafflecap_8_8_0[14|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1056 vcm adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|25]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1057 adc_array_wafflecap_8_8_0[6|4]/adc_array_circuit_150n_0/vint1 col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1058 adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/vdrv row_n[6] adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1059 vcm adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|3]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1060 adc_array_wafflecap_8_8_0[2|5]/adc_array_circuit_150n_0/vint1 col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1061 VSS row_n[11] adc_array_wafflecap_8_8_0[10|21]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1062 vcm adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|15]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1063 VDD rowon_n[0] adc_array_wafflecap_8_8_1[5]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1064 adc_array_wafflecap_8_8_0[12|5]/adc_array_circuit_150n_0/vint2 rowon_n[13] adc_array_wafflecap_8_8_0[12|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1065 adc_array_wafflecap_8_8_0[12|15]/adc_array_circuit_150n_0/vint2 rowon_n[13] adc_array_wafflecap_8_8_0[12|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1066 VDD sample adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1067 adc_array_wafflecap_8_8_0[0|29]/adc_array_circuit_150n_0/vdrv row_n[1] adc_array_wafflecap_8_8_0[0|29]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1068 vcm VSS adc_array_wafflecap_8_Dummy_4[13]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1069 adc_array_wafflecap_8_8_0[8|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1070 VDD rowon_n[6] adc_array_wafflecap_8_8_0[5|18]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1071 adc_array_wafflecap_8_8_1[26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1072 vcm VSS adc_array_wafflecap_8_Dummy_4[3]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1073 adc_array_wafflecap_8_8_0[5|7]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|7]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1074 adc_array_wafflecap_8_8_0[5|16]/adc_array_circuit_150n_0/vint1 col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1075 vcm adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[13]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1076 adc_array_wafflecap_8_8_0[0|15]/adc_array_circuit_150n_0/vint1 col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1077 adc_array_wafflecap_8_8_0[1|8]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|8]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1078 VDD rowon_n[13] adc_array_wafflecap_8_8_0[12|20]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1079 adc_array_wafflecap_8_8_0[5|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1080 adc_array_wafflecap_8_8_0[1|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1081 VDD rowon_n[12] adc_array_wafflecap_8_8_0[11|1]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1082 VDD rowon_n[12] adc_array_wafflecap_8_8_0[11|11]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1083 adc_array_wafflecap_8_8_0[8|21]/adc_array_circuit_150n_0/vint1 col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1084 VDD rowon_n[11] adc_array_wafflecap_8_8_0[10|15]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1085 VDD rowon_n[11] adc_array_wafflecap_8_8_0[10|5]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1086 adc_array_wafflecap_8_8_0[4|20]/adc_array_circuit_150n_0/vint2 rowon_n[5] adc_array_wafflecap_8_8_0[4|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1087 adc_array_wafflecap_8_8_0[0|21]/adc_array_circuit_150n_0/vint2 rowon_n[1] adc_array_wafflecap_8_8_0[0|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1088 adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/vint2 VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1089 adc_array_wafflecap_8_8_0[8|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1090 VSS row_n[15] adc_array_wafflecap_8_8_0[14|9]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1091 VDD rowon_n[4] adc_array_wafflecap_8_8_0[3|23]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1092 adc_array_wafflecap_8_8_0[0|0]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|0]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1093 adc_array_wafflecap_8_8_0[10|10]/adc_array_circuit_150n_0/vint2 col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1094 adc_array_wafflecap_8_8_0[3|12]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|12]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1095 adc_array_wafflecap_8_8_0[10|0]/adc_array_circuit_150n_0/vint2 col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1096 VDD sample adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1097 VDD VSS adc_array_wafflecap_8_Dummy_2[4]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1098 adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/vdrv row_n[13] adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1099 adc_array_wafflecap_8_8_0[12|9]/adc_array_circuit_150n_0/vint1 col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1100 adc_array_wafflecap_8_8_0[9|6]/adc_array_circuit_150n_0/vdrv row_n[10] adc_array_wafflecap_8_8_0[9|6]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1101 adc_array_wafflecap_8_8_0[3|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1102 adc_array_wafflecap_8_8_0[2|25]/adc_array_circuit_150n_0/vint2 rowon_n[3] adc_array_wafflecap_8_8_0[2|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1103 vcm adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1104 adc_array_wafflecap_8_8_0[12|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1105 adc_array_wafflecap_8_8_0[12|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1106 adc_array_wafflecap_8_8_0[9|23]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|23]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1107 adc_array_wafflecap_8_8_0[8|0]/adc_array_circuit_150n_0/vdrv row_n[9] adc_array_wafflecap_8_8_0[8|0]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1108 adc_array_wafflecap_8_8_0[8|10]/adc_array_circuit_150n_0/vdrv row_n[9] adc_array_wafflecap_8_8_0[8|10]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1109 adc_array_wafflecap_8_Dummy_8[3]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_8[3]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1110 adc_array_wafflecap_8_8_0[11|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1111 vcm adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|9]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1112 adc_array_wafflecap_8_8_0[11|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1113 VSS sample_n adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1114 adc_array_wafflecap_8_8_0[3|9]/adc_array_circuit_150n_0/vint2 col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1115 adc_array_wafflecap_8_8_0[4|20]/adc_array_circuit_150n_0/vdrv row_n[5] adc_array_wafflecap_8_8_0[4|20]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1116 adc_array_wafflecap_8_8_1[23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_1[23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1117 VDD rowon_n[1] adc_array_wafflecap_8_8_0[0|25]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1118 vcm adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|28]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1119 adc_array_wafflecap_8_8_0[4|21]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|21]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1120 adc_array_wafflecap_8_8_0[4|30]/adc_array_circuit_150n_0/vint1 col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1121 adc_array_wafflecap_8_Dummy_8[1]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_8[1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1122 vcm adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|29]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1123 adc_array_wafflecap_8_8_0[2|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1124 adc_array_wafflecap_8_Dummy_4[19]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1125 adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/vint2 rowon_n[15] adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1126 adc_array_wafflecap_8_8_0[5|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1127 adc_array_wafflecap_8_8_0[1|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1128 adc_array_wafflecap_8_8_0[14|9]/adc_array_circuit_150n_0/vint2 rowon_n[15] adc_array_wafflecap_8_8_0[14|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1129 VSS row_n[12] adc_array_wafflecap_8_8_0[11|19]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1130 adc_array_wafflecap_8_8_0[13|13]/adc_array_circuit_150n_0/vint2 rowon_n[14] adc_array_wafflecap_8_8_0[13|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1131 VSS row_n[11] adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1132 adc_array_wafflecap_8_8_0[7|29]/adc_array_circuit_150n_0/vint2 col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1133 adc_array_wafflecap_8_8_1[27]/adc_array_circuit_150n_0/vint1 col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1134 adc_array_wafflecap_8_8_0[13|3]/adc_array_circuit_150n_0/vint2 rowon_n[14] adc_array_wafflecap_8_8_0[13|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1135 adc_array_wafflecap_8_8_1[22]/adc_array_circuit_150n_0/vint2 col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1136 adc_array_wafflecap_8_8_0[0|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1137 adc_array_wafflecap_8_8_0[2|1]/adc_array_circuit_150n_0/vint2 col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1138 VDD rowon_n[14] adc_array_wafflecap_8_8_0[13|18]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1139 adc_array_wafflecap_8_8_0[12|15]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|15]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1140 adc_array_wafflecap_8_8_0[5|13]/adc_array_circuit_150n_0/vint2 col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1141 adc_array_wafflecap_8_8_0[1|14]/adc_array_circuit_150n_0/vint2 col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1142 adc_array_wafflecap_8_8_0[12|5]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|5]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1143 VDD rowon_n[13] adc_array_wafflecap_8_8_0[12|9]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1144 VDD rowon_n[13] adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1145 adc_array_wafflecap_8_8_0[11|24]/adc_array_circuit_150n_0/vdrv row_n[12] adc_array_wafflecap_8_8_0[11|24]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1146 adc_array_wafflecap_8_8_0[9|28]/adc_array_circuit_150n_0/vint1 col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1147 adc_array_wafflecap_8_8_0[2|25]/adc_array_circuit_150n_0/vdrv row_n[3] adc_array_wafflecap_8_8_0[2|25]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1148 adc_array_wafflecap_8_8_0[5|3]/adc_array_circuit_150n_0/vdrv row_n[6] adc_array_wafflecap_8_8_0[5|3]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1149 adc_array_wafflecap_8_8_0[4|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1150 adc_array_wafflecap_8_8_0[2|26]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|26]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1151 adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/vint1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1152 adc_array_wafflecap_8_8_0[5|4]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|4]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1153 adc_array_wafflecap_8_Dummy_4[31]/adc_array_circuit_150n_0/vint2 col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1154 adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1155 adc_array_wafflecap_8_8_0[0|1]/adc_array_circuit_150n_0/vdrv row_n[1] adc_array_wafflecap_8_8_0[0|1]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1156 adc_array_wafflecap_8_8_0[2|7]/adc_array_circuit_150n_0/vint2 rowon_n[3] adc_array_wafflecap_8_8_0[2|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1157 VSS VDD adc_array_wafflecap_8_Dummy_4[8]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1158 adc_array_wafflecap_8_8_0[2|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1159 adc_array_wafflecap_8_Dummy_1[3]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1160 adc_array_wafflecap_8_8_0[4|5]/adc_array_circuit_150n_0/vint2 col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1161 adc_array_wafflecap_8_8_0[1|14]/adc_array_circuit_150n_0/vdrv row_n[2] adc_array_wafflecap_8_8_0[1|14]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1162 adc_array_wafflecap_8_Dummy_4[18]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[18]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1163 adc_array_wafflecap_8_8_0[14|26]/adc_array_circuit_150n_0/vdrv row_n[15] adc_array_wafflecap_8_8_0[14|26]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1164 adc_array_wafflecap_8_8_0[11|8]/adc_array_circuit_150n_0/vint2 col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1165 VDD rowon_n[6] adc_array_wafflecap_8_8_0[5|9]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1166 adc_array_wafflecap_8_8_0[13|30]/adc_array_circuit_150n_0/vdrv row_n[14] adc_array_wafflecap_8_8_0[13|30]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1167 vcm adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|30]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1168 VSS row_n[4] adc_array_wafflecap_8_8_0[3|19]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1169 adc_array_wafflecap_8_8_0[3|29]/adc_array_circuit_150n_0/vint2 rowon_n[4] adc_array_wafflecap_8_8_0[3|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1170 VDD rowon_n[1] adc_array_wafflecap_8_8_0[0|7]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1171 adc_array_wafflecap_8_8_0[14|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1172 adc_array_wafflecap_8_8_0[13|7]/adc_array_circuit_150n_0/vint1 col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1173 vcm adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|29]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1174 adc_array_wafflecap_8_8_0[7|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1175 adc_array_wafflecap_8_8_0[3|17]/adc_array_circuit_150n_0/vint2 col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1176 adc_array_wafflecap_8_8_0[4|11]/adc_array_circuit_150n_0/vint2 rowon_n[5] adc_array_wafflecap_8_8_0[4|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1177 adc_array_wafflecap_8_8_0[0|12]/adc_array_circuit_150n_0/vint2 rowon_n[1] adc_array_wafflecap_8_8_0[0|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1178 adc_array_wafflecap_8_8_0[0|30]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|30]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1179 adc_array_wafflecap_8_8_0[13|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1180 adc_array_wafflecap_8_8_0[10|21]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|21]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1181 adc_array_wafflecap_8_8_0[6|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1182 adc_array_wafflecap_8_8_0[0|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1183 VDD rowon_n[5] adc_array_wafflecap_8_8_0[4|1]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1184 VSS row_n[3] adc_array_wafflecap_8_8_0[2|8]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1185 VDD rowon_n[4] adc_array_wafflecap_8_8_0[3|14]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1186 adc_array_wafflecap_8_8_0[9|30]/adc_array_circuit_150n_0/vint2 rowon_n[10] adc_array_wafflecap_8_8_0[9|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1187 adc_array_wafflecap_8_8_0[6|5]/adc_array_circuit_150n_0/vint2 rowon_n[7] adc_array_wafflecap_8_8_0[6|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1188 adc_array_wafflecap_8_8_0[4|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1189 adc_array_wafflecap_8_8_0[0|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1190 adc_array_wafflecap_8_8_0[9|8]/adc_array_circuit_150n_0/vint2 rowon_n[10] adc_array_wafflecap_8_8_0[9|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1191 vcm adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|8]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1192 adc_array_wafflecap_8_8_1[18]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[18]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1193 VSS row_n[2] adc_array_wafflecap_8_8_0[1|24]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1194 adc_array_wafflecap_8_8_0[6|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1195 adc_array_wafflecap_8_8_0[5|10]/adc_array_circuit_150n_0/vint1 col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1196 VDD VSS adc_array_wafflecap_8_Dummy_1[3]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1197 adc_array_wafflecap_8_Dummy_4[8]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1198 adc_array_wafflecap_8_Dummy_4[30]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1199 adc_array_wafflecap_8_8_1[3]/adc_array_circuit_150n_0/vint2 rowon_n[0] adc_array_wafflecap_8_8_1[3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1200 VSS row_n[12] adc_array_wafflecap_8_8_0[11|30]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1201 adc_array_wafflecap_8_8_0[0|8]/adc_array_circuit_150n_0/vint1 col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1202 adc_array_wafflecap_8_8_0[2|16]/adc_array_circuit_150n_0/vint2 rowon_n[3] adc_array_wafflecap_8_8_0[2|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1203 adc_array_wafflecap_8_8_0[4|26]/adc_array_circuit_150n_0/vint2 col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1204 adc_array_wafflecap_8_8_0[14|9]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|9]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1205 VDD rowon_n[8] adc_array_wafflecap_8_8_0[7|8]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1206 VDD rowon_n[8] adc_array_wafflecap_8_8_0[7|30]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1207 VDD rowon_n[3] adc_array_wafflecap_8_8_0[2|6]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1208 VSS row_n[1] adc_array_wafflecap_8_8_0[0|13]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1209 VDD sample_n adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1210 VDD rowon_n[7] adc_array_wafflecap_8_8_0[6|5]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1211 VSS row_n[5] adc_array_wafflecap_8_8_0[4|12]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1212 vcm VSS adc_array_wafflecap_8_Dummy_2[6]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1213 vcm adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|22]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1214 adc_array_wafflecap_8_Dummy_4[26]/adc_array_circuit_150n_0/vint1 col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1215 adc_array_wafflecap_8_8_0[13|13]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|13]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1216 VDD rowon_n[14] adc_array_wafflecap_8_8_0[13|29]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1217 adc_array_wafflecap_8_8_0[11|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1218 adc_array_wafflecap_8_8_0[9|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1219 vcm adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|0]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1220 adc_array_wafflecap_8_8_0[3|29]/adc_array_circuit_150n_0/vdrv row_n[4] adc_array_wafflecap_8_8_0[3|29]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1221 vcm adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|1]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1222 adc_array_wafflecap_8_8_0[1|24]/adc_array_circuit_150n_0/vint1 col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1223 adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1224 adc_array_wafflecap_8_8_0[13|3]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|3]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1225 VDD rowon_n[14] adc_array_wafflecap_8_8_0[13|7]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1226 adc_array_wafflecap_8_8_0[4|2]/adc_array_circuit_150n_0/vint1 col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1227 adc_array_wafflecap_8_8_0[4|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1228 adc_array_wafflecap_8_8_0[3|15]/adc_array_circuit_150n_0/vint1 col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1229 VDD rowon_n[1] adc_array_wafflecap_8_8_0[0|16]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1230 VSS row_n[11] adc_array_wafflecap_8_8_0[10|6]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1231 adc_array_wafflecap_8_Dummy_7/adc_array_circuit_150n_0/vint1 col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1232 adc_array_wafflecap_8_Dummy_1[4]/adc_array_circuit_150n_0/vint1 col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1233 VSS row_n[0] adc_array_wafflecap_8_8_1[4]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1234 adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/vint2 col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1235 VSS VDD adc_array_wafflecap_8_Dummy_4[19]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1236 adc_array_wafflecap_8_8_0[7|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1237 vcm adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|23]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1238 adc_array_wafflecap_8_8_0[12|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1239 adc_array_wafflecap_8_8_0[11|19]/adc_array_circuit_150n_0/vint2 col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1240 vcm adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|5]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1241 adc_array_wafflecap_8_Dummy_2[2]/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_2[2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1242 adc_array_wafflecap_8_8_0[2|18]/adc_array_circuit_150n_0/vint2 rowon_n[3] adc_array_wafflecap_8_8_0[2|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1243 adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1244 adc_array_wafflecap_8_8_0[9|15]/adc_array_circuit_150n_0/vdrv row_n[10] adc_array_wafflecap_8_8_0[9|15]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1245 adc_array_wafflecap_8_8_0[9|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1246 adc_array_wafflecap_8_8_0[8|6]/adc_array_circuit_150n_0/vint1 col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1247 adc_array_wafflecap_8_Dummy_8[5]/adc_array_circuit_150n_0/vint2 col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1248 adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1249 adc_array_wafflecap_8_8_0[9|5]/adc_array_circuit_150n_0/vdrv row_n[10] adc_array_wafflecap_8_8_0[9|5]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1250 vcm adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|28]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1251 VSS VSS adc_array_wafflecap_8_Dummy_2[0]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1252 VSS row_n[3] adc_array_wafflecap_8_8_0[2|16]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1253 adc_array_wafflecap_8_8_0[14|17]/adc_array_circuit_150n_0/vint2 col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1254 VDD rowon_n[6] adc_array_wafflecap_8_8_0[5|20]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1255 adc_array_wafflecap_8_8_1[28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1256 adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/vdrv row_n[1] adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1257 adc_array_wafflecap_8_Dummy_4[5]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[5]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1258 adc_array_wafflecap_8_Dummy_4[15]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[15]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1259 adc_array_wafflecap_8_8_0[13|18]/adc_array_circuit_150n_0/vint1 col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1260 vcm adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|4]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1261 vcm adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|14]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1262 adc_array_wafflecap_8_8_0[7|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1263 vcm adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[15]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1264 adc_array_wafflecap_8_8_0[1|10]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|10]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1265 VDD rowon_n[1] adc_array_wafflecap_8_8_0[0|18]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1266 adc_array_wafflecap_8_8_0[0|23]/adc_array_circuit_150n_0/vint2 rowon_n[1] adc_array_wafflecap_8_8_0[0|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1267 adc_array_wafflecap_8_8_0[0|16]/adc_array_circuit_150n_0/vint1 col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1268 adc_array_wafflecap_8_8_0[1|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1269 adc_array_wafflecap_8_8_0[12|17]/adc_array_circuit_150n_0/vdrv row_n[13] adc_array_wafflecap_8_8_0[12|17]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1270 VSS row_n[13] adc_array_wafflecap_8_8_0[12|24]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1271 adc_array_wafflecap_8_8_0[10|28]/adc_array_circuit_150n_0/vint2 rowon_n[11] adc_array_wafflecap_8_8_0[10|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1272 adc_array_wafflecap_8_8_0[9|21]/adc_array_circuit_150n_0/vint2 col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1273 VSS row_n[7] adc_array_wafflecap_8_8_0[6|27]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1274 adc_array_wafflecap_8_8_0[5|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1275 adc_array_wafflecap_8_8_0[8|25]/adc_array_circuit_150n_0/vint2 col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1276 VDD rowon_n[4] adc_array_wafflecap_8_8_0[3|25]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1277 adc_array_wafflecap_8_8_0[0|2]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|2]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1278 VDD rowon_n[15] adc_array_wafflecap_8_8_0[14|23]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1279 adc_array_wafflecap_8_8_0[12|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1280 adc_array_wafflecap_8_8_0[12|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1281 adc_array_wafflecap_8_8_0[11|20]/adc_array_circuit_150n_0/vint1 col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1282 adc_array_wafflecap_8_8_0[9|8]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|8]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1283 VSS row_n[8] adc_array_wafflecap_8_8_0[7|5]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1284 VSS row_n[8] adc_array_wafflecap_8_8_0[7|15]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1285 adc_array_wafflecap_8_8_0[10|24]/adc_array_circuit_150n_0/vint1 col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1286 adc_array_wafflecap_8_8_0[7|21]/adc_array_circuit_150n_0/vdrv row_n[8] adc_array_wafflecap_8_8_0[7|21]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1287 adc_array_wafflecap_8_8_0[5|6]/adc_array_circuit_150n_0/vint2 col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1288 VDD VSS adc_array_wafflecap_8_Dummy_2[6]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1289 VDD rowon_n[9] adc_array_wafflecap_8_8_0[8|28]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1290 adc_array_wafflecap_8_8_0[2|28]/adc_array_circuit_150n_0/vint1 col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1291 adc_array_wafflecap_8_8_0[0|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1292 VSS VDD adc_array_wafflecap_8_Dummy_4[27]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1293 adc_array_wafflecap_8_8_0[6|27]/adc_array_circuit_150n_0/vint1 col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1294 adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1295 adc_array_wafflecap_8_8_0[10|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1296 adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1297 adc_array_wafflecap_8_8_0[3|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1298 adc_array_wafflecap_8_8_0[11|27]/adc_array_circuit_150n_0/vint2 col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1299 adc_array_wafflecap_8_8_0[12|13]/adc_array_circuit_150n_0/vint2 col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1300 VSS row_n[11] adc_array_wafflecap_8_8_0[10|17]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1301 adc_array_wafflecap_8_8_0[12|3]/adc_array_circuit_150n_0/vint2 col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1302 adc_array_wafflecap_8_8_0[7|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1303 adc_array_wafflecap_8_Dummy_4[23]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[23]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1304 adc_array_wafflecap_8_8_0[13|26]/adc_array_circuit_150n_0/vint1 col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1305 vcm adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|22]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1306 adc_array_wafflecap_8_8_0[3|11]/adc_array_circuit_150n_0/vint2 col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1307 vcm adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|30]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1308 adc_array_wafflecap_8_8_0[4|22]/adc_array_circuit_150n_0/vdrv row_n[5] adc_array_wafflecap_8_8_0[4|22]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1309 adc_array_wafflecap_8_8_0[4|23]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|23]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1310 adc_array_wafflecap_8_Dummy_8[3]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_8[3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1311 adc_array_wafflecap_8_8_1[25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_1[25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1312 adc_array_wafflecap_8_8_0[0|24]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|24]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1313 vcm adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1314 vcm VSS adc_array_wafflecap_8_Dummy_4[22]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1315 adc_array_wafflecap_8_8_0[14|12]/adc_array_circuit_150n_0/vint1 col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1316 adc_array_wafflecap_8_8_0[11|9]/adc_array_circuit_150n_0/vdrv row_n[12] adc_array_wafflecap_8_8_0[11|9]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1317 adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/vint1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1318 adc_array_wafflecap_8_8_0[3|1]/adc_array_circuit_150n_0/vdrv row_n[4] adc_array_wafflecap_8_8_0[3|1]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1319 adc_array_wafflecap_8_8_0[2|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1320 adc_array_wafflecap_8_8_0[14|2]/adc_array_circuit_150n_0/vint1 col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1321 adc_array_wafflecap_8_8_0[6|14]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|14]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1322 adc_array_wafflecap_8_8_0[5|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1323 adc_array_wafflecap_8_8_1[19]/adc_array_circuit_150n_0/vdrv row_n[0] adc_array_wafflecap_8_8_1[19]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1324 adc_array_wafflecap_8_8_0[10|3]/adc_array_circuit_150n_0/vdrv row_n[11] adc_array_wafflecap_8_8_0[10|3]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1325 adc_array_wafflecap_8_8_0[10|13]/adc_array_circuit_150n_0/vdrv row_n[11] adc_array_wafflecap_8_8_0[10|13]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1326 adc_array_wafflecap_8_8_0[8|17]/adc_array_circuit_150n_0/vint1 col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1327 adc_array_wafflecap_8_8_0[8|24]/adc_array_circuit_150n_0/vint2 rowon_n[9] adc_array_wafflecap_8_8_0[8|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1328 adc_array_wafflecap_8_8_0[7|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1329 adc_array_wafflecap_8_8_0[7|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1330 adc_array_wafflecap_8_Dummy_0[0]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_0[0]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1331 adc_array_wafflecap_8_8_1[29]/adc_array_circuit_150n_0/vint1 col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1332 adc_array_wafflecap_8_8_0[9|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1333 adc_array_wafflecap_8_8_0[13|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1334 adc_array_wafflecap_8_8_1[24]/adc_array_circuit_150n_0/vint2 col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1335 adc_array_wafflecap_8_8_0[0|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1336 adc_array_wafflecap_8_8_0[13|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1337 vcm adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|19]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1338 adc_array_wafflecap_8_Dummy_8[2]/adc_array_circuit_150n_0/vint2 col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1339 adc_array_wafflecap_8_8_0[2|3]/adc_array_circuit_150n_0/vint2 col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1340 adc_array_wafflecap_8_8_0[5|15]/adc_array_circuit_150n_0/vint2 col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1341 VDD rowon_n[4] adc_array_wafflecap_8_8_0[3|7]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1342 adc_array_wafflecap_8_8_0[5|5]/adc_array_circuit_150n_0/vdrv row_n[6] adc_array_wafflecap_8_8_0[5|5]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1343 adc_array_wafflecap_8_8_0[5|6]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|6]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1344 adc_array_wafflecap_8_8_0[5|26]/adc_array_circuit_150n_0/vint2 rowon_n[6] adc_array_wafflecap_8_8_0[5|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1345 adc_array_wafflecap_8_8_0[1|27]/adc_array_circuit_150n_0/vint2 rowon_n[2] adc_array_wafflecap_8_8_0[1|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1346 VSS row_n[14] adc_array_wafflecap_8_8_0[13|22]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1347 adc_array_wafflecap_8_8_0[7|5]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|5]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1348 adc_array_wafflecap_8_8_0[7|15]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|15]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1349 adc_array_wafflecap_8_Dummy_4[17]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1350 adc_array_wafflecap_8_8_0[14|28]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|28]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1351 adc_array_wafflecap_8_8_0[11|26]/adc_array_circuit_150n_0/vint2 rowon_n[12] adc_array_wafflecap_8_8_0[11|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1352 adc_array_wafflecap_8_Dummy_3[3]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_3[3]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1353 adc_array_wafflecap_8_Dummy_4[7]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1354 adc_array_wafflecap_8_8_0[10|17]/adc_array_circuit_150n_0/vint2 rowon_n[11] adc_array_wafflecap_8_8_0[10|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1355 adc_array_wafflecap_8_8_0[2|27]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|27]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1356 adc_array_wafflecap_8_8_1[0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1357 adc_array_wafflecap_8_8_0[0|3]/adc_array_circuit_150n_0/vdrv row_n[1] adc_array_wafflecap_8_8_0[0|3]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1358 adc_array_wafflecap_8_8_0[2|9]/adc_array_circuit_150n_0/vint2 rowon_n[3] adc_array_wafflecap_8_8_0[2|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1359 adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1360 adc_array_wafflecap_8_Dummy_1[5]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1361 VDD VDD adc_array_wafflecap_8_Dummy_4[22]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1362 adc_array_wafflecap_8_8_0[13|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1363 VSS row_n[9] adc_array_wafflecap_8_8_0[8|13]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1364 VDD rowon_n[15] adc_array_wafflecap_8_8_0[14|12]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1365 adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1366 adc_array_wafflecap_8_8_0[9|19]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|19]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1367 VSS row_n[9] adc_array_wafflecap_8_8_0[8|3]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1368 VDD rowon_n[6] adc_array_wafflecap_8_8_0[5|11]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1369 VDD rowon_n[15] adc_array_wafflecap_8_8_0[14|2]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1370 VDD rowon_n[2] adc_array_wafflecap_8_8_0[1|27]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1371 VDD rowon_n[14] adc_array_wafflecap_8_8_0[13|16]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1372 VDD rowon_n[9] adc_array_wafflecap_8_8_0[8|17]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1373 adc_array_wafflecap_8_8_0[3|8]/adc_array_circuit_150n_0/vint1 col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1374 VSS row_n[4] adc_array_wafflecap_8_8_0[3|21]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1375 adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/vint2 rowon_n[4] adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1376 VDD rowon_n[14] adc_array_wafflecap_8_8_0[13|6]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1377 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X1378 VDD rowon_n[1] adc_array_wafflecap_8_8_0[0|9]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1379 adc_array_wafflecap_8_8_0[7|12]/adc_array_circuit_150n_0/vint2 col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1380 adc_array_wafflecap_8_8_0[7|2]/adc_array_circuit_150n_0/vint2 col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1381 adc_array_wafflecap_8_8_0[6|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1382 adc_array_wafflecap_8_8_0[4|13]/adc_array_circuit_150n_0/vint2 rowon_n[5] adc_array_wafflecap_8_8_0[4|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1383 adc_array_wafflecap_8_8_0[0|14]/adc_array_circuit_150n_0/vint2 rowon_n[1] adc_array_wafflecap_8_8_0[0|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1384 adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1385 adc_array_wafflecap_8_8_0[14|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1386 adc_array_wafflecap_8_8_0[13|1]/adc_array_circuit_150n_0/vint2 col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1387 adc_array_wafflecap_8_8_0[13|11]/adc_array_circuit_150n_0/vint2 col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1388 VDD rowon_n[5] adc_array_wafflecap_8_8_0[4|3]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1389 VSS row_n[3] adc_array_wafflecap_8_8_0[2|10]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1390 adc_array_wafflecap_8_8_0[9|11]/adc_array_circuit_150n_0/vint1 col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1391 adc_array_wafflecap_8_8_0[8|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1392 VDD rowon_n[4] adc_array_wafflecap_8_8_0[3|16]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1393 adc_array_wafflecap_8_8_1[22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1394 adc_array_wafflecap_8_8_0[0|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1395 vcm adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|20]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1396 vcm adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|20]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1397 adc_array_wafflecap_8_8_0[9|1]/adc_array_circuit_150n_0/vint1 col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1398 adc_array_wafflecap_8_8_0[5|26]/adc_array_circuit_150n_0/vdrv row_n[6] adc_array_wafflecap_8_8_0[5|26]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1399 adc_array_wafflecap_8_8_0[4|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1400 adc_array_wafflecap_8_8_0[2|0]/adc_array_circuit_150n_0/vint1 col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1401 vcm adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|10]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1402 adc_array_wafflecap_8_8_0[5|12]/adc_array_circuit_150n_0/vint1 col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1403 VDD rowon_n[0] adc_array_wafflecap_8_8_1[0]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1404 adc_array_wafflecap_8_Dummy_4[1]/adc_array_circuit_150n_0/vint1 col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1405 adc_array_wafflecap_8_Dummy_4[11]/adc_array_circuit_150n_0/vint1 col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1406 adc_array_wafflecap_8_8_0[9|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1407 adc_array_wafflecap_8_8_0[9|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1408 adc_array_wafflecap_8_8_0[5|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1409 VDD VSS adc_array_wafflecap_8_Dummy_1[5]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1410 adc_array_wafflecap_8_8_0[8|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1411 adc_array_wafflecap_8_8_1[5]/adc_array_circuit_150n_0/vint2 rowon_n[0] adc_array_wafflecap_8_8_1[5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1412 adc_array_wafflecap_8_8_0[12|24]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|24]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1413 adc_array_wafflecap_8_8_0[10|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1414 adc_array_wafflecap_8_8_0[8|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1415 vcm adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[8]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1416 adc_array_wafflecap_8_8_0[0|10]/adc_array_circuit_150n_0/vint1 col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1417 adc_array_wafflecap_8_8_0[4|28]/adc_array_circuit_150n_0/vint2 col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1418 adc_array_wafflecap_8_8_0[0|29]/adc_array_circuit_150n_0/vint2 col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1419 VSS row_n[5] adc_array_wafflecap_8_8_0[4|14]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1420 VSS row_n[1] adc_array_wafflecap_8_8_0[0|15]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1421 adc_array_wafflecap_8_8_0[12|20]/adc_array_circuit_150n_0/vint2 rowon_n[13] adc_array_wafflecap_8_8_0[12|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1422 adc_array_wafflecap_8_8_0[6|19]/adc_array_circuit_150n_0/vint2 col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1423 vcm VSS adc_array_wafflecap_8_Dummy_3[0]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1424 vcm adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|2]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1425 adc_array_wafflecap_8_8_0[4|4]/adc_array_circuit_150n_0/vint1 col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1426 adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/vdrv row_n[4] adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1427 vcm adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|3]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1428 vcm adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|8]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1429 adc_array_wafflecap_8_8_0[9|27]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|27]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1430 VSS row_n[9] adc_array_wafflecap_8_8_0[8|21]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1431 adc_array_wafflecap_8_8_0[4|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1432 adc_array_wafflecap_8_8_0[10|5]/adc_array_circuit_150n_0/vint2 rowon_n[11] adc_array_wafflecap_8_8_0[10|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1433 adc_array_wafflecap_8_8_0[10|15]/adc_array_circuit_150n_0/vint2 rowon_n[11] adc_array_wafflecap_8_8_0[10|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1434 VDD sample adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1435 adc_array_wafflecap_8_8_0[8|13]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|13]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1436 adc_array_wafflecap_8_Dummy_3[4]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_3[4]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1437 vcm adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|2]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1438 vcm adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|12]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1439 adc_array_wafflecap_8_8_0[8|3]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|3]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1440 VDD rowon_n[4] adc_array_wafflecap_8_8_0[3|18]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1441 adc_array_wafflecap_8_8_1[1]/adc_array_circuit_150n_0/vint1 col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1442 adc_array_wafflecap_8_8_0[3|7]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|7]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1443 adc_array_wafflecap_8_8_0[3|16]/adc_array_circuit_150n_0/vint1 col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1444 adc_array_wafflecap_8_Dummy_1[6]/adc_array_circuit_150n_0/vint1 col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1445 VDD rowon_n[11] adc_array_wafflecap_8_8_0[10|20]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1446 adc_array_wafflecap_8_8_0[3|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1447 VDD rowon_n[10] adc_array_wafflecap_8_8_0[9|1]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1448 VDD rowon_n[10] adc_array_wafflecap_8_8_0[9|11]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1449 adc_array_wafflecap_8_8_0[6|19]/adc_array_circuit_150n_0/vdrv row_n[7] adc_array_wafflecap_8_8_0[6|19]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1450 adc_array_wafflecap_8_Dummy_4[17]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[17]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1451 VDD rowon_n[9] adc_array_wafflecap_8_8_0[8|15]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1452 adc_array_wafflecap_8_Dummy_4[7]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[7]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1453 VDD VDD adc_array_wafflecap_8_Dummy_4[33]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1454 VDD rowon_n[9] adc_array_wafflecap_8_8_0[8|5]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1455 adc_array_wafflecap_8_Dummy_2[4]/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_2[4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1456 adc_array_wafflecap_8_8_0[2|20]/adc_array_circuit_150n_0/vint2 rowon_n[3] adc_array_wafflecap_8_8_0[2|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1457 adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/vint2 VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1458 VSS row_n[13] adc_array_wafflecap_8_8_0[12|9]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1459 adc_array_wafflecap_8_8_0[9|6]/adc_array_circuit_150n_0/vint2 col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1460 adc_array_wafflecap_8_Dummy_0[1]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_0[1]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1461 adc_array_wafflecap_8_8_1[30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1462 adc_array_wafflecap_8_8_0[8|10]/adc_array_circuit_150n_0/vint2 col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1463 adc_array_wafflecap_8_8_0[5|17]/adc_array_circuit_150n_0/vint2 rowon_n[6] adc_array_wafflecap_8_8_0[5|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1464 vcm adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|24]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1465 adc_array_wafflecap_8_8_0[1|12]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|12]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1466 adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/vint1 col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1467 adc_array_wafflecap_8_8_0[11|28]/adc_array_circuit_150n_0/vdrv row_n[12] adc_array_wafflecap_8_8_0[11|28]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1468 adc_array_wafflecap_8_8_0[8|0]/adc_array_circuit_150n_0/vint2 col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1469 adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/vdrv row_n[11] adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1470 adc_array_wafflecap_8_8_1[18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_1[18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1471 VDD rowon_n[1] adc_array_wafflecap_8_8_0[0|20]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1472 adc_array_wafflecap_8_8_0[14|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1473 adc_array_wafflecap_8_8_0[10|9]/adc_array_circuit_150n_0/vint1 col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1474 adc_array_wafflecap_8_8_0[7|6]/adc_array_circuit_150n_0/vdrv row_n[8] adc_array_wafflecap_8_8_0[7|6]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1475 adc_array_wafflecap_8_8_0[5|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1476 vcm adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[16]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1477 adc_array_wafflecap_8_8_0[0|25]/adc_array_circuit_150n_0/vint2 rowon_n[1] adc_array_wafflecap_8_8_0[0|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1478 adc_array_wafflecap_8_8_0[1|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1479 vcm adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1480 VSS row_n[7] adc_array_wafflecap_8_8_0[6|29]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1481 adc_array_wafflecap_8_8_0[10|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1482 adc_array_wafflecap_8_8_0[10|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1483 VSS row_n[0] adc_array_wafflecap_8_8_1[27]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1484 adc_array_wafflecap_8_8_0[5|8]/adc_array_circuit_150n_0/vint2 col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1485 adc_array_wafflecap_8_8_0[1|9]/adc_array_circuit_150n_0/vint2 col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1486 VSS row_n[6] adc_array_wafflecap_8_8_0[5|18]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1487 adc_array_wafflecap_8_8_0[2|20]/adc_array_circuit_150n_0/vdrv row_n[3] adc_array_wafflecap_8_8_0[2|20]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1488 VDD VSS adc_array_wafflecap_8_Dummy_3[0]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1489 adc_array_wafflecap_8_Dummy_4[8]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[8]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1490 adc_array_wafflecap_8_8_0[13|18]/adc_array_circuit_150n_0/vint2 rowon_n[14] adc_array_wafflecap_8_8_0[13|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1491 vcm adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|7]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1492 adc_array_wafflecap_8_8_0[7|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1493 adc_array_wafflecap_8_8_0[7|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1494 adc_array_wafflecap_8_8_0[6|29]/adc_array_circuit_150n_0/vint1 col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1495 adc_array_wafflecap_8_8_0[4|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1496 vcm adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|28]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1497 adc_array_wafflecap_8_8_0[2|21]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|21]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1498 adc_array_wafflecap_8_8_0[2|30]/adc_array_circuit_150n_0/vint1 col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1499 adc_array_wafflecap_8_8_0[0|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1500 adc_array_wafflecap_8_8_0[12|9]/adc_array_circuit_150n_0/vint2 rowon_n[13] adc_array_wafflecap_8_8_0[12|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1501 adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/vint2 rowon_n[13] adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1502 VSS row_n[10] adc_array_wafflecap_8_8_0[9|28]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1503 VDD sample_n adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1504 adc_array_wafflecap_8_8_0[3|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1505 vcm adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|19]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1506 adc_array_wafflecap_8_8_0[11|13]/adc_array_circuit_150n_0/vint2 rowon_n[12] adc_array_wafflecap_8_8_0[11|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1507 VSS row_n[9] adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1508 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.64e+07u l=1.6e+07u
X1509 adc_array_wafflecap_8_8_0[11|3]/adc_array_circuit_150n_0/vint2 rowon_n[12] adc_array_wafflecap_8_8_0[11|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1510 adc_array_wafflecap_8_Dummy_8[5]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1511 adc_array_wafflecap_8_8_0[14|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1512 adc_array_wafflecap_8_8_0[14|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1513 VDD rowon_n[12] adc_array_wafflecap_8_8_0[11|27]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1514 adc_array_wafflecap_8_8_0[4|0]/adc_array_circuit_150n_0/vint2 col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1515 adc_array_wafflecap_8_8_0[0|1]/adc_array_circuit_150n_0/vint2 col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1516 adc_array_wafflecap_8_8_0[1|9]/adc_array_circuit_150n_0/vdrv row_n[2] adc_array_wafflecap_8_8_0[1|9]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1517 adc_array_wafflecap_8_8_0[10|15]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|15]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1518 adc_array_wafflecap_8_8_0[3|13]/adc_array_circuit_150n_0/vint2 col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1519 adc_array_wafflecap_8_8_0[10|5]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|5]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1520 VDD rowon_n[11] adc_array_wafflecap_8_8_0[10|9]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1521 VDD rowon_n[11] adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1522 adc_array_wafflecap_8_8_0[9|24]/adc_array_circuit_150n_0/vdrv row_n[10] adc_array_wafflecap_8_8_0[9|24]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1523 adc_array_wafflecap_8_8_0[7|28]/adc_array_circuit_150n_0/vint1 col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1524 vcm adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1525 adc_array_wafflecap_8_8_0[4|25]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|25]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1526 adc_array_wafflecap_8_8_0[3|3]/adc_array_circuit_150n_0/vdrv row_n[4] adc_array_wafflecap_8_8_0[3|3]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1527 adc_array_wafflecap_8_8_0[0|26]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|26]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1528 adc_array_wafflecap_8_8_0[2|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1529 adc_array_wafflecap_8_8_0[14|26]/adc_array_circuit_150n_0/vint2 col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1530 adc_array_wafflecap_8_8_0[3|4]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|4]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1531 adc_array_wafflecap_8_8_0[13|30]/adc_array_circuit_150n_0/vint2 col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1532 adc_array_wafflecap_8_8_0[6|16]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|16]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1533 adc_array_wafflecap_8_8_1[21]/adc_array_circuit_150n_0/vdrv row_n[0] adc_array_wafflecap_8_8_1[21]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1534 adc_array_wafflecap_8_1_1/adc_array_circuit_150n_0/vdrv en_C0_n adc_array_wafflecap_8_1_1/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1535 adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/vint1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1536 adc_array_wafflecap_8_8_0[0|7]/adc_array_circuit_150n_0/vint2 rowon_n[1] adc_array_wafflecap_8_8_0[0|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1537 VSS row_n[14] adc_array_wafflecap_8_8_0[13|7]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1538 adc_array_wafflecap_8_8_0[4|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1539 adc_array_wafflecap_8_8_0[0|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1540 adc_array_wafflecap_8_8_0[2|5]/adc_array_circuit_150n_0/vint2 col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1541 adc_array_wafflecap_8_Dummy_4[30]/adc_array_circuit_150n_0/vint1 col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1542 adc_array_wafflecap_8_8_0[13|17]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|17]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1543 adc_array_wafflecap_8_8_0[12|26]/adc_array_circuit_150n_0/vdrv row_n[13] adc_array_wafflecap_8_8_0[12|26]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1544 adc_array_wafflecap_8_8_0[9|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1545 VDD rowon_n[4] adc_array_wafflecap_8_8_0[3|9]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1546 adc_array_wafflecap_8_8_0[6|0]/adc_array_circuit_150n_0/vint2 rowon_n[7] adc_array_wafflecap_8_8_0[6|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1547 VSS row_n[2] adc_array_wafflecap_8_8_0[1|19]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1548 adc_array_wafflecap_8_Dummy_4[29]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1549 adc_array_wafflecap_8_8_0[5|28]/adc_array_circuit_150n_0/vint2 rowon_n[6] adc_array_wafflecap_8_8_0[5|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1550 VDD VSS adc_array_wafflecap_8_Dummy_8[5]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1551 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X1552 adc_array_wafflecap_8_8_0[1|29]/adc_array_circuit_150n_0/vint2 rowon_n[2] adc_array_wafflecap_8_8_0[1|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1553 adc_array_wafflecap_8_8_0[12|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1554 vcm adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|29]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1555 adc_array_wafflecap_8_8_0[1|17]/adc_array_circuit_150n_0/vint2 col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1556 adc_array_wafflecap_8_Dummy_3[5]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_3[5]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1557 adc_array_wafflecap_8_Dummy_1[3]/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_1[3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1558 adc_array_wafflecap_8_8_0[0|5]/adc_array_circuit_150n_0/vdrv row_n[1] adc_array_wafflecap_8_8_0[0|5]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1559 adc_array_wafflecap_8_8_0[2|11]/adc_array_circuit_150n_0/vint2 rowon_n[3] adc_array_wafflecap_8_8_0[2|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1560 adc_array_wafflecap_8_8_0[11|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1561 adc_array_wafflecap_8_2_0/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1562 VDD rowon_n[3] adc_array_wafflecap_8_8_0[2|1]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1563 VSS row_n[1] adc_array_wafflecap_8_8_0[0|8]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1564 vcm adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|27]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1565 VDD rowon_n[7] adc_array_wafflecap_8_8_0[6|0]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1566 VSS row_n[5] adc_array_wafflecap_8_8_0[4|7]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1567 VSS sample adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1568 adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1569 adc_array_wafflecap_8_8_0[7|30]/adc_array_circuit_150n_0/vint2 rowon_n[8] adc_array_wafflecap_8_8_0[7|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1570 VDD rowon_n[6] adc_array_wafflecap_8_8_0[5|13]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1571 adc_array_wafflecap_8_Dummy_3[3]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_3[3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1572 VDD rowon_n[2] adc_array_wafflecap_8_8_0[1|29]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1573 adc_array_wafflecap_8_8_0[1|19]/adc_array_circuit_150n_0/vint1 col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1574 adc_array_wafflecap_8_8_0[2|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1575 adc_array_wafflecap_8_8_0[8|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1576 adc_array_wafflecap_8_8_0[7|8]/adc_array_circuit_150n_0/vint2 rowon_n[8] adc_array_wafflecap_8_8_0[7|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1577 adc_array_wafflecap_8_8_0[1|17]/adc_array_circuit_150n_0/vdrv row_n[2] adc_array_wafflecap_8_8_0[1|17]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1578 VSS VDD adc_array_wafflecap_8_Dummy_4[26]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1579 adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1580 VSS row_n[7] adc_array_wafflecap_8_8_0[6|1]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1581 adc_array_wafflecap_8_8_0[3|10]/adc_array_circuit_150n_0/vint1 col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1582 VDD rowon_n[1] adc_array_wafflecap_8_8_0[0|11]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1583 adc_array_wafflecap_8_Dummy_4[19]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[19]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1584 adc_array_wafflecap_8_8_0[13|7]/adc_array_circuit_150n_0/vint2 rowon_n[14] adc_array_wafflecap_8_8_0[13|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1585 adc_array_wafflecap_8_8_0[13|29]/adc_array_circuit_150n_0/vint2 rowon_n[14] adc_array_wafflecap_8_8_0[13|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1586 vcm adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|18]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1587 VDD rowon_n[12] adc_array_wafflecap_8_8_0[11|25]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1588 adc_array_wafflecap_8_4_0/adc_array_circuit_150n_0/vint1 en_n_bit[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1589 adc_array_wafflecap_8_8_0[0|16]/adc_array_circuit_150n_0/vint2 rowon_n[1] adc_array_wafflecap_8_8_0[0|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1590 adc_array_wafflecap_8_8_0[6|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1591 adc_array_wafflecap_8_8_0[4|15]/adc_array_circuit_150n_0/vint2 rowon_n[5] adc_array_wafflecap_8_8_0[4|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1592 VSS row_n[0] adc_array_wafflecap_8_Dummy_7/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1593 adc_array_wafflecap_8_8_0[2|26]/adc_array_circuit_150n_0/vint2 col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1594 adc_array_wafflecap_8_Dummy_4[13]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1595 adc_array_wafflecap_8_8_0[12|9]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|9]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1596 VSS VSS adc_array_wafflecap_8_Dummy_1[4]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1597 adc_array_wafflecap_8_Dummy_4[3]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1598 VDD sample_n adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1599 VDD rowon_n[5] adc_array_wafflecap_8_8_0[4|5]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1600 vcm adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|22]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1601 VSS row_n[3] adc_array_wafflecap_8_8_0[2|12]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1602 adc_array_wafflecap_8_8_0[13|25]/adc_array_circuit_150n_0/vint1 col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1603 adc_array_wafflecap_8_8_0[11|13]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|13]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1604 adc_array_wafflecap_8_8_0[7|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1605 adc_array_wafflecap_8_8_0[5|28]/adc_array_circuit_150n_0/vdrv row_n[6] adc_array_wafflecap_8_8_0[5|28]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1606 adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1607 vcm adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|0]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1608 adc_array_wafflecap_8_8_1[24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1609 adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1610 adc_array_wafflecap_8_8_0[11|3]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|3]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1611 adc_array_wafflecap_8_8_0[6|1]/adc_array_circuit_150n_0/vint1 col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1612 adc_array_wafflecap_8_8_0[5|29]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|29]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1613 adc_array_wafflecap_8_8_0[2|2]/adc_array_circuit_150n_0/vint1 col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1614 adc_array_wafflecap_8_8_0[2|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1615 VDD rowon_n[0] adc_array_wafflecap_8_8_1[2]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1616 vcm adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|12]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1617 adc_array_wafflecap_8_8_0[5|14]/adc_array_circuit_150n_0/vint1 col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1618 adc_array_wafflecap_8_8_0[5|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1619 VDD en_n_bit[1] adc_array_wafflecap_8_2_0/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1620 adc_array_wafflecap_8_8_0[9|15]/adc_array_circuit_150n_0/vint2 col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1621 VSS row_n[9] adc_array_wafflecap_8_8_0[8|6]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1622 adc_array_wafflecap_8_8_0[0|26]/adc_array_circuit_150n_0/vdrv row_n[1] adc_array_wafflecap_8_8_0[0|26]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1623 adc_array_wafflecap_8_8_0[9|5]/adc_array_circuit_150n_0/vint2 col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1624 adc_array_wafflecap_8_8_0[0|12]/adc_array_circuit_150n_0/vint1 col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1625 adc_array_wafflecap_8_8_0[4|30]/adc_array_circuit_150n_0/vint2 col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1626 vcm adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[10]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1627 adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/vint2 col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1628 adc_array_wafflecap_8_Dummy_4[5]/adc_array_circuit_150n_0/vint2 col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1629 adc_array_wafflecap_8_Dummy_4[15]/adc_array_circuit_150n_0/vint2 col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1630 VSS row_n[14] adc_array_wafflecap_8_8_0[13|18]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1631 VSS row_n[7] adc_array_wafflecap_8_8_0[6|23]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1632 adc_array_wafflecap_8_8_0[11|14]/adc_array_circuit_150n_0/vint1 col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1633 adc_array_wafflecap_8_8_0[7|24]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|24]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1634 adc_array_wafflecap_8_Dummy_4[27]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1635 vcm adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|23]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1636 adc_array_wafflecap_8_8_0[11|4]/adc_array_circuit_150n_0/vint1 col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1637 adc_array_wafflecap_8_8_0[10|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1638 adc_array_wafflecap_8_8_0[0|18]/adc_array_circuit_150n_0/vint2 rowon_n[1] adc_array_wafflecap_8_8_0[0|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1639 vcm adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|5]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1640 adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1641 adc_array_wafflecap_8_8_0[7|15]/adc_array_circuit_150n_0/vdrv row_n[8] adc_array_wafflecap_8_8_0[7|15]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1642 adc_array_wafflecap_8_8_0[7|5]/adc_array_circuit_150n_0/vdrv row_n[8] adc_array_wafflecap_8_8_0[7|5]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1643 VSS row_n[1] adc_array_wafflecap_8_8_0[0|16]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1644 adc_array_wafflecap_8_8_0[12|17]/adc_array_circuit_150n_0/vint2 col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1645 VDD rowon_n[4] adc_array_wafflecap_8_8_0[3|20]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1646 adc_array_wafflecap_8_8_1[3]/adc_array_circuit_150n_0/vint1 col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1647 adc_array_wafflecap_8_8_0[13|4]/adc_array_circuit_150n_0/vdrv row_n[14] adc_array_wafflecap_8_8_0[13|4]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1648 adc_array_wafflecap_8_8_0[13|14]/adc_array_circuit_150n_0/vdrv row_n[14] adc_array_wafflecap_8_8_0[13|14]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1649 vcm adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|4]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1650 vcm adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|14]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1651 adc_array_wafflecap_8_8_0[6|23]/adc_array_circuit_150n_0/vint1 col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1652 VDD VSS adc_array_wafflecap_8_Dummy_2[1]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1653 adc_array_wafflecap_8_8_0[14|16]/adc_array_circuit_150n_0/vint1 col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1654 adc_array_wafflecap_8_8_0[14|23]/adc_array_circuit_150n_0/vint2 rowon_n[15] adc_array_wafflecap_8_8_0[14|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1655 adc_array_wafflecap_8_2_0/adc_array_circuit_150n_0/vint1 en_n_bit[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1656 adc_array_wafflecap_8_Dummy_2[6]/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_2[6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1657 adc_array_wafflecap_8_8_0[10|17]/adc_array_circuit_150n_0/vdrv row_n[11] adc_array_wafflecap_8_8_0[10|17]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1658 VSS row_n[11] adc_array_wafflecap_8_8_0[10|24]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1659 adc_array_wafflecap_8_8_0[8|28]/adc_array_circuit_150n_0/vint2 rowon_n[9] adc_array_wafflecap_8_8_0[8|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1660 adc_array_wafflecap_8_8_0[7|21]/adc_array_circuit_150n_0/vint2 col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1661 adc_array_wafflecap_8_8_0[3|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1662 vcm VSS adc_array_wafflecap_8_Dummy_4[16]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1663 adc_array_wafflecap_8_Dummy_8[0]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_8[0]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1664 vcm VSS adc_array_wafflecap_8_Dummy_4[6]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1665 vcm adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|26]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1666 VDD rowon_n[13] adc_array_wafflecap_8_8_0[12|23]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1667 adc_array_wafflecap_8_8_0[10|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1668 adc_array_wafflecap_8_8_0[10|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1669 adc_array_wafflecap_8_8_0[9|20]/adc_array_circuit_150n_0/vint1 col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1670 VDD rowon_n[12] adc_array_wafflecap_8_8_0[11|4]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1671 VDD rowon_n[12] adc_array_wafflecap_8_8_0[11|14]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1672 adc_array_wafflecap_8_8_0[8|24]/adc_array_circuit_150n_0/vint1 col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1673 adc_array_wafflecap_8_8_0[3|6]/adc_array_circuit_150n_0/vint2 col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1674 adc_array_wafflecap_8_Dummy_0[1]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_0[1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1675 adc_array_wafflecap_8_8_1[20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_1[20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1676 adc_array_wafflecap_8_Dummy_4[23]/adc_array_circuit_150n_0/vint2 col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1677 VSS row_n[14] adc_array_wafflecap_8_8_0[13|26]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1678 adc_array_wafflecap_8_8_0[4|27]/adc_array_circuit_150n_0/vint1 col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1679 adc_array_wafflecap_8_8_0[4|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1680 adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1681 adc_array_wafflecap_8_8_0[8|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1682 adc_array_wafflecap_8_8_0[6|9]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|9]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1683 VSS row_n[7] adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1684 adc_array_wafflecap_8_8_0[5|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1685 adc_array_wafflecap_8_8_0[1|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1686 VSS row_n[15] adc_array_wafflecap_8_8_0[14|12]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1687 VSS row_n[15] adc_array_wafflecap_8_8_0[14|2]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1688 adc_array_wafflecap_8_8_0[10|13]/adc_array_circuit_150n_0/vint2 col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1689 VSS row_n[9] adc_array_wafflecap_8_8_0[8|17]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1690 VSS row_n[0] adc_array_wafflecap_8_8_1[29]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1691 adc_array_wafflecap_8_8_1[19]/adc_array_circuit_150n_0/vint2 col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1692 adc_array_wafflecap_8_8_0[10|3]/adc_array_circuit_150n_0/vint2 col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1693 adc_array_wafflecap_8_8_0[5|22]/adc_array_circuit_150n_0/vint2 rowon_n[6] adc_array_wafflecap_8_8_0[5|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1694 adc_array_wafflecap_8_Dummy_0[0]/adc_array_circuit_150n_0/vint2 VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1695 adc_array_wafflecap_8_8_0[13|22]/adc_array_circuit_150n_0/vdrv row_n[14] adc_array_wafflecap_8_8_0[13|22]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1696 vcm adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|22]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1697 adc_array_wafflecap_8_8_0[5|10]/adc_array_circuit_150n_0/vint2 col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1698 adc_array_wafflecap_8_8_0[1|11]/adc_array_circuit_150n_0/vint2 col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1699 vcm adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|30]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1700 adc_array_wafflecap_8_8_0[2|22]/adc_array_circuit_150n_0/vdrv row_n[3] adc_array_wafflecap_8_8_0[2|22]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1701 adc_array_wafflecap_8_8_0[2|23]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|23]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1702 adc_array_wafflecap_8_1_0/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_1_0/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1703 vcm adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|21]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1704 adc_array_wafflecap_8_8_0[12|12]/adc_array_circuit_150n_0/vint1 col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1705 adc_array_wafflecap_8_8_0[9|9]/adc_array_circuit_150n_0/vdrv row_n[10] adc_array_wafflecap_8_8_0[9|9]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1706 adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/vint1 col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1707 adc_array_wafflecap_8_8_0[5|0]/adc_array_circuit_150n_0/vdrv row_n[6] adc_array_wafflecap_8_8_0[5|0]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1708 adc_array_wafflecap_8_8_0[5|1]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|1]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1709 adc_array_wafflecap_8_8_0[0|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1710 adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/vint1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1711 adc_array_wafflecap_8_8_0[12|2]/adc_array_circuit_150n_0/vint1 col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1712 adc_array_wafflecap_8_8_0[3|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1713 adc_array_wafflecap_8_8_0[9|26]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|26]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1714 adc_array_wafflecap_8_8_0[8|3]/adc_array_circuit_150n_0/vdrv row_n[9] adc_array_wafflecap_8_8_0[8|3]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1715 adc_array_wafflecap_8_8_0[8|13]/adc_array_circuit_150n_0/vdrv row_n[9] adc_array_wafflecap_8_8_0[8|13]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1716 adc_array_wafflecap_8_8_0[11|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1717 adc_array_wafflecap_8_Dummy_1[0]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1718 adc_array_wafflecap_8_8_0[1|11]/adc_array_circuit_150n_0/vdrv row_n[2] adc_array_wafflecap_8_8_0[1|11]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1719 adc_array_wafflecap_8_8_0[11|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1720 adc_array_wafflecap_8_8_0[4|2]/adc_array_circuit_150n_0/vint2 col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1721 adc_array_wafflecap_8_8_0[0|3]/adc_array_circuit_150n_0/vint2 col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1722 vcm adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|19]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1723 adc_array_wafflecap_8_8_0[3|15]/adc_array_circuit_150n_0/vint2 col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1724 adc_array_wafflecap_8_Dummy_4[22]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1725 adc_array_wafflecap_8_8_0[3|5]/adc_array_circuit_150n_0/vdrv row_n[4] adc_array_wafflecap_8_8_0[3|5]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1726 adc_array_wafflecap_8_8_0[3|6]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|6]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1727 adc_array_wafflecap_8_8_0[3|26]/adc_array_circuit_150n_0/vint2 rowon_n[4] adc_array_wafflecap_8_8_0[3|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1728 adc_array_wafflecap_8_8_0[14|2]/adc_array_circuit_150n_0/vint2 rowon_n[15] adc_array_wafflecap_8_8_0[14|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1729 adc_array_wafflecap_8_8_0[14|12]/adc_array_circuit_150n_0/vint2 rowon_n[15] adc_array_wafflecap_8_8_0[14|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1730 VSS row_n[12] adc_array_wafflecap_8_8_0[11|22]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1731 adc_array_wafflecap_8_Dummy_4[32]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1732 adc_array_wafflecap_8_8_0[13|16]/adc_array_circuit_150n_0/vint2 rowon_n[14] adc_array_wafflecap_8_8_0[13|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1733 adc_array_wafflecap_8_8_0[12|28]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|28]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1734 adc_array_wafflecap_8_Dummy_8[1]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_8[1]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1735 adc_array_wafflecap_8_8_0[13|6]/adc_array_circuit_150n_0/vint2 rowon_n[14] adc_array_wafflecap_8_8_0[13|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1736 adc_array_wafflecap_8_8_0[8|17]/adc_array_circuit_150n_0/vint2 rowon_n[9] adc_array_wafflecap_8_8_0[8|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1737 adc_array_wafflecap_8_8_0[6|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1738 adc_array_wafflecap_8_8_0[4|8]/adc_array_circuit_150n_0/vint2 rowon_n[5] adc_array_wafflecap_8_8_0[4|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1739 adc_array_wafflecap_8_8_0[0|9]/adc_array_circuit_150n_0/vint2 rowon_n[1] adc_array_wafflecap_8_8_0[0|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1740 adc_array_wafflecap_8_8_0[0|27]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|27]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1741 adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1742 adc_array_wafflecap_8_8_0[4|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1743 VDD rowon_n[14] adc_array_wafflecap_8_8_0[13|21]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1744 adc_array_wafflecap_8_8_0[11|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1745 adc_array_wafflecap_8_8_0[6|17]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|17]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1746 VDD rowon_n[13] adc_array_wafflecap_8_8_0[12|12]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1747 adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1748 VDD rowon_n[4] adc_array_wafflecap_8_8_0[3|11]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1749 VDD rowon_n[13] adc_array_wafflecap_8_8_0[12|2]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1750 VSS row_n[2] adc_array_wafflecap_8_8_0[1|21]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1751 adc_array_wafflecap_8_8_0[8|17]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|17]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1752 adc_array_wafflecap_8_8_0[5|7]/adc_array_circuit_150n_0/vint1 col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1753 VDD VSS adc_array_wafflecap_8_Dummy_1[0]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1754 adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/vint2 rowon_n[2] adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1755 VSS row_n[10] adc_array_wafflecap_8_8_0[9|1]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1756 VSS row_n[10] adc_array_wafflecap_8_8_0[9|11]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1757 adc_array_wafflecap_8_8_0[5|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1758 adc_array_wafflecap_8_8_0[5|30]/adc_array_circuit_150n_0/vint2 rowon_n[6] adc_array_wafflecap_8_8_0[5|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1759 adc_array_wafflecap_8_8_0[4|24]/adc_array_circuit_150n_0/vint2 col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1760 adc_array_wafflecap_8_Dummy_6/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_6/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1761 adc_array_wafflecap_8_8_1[0]/adc_array_circuit_150n_0/vint2 rowon_n[0] adc_array_wafflecap_8_8_1[0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1762 VSS VDD adc_array_wafflecap_8_Dummy_4[11]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1763 adc_array_wafflecap_8_Dummy_1[5]/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_1[5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1764 adc_array_wafflecap_8_8_0[2|13]/adc_array_circuit_150n_0/vint2 rowon_n[3] adc_array_wafflecap_8_8_0[2|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1765 VSS VDD adc_array_wafflecap_8_Dummy_4[1]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1766 adc_array_wafflecap_8_8_0[7|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1767 adc_array_wafflecap_8_8_0[14|29]/adc_array_circuit_150n_0/vdrv row_n[15] adc_array_wafflecap_8_8_0[14|29]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1768 adc_array_wafflecap_8_8_0[12|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1769 adc_array_wafflecap_8_8_0[11|1]/adc_array_circuit_150n_0/vint2 col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1770 adc_array_wafflecap_8_8_0[11|11]/adc_array_circuit_150n_0/vint2 col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1771 VSS row_n[5] adc_array_wafflecap_8_8_0[4|9]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1772 VDD rowon_n[3] adc_array_wafflecap_8_8_0[2|3]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1773 analog_in sw_n ctop VDD sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=5.9e+11p ps=3.18e+06u w=1e+06u l=1e+06u
X1774 VSS row_n[1] adc_array_wafflecap_8_8_0[0|10]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1775 adc_array_wafflecap_8_8_0[7|11]/adc_array_circuit_150n_0/vint1 col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1776 VDD rowon_n[6] adc_array_wafflecap_8_8_0[5|15]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1777 adc_array_wafflecap_8_Dummy_3[5]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_3[5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1778 vcm VSS adc_array_wafflecap_8_Dummy_2[3]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1779 adc_array_wafflecap_8_8_0[1|21]/adc_array_circuit_150n_0/vint1 col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1780 vcm adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|20]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1781 adc_array_wafflecap_8_8_0[7|1]/adc_array_circuit_150n_0/vint1 col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1782 adc_array_wafflecap_8_8_0[3|26]/adc_array_circuit_150n_0/vdrv row_n[4] adc_array_wafflecap_8_8_0[3|26]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1783 VDD rowon_n[2] adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1784 adc_array_wafflecap_8_8_0[2|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1785 adc_array_wafflecap_8_8_0[4|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1786 adc_array_wafflecap_8_8_0[3|12]/adc_array_circuit_150n_0/vint1 col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1787 adc_array_wafflecap_8_8_0[14|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1788 adc_array_wafflecap_8_8_0[13|0]/adc_array_circuit_150n_0/vint1 col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1789 adc_array_wafflecap_8_8_0[13|10]/adc_array_circuit_150n_0/vint1 col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1790 adc_array_wafflecap_8_8_0[7|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1791 adc_array_wafflecap_8_8_0[7|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1792 adc_array_wafflecap_8_8_0[3|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1793 VDD rowon_n[1] adc_array_wafflecap_8_8_0[0|13]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1794 adc_array_wafflecap_8_8_0[10|24]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|24]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1795 adc_array_wafflecap_8_Dummy_1[1]/adc_array_circuit_150n_0/vint1 col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1796 adc_array_wafflecap_8_Dummy_3[4]/adc_array_circuit_150n_0/vint2 col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1797 VSS row_n[0] adc_array_wafflecap_8_8_1[1]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1798 adc_array_wafflecap_8_8_0[2|28]/adc_array_circuit_150n_0/vint2 col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1799 VSS VSS adc_array_wafflecap_8_Dummy_1[6]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1800 VSS row_n[3] adc_array_wafflecap_8_8_0[2|14]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1801 adc_array_wafflecap_8_8_0[10|20]/adc_array_circuit_150n_0/vint2 rowon_n[11] adc_array_wafflecap_8_8_0[10|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1802 adc_array_wafflecap_8_8_0[9|1]/adc_array_circuit_150n_0/vint2 rowon_n[10] adc_array_wafflecap_8_8_0[9|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1803 adc_array_wafflecap_8_8_0[9|11]/adc_array_circuit_150n_0/vint2 rowon_n[10] adc_array_wafflecap_8_8_0[9|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1804 adc_array_wafflecap_8_8_0[5|30]/adc_array_circuit_150n_0/vdrv row_n[6] adc_array_wafflecap_8_8_0[5|30]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1805 adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1806 vcm adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|2]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1807 adc_array_wafflecap_8_8_0[2|4]/adc_array_circuit_150n_0/vint1 col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1808 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X1809 adc_array_wafflecap_8_Dummy_4[12]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1810 vcm adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|8]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1811 VDD sample_n adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1812 adc_array_wafflecap_8_8_0[7|9]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|9]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1813 adc_array_wafflecap_8_8_0[2|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1814 VDD rowon_n[0] adc_array_wafflecap_8_8_1[4]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1815 adc_array_wafflecap_8_Dummy_4[2]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1816 adc_array_wafflecap_8_Dummy_4[33]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[33]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1817 adc_array_wafflecap_8_8_0[8|5]/adc_array_circuit_150n_0/vint2 rowon_n[9] adc_array_wafflecap_8_8_0[8|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1818 adc_array_wafflecap_8_8_0[8|15]/adc_array_circuit_150n_0/vint2 rowon_n[9] adc_array_wafflecap_8_8_0[8|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1819 adc_array_wafflecap_8_8_0[0|28]/adc_array_circuit_150n_0/vdrv row_n[1] adc_array_wafflecap_8_8_0[0|28]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1820 vcm adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|2]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1821 vcm adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|12]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1822 vcm adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[12]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1823 adc_array_wafflecap_8_8_0[0|14]/adc_array_circuit_150n_0/vint1 col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1824 adc_array_wafflecap_8_8_0[1|7]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|7]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1825 VDD rowon_n[9] adc_array_wafflecap_8_8_0[8|20]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1826 VSS row_n[7] adc_array_wafflecap_8_8_0[6|25]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1827 adc_array_wafflecap_8_8_0[4|19]/adc_array_circuit_150n_0/vdrv row_n[5] adc_array_wafflecap_8_8_0[4|19]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1828 adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/vint2 VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1829 adc_array_wafflecap_8_8_0[1|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1830 VDD rowon_n[8] adc_array_wafflecap_8_8_0[7|1]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1831 VDD rowon_n[8] adc_array_wafflecap_8_8_0[7|11]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1832 VSS row_n[15] adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1833 adc_array_wafflecap_8_8_0[13|16]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|16]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1834 VDD rowon_n[14] adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1835 adc_array_wafflecap_8_8_0[13|6]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|6]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1836 adc_array_wafflecap_8_8_0[0|20]/adc_array_circuit_150n_0/vint2 rowon_n[1] adc_array_wafflecap_8_8_0[0|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1837 adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/vint2 VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1838 VSS row_n[11] adc_array_wafflecap_8_8_0[10|9]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1839 adc_array_wafflecap_8_8_0[7|6]/adc_array_circuit_150n_0/vint2 col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1840 adc_array_wafflecap_8_8_0[6|25]/adc_array_circuit_150n_0/vint1 col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1841 adc_array_wafflecap_8_8_0[3|17]/adc_array_circuit_150n_0/vint2 rowon_n[4] adc_array_wafflecap_8_8_0[3|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1842 vcm adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|24]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1843 adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/vint1 col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1844 adc_array_wafflecap_8_8_0[9|28]/adc_array_circuit_150n_0/vdrv row_n[10] adc_array_wafflecap_8_8_0[9|28]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1845 VDD VSS adc_array_wafflecap_8_Dummy_2[3]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1846 adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/vdrv row_n[9] adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1847 vcm adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|26]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1848 adc_array_wafflecap_8_8_0[12|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1849 adc_array_wafflecap_8_8_0[9|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1850 adc_array_wafflecap_8_8_0[8|9]/adc_array_circuit_150n_0/vint1 col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1851 adc_array_wafflecap_8_8_0[3|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1852 adc_array_wafflecap_8_Dummy_3[0]/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_3[0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1853 vcm adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1854 adc_array_wafflecap_8_Dummy_4[8]/adc_array_circuit_150n_0/vint2 col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1855 adc_array_wafflecap_8_8_0[8|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1856 adc_array_wafflecap_8_8_0[3|8]/adc_array_circuit_150n_0/vint2 col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1857 VSS row_n[4] adc_array_wafflecap_8_8_0[3|18]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1858 adc_array_wafflecap_8_8_0[13|7]/adc_array_circuit_150n_0/vdrv row_n[14] adc_array_wafflecap_8_8_0[13|7]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1859 adc_array_wafflecap_8_8_0[11|18]/adc_array_circuit_150n_0/vint2 rowon_n[12] adc_array_wafflecap_8_8_0[11|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1860 vcm adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|7]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1861 vcm adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|27]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1862 adc_array_wafflecap_8_8_0[4|20]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|20]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1863 adc_array_wafflecap_8_8_0[4|29]/adc_array_circuit_150n_0/vint1 col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1864 adc_array_wafflecap_8_Dummy_8[0]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_8[0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1865 adc_array_wafflecap_8_8_0[0|21]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|21]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1866 vcm adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|28]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1867 adc_array_wafflecap_8_8_0[2|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1868 adc_array_wafflecap_8_8_0[14|20]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|20]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1869 adc_array_wafflecap_8_8_0[10|9]/adc_array_circuit_150n_0/vint2 rowon_n[11] adc_array_wafflecap_8_8_0[10|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1870 adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/vint2 rowon_n[11] adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1871 adc_array_wafflecap_8_8_0[9|24]/adc_array_circuit_150n_0/vint2 col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1872 VSS row_n[8] adc_array_wafflecap_8_8_0[7|28]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1873 adc_array_wafflecap_8_8_0[4|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1874 VDD sample_n adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1875 adc_array_wafflecap_8_8_0[1|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1876 adc_array_wafflecap_8_8_0[6|11]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|11]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1877 vcm adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|19]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1878 adc_array_wafflecap_8_8_1[26]/adc_array_circuit_150n_0/vint1 col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1879 adc_array_wafflecap_8_8_1[21]/adc_array_circuit_150n_0/vint2 col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1880 adc_array_wafflecap_8_8_0[12|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1881 adc_array_wafflecap_8_8_0[12|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1882 adc_array_wafflecap_8_8_0[11|23]/adc_array_circuit_150n_0/vint1 col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1883 adc_array_wafflecap_8_8_0[9|1]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|1]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1884 adc_array_wafflecap_8_8_0[9|11]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|11]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1885 VDD rowon_n[10] adc_array_wafflecap_8_8_0[9|27]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1886 VSS row_n[0] adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1887 adc_array_wafflecap_8_1_1/adc_array_circuit_150n_0/vint2 en_C0_n VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1888 adc_array_wafflecap_8_8_0[2|0]/adc_array_circuit_150n_0/vint2 col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1889 adc_array_wafflecap_8_8_0[5|24]/adc_array_circuit_150n_0/vint2 rowon_n[6] adc_array_wafflecap_8_8_0[5|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1890 adc_array_wafflecap_8_8_0[1|13]/adc_array_circuit_150n_0/vint2 col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1891 VDD rowon_n[9] adc_array_wafflecap_8_8_0[8|9]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1892 VDD rowon_n[9] adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1893 adc_array_wafflecap_8_8_0[7|24]/adc_array_circuit_150n_0/vdrv row_n[8] adc_array_wafflecap_8_8_0[7|24]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1894 adc_array_wafflecap_8_8_0[5|12]/adc_array_circuit_150n_0/vint2 col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1895 VSS VDD adc_array_wafflecap_8_Dummy_4[30]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1896 vcm adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1897 adc_array_wafflecap_8_8_0[2|25]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|25]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1898 adc_array_wafflecap_8_Dummy_3[1]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_3[1]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1899 adc_array_wafflecap_8_8_0[0|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1900 adc_array_wafflecap_8_8_0[12|26]/adc_array_circuit_150n_0/vint2 col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1901 adc_array_wafflecap_8_8_0[5|2]/adc_array_circuit_150n_0/vdrv row_n[6] adc_array_wafflecap_8_8_0[5|2]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1902 adc_array_wafflecap_8_8_0[5|3]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|3]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1903 adc_array_wafflecap_8_8_0[1|4]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|4]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1904 adc_array_wafflecap_8_8_0[11|30]/adc_array_circuit_150n_0/vint2 col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1905 adc_array_wafflecap_8_Dummy_8[5]/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_8[5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1906 adc_array_wafflecap_8_8_0[0|0]/adc_array_circuit_150n_0/vdrv row_n[1] adc_array_wafflecap_8_8_0[0|0]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1907 VSS row_n[12] adc_array_wafflecap_8_8_0[11|7]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1908 adc_array_wafflecap_8_Dummy_1[2]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1909 adc_array_wafflecap_8_8_0[2|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1910 adc_array_wafflecap_8_8_0[0|5]/adc_array_circuit_150n_0/vint2 col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1911 adc_array_wafflecap_8_8_0[1|13]/adc_array_circuit_150n_0/vdrv row_n[2] adc_array_wafflecap_8_8_0[1|13]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1912 adc_array_wafflecap_8_Dummy_4[26]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[26]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1913 adc_array_wafflecap_8_8_0[13|29]/adc_array_circuit_150n_0/vint1 col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1914 adc_array_wafflecap_8_8_0[11|17]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|17]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1915 adc_array_wafflecap_8_8_0[10|26]/adc_array_circuit_150n_0/vdrv row_n[11] adc_array_wafflecap_8_8_0[10|26]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1916 vcm adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|25]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1917 adc_array_wafflecap_8_8_0[7|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1918 VDD rowon_n[6] adc_array_wafflecap_8_8_0[5|8]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1919 vcm VSS adc_array_wafflecap_8_Dummy_4[25]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1920 adc_array_wafflecap_8_8_0[14|15]/adc_array_circuit_150n_0/vint1 col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1921 adc_array_wafflecap_8_8_0[14|5]/adc_array_circuit_150n_0/vint1 col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1922 adc_array_wafflecap_8_8_0[13|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1923 adc_array_wafflecap_8_8_0[3|28]/adc_array_circuit_150n_0/vint2 rowon_n[4] adc_array_wafflecap_8_8_0[3|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1924 adc_array_wafflecap_8_8_0[10|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1925 adc_array_wafflecap_8_Dummy_8[3]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_8[3]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1926 adc_array_wafflecap_8_8_0[0|11]/adc_array_circuit_150n_0/vint2 rowon_n[1] adc_array_wafflecap_8_8_0[0|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1927 adc_array_wafflecap_8_Dummy_4[19]/adc_array_circuit_150n_0/vint2 col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1928 adc_array_wafflecap_8_8_0[6|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1929 adc_array_wafflecap_8_8_0[5|24]/adc_array_circuit_150n_0/vdrv row_n[6] adc_array_wafflecap_8_8_0[5|24]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1930 adc_array_wafflecap_8_8_0[4|10]/adc_array_circuit_150n_0/vint2 rowon_n[5] adc_array_wafflecap_8_8_0[4|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1931 adc_array_wafflecap_8_8_0[7|28]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|28]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1932 VSS en_n_bit[2] adc_array_wafflecap_8_4_0/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1933 vcm adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|27]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1934 VDD rowon_n[5] adc_array_wafflecap_8_8_0[4|0]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1935 VSS row_n[3] adc_array_wafflecap_8_8_0[2|7]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1936 VSS sample adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1937 VDD rowon_n[4] adc_array_wafflecap_8_8_0[3|13]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1938 adc_array_wafflecap_8_8_1[19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1939 adc_array_wafflecap_8_8_0[0|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1940 VSS row_n[14] adc_array_wafflecap_8_8_0[13|25]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1941 vcm adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|7]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1942 adc_array_wafflecap_8_8_0[6|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1943 adc_array_wafflecap_8_8_0[5|9]/adc_array_circuit_150n_0/vint1 col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1944 adc_array_wafflecap_8_8_0[5|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1945 VDD VSS adc_array_wafflecap_8_Dummy_1[2]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1946 adc_array_wafflecap_8_8_1[17]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[17]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1947 adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1948 adc_array_wafflecap_8_8_0[13|18]/adc_array_circuit_150n_0/vdrv row_n[14] adc_array_wafflecap_8_8_0[13|18]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1949 adc_array_wafflecap_8_8_0[11|7]/adc_array_circuit_150n_0/vint2 rowon_n[12] adc_array_wafflecap_8_8_0[11|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1950 adc_array_wafflecap_8_8_0[11|29]/adc_array_circuit_150n_0/vint2 rowon_n[12] adc_array_wafflecap_8_8_0[11|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1951 vcm adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|18]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1952 adc_array_wafflecap_8_8_1[2]/adc_array_circuit_150n_0/vint2 rowon_n[0] adc_array_wafflecap_8_8_1[2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1953 VDD rowon_n[10] adc_array_wafflecap_8_8_0[9|25]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1954 adc_array_wafflecap_8_2_0/adc_array_circuit_150n_0/vint2 en_n_bit[1] adc_array_wafflecap_8_2_0/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1955 adc_array_wafflecap_8_8_0[0|7]/adc_array_circuit_150n_0/vint1 col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1956 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.64e+07u l=1.6e+07u
X1957 adc_array_wafflecap_8_8_0[14|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1958 adc_array_wafflecap_8_8_0[0|26]/adc_array_circuit_150n_0/vint2 col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1959 adc_array_wafflecap_8_8_0[2|15]/adc_array_circuit_150n_0/vint2 rowon_n[3] adc_array_wafflecap_8_8_0[2|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1960 VDD VDD adc_array_wafflecap_8_Dummy_4[25]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1961 adc_array_wafflecap_8_8_0[13|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1962 adc_array_wafflecap_8_8_0[10|9]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|9]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1963 adc_array_wafflecap_8_8_0[13|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1964 VDD sample_n adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1965 adc_array_wafflecap_8_8_0[6|16]/adc_array_circuit_150n_0/vint2 col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1966 VSS row_n[5] adc_array_wafflecap_8_8_0[4|11]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1967 VDD rowon_n[3] adc_array_wafflecap_8_8_0[2|5]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1968 vcm VSS adc_array_wafflecap_8_Dummy_2[5]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1969 VSS row_n[1] adc_array_wafflecap_8_8_0[0|12]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1970 adc_array_wafflecap_8_8_0[3|28]/adc_array_circuit_150n_0/vdrv row_n[4] adc_array_wafflecap_8_8_0[3|28]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1971 adc_array_wafflecap_8_Dummy_6/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_6/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1972 vcm adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|0]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1973 adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1974 adc_array_wafflecap_8_8_0[4|1]/adc_array_circuit_150n_0/vint1 col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1975 adc_array_wafflecap_8_8_0[4|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1976 adc_array_wafflecap_8_8_0[3|29]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|29]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1977 adc_array_wafflecap_8_8_0[0|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1978 adc_array_wafflecap_8_8_0[3|14]/adc_array_circuit_150n_0/vint1 col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1979 adc_array_wafflecap_8_8_0[3|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1980 VDD rowon_n[1] adc_array_wafflecap_8_8_0[0|15]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1981 adc_array_wafflecap_8_8_0[11|20]/adc_array_circuit_150n_0/vdrv row_n[12] adc_array_wafflecap_8_8_0[11|20]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1982 adc_array_wafflecap_8_8_0[7|15]/adc_array_circuit_150n_0/vint2 col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1983 VSS sample adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1984 adc_array_wafflecap_8_Dummy_3[1]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_3[1]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1985 adc_array_wafflecap_8_8_0[7|5]/adc_array_circuit_150n_0/vint2 col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1986 adc_array_wafflecap_8_Dummy_1[3]/adc_array_circuit_150n_0/vint1 col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1987 adc_array_wafflecap_8_8_0[2|30]/adc_array_circuit_150n_0/vint2 col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1988 adc_array_wafflecap_8_8_0[14|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1989 adc_array_wafflecap_8_8_0[13|4]/adc_array_circuit_150n_0/vint2 col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1990 adc_array_wafflecap_8_8_0[13|14]/adc_array_circuit_150n_0/vint2 col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1991 VSS row_n[12] adc_array_wafflecap_8_8_0[11|18]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1992 adc_array_wafflecap_8_8_0[6|16]/adc_array_circuit_150n_0/vdrv row_n[7] adc_array_wafflecap_8_8_0[6|16]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1993 VSS row_n[0] adc_array_wafflecap_8_8_1[3]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1994 adc_array_wafflecap_8_8_0[9|14]/adc_array_circuit_150n_0/vint1 col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1995 adc_array_wafflecap_8_8_0[13|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1996 vcm adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|23]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1997 adc_array_wafflecap_8_8_0[9|4]/adc_array_circuit_150n_0/vint1 col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1998 adc_array_wafflecap_8_8_0[8|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1999 adc_array_wafflecap_8_Dummy_2[1]/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_2[1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2000 VSS row_n[15] adc_array_wafflecap_8_8_0[14|16]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2001 adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2002 adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/vdrv row_n[6] adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2003 adc_array_wafflecap_8_Dummy_4[4]/adc_array_circuit_150n_0/vint1 col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2004 adc_array_wafflecap_8_Dummy_4[14]/adc_array_circuit_150n_0/vint1 col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2005 adc_array_wafflecap_8_8_0[9|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2006 adc_array_wafflecap_8_8_0[9|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2007 VSS en_n_bit[1] adc_array_wafflecap_8_2_0/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2008 adc_array_wafflecap_8_8_0[10|17]/adc_array_circuit_150n_0/vint2 col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2009 adc_array_wafflecap_8_8_0[0|30]/adc_array_circuit_150n_0/vdrv row_n[1] adc_array_wafflecap_8_8_0[0|30]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2010 vcm adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|21]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2011 adc_array_wafflecap_8_8_0[4|23]/adc_array_circuit_150n_0/vint1 col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2012 vcm adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[14]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2013 adc_array_wafflecap_8_8_0[14|2]/adc_array_circuit_150n_0/vdrv row_n[15] adc_array_wafflecap_8_8_0[14|2]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2014 adc_array_wafflecap_8_8_0[14|12]/adc_array_circuit_150n_0/vdrv row_n[15] adc_array_wafflecap_8_8_0[14|12]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2015 adc_array_wafflecap_8_8_0[12|16]/adc_array_circuit_150n_0/vint1 col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2016 adc_array_wafflecap_8_8_0[12|23]/adc_array_circuit_150n_0/vint2 rowon_n[13] adc_array_wafflecap_8_8_0[12|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2017 VSS row_n[10] adc_array_wafflecap_8_8_0[9|20]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2018 vcm adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|11]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2019 adc_array_wafflecap_8_8_0[9|30]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|30]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2020 adc_array_wafflecap_8_8_0[8|17]/adc_array_circuit_150n_0/vdrv row_n[9] adc_array_wafflecap_8_8_0[8|17]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2021 VSS row_n[9] adc_array_wafflecap_8_8_0[8|24]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2022 VSS row_n[7] adc_array_wafflecap_8_8_0[6|26]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2023 adc_array_wafflecap_8_8_1[18]/adc_array_circuit_150n_0/vdrv row_n[0] adc_array_wafflecap_8_8_1[18]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2024 adc_array_wafflecap_8_8_0[1|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2025 vcm adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|1]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2026 adc_array_wafflecap_8_8_0[8|16]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|16]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2027 vcm adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|15]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2028 VDD rowon_n[12] adc_array_wafflecap_8_8_0[11|19]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2029 adc_array_wafflecap_8_8_0[9|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2030 adc_array_wafflecap_8_8_0[8|6]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|6]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2031 adc_array_wafflecap_8_Dummy_4[30]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[30]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2032 vcm adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|5]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2033 vcm adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|26]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2034 VDD rowon_n[11] adc_array_wafflecap_8_8_0[10|23]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2035 adc_array_wafflecap_8_8_0[7|20]/adc_array_circuit_150n_0/vint1 col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2036 vcm adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|4]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2037 VDD rowon_n[10] adc_array_wafflecap_8_8_0[9|4]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2038 VDD rowon_n[10] adc_array_wafflecap_8_8_0[9|14]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2039 adc_array_wafflecap_8_8_0[1|6]/adc_array_circuit_150n_0/vint2 col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2040 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X2041 adc_array_wafflecap_8_8_0[13|22]/adc_array_circuit_150n_0/vint2 col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2042 VSS row_n[12] adc_array_wafflecap_8_8_0[11|26]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2043 adc_array_wafflecap_8_8_0[6|26]/adc_array_circuit_150n_0/vint1 col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2044 adc_array_wafflecap_8_8_0[2|27]/adc_array_circuit_150n_0/vint1 col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2045 adc_array_wafflecap_8_8_0[2|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2046 adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2047 adc_array_wafflecap_8_8_0[3|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2048 VSS row_n[13] adc_array_wafflecap_8_8_0[12|12]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2049 adc_array_wafflecap_8_8_0[9|9]/adc_array_circuit_150n_0/vint2 col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2050 VSS row_n[13] adc_array_wafflecap_8_8_0[12|2]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2051 adc_array_wafflecap_8_Dummy_4[22]/adc_array_circuit_150n_0/vint1 col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2052 adc_array_wafflecap_8_8_0[9|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2053 adc_array_wafflecap_8_8_0[8|13]/adc_array_circuit_150n_0/vint2 col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2054 adc_array_wafflecap_8_8_0[1|6]/adc_array_circuit_150n_0/vdrv row_n[2] adc_array_wafflecap_8_8_0[1|6]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2055 adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/vdrv row_n[12] adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2056 adc_array_wafflecap_8_8_0[8|3]/adc_array_circuit_150n_0/vint2 col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2057 adc_array_wafflecap_8_8_0[3|22]/adc_array_circuit_150n_0/vint2 rowon_n[4] adc_array_wafflecap_8_8_0[3|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2058 adc_array_wafflecap_8_8_0[11|8]/adc_array_circuit_150n_0/vint1 col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2059 adc_array_wafflecap_8_8_0[3|10]/adc_array_circuit_150n_0/vint2 col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2060 adc_array_wafflecap_8_Dummy_4[21]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2061 adc_array_wafflecap_8_8_0[0|23]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|23]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2062 vcm adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|30]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2063 vcm adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|21]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2064 adc_array_wafflecap_8_8_0[10|12]/adc_array_circuit_150n_0/vint1 col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2065 adc_array_wafflecap_8_8_0[7|9]/adc_array_circuit_150n_0/vdrv row_n[8] adc_array_wafflecap_8_8_0[7|9]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2066 adc_array_wafflecap_8_8_0[4|22]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|22]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2067 adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/vint1 col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2068 adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2069 adc_array_wafflecap_8_8_0[3|0]/adc_array_circuit_150n_0/vdrv row_n[4] adc_array_wafflecap_8_8_0[3|0]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2070 adc_array_wafflecap_8_8_0[3|1]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|1]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2071 adc_array_wafflecap_8_Dummy_8[2]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_8[2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2072 adc_array_wafflecap_8_8_0[10|2]/adc_array_circuit_150n_0/vint1 col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2073 adc_array_wafflecap_8_8_0[1|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2074 adc_array_wafflecap_8_8_0[6|13]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|13]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2075 adc_array_wafflecap_8_8_1[28]/adc_array_circuit_150n_0/vint1 col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2076 adc_array_wafflecap_8_8_0[4|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2077 vcm adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|18]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2078 adc_array_wafflecap_8_Dummy_8[1]/adc_array_circuit_150n_0/vint2 col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2079 vcm adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|19]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2080 adc_array_wafflecap_8_8_0[2|2]/adc_array_circuit_150n_0/vint2 col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2081 adc_array_wafflecap_8_8_0[1|15]/adc_array_circuit_150n_0/vint2 col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2082 adc_array_wafflecap_8_Dummy_4[11]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[11]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2083 adc_array_wafflecap_8_8_0[7|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2084 adc_array_wafflecap_8_8_0[7|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2085 adc_array_wafflecap_8_Dummy_4[1]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[1]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2086 adc_array_wafflecap_8_8_0[14|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2087 adc_array_wafflecap_8_8_0[13|21]/adc_array_circuit_150n_0/vint2 rowon_n[14] adc_array_wafflecap_8_8_0[13|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2088 vcm adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|0]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2089 vcm adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|10]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2090 adc_array_wafflecap_8_8_0[1|26]/adc_array_circuit_150n_0/vint2 rowon_n[2] adc_array_wafflecap_8_8_0[1|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2091 adc_array_wafflecap_8_8_0[1|6]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|6]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2092 adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2093 adc_array_wafflecap_8_8_0[12|2]/adc_array_circuit_150n_0/vint2 rowon_n[13] adc_array_wafflecap_8_8_0[12|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2094 adc_array_wafflecap_8_8_0[12|12]/adc_array_circuit_150n_0/vint2 rowon_n[13] adc_array_wafflecap_8_8_0[12|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2095 adc_array_wafflecap_8_8_0[5|5]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|5]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2096 vcm VSS adc_array_wafflecap_8_Dummy_4[0]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2097 vcm VSS adc_array_wafflecap_8_Dummy_4[10]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2098 adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2099 adc_array_wafflecap_8_8_0[11|16]/adc_array_circuit_150n_0/vint2 rowon_n[12] adc_array_wafflecap_8_8_0[11|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2100 adc_array_wafflecap_8_8_0[10|28]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|28]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2101 adc_array_wafflecap_8_Dummy_3[2]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_3[2]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2102 adc_array_wafflecap_8_8_0[11|6]/adc_array_circuit_150n_0/vint2 rowon_n[12] adc_array_wafflecap_8_8_0[11|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2103 adc_array_wafflecap_8_Dummy_1[0]/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_1[0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2104 adc_array_wafflecap_8_8_0[0|2]/adc_array_circuit_150n_0/vdrv row_n[1] adc_array_wafflecap_8_8_0[0|2]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2105 adc_array_wafflecap_8_8_0[2|8]/adc_array_circuit_150n_0/vint2 rowon_n[3] adc_array_wafflecap_8_8_0[2|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2106 adc_array_wafflecap_8_8_0[9|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2107 adc_array_wafflecap_8_8_0[2|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2108 adc_array_wafflecap_8_8_0[5|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2109 adc_array_wafflecap_8_8_0[1|15]/adc_array_circuit_150n_0/vdrv row_n[2] adc_array_wafflecap_8_8_0[1|15]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2110 VDD rowon_n[11] adc_array_wafflecap_8_8_0[10|12]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2111 VDD rowon_n[6] adc_array_wafflecap_8_8_0[5|10]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2112 VDD rowon_n[11] adc_array_wafflecap_8_8_0[10|2]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2113 VDD rowon_n[2] adc_array_wafflecap_8_8_0[1|26]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2114 adc_array_wafflecap_8_8_0[14|29]/adc_array_circuit_150n_0/vint2 col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2115 adc_array_wafflecap_8_8_0[3|7]/adc_array_circuit_150n_0/vint1 col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2116 VSS row_n[8] adc_array_wafflecap_8_8_0[7|1]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2117 VSS row_n[8] adc_array_wafflecap_8_8_0[7|11]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2118 adc_array_wafflecap_8_8_0[3|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2119 adc_array_wafflecap_8_8_0[3|30]/adc_array_circuit_150n_0/vint2 rowon_n[4] adc_array_wafflecap_8_8_0[3|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2120 VDD rowon_n[1] adc_array_wafflecap_8_8_0[0|8]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2121 adc_array_wafflecap_8_8_0[2|24]/adc_array_circuit_150n_0/vint2 col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2122 VSS row_n[14] adc_array_wafflecap_8_8_0[13|10]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2123 adc_array_wafflecap_8_8_0[0|13]/adc_array_circuit_150n_0/vint2 rowon_n[1] adc_array_wafflecap_8_8_0[0|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2124 VSS row_n[14] adc_array_wafflecap_8_8_0[13|0]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2125 adc_array_wafflecap_8_Dummy_4[33]/adc_array_circuit_150n_0/vint1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2126 adc_array_wafflecap_8_8_0[12|29]/adc_array_circuit_150n_0/vdrv row_n[13] adc_array_wafflecap_8_8_0[12|29]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2127 adc_array_wafflecap_8_8_0[10|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2128 adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2129 VSS VSS adc_array_wafflecap_8_Dummy_1[1]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2130 VSS row_n[3] adc_array_wafflecap_8_8_0[2|9]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2131 VDD rowon_n[4] adc_array_wafflecap_8_8_0[3|15]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2132 adc_array_wafflecap_8_8_0[0|24]/adc_array_circuit_150n_0/vdrv row_n[1] adc_array_wafflecap_8_8_0[0|24]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2133 adc_array_wafflecap_8_8_1[21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2134 adc_array_wafflecap_8_8_0[0|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2135 adc_array_wafflecap_8_8_0[5|11]/adc_array_circuit_150n_0/vint1 col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2136 adc_array_wafflecap_8_8_0[2|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2137 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X2138 VDD rowon_n[0] adc_array_wafflecap_8_Dummy_7/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2139 adc_array_wafflecap_8_8_0[12|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2140 adc_array_wafflecap_8_8_0[5|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2141 VDD VSS adc_array_wafflecap_8_Dummy_1[4]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2142 adc_array_wafflecap_8_8_0[1|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2143 adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n sample VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2144 adc_array_wafflecap_8_8_1[4]/adc_array_circuit_150n_0/vint2 rowon_n[0] adc_array_wafflecap_8_8_1[4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2145 vcm adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[7]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2146 adc_array_wafflecap_8_8_0[0|9]/adc_array_circuit_150n_0/vint1 col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2147 VSS row_n[7] adc_array_wafflecap_8_8_0[6|20]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2148 adc_array_wafflecap_8_8_0[4|27]/adc_array_circuit_150n_0/vint2 col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2149 adc_array_wafflecap_8_8_1[17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_1[17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2150 adc_array_wafflecap_8_8_0[0|28]/adc_array_circuit_150n_0/vint2 col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2151 vcm adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|30]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2152 VSS row_n[1] adc_array_wafflecap_8_8_0[0|14]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2153 adc_array_wafflecap_8_8_0[14|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2154 adc_array_wafflecap_8_8_0[8|20]/adc_array_circuit_150n_0/vint2 rowon_n[9] adc_array_wafflecap_8_8_0[8|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2155 adc_array_wafflecap_8_8_0[6|18]/adc_array_circuit_150n_0/vint2 col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2156 adc_array_wafflecap_8_8_0[8|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2157 adc_array_wafflecap_8_8_0[7|1]/adc_array_circuit_150n_0/vint2 rowon_n[8] adc_array_wafflecap_8_8_0[7|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2158 adc_array_wafflecap_8_8_0[7|11]/adc_array_circuit_150n_0/vint2 rowon_n[8] adc_array_wafflecap_8_8_0[7|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2159 adc_array_wafflecap_8_8_0[3|30]/adc_array_circuit_150n_0/vdrv row_n[4] adc_array_wafflecap_8_8_0[3|30]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2160 adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2161 vcm adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|2]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2162 adc_array_wafflecap_8_8_0[13|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2163 vcm adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|8]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2164 adc_array_wafflecap_8_8_0[8|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2165 adc_array_wafflecap_8_8_0[4|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2166 adc_array_wafflecap_8_8_0[0|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2167 adc_array_wafflecap_8_8_0[13|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2168 adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/vint2 rowon_n[14] adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2169 adc_array_wafflecap_8_Dummy_3[3]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_3[3]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2170 adc_array_wafflecap_8_8_0[9|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2171 adc_array_wafflecap_8_8_1[0]/adc_array_circuit_150n_0/vint1 col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2172 adc_array_wafflecap_8_8_0[9|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2173 adc_array_wafflecap_8_8_0[6|20]/adc_array_circuit_150n_0/vint1 col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2174 adc_array_wafflecap_8_Dummy_1[5]/adc_array_circuit_150n_0/vint1 col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2175 adc_array_wafflecap_8_Dummy_4[16]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2176 adc_array_wafflecap_8_8_0[2|19]/adc_array_circuit_150n_0/vdrv row_n[3] adc_array_wafflecap_8_8_0[2|19]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2177 VSS sample adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2178 adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/vint2 VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2179 adc_array_wafflecap_8_Dummy_4[6]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2180 adc_array_wafflecap_8_8_0[6|18]/adc_array_circuit_150n_0/vdrv row_n[7] adc_array_wafflecap_8_8_0[6|18]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2181 VSS row_n[13] adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2182 adc_array_wafflecap_8_8_0[11|16]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|16]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2183 adc_array_wafflecap_8_8_0[9|28]/adc_array_circuit_150n_0/vint2 col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2184 adc_array_wafflecap_8_8_0[11|6]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|6]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2185 adc_array_wafflecap_8_Dummy_2[3]/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_2[3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2186 adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/vint2 VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2187 VSS row_n[9] adc_array_wafflecap_8_8_0[8|9]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2188 VDD rowon_n[15] adc_array_wafflecap_8_8_0[14|8]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2189 VDD rowon_n[15] adc_array_wafflecap_8_8_0[14|30]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2190 adc_array_wafflecap_8_8_0[11|27]/adc_array_circuit_150n_0/vint1 col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2191 adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/vdrv row_n[1] adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2192 vcm adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|23]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2193 adc_array_wafflecap_8_8_0[4|25]/adc_array_circuit_150n_0/vint1 col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2194 vcm adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|24]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2195 adc_array_wafflecap_8_8_0[1|17]/adc_array_circuit_150n_0/vint2 rowon_n[2] adc_array_wafflecap_8_8_0[1|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2196 adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/vint1 col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2197 adc_array_wafflecap_8_8_0[7|28]/adc_array_circuit_150n_0/vdrv row_n[8] adc_array_wafflecap_8_8_0[7|28]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2198 vcm adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|26]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2199 adc_array_wafflecap_8_8_0[10|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2200 adc_array_wafflecap_8_8_1[22]/adc_array_circuit_150n_0/vint1 col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2201 adc_array_wafflecap_8_8_0[1|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2202 adc_array_wafflecap_8_8_0[13|7]/adc_array_circuit_150n_0/vint2 col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2203 VDD rowon_n[2] adc_array_wafflecap_8_8_0[1|17]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2204 VSS row_n[0] adc_array_wafflecap_8_8_1[26]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2205 vcm adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|6]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2206 adc_array_wafflecap_8_8_0[5|19]/adc_array_circuit_150n_0/vint2 rowon_n[6] adc_array_wafflecap_8_8_0[5|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2207 adc_array_wafflecap_8_8_0[1|8]/adc_array_circuit_150n_0/vint2 col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2208 adc_array_wafflecap_8_Dummy_4[7]/adc_array_circuit_150n_0/vint1 col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2209 vcm VSS adc_array_wafflecap_8_Dummy_4[29]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2210 adc_array_wafflecap_8_8_0[11|16]/adc_array_circuit_150n_0/vdrv row_n[12] adc_array_wafflecap_8_8_0[11|16]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2211 adc_array_wafflecap_8_8_0[9|27]/adc_array_circuit_150n_0/vint2 rowon_n[10] adc_array_wafflecap_8_8_0[9|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2212 adc_array_wafflecap_8_8_0[5|7]/adc_array_circuit_150n_0/vint2 col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2213 VSS row_n[6] adc_array_wafflecap_8_8_0[5|17]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2214 VSS row_n[2] adc_array_wafflecap_8_8_0[1|18]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2215 vcm adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|27]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2216 adc_array_wafflecap_8_8_0[2|20]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|20]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2217 adc_array_wafflecap_8_8_0[2|29]/adc_array_circuit_150n_0/vint1 col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2218 adc_array_wafflecap_8_Dummy_2[4]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_2[4]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2219 adc_array_wafflecap_8_8_0[0|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2220 adc_array_wafflecap_8_8_0[12|20]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|20]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2221 adc_array_wafflecap_8_8_0[8|9]/adc_array_circuit_150n_0/vint2 rowon_n[9] adc_array_wafflecap_8_8_0[8|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2222 adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/vint2 rowon_n[9] adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2223 adc_array_wafflecap_8_8_0[7|24]/adc_array_circuit_150n_0/vint2 col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2224 adc_array_wafflecap_8_8_0[2|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2225 VDD sample_n adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2226 adc_array_wafflecap_8_8_0[14|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2227 vcm adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|19]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2228 adc_array_wafflecap_8_8_0[10|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2229 adc_array_wafflecap_8_8_0[10|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2230 adc_array_wafflecap_8_8_0[9|23]/adc_array_circuit_150n_0/vint1 col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2231 VDD rowon_n[8] adc_array_wafflecap_8_8_0[7|27]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2232 adc_array_wafflecap_8_8_0[0|0]/adc_array_circuit_150n_0/vint2 col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2233 adc_array_wafflecap_8_8_0[1|8]/adc_array_circuit_150n_0/vdrv row_n[2] adc_array_wafflecap_8_8_0[1|8]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2234 adc_array_wafflecap_8_8_0[3|24]/adc_array_circuit_150n_0/vint2 rowon_n[4] adc_array_wafflecap_8_8_0[3|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2235 adc_array_wafflecap_8_8_0[1|18]/adc_array_circuit_150n_0/vint1 col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2236 adc_array_wafflecap_8_8_0[3|12]/adc_array_circuit_150n_0/vint2 col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2237 adc_array_wafflecap_8_Dummy_4[26]/adc_array_circuit_150n_0/vint2 col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2238 VSS row_n[14] adc_array_wafflecap_8_8_0[13|29]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2239 adc_array_wafflecap_8_8_0[10|26]/adc_array_circuit_150n_0/vint2 col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2240 adc_array_wafflecap_8_Dummy_8[4]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_8[4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2241 adc_array_wafflecap_8_8_0[0|25]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|25]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2242 vcm adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2243 adc_array_wafflecap_8_8_0[3|2]/adc_array_circuit_150n_0/vdrv row_n[4] adc_array_wafflecap_8_8_0[3|2]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2244 adc_array_wafflecap_8_8_0[3|3]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|3]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2245 VSS row_n[15] adc_array_wafflecap_8_8_0[14|15]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2246 adc_array_wafflecap_8_8_0[6|15]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|15]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2247 VSS row_n[15] adc_array_wafflecap_8_8_0[14|5]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2248 adc_array_wafflecap_8_Dummy_0[1]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_0[1]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2249 adc_array_wafflecap_8_8_1[30]/adc_array_circuit_150n_0/vint1 col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2250 adc_array_wafflecap_8_Dummy_4[13]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[13]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2251 VDD VDD adc_array_wafflecap_8_Dummy_4[29]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2252 adc_array_wafflecap_8_8_0[14|21]/adc_array_circuit_150n_0/vdrv row_n[15] adc_array_wafflecap_8_8_0[14|21]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2253 adc_array_wafflecap_8_8_0[4|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2254 adc_array_wafflecap_8_8_0[0|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2255 adc_array_wafflecap_8_Dummy_4[3]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[3]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2256 adc_array_wafflecap_8_Dummy_8[3]/adc_array_circuit_150n_0/vint2 col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2257 adc_array_wafflecap_8_8_1[13]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[13]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2258 adc_array_wafflecap_8_8_0[13|25]/adc_array_circuit_150n_0/vdrv row_n[14] adc_array_wafflecap_8_8_0[13|25]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2259 adc_array_wafflecap_8_8_0[8|26]/adc_array_circuit_150n_0/vdrv row_n[9] adc_array_wafflecap_8_8_0[8|26]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2260 vcm adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|25]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2261 adc_array_wafflecap_8_8_0[6|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2262 VDD rowon_n[4] adc_array_wafflecap_8_8_0[3|8]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2263 vcm adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|24]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2264 adc_array_wafflecap_8_8_0[12|15]/adc_array_circuit_150n_0/vint1 col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2265 adc_array_wafflecap_8_8_0[12|5]/adc_array_circuit_150n_0/vint1 col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2266 adc_array_wafflecap_8_8_0[11|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2267 adc_array_wafflecap_8_8_0[4|21]/adc_array_circuit_150n_0/vint2 col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2268 adc_array_wafflecap_8_8_0[1|28]/adc_array_circuit_150n_0/vint2 rowon_n[2] adc_array_wafflecap_8_8_0[1|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2269 adc_array_wafflecap_8_Dummy_1[2]/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_1[2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2270 adc_array_wafflecap_8_8_0[13|18]/adc_array_circuit_150n_0/vint2 col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2271 adc_array_wafflecap_8_8_0[3|24]/adc_array_circuit_150n_0/vdrv row_n[4] adc_array_wafflecap_8_8_0[3|24]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2272 adc_array_wafflecap_8_8_0[2|10]/adc_array_circuit_150n_0/vint2 rowon_n[3] adc_array_wafflecap_8_8_0[2|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2273 adc_array_wafflecap_8_8_0[9|25]/adc_array_circuit_150n_0/vint2 rowon_n[10] adc_array_wafflecap_8_8_0[9|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2274 adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2275 adc_array_wafflecap_8_8_0[5|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2276 vcm adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|27]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2277 VSS row_n[5] adc_array_wafflecap_8_8_0[4|6]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2278 VDD rowon_n[3] adc_array_wafflecap_8_8_0[2|0]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2279 VSS row_n[1] adc_array_wafflecap_8_8_0[0|7]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2280 VSS sample adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2281 adc_array_wafflecap_8_Dummy_3[2]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_3[2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2282 VDD rowon_n[2] adc_array_wafflecap_8_8_0[1|28]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2283 adc_array_wafflecap_8_Dummy_4[18]/adc_array_circuit_150n_0/vint1 col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2284 adc_array_wafflecap_8_Dummy_4[25]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2285 adc_array_wafflecap_8_8_0[14|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2286 adc_array_wafflecap_8_8_0[14|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2287 adc_array_wafflecap_8_8_0[9|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2288 VSS row_n[12] adc_array_wafflecap_8_8_0[11|25]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2289 adc_array_wafflecap_8_8_0[3|9]/adc_array_circuit_150n_0/vint1 col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2290 adc_array_wafflecap_8_8_0[3|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2291 VDD rowon_n[1] adc_array_wafflecap_8_8_0[0|10]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2292 adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2293 adc_array_wafflecap_8_8_0[5|4]/adc_array_circuit_150n_0/vint2 col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2294 VDD rowon_n[8] adc_array_wafflecap_8_8_0[7|25]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2295 adc_array_wafflecap_8_Dummy_8[5]/adc_array_circuit_150n_0/vint1 col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2296 adc_array_wafflecap_8_8_0[12|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2297 adc_array_wafflecap_8_Dummy_3[1]/adc_array_circuit_150n_0/vint2 col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2298 adc_array_wafflecap_8_8_0[0|15]/adc_array_circuit_150n_0/vint2 rowon_n[1] adc_array_wafflecap_8_8_0[0|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2299 VDD rowon_n[14] adc_array_wafflecap_8_8_0[13|24]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2300 adc_array_wafflecap_8_8_0[11|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2301 adc_array_wafflecap_8_8_0[11|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2302 VSS VSS adc_array_wafflecap_8_Dummy_1[3]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2303 VSS row_n[3] adc_array_wafflecap_8_8_0[2|11]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2304 adc_array_wafflecap_8_8_1[23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2305 adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2306 adc_array_wafflecap_8_8_0[5|27]/adc_array_circuit_150n_0/vdrv row_n[6] adc_array_wafflecap_8_8_0[5|27]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2307 adc_array_wafflecap_8_8_0[5|28]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|28]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2308 adc_array_wafflecap_8_8_0[2|1]/adc_array_circuit_150n_0/vint1 col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2309 adc_array_wafflecap_8_8_0[2|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2310 adc_array_wafflecap_8_Dummy_8[1]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2311 adc_array_wafflecap_8_8_0[1|29]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|29]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2312 VSS row_n[10] adc_array_wafflecap_8_8_0[9|4]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2313 VSS row_n[10] adc_array_wafflecap_8_8_0[9|14]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2314 VDD VSS adc_array_wafflecap_8_Dummy_1[6]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2315 adc_array_wafflecap_8_8_0[1|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2316 adc_array_wafflecap_8_8_0[9|20]/adc_array_circuit_150n_0/vdrv row_n[10] adc_array_wafflecap_8_8_0[9|20]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2317 adc_array_wafflecap_8_8_0[5|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2318 VSS VDD adc_array_wafflecap_8_Dummy_4[14]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2319 VSS VDD adc_array_wafflecap_8_Dummy_4[4]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2320 adc_array_wafflecap_8_8_0[7|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2321 vcm adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[9]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2322 adc_array_wafflecap_8_8_0[0|30]/adc_array_circuit_150n_0/vint2 col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2323 adc_array_wafflecap_8_8_0[0|11]/adc_array_circuit_150n_0/vint1 col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2324 adc_array_wafflecap_8_8_0[12|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2325 adc_array_wafflecap_8_8_0[11|4]/adc_array_circuit_150n_0/vint2 col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2326 adc_array_wafflecap_8_8_0[11|14]/adc_array_circuit_150n_0/vint2 col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2327 VSS row_n[7] adc_array_wafflecap_8_8_0[6|22]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2328 adc_array_wafflecap_8_8_0[4|16]/adc_array_circuit_150n_0/vdrv row_n[5] adc_array_wafflecap_8_8_0[4|16]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2329 VDD VDD adc_array_wafflecap_8_Dummy_4[18]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2330 adc_array_wafflecap_8_8_0[7|14]/adc_array_circuit_150n_0/vint1 col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2331 adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/vint2 rowon_n[7] adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2332 adc_array_wafflecap_8_8_0[11|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2333 vcm adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|23]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2334 adc_array_wafflecap_8_8_0[7|4]/adc_array_circuit_150n_0/vint1 col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2335 adc_array_wafflecap_8_8_0[4|2]/adc_array_circuit_150n_0/vint2 rowon_n[5] adc_array_wafflecap_8_8_0[4|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2336 adc_array_wafflecap_8_8_0[14|12]/adc_array_circuit_150n_0/vint2 col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2337 VSS row_n[13] adc_array_wafflecap_8_8_0[12|16]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2338 adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/vdrv row_n[4] adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2339 adc_array_wafflecap_8_8_0[14|2]/adc_array_circuit_150n_0/vint2 col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2340 adc_array_wafflecap_8_8_0[13|3]/adc_array_circuit_150n_0/vint1 col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2341 adc_array_wafflecap_8_8_0[13|13]/adc_array_circuit_150n_0/vint1 col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2342 adc_array_wafflecap_8_8_0[7|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2343 adc_array_wafflecap_8_8_0[7|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2344 adc_array_wafflecap_8_8_0[4|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2345 adc_array_wafflecap_8_8_0[8|17]/adc_array_circuit_150n_0/vint2 col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2346 adc_array_wafflecap_8_Dummy_3[5]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_3[5]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2347 adc_array_wafflecap_8_8_1[18]/adc_array_circuit_150n_0/vint2 col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2348 vcm adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|21]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2349 adc_array_wafflecap_8_8_0[2|23]/adc_array_circuit_150n_0/vint1 col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2350 VSS sample_n adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2351 adc_array_wafflecap_8_8_0[6|22]/adc_array_circuit_150n_0/vint1 col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2352 VDD rowon_n[7] adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2353 adc_array_wafflecap_8_8_0[12|2]/adc_array_circuit_150n_0/vdrv row_n[13] adc_array_wafflecap_8_8_0[12|2]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2354 adc_array_wafflecap_8_8_0[12|12]/adc_array_circuit_150n_0/vdrv row_n[13] adc_array_wafflecap_8_8_0[12|12]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2355 adc_array_wafflecap_8_8_0[10|16]/adc_array_circuit_150n_0/vint1 col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2356 adc_array_wafflecap_8_8_0[10|23]/adc_array_circuit_150n_0/vint2 rowon_n[11] adc_array_wafflecap_8_8_0[10|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2357 VSS row_n[8] adc_array_wafflecap_8_8_0[7|20]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2358 adc_array_wafflecap_8_8_0[9|14]/adc_array_circuit_150n_0/vint2 rowon_n[10] adc_array_wafflecap_8_8_0[9|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2359 adc_array_wafflecap_8_Dummy_4[15]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2360 vcm adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|11]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2361 adc_array_wafflecap_8_8_0[9|4]/adc_array_circuit_150n_0/vint2 rowon_n[10] adc_array_wafflecap_8_8_0[9|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2362 adc_array_wafflecap_8_Dummy_4[5]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2363 vcm adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|1]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2364 vcm adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|15]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2365 VDD rowon_n[10] adc_array_wafflecap_8_8_0[9|19]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2366 VSS row_n[5] adc_array_wafflecap_8_8_0[4|3]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2367 adc_array_wafflecap_8_8_0[13|29]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|29]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2368 vcm adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|5]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2369 vcm adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|25]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2370 vcm adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|26]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2371 VDD rowon_n[9] adc_array_wafflecap_8_8_0[8|23]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2372 VSS VDD adc_array_wafflecap_8_Dummy_4[22]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2373 VDD rowon_n[8] adc_array_wafflecap_8_8_0[7|4]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2374 VDD rowon_n[8] adc_array_wafflecap_8_8_0[7|14]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2375 adc_array_wafflecap_8_8_1[24]/adc_array_circuit_150n_0/vint1 col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2376 adc_array_wafflecap_8_8_0[11|22]/adc_array_circuit_150n_0/vint2 col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2377 adc_array_wafflecap_8_8_0[4|26]/adc_array_circuit_150n_0/vint1 col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2378 adc_array_wafflecap_8_8_0[4|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2379 adc_array_wafflecap_8_Dummy_0[0]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_0[0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2380 adc_array_wafflecap_8_8_0[0|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2381 adc_array_wafflecap_8_8_0[1|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2382 VSS row_n[11] adc_array_wafflecap_8_8_0[10|12]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2383 adc_array_wafflecap_8_8_0[7|9]/adc_array_circuit_150n_0/vint2 col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2384 adc_array_wafflecap_8_8_0[6|8]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|8]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2385 adc_array_wafflecap_8_8_0[6|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2386 vcm adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|14]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2387 VSS row_n[11] adc_array_wafflecap_8_8_0[10|2]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2388 adc_array_wafflecap_8_8_0[13|21]/adc_array_circuit_150n_0/vint1 col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2389 adc_array_wafflecap_8_8_0[7|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2390 VDD VDD adc_array_wafflecap_8_Dummy_4[16]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2391 adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/vdrv row_n[10] adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2392 adc_array_wafflecap_8_8_0[5|21]/adc_array_circuit_150n_0/vint2 rowon_n[6] adc_array_wafflecap_8_8_0[5|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2393 VSS row_n[0] adc_array_wafflecap_8_8_1[28]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2394 adc_array_wafflecap_8_8_0[1|22]/adc_array_circuit_150n_0/vint2 rowon_n[2] adc_array_wafflecap_8_8_0[1|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2395 VDD VDD adc_array_wafflecap_8_Dummy_4[6]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2396 adc_array_wafflecap_8_8_0[13|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2397 adc_array_wafflecap_8_8_0[9|8]/adc_array_circuit_150n_0/vint1 col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2398 adc_array_wafflecap_8_8_0[1|10]/adc_array_circuit_150n_0/vint2 col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2399 adc_array_wafflecap_8_Dummy_2[6]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_2[6]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2400 adc_array_wafflecap_8_8_0[9|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2401 adc_array_wafflecap_8_8_0[8|12]/adc_array_circuit_150n_0/vint1 col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2402 adc_array_wafflecap_8_8_0[2|22]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|22]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2403 adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/vint1 col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2404 adc_array_wafflecap_8_8_0[1|1]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|1]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2405 adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2406 adc_array_wafflecap_8_8_0[8|2]/adc_array_circuit_150n_0/vint1 col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2407 adc_array_wafflecap_8_8_0[5|0]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|0]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2408 adc_array_wafflecap_8_Dummy_4[1]/adc_array_circuit_150n_0/vint2 col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2409 adc_array_wafflecap_8_Dummy_4[11]/adc_array_circuit_150n_0/vint2 col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2410 adc_array_wafflecap_8_8_0[7|20]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|20]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2411 adc_array_wafflecap_8_8_0[2|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2412 VDD rowon_n[2] adc_array_wafflecap_8_8_0[1|22]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2413 vcm VSS adc_array_wafflecap_8_Dummy_2[2]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2414 adc_array_wafflecap_8_8_0[0|2]/adc_array_circuit_150n_0/vint2 col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2415 adc_array_wafflecap_8_8_0[1|10]/adc_array_circuit_150n_0/vdrv row_n[2] adc_array_wafflecap_8_8_0[1|10]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2416 vcm adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|18]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2417 adc_array_wafflecap_8_8_0[14|6]/adc_array_circuit_150n_0/vdrv row_n[15] adc_array_wafflecap_8_8_0[14|6]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2418 adc_array_wafflecap_8_8_0[13|10]/adc_array_circuit_150n_0/vdrv row_n[14] adc_array_wafflecap_8_8_0[13|10]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2419 adc_array_wafflecap_8_8_0[11|21]/adc_array_circuit_150n_0/vint2 rowon_n[12] adc_array_wafflecap_8_8_0[11|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2420 vcm adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|10]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2421 adc_array_wafflecap_8_8_0[14|23]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|23]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2422 adc_array_wafflecap_8_8_0[13|0]/adc_array_circuit_150n_0/vdrv row_n[14] adc_array_wafflecap_8_8_0[13|0]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2423 adc_array_wafflecap_8_8_0[12|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2424 vcm adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|0]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2425 adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2426 adc_array_wafflecap_8_8_0[10|2]/adc_array_circuit_150n_0/vint2 rowon_n[11] adc_array_wafflecap_8_8_0[10|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2427 adc_array_wafflecap_8_8_0[10|12]/adc_array_circuit_150n_0/vint2 rowon_n[11] adc_array_wafflecap_8_8_0[10|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2428 adc_array_wafflecap_8_8_0[3|5]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|5]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2429 VSS sample_n adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2430 vcm adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|9]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2431 adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2432 adc_array_wafflecap_8_Dummy_8[0]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_8[0]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2433 adc_array_wafflecap_8_8_0[0|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2434 adc_array_wafflecap_8_8_0[0|8]/adc_array_circuit_150n_0/vint2 rowon_n[1] adc_array_wafflecap_8_8_0[0|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2435 adc_array_wafflecap_8_8_0[9|4]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|4]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2436 adc_array_wafflecap_8_8_0[9|14]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|14]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2437 vcm adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|29]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2438 adc_array_wafflecap_8_8_0[5|21]/adc_array_circuit_150n_0/vdrv row_n[6] adc_array_wafflecap_8_8_0[5|21]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2439 adc_array_wafflecap_8_8_0[4|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2440 ctop sw analog_in VSS sky130_fd_pr__nfet_01v8 ad=1.45e+11p pd=1.58e+06u as=2.9e+11p ps=3.16e+06u w=500000u l=500000u
X2441 adc_array_wafflecap_8_8_0[3|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2442 adc_array_wafflecap_8_8_1[15]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[15]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2443 VDD rowon_n[9] adc_array_wafflecap_8_8_0[8|12]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2444 adc_array_wafflecap_8_8_0[6|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2445 VDD rowon_n[4] adc_array_wafflecap_8_8_0[3|10]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2446 VDD rowon_n[9] adc_array_wafflecap_8_8_0[8|2]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2447 VSS VDD adc_array_wafflecap_8_Dummy_4[33]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2448 adc_array_wafflecap_8_8_0[12|29]/adc_array_circuit_150n_0/vint2 col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2449 adc_array_wafflecap_8_8_0[5|6]/adc_array_circuit_150n_0/vint1 col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2450 adc_array_wafflecap_8_8_0[1|30]/adc_array_circuit_150n_0/vint2 rowon_n[2] adc_array_wafflecap_8_8_0[1|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2451 adc_array_wafflecap_8_8_0[5|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2452 adc_array_wafflecap_8_8_0[4|23]/adc_array_circuit_150n_0/vint2 col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2453 VDD en_n_bit[2] adc_array_wafflecap_8_4_0/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2454 adc_array_wafflecap_8_8_0[0|24]/adc_array_circuit_150n_0/vint2 col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2455 adc_array_wafflecap_8_8_0[1|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2456 VDD rowon_n[12] adc_array_wafflecap_8_8_0[11|0]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2457 VDD rowon_n[12] adc_array_wafflecap_8_8_0[11|10]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2458 adc_array_wafflecap_8_Dummy_7/adc_array_circuit_150n_0/vint2 rowon_n[0] adc_array_wafflecap_8_Dummy_7/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2459 VSS row_n[12] adc_array_wafflecap_8_8_0[11|0]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2460 VSS row_n[12] adc_array_wafflecap_8_8_0[11|10]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2461 adc_array_wafflecap_8_8_0[6|14]/adc_array_circuit_150n_0/vint2 col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2462 adc_array_wafflecap_8_Dummy_1[4]/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_1[4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2463 adc_array_wafflecap_8_8_0[14|28]/adc_array_circuit_150n_0/vint1 col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2464 adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/vint1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2465 adc_array_wafflecap_8_8_0[10|29]/adc_array_circuit_150n_0/vdrv row_n[11] adc_array_wafflecap_8_8_0[10|29]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2466 adc_array_wafflecap_8_8_0[8|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2467 adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2468 VSS row_n[1] adc_array_wafflecap_8_8_0[0|9]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2469 adc_array_wafflecap_8_1_0/adc_array_circuit_150n_0/vdrv en_n_bit[0] adc_array_wafflecap_8_1_0/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2470 adc_array_wafflecap_8_Dummy_3[4]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_3[4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2471 VDD rowon_n[2] adc_array_wafflecap_8_8_0[1|30]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2472 adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2473 adc_array_wafflecap_8_8_0[3|11]/adc_array_circuit_150n_0/vint1 col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2474 adc_array_wafflecap_8_8_0[0|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2475 adc_array_wafflecap_8_8_0[10|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2476 adc_array_wafflecap_8_8_0[3|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2477 adc_array_wafflecap_8_8_0[6|14]/adc_array_circuit_150n_0/vdrv row_n[7] adc_array_wafflecap_8_8_0[6|14]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2478 adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n sample VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2479 adc_array_wafflecap_8_Dummy_1[0]/adc_array_circuit_150n_0/vint1 col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2480 adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2481 adc_array_wafflecap_8_Dummy_3[3]/adc_array_circuit_150n_0/vint2 col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2482 VSS row_n[0] adc_array_wafflecap_8_8_1[0]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2483 adc_array_wafflecap_8_8_0[2|27]/adc_array_circuit_150n_0/vint2 col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2484 vcm adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|30]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2485 VSS VSS adc_array_wafflecap_8_Dummy_1[5]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2486 adc_array_wafflecap_8_8_0[12|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2487 adc_array_wafflecap_8_8_0[9|22]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|22]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2488 adc_array_wafflecap_8_8_0[7|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2489 adc_array_wafflecap_8_8_1[25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2490 adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2491 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.64e+07u l=1.6e+07u
X2492 adc_array_wafflecap_8_Dummy_4[22]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[22]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2493 adc_array_wafflecap_8_8_0[11|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2494 vcm adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|8]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2495 adc_array_wafflecap_8_8_0[5|30]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|30]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2496 adc_array_wafflecap_8_8_0[5|12]/adc_array_circuit_150n_0/vint2 rowon_n[6] adc_array_wafflecap_8_8_0[5|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2497 adc_array_wafflecap_8_8_0[2|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2498 adc_array_wafflecap_8_Dummy_8[3]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2499 adc_array_wafflecap_8_8_0[11|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2500 adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/vint2 rowon_n[12] adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2501 adc_array_wafflecap_8_8_0[5|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2502 VDD rowon_n[6] adc_array_wafflecap_8_8_0[5|2]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2503 adc_array_wafflecap_8_8_0[0|27]/adc_array_circuit_150n_0/vdrv row_n[1] adc_array_wafflecap_8_8_0[0|27]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2504 adc_array_wafflecap_8_8_0[4|20]/adc_array_circuit_150n_0/vint1 col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2505 adc_array_wafflecap_8_8_0[14|8]/adc_array_circuit_150n_0/vint2 rowon_n[15] adc_array_wafflecap_8_8_0[14|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2506 adc_array_wafflecap_8_8_0[14|30]/adc_array_circuit_150n_0/vint2 rowon_n[15] adc_array_wafflecap_8_8_0[14|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2507 adc_array_wafflecap_8_8_0[13|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2508 adc_array_wafflecap_8_8_0[5|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2509 vcm adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[11]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2510 VSS sample adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2511 adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/vint2 VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2512 adc_array_wafflecap_8_8_0[13|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2513 VSS row_n[7] adc_array_wafflecap_8_8_0[6|24]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2514 adc_array_wafflecap_8_8_0[4|18]/adc_array_circuit_150n_0/vdrv row_n[5] adc_array_wafflecap_8_8_0[4|18]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2515 adc_array_wafflecap_8_8_0[4|19]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|19]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2516 VSS row_n[11] adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2517 adc_array_wafflecap_8_8_0[7|28]/adc_array_circuit_150n_0/vint2 col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2518 adc_array_wafflecap_8_8_0[4|4]/adc_array_circuit_150n_0/vint2 rowon_n[5] adc_array_wafflecap_8_8_0[4|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2519 adc_array_wafflecap_8_8_1[15]/adc_array_circuit_150n_0/vdrv row_n[0] adc_array_wafflecap_8_8_1[15]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2520 VSS row_n[0] adc_array_wafflecap_8_8_1[22]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2521 VDD rowon_n[13] adc_array_wafflecap_8_8_0[12|8]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2522 VDD rowon_n[13] adc_array_wafflecap_8_8_0[12|30]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2523 adc_array_wafflecap_8_8_0[11|23]/adc_array_circuit_150n_0/vdrv row_n[12] adc_array_wafflecap_8_8_0[11|23]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2524 adc_array_wafflecap_8_8_0[9|27]/adc_array_circuit_150n_0/vint1 col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2525 VSS row_n[6] adc_array_wafflecap_8_8_0[5|13]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2526 adc_array_wafflecap_8_Dummy_6/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_6/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2527 adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/vint1 col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2528 adc_array_wafflecap_8_8_0[6|24]/adc_array_circuit_150n_0/vint1 col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2529 vcm adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|23]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2530 adc_array_wafflecap_8_8_0[2|25]/adc_array_circuit_150n_0/vint1 col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2531 adc_array_wafflecap_8_8_0[14|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2532 vcm adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|1]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2533 adc_array_wafflecap_8_8_0[5|3]/adc_array_circuit_150n_0/vint1 col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2534 vcm adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|26]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2535 adc_array_wafflecap_8_8_0[8|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2536 VSS VDD adc_array_wafflecap_8_Dummy_4[7]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2537 adc_array_wafflecap_8_8_0[11|7]/adc_array_circuit_150n_0/vint2 col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2538 VSS row_n[5] adc_array_wafflecap_8_8_0[4|5]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2539 adc_array_wafflecap_8_8_0[3|19]/adc_array_circuit_150n_0/vint2 rowon_n[4] adc_array_wafflecap_8_8_0[3|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2540 adc_array_wafflecap_8_8_0[14|15]/adc_array_circuit_150n_0/vdrv row_n[15] adc_array_wafflecap_8_8_0[14|15]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2541 adc_array_wafflecap_8_8_0[14|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2542 adc_array_wafflecap_8_8_0[13|6]/adc_array_circuit_150n_0/vint1 col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2543 vcm adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|28]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2544 adc_array_wafflecap_8_8_0[9|16]/adc_array_circuit_150n_0/vdrv row_n[10] adc_array_wafflecap_8_8_0[9|16]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2545 VSS row_n[10] adc_array_wafflecap_8_8_0[9|23]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2546 adc_array_wafflecap_8_8_0[8|29]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|29]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2547 adc_array_wafflecap_8_8_0[7|27]/adc_array_circuit_150n_0/vint2 rowon_n[8] adc_array_wafflecap_8_8_0[7|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2548 adc_array_wafflecap_8_8_0[3|7]/adc_array_circuit_150n_0/vint2 col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2549 VSS row_n[4] adc_array_wafflecap_8_8_0[3|17]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2550 adc_array_wafflecap_8_8_0[14|5]/adc_array_circuit_150n_0/vdrv row_n[15] adc_array_wafflecap_8_8_0[14|5]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2551 adc_array_wafflecap_8_1_1/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_1_1/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2552 adc_array_wafflecap_8_8_0[0|20]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|20]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2553 vcm adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|27]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2554 vcm adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|14]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2555 adc_array_wafflecap_8_8_0[10|20]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|20]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2556 adc_array_wafflecap_8_8_0[4|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2557 adc_array_wafflecap_8_8_0[0|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2558 vcm adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|4]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2559 adc_array_wafflecap_8_8_0[12|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2560 adc_array_wafflecap_8_8_0[6|10]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|10]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2561 VDD rowon_n[12] adc_array_wafflecap_8_8_0[11|22]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2562 adc_array_wafflecap_8_8_0[9|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2563 vcm adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|19]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2564 vcm adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|16]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2565 adc_array_wafflecap_8_8_1[25]/adc_array_circuit_150n_0/vint1 col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2566 adc_array_wafflecap_8_8_0[9|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2567 adc_array_wafflecap_8_8_0[7|23]/adc_array_circuit_150n_0/vint1 col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2568 VSS row_n[0] adc_array_wafflecap_8_8_1[30]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2569 adc_array_wafflecap_8_Dummy_0[1]/adc_array_circuit_150n_0/vint2 col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2570 adc_array_wafflecap_8_8_1[8]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[8]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2571 adc_array_wafflecap_8_8_0[14|21]/adc_array_circuit_150n_0/vint2 col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2572 adc_array_wafflecap_8_8_0[6|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2573 adc_array_wafflecap_8_8_0[5|23]/adc_array_circuit_150n_0/vint2 rowon_n[6] adc_array_wafflecap_8_8_0[5|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2574 adc_array_wafflecap_8_8_0[1|24]/adc_array_circuit_150n_0/vint2 rowon_n[2] adc_array_wafflecap_8_8_0[1|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2575 adc_array_wafflecap_8_Dummy_4[29]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2576 adc_array_wafflecap_8_8_0[1|12]/adc_array_circuit_150n_0/vint2 col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2577 adc_array_wafflecap_8_8_0[13|25]/adc_array_circuit_150n_0/vint2 col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2578 VSS row_n[12] adc_array_wafflecap_8_8_0[11|29]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2579 adc_array_wafflecap_8_8_0[8|26]/adc_array_circuit_150n_0/vint2 col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2580 adc_array_wafflecap_8_Dummy_3[0]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_3[0]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2581 adc_array_wafflecap_8_8_0[5|2]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|2]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2582 adc_array_wafflecap_8_8_0[1|3]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|3]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2583 adc_array_wafflecap_8_8_0[14|8]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|8]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2584 VSS row_n[13] adc_array_wafflecap_8_8_0[12|15]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2585 VSS row_n[13] adc_array_wafflecap_8_8_0[12|5]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2586 adc_array_wafflecap_8_Dummy_4[25]/adc_array_circuit_150n_0/vint1 col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2587 adc_array_wafflecap_8_8_0[13|12]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|12]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2588 VDD rowon_n[14] adc_array_wafflecap_8_8_0[13|28]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2589 adc_array_wafflecap_8_8_0[12|21]/adc_array_circuit_150n_0/vdrv row_n[13] adc_array_wafflecap_8_8_0[12|21]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2590 adc_array_wafflecap_8_8_0[9|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2591 adc_array_wafflecap_8_Dummy_2[6]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_2[6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2592 VDD rowon_n[2] adc_array_wafflecap_8_8_0[1|24]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2593 adc_array_wafflecap_8_8_0[2|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2594 adc_array_wafflecap_8_8_0[13|2]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|2]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2595 adc_array_wafflecap_8_8_0[5|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2596 adc_array_wafflecap_8_8_0[1|12]/adc_array_circuit_150n_0/vdrv row_n[2] adc_array_wafflecap_8_8_0[1|12]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2597 adc_array_wafflecap_8_Dummy_4[24]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2598 vcm adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|24]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2599 adc_array_wafflecap_8_8_0[10|15]/adc_array_circuit_150n_0/vint1 col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2600 adc_array_wafflecap_8_8_0[10|5]/adc_array_circuit_150n_0/vint1 col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2601 adc_array_wafflecap_8_8_0[2|21]/adc_array_circuit_150n_0/vint2 col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2602 VSS VDD adc_array_wafflecap_8_Dummy_4[18]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2603 adc_array_wafflecap_8_8_0[7|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2604 vcm adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|22]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2605 adc_array_wafflecap_8_8_0[11|18]/adc_array_circuit_150n_0/vint2 col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2606 adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2607 adc_array_wafflecap_8_8_0[5|23]/adc_array_circuit_150n_0/vdrv row_n[6] adc_array_wafflecap_8_8_0[5|23]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2608 adc_array_wafflecap_8_8_0[4|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2609 adc_array_wafflecap_8_8_0[0|10]/adc_array_circuit_150n_0/vint2 rowon_n[1] adc_array_wafflecap_8_8_0[0|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2610 adc_array_wafflecap_8_8_0[7|25]/adc_array_circuit_150n_0/vint2 rowon_n[8] adc_array_wafflecap_8_8_0[7|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2611 vcm adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2612 adc_array_wafflecap_8_8_0[5|24]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|24]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2613 adc_array_wafflecap_8_8_0[3|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2614 vcm adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|27]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2615 VSS VSS adc_array_wafflecap_8_Dummy_8[5]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2616 VSS row_n[3] adc_array_wafflecap_8_8_0[2|6]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2617 VSS sample adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2618 adc_array_wafflecap_8_8_1[18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2619 adc_array_wafflecap_8_8_0[0|21]/adc_array_circuit_150n_0/vdrv row_n[1] adc_array_wafflecap_8_8_0[0|21]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2620 adc_array_wafflecap_8_Dummy_4[4]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[4]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2621 adc_array_wafflecap_8_Dummy_4[14]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[14]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2622 adc_array_wafflecap_8_8_0[14|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2623 adc_array_wafflecap_8_8_0[13|17]/adc_array_circuit_150n_0/vint1 col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2624 adc_array_wafflecap_8_8_0[13|24]/adc_array_circuit_150n_0/vint2 rowon_n[14] adc_array_wafflecap_8_8_0[13|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2625 adc_array_wafflecap_8_8_0[12|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2626 adc_array_wafflecap_8_8_0[12|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2627 vcm adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|3]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2628 vcm adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|13]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2629 adc_array_wafflecap_8_8_0[7|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2630 adc_array_wafflecap_8_8_0[4|25]/adc_array_circuit_150n_0/vint2 col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2631 VDD VSS adc_array_wafflecap_8_Dummy_1[1]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2632 adc_array_wafflecap_8_8_1[16]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[16]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2633 adc_array_wafflecap_8_8_0[1|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2634 adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2635 adc_array_wafflecap_8_8_0[5|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2636 adc_array_wafflecap_8_8_0[3|4]/adc_array_circuit_150n_0/vint2 col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2637 adc_array_wafflecap_8_8_0[10|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2638 adc_array_wafflecap_8_Dummy_1[6]/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_1[6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2639 adc_array_wafflecap_8_8_0[0|6]/adc_array_circuit_150n_0/vint1 col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2640 adc_array_wafflecap_8_8_0[9|20]/adc_array_circuit_150n_0/vint2 col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2641 adc_array_wafflecap_8_8_0[6|27]/adc_array_circuit_150n_0/vint2 rowon_n[7] adc_array_wafflecap_8_8_0[6|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2642 VSS row_n[1] adc_array_wafflecap_8_8_0[0|11]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2643 adc_array_wafflecap_8_8_0[3|27]/adc_array_circuit_150n_0/vdrv row_n[4] adc_array_wafflecap_8_8_0[3|27]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2644 adc_array_wafflecap_8_Dummy_4[18]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2645 adc_array_wafflecap_8_8_0[3|28]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|28]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2646 adc_array_wafflecap_8_8_0[0|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2647 adc_array_wafflecap_8_8_0[11|19]/adc_array_circuit_150n_0/vint1 col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2648 adc_array_wafflecap_8_8_0[9|7]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|7]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2649 VSS row_n[8] adc_array_wafflecap_8_8_0[7|4]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2650 VSS row_n[8] adc_array_wafflecap_8_8_0[7|14]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2651 adc_array_wafflecap_8_8_0[4|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2652 adc_array_wafflecap_8_8_0[7|20]/adc_array_circuit_150n_0/vdrv row_n[8] adc_array_wafflecap_8_8_0[7|20]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2653 adc_array_wafflecap_8_8_0[3|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2654 VSS row_n[14] adc_array_wafflecap_8_8_0[13|13]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2655 adc_array_wafflecap_8_8_0[14|19]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|19]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2656 VSS row_n[14] adc_array_wafflecap_8_8_0[13|3]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2657 VDD rowon_n[7] adc_array_wafflecap_8_8_0[6|27]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2658 adc_array_wafflecap_8_Dummy_1[2]/adc_array_circuit_150n_0/vint1 col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2659 adc_array_wafflecap_8_Dummy_3[5]/adc_array_circuit_150n_0/vint2 col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2660 adc_array_wafflecap_8_8_0[10|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2661 adc_array_wafflecap_8_8_0[2|16]/adc_array_circuit_150n_0/vdrv row_n[3] adc_array_wafflecap_8_8_0[2|16]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2662 VDD rowon_n[14] adc_array_wafflecap_8_8_0[13|17]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2663 adc_array_wafflecap_8_8_0[2|2]/adc_array_circuit_150n_0/vint2 rowon_n[3] adc_array_wafflecap_8_8_0[2|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2664 adc_array_wafflecap_8_8_0[12|12]/adc_array_circuit_150n_0/vint2 col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2665 VSS row_n[11] adc_array_wafflecap_8_8_0[10|16]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2666 adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2667 adc_array_wafflecap_8_8_0[12|2]/adc_array_circuit_150n_0/vint2 col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2668 adc_array_wafflecap_8_8_0[5|14]/adc_array_circuit_150n_0/vint2 rowon_n[6] adc_array_wafflecap_8_8_0[5|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2669 adc_array_wafflecap_8_8_0[2|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2670 VDD rowon_n[6] adc_array_wafflecap_8_8_0[5|4]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2671 vcm adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|20]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2672 vcm adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|21]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2673 vcm VSS adc_array_wafflecap_8_Dummy_4[21]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2674 adc_array_wafflecap_8_8_0[14|11]/adc_array_circuit_150n_0/vint1 col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2675 adc_array_wafflecap_8_8_0[11|8]/adc_array_circuit_150n_0/vdrv row_n[12] adc_array_wafflecap_8_8_0[11|8]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2676 adc_array_wafflecap_8_8_0[9|19]/adc_array_circuit_150n_0/vint2 rowon_n[10] adc_array_wafflecap_8_8_0[9|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2677 adc_array_wafflecap_8_8_0[5|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2678 adc_array_wafflecap_8_8_0[4|22]/adc_array_circuit_150n_0/vint1 col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2679 adc_array_wafflecap_8_8_0[4|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2680 VDD rowon_n[5] adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2681 adc_array_wafflecap_8_8_0[14|1]/adc_array_circuit_150n_0/vint1 col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2682 VDD rowon_n[1] adc_array_wafflecap_8_8_0[0|2]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2683 adc_array_wafflecap_8_8_0[14|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2684 adc_array_wafflecap_8_8_0[10|2]/adc_array_circuit_150n_0/vdrv row_n[11] adc_array_wafflecap_8_8_0[10|2]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2685 adc_array_wafflecap_8_8_0[10|12]/adc_array_circuit_150n_0/vdrv row_n[11] adc_array_wafflecap_8_8_0[10|12]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2686 adc_array_wafflecap_8_8_0[9|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2687 adc_array_wafflecap_8_8_0[8|16]/adc_array_circuit_150n_0/vint1 col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2688 adc_array_wafflecap_8_8_0[8|23]/adc_array_circuit_150n_0/vint2 rowon_n[9] adc_array_wafflecap_8_8_0[8|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2689 adc_array_wafflecap_8_8_1[19]/adc_array_circuit_150n_0/vint1 col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2690 adc_array_wafflecap_8_8_0[14|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2691 adc_array_wafflecap_8_8_0[7|4]/adc_array_circuit_150n_0/vint2 rowon_n[8] adc_array_wafflecap_8_8_0[7|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2692 adc_array_wafflecap_8_8_0[7|14]/adc_array_circuit_150n_0/vint2 rowon_n[8] adc_array_wafflecap_8_8_0[7|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2693 adc_array_wafflecap_8_8_0[13|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2694 vcm adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|11]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2695 adc_array_wafflecap_8_8_0[8|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2696 adc_array_wafflecap_8_8_0[8|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2697 adc_array_wafflecap_8_8_0[4|6]/adc_array_circuit_150n_0/vint2 rowon_n[5] adc_array_wafflecap_8_8_0[4|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2698 VSS row_n[0] adc_array_wafflecap_8_8_1[24]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2699 adc_array_wafflecap_8_8_1[17]/adc_array_circuit_150n_0/vdrv row_n[0] adc_array_wafflecap_8_8_1[17]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2700 adc_array_wafflecap_8_Dummy_4[29]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2701 adc_array_wafflecap_8_8_0[13|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2702 vcm adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|1]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2703 adc_array_wafflecap_8_8_0[5|29]/adc_array_circuit_150n_0/vint2 col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2704 vcm adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|9]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2705 VDD rowon_n[8] adc_array_wafflecap_8_8_0[7|19]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2706 VSS row_n[3] adc_array_wafflecap_8_8_0[2|3]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2707 adc_array_wafflecap_8_8_0[11|29]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|29]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2708 VSS row_n[6] adc_array_wafflecap_8_8_0[5|15]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2709 vcm adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|25]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2710 VSS row_n[14] adc_array_wafflecap_8_8_0[13|21]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2711 vcm adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|3]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2712 adc_array_wafflecap_8_8_0[5|5]/adc_array_circuit_150n_0/vint1 col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2713 adc_array_wafflecap_8_Dummy_4[16]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2714 adc_array_wafflecap_8_8_0[14|27]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|27]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2715 adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/vint2 col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2716 adc_array_wafflecap_8_Dummy_4[6]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2717 VDD sample adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2718 adc_array_wafflecap_8_8_0[2|26]/adc_array_circuit_150n_0/vint1 col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2719 adc_array_wafflecap_8_8_0[2|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2720 adc_array_wafflecap_8_Dummy_3[3]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2721 adc_array_wafflecap_8_8_0[0|3]/adc_array_circuit_150n_0/vint1 col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2722 VSS row_n[10] adc_array_wafflecap_8_8_0[9|8]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2723 VDD VDD adc_array_wafflecap_8_Dummy_4[21]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2724 VSS row_n[9] adc_array_wafflecap_8_8_0[8|12]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2725 vcm adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|14]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2726 VDD rowon_n[15] adc_array_wafflecap_8_8_0[14|11]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2727 adc_array_wafflecap_8_8_0[11|30]/adc_array_circuit_150n_0/vint1 col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2728 adc_array_wafflecap_8_8_0[9|18]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|18]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2729 VSS row_n[9] adc_array_wafflecap_8_8_0[8|2]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2730 VDD rowon_n[15] adc_array_wafflecap_8_8_0[14|1]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2731 VDD rowon_n[14] adc_array_wafflecap_8_8_0[13|15]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2732 adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/vdrv row_n[8] adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2733 adc_array_wafflecap_8_8_0[3|21]/adc_array_circuit_150n_0/vint2 rowon_n[4] adc_array_wafflecap_8_8_0[3|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2734 VDD rowon_n[14] adc_array_wafflecap_8_8_0[13|5]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2735 adc_array_wafflecap_8_8_0[11|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2736 adc_array_wafflecap_8_8_0[7|8]/adc_array_circuit_150n_0/vint1 col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2737 adc_array_wafflecap_8_8_0[0|22]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|22]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2738 adc_array_wafflecap_8_8_0[14|6]/adc_array_circuit_150n_0/vint2 col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2739 adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2740 adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2741 adc_array_wafflecap_8_8_0[3|0]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|0]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2742 adc_array_wafflecap_8_8_0[13|0]/adc_array_circuit_150n_0/vint2 col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2743 adc_array_wafflecap_8_8_0[13|10]/adc_array_circuit_150n_0/vint2 col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2744 adc_array_wafflecap_8_8_0[6|12]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|12]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2745 adc_array_wafflecap_8_8_0[0|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2746 adc_array_wafflecap_8_Dummy_4[33]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[33]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2747 vcm adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2748 adc_array_wafflecap_8_8_0[4|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2749 vcm adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|17]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2750 adc_array_wafflecap_8_Dummy_8[0]/adc_array_circuit_150n_0/vint2 col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2751 adc_array_wafflecap_8_8_1[10]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[10]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2752 vcm adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|18]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2753 adc_array_wafflecap_8_Dummy_4[0]/adc_array_circuit_150n_0/vint1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2754 adc_array_wafflecap_8_Dummy_4[10]/adc_array_circuit_150n_0/vint1 col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2755 vcm VSS adc_array_wafflecap_8_Dummy_4[32]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2756 adc_array_wafflecap_8_8_0[12|6]/adc_array_circuit_150n_0/vdrv row_n[13] adc_array_wafflecap_8_8_0[12|6]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2757 adc_array_wafflecap_8_8_0[11|19]/adc_array_circuit_150n_0/vdrv row_n[12] adc_array_wafflecap_8_8_0[11|19]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2758 adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2759 adc_array_wafflecap_8_8_0[9|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2760 adc_array_wafflecap_8_8_0[6|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2761 adc_array_wafflecap_8_8_0[5|25]/adc_array_circuit_150n_0/vint2 rowon_n[6] adc_array_wafflecap_8_8_0[5|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2762 adc_array_wafflecap_8_Dummy_4[27]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2763 adc_array_wafflecap_8_Dummy_4[9]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2764 adc_array_wafflecap_8_8_0[12|23]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|23]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2765 adc_array_wafflecap_8_8_0[10|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2766 adc_array_wafflecap_8_8_0[8|12]/adc_array_circuit_150n_0/vint2 rowon_n[9] adc_array_wafflecap_8_8_0[8|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2767 adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2768 adc_array_wafflecap_8_8_0[8|2]/adc_array_circuit_150n_0/vint2 rowon_n[9] adc_array_wafflecap_8_8_0[8|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2769 adc_array_wafflecap_8_8_0[1|5]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|5]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2770 VSS sample_n adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2771 vcm adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|9]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2772 VSS row_n[5] adc_array_wafflecap_8_8_0[4|28]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2773 adc_array_wafflecap_8_8_0[6|9]/adc_array_circuit_150n_0/vint2 col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2774 adc_array_wafflecap_8_4_0/adc_array_circuit_150n_0/vint2 en_n_bit[2] adc_array_wafflecap_8_4_0/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2775 adc_array_wafflecap_8_Dummy_3[0]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_3[0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2776 adc_array_wafflecap_8_8_0[3|21]/adc_array_circuit_150n_0/vdrv row_n[4] adc_array_wafflecap_8_8_0[3|21]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2777 adc_array_wafflecap_8_8_0[2|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2778 vcm adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|7]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2779 adc_array_wafflecap_8_8_0[5|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2780 adc_array_wafflecap_8_8_0[1|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2781 VSS row_n[15] adc_array_wafflecap_8_8_0[14|28]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2782 adc_array_wafflecap_8_8_0[8|12]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|12]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2783 adc_array_wafflecap_8_8_0[8|2]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|2]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2784 VSS row_n[14] adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2785 adc_array_wafflecap_8_8_0[10|29]/adc_array_circuit_150n_0/vint2 col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2786 adc_array_wafflecap_8_8_0[3|6]/adc_array_circuit_150n_0/vint1 col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2787 adc_array_wafflecap_8_1_0/adc_array_circuit_150n_0/vint2 en_n_bit[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2788 adc_array_wafflecap_8_8_0[6|9]/adc_array_circuit_150n_0/vdrv row_n[7] adc_array_wafflecap_8_8_0[6|9]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2789 adc_array_wafflecap_8_8_0[3|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2790 adc_array_wafflecap_8_8_0[2|23]/adc_array_circuit_150n_0/vint2 col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2791 VDD rowon_n[10] adc_array_wafflecap_8_8_0[9|0]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2792 VDD rowon_n[10] adc_array_wafflecap_8_8_0[9|10]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2793 adc_array_wafflecap_8_8_0[5|1]/adc_array_circuit_150n_0/vint2 col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2794 adc_array_wafflecap_8_Dummy_4[16]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[16]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2795 VDD VDD adc_array_wafflecap_8_Dummy_4[32]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2796 adc_array_wafflecap_8_8_0[14|24]/adc_array_circuit_150n_0/vdrv row_n[15] adc_array_wafflecap_8_8_0[14|24]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2797 adc_array_wafflecap_8_Dummy_4[6]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[6]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2798 VDD VDD adc_array_wafflecap_8_Dummy_4[10]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2799 adc_array_wafflecap_8_8_0[12|28]/adc_array_circuit_150n_0/vint1 col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2800 adc_array_wafflecap_8_8_0[5|25]/adc_array_circuit_150n_0/vdrv row_n[6] adc_array_wafflecap_8_8_0[5|25]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2801 adc_array_wafflecap_8_8_0[5|26]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|26]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2802 VDD VDD adc_array_wafflecap_8_Dummy_4[0]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2803 adc_array_wafflecap_8_8_0[8|29]/adc_array_circuit_150n_0/vdrv row_n[9] adc_array_wafflecap_8_8_0[8|29]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2804 VSS VSS adc_array_wafflecap_8_Dummy_1[0]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2805 adc_array_wafflecap_8_8_0[0|23]/adc_array_circuit_150n_0/vdrv row_n[1] adc_array_wafflecap_8_8_0[0|23]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2806 adc_array_wafflecap_8_8_1[20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2807 adc_array_wafflecap_8_8_0[5|7]/adc_array_circuit_150n_0/vint2 rowon_n[6] adc_array_wafflecap_8_8_0[5|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2808 adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2809 adc_array_wafflecap_8_Dummy_0[1]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2810 adc_array_wafflecap_8_8_0[11|27]/adc_array_circuit_150n_0/vdrv row_n[12] adc_array_wafflecap_8_8_0[11|27]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2811 adc_array_wafflecap_8_8_0[5|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2812 adc_array_wafflecap_8_8_0[4|14]/adc_array_circuit_150n_0/vdrv row_n[5] adc_array_wafflecap_8_8_0[4|14]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2813 adc_array_wafflecap_8_8_0[1|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2814 adc_array_wafflecap_8_8_0[14|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2815 adc_array_wafflecap_8_8_1[16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_1[16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2816 vcm adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[6]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2817 adc_array_wafflecap_8_8_0[0|27]/adc_array_circuit_150n_0/vint2 col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2818 vcm adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|30]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2819 VSS row_n[7] adc_array_wafflecap_8_8_0[6|19]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2820 adc_array_wafflecap_8_8_0[6|29]/adc_array_circuit_150n_0/vint2 rowon_n[7] adc_array_wafflecap_8_8_0[6|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2821 adc_array_wafflecap_8_8_0[10|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2822 adc_array_wafflecap_8_8_0[6|17]/adc_array_circuit_150n_0/vint2 col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2823 adc_array_wafflecap_8_8_0[13|21]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|21]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2824 adc_array_wafflecap_8_8_0[3|30]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|30]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2825 adc_array_wafflecap_8_8_0[3|12]/adc_array_circuit_150n_0/vint2 rowon_n[4] adc_array_wafflecap_8_8_0[3|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2826 adc_array_wafflecap_8_8_0[0|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2827 adc_array_wafflecap_8_8_0[3|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2828 adc_array_wafflecap_8_8_1[15]/adc_array_circuit_150n_0/vint2 col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2829 VSS row_n[6] adc_array_wafflecap_8_8_0[5|8]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2830 VDD rowon_n[4] adc_array_wafflecap_8_8_0[3|2]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2831 adc_array_wafflecap_8_Dummy_3[2]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_3[2]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2832 adc_array_wafflecap_8_8_0[6|19]/adc_array_circuit_150n_0/vint1 col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2833 adc_array_wafflecap_8_8_0[2|20]/adc_array_circuit_150n_0/vint1 col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2834 adc_array_wafflecap_8_8_0[12|8]/adc_array_circuit_150n_0/vint2 rowon_n[13] adc_array_wafflecap_8_8_0[12|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2835 adc_array_wafflecap_8_8_0[12|30]/adc_array_circuit_150n_0/vint2 rowon_n[13] adc_array_wafflecap_8_8_0[12|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2836 adc_array_wafflecap_8_8_0[11|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2837 VSS row_n[10] adc_array_wafflecap_8_8_0[9|27]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2838 VDD rowon_n[7] adc_array_wafflecap_8_8_0[6|29]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2839 adc_array_wafflecap_8_8_0[3|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2840 adc_array_wafflecap_8_Dummy_6/adc_array_circuit_150n_0/vint2 VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2841 adc_array_wafflecap_8_8_0[11|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2842 adc_array_wafflecap_8_8_0[6|17]/adc_array_circuit_150n_0/vdrv row_n[7] adc_array_wafflecap_8_8_0[6|17]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2843 adc_array_wafflecap_8_8_0[2|18]/adc_array_circuit_150n_0/vdrv row_n[3] adc_array_wafflecap_8_8_0[2|18]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2844 adc_array_wafflecap_8_8_0[2|19]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|19]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2845 vcm adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|18]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2846 VSS row_n[9] adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2847 adc_array_wafflecap_8_8_0[2|4]/adc_array_circuit_150n_0/vint2 rowon_n[3] adc_array_wafflecap_8_8_0[2|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2848 VDD rowon_n[12] adc_array_wafflecap_8_8_0[11|26]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2849 adc_array_wafflecap_8_8_0[5|16]/adc_array_circuit_150n_0/vint2 rowon_n[6] adc_array_wafflecap_8_8_0[5|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2850 VSS row_n[5] adc_array_wafflecap_8_8_0[4|0]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2851 VDD rowon_n[11] adc_array_wafflecap_8_8_0[10|8]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2852 VDD rowon_n[11] adc_array_wafflecap_8_8_0[10|30]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2853 adc_array_wafflecap_8_8_0[9|23]/adc_array_circuit_150n_0/vdrv row_n[10] adc_array_wafflecap_8_8_0[9|23]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2854 adc_array_wafflecap_8_8_0[7|27]/adc_array_circuit_150n_0/vint1 col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2855 VDD rowon_n[6] adc_array_wafflecap_8_8_0[5|6]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2856 VSS row_n[4] adc_array_wafflecap_8_8_0[3|13]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2857 vcm adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|22]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2858 adc_array_wafflecap_8_8_0[4|24]/adc_array_circuit_150n_0/vint1 col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2859 vcm adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|23]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2860 adc_array_wafflecap_8_8_0[12|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2861 adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2862 adc_array_wafflecap_8_8_0[4|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2863 adc_array_wafflecap_8_8_0[3|3]/adc_array_circuit_150n_0/vint1 col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2864 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X2865 VDD rowon_n[1] adc_array_wafflecap_8_8_0[0|4]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2866 vcm adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|26]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2867 adc_array_wafflecap_8_8_1[21]/adc_array_circuit_150n_0/vint1 col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2868 adc_array_wafflecap_8_8_0[14|15]/adc_array_circuit_150n_0/vint2 col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2869 VSS row_n[14] adc_array_wafflecap_8_8_0[13|6]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2870 adc_array_wafflecap_8_8_0[9|16]/adc_array_circuit_150n_0/vint2 col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2871 VDD rowon_n[0] adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2872 adc_array_wafflecap_8_8_0[14|5]/adc_array_circuit_150n_0/vint2 col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2873 adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/vint2 col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2874 vcm adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|11]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2875 VSS row_n[3] adc_array_wafflecap_8_8_0[2|5]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2876 VSS row_n[0] adc_array_wafflecap_8_8_1[25]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2877 adc_array_wafflecap_8_Dummy_4[28]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2878 vcm adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|5]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2879 adc_array_wafflecap_8_8_0[5|18]/adc_array_circuit_150n_0/vint2 rowon_n[6] adc_array_wafflecap_8_8_0[5|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2880 adc_array_wafflecap_8_8_0[1|19]/adc_array_circuit_150n_0/vint2 rowon_n[2] adc_array_wafflecap_8_8_0[1|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2881 adc_array_wafflecap_8_8_0[12|5]/adc_array_circuit_150n_0/vdrv row_n[13] adc_array_wafflecap_8_8_0[12|5]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2882 adc_array_wafflecap_8_8_0[12|15]/adc_array_circuit_150n_0/vdrv row_n[13] adc_array_wafflecap_8_8_0[12|15]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2883 adc_array_wafflecap_8_8_0[12|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2884 vcm adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|28]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2885 adc_array_wafflecap_8_8_0[7|16]/adc_array_circuit_150n_0/vdrv row_n[8] adc_array_wafflecap_8_8_0[7|16]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2886 VSS row_n[8] adc_array_wafflecap_8_8_0[7|23]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2887 VSS row_n[2] adc_array_wafflecap_8_8_0[1|17]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2888 adc_array_wafflecap_8_8_0[1|7]/adc_array_circuit_150n_0/vint2 col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2889 VSS row_n[6] adc_array_wafflecap_8_8_0[5|16]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2890 adc_array_wafflecap_8_Dummy_2[3]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_2[3]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2891 vcm adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|14]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2892 adc_array_wafflecap_8_8_0[2|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2893 adc_array_wafflecap_8_Dummy_3[5]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2894 vcm adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[3]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2895 adc_array_wafflecap_8_8_0[0|5]/adc_array_circuit_150n_0/vint1 col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2896 vcm adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|4]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2897 adc_array_wafflecap_8_8_0[10|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2898 VDD rowon_n[10] adc_array_wafflecap_8_8_0[9|22]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2899 vcm adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|16]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2900 VDD rowon_n[2] adc_array_wafflecap_8_8_0[1|19]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2901 adc_array_wafflecap_8_8_0[1|7]/adc_array_circuit_150n_0/vdrv row_n[2] adc_array_wafflecap_8_8_0[1|7]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2902 VSS VDD adc_array_wafflecap_8_Dummy_4[25]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2903 adc_array_wafflecap_8_8_0[12|21]/adc_array_circuit_150n_0/vint2 col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2904 adc_array_wafflecap_8_8_0[3|23]/adc_array_circuit_150n_0/vint2 rowon_n[4] adc_array_wafflecap_8_8_0[3|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2905 adc_array_wafflecap_8_8_0[1|17]/adc_array_circuit_150n_0/vint1 col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2906 adc_array_wafflecap_8_Dummy_4[18]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[18]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2907 adc_array_wafflecap_8_8_0[13|28]/adc_array_circuit_150n_0/vint2 rowon_n[14] adc_array_wafflecap_8_8_0[13|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2908 vcm adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|17]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2909 adc_array_wafflecap_8_8_0[11|25]/adc_array_circuit_150n_0/vint2 col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2910 adc_array_wafflecap_8_8_0[3|2]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|2]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2911 adc_array_wafflecap_8_Dummy_4[12]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2912 adc_array_wafflecap_8_8_0[14|20]/adc_array_circuit_150n_0/vint1 col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2913 adc_array_wafflecap_8_8_0[12|8]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|8]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2914 VSS row_n[11] adc_array_wafflecap_8_8_0[10|15]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2915 adc_array_wafflecap_8_Dummy_4[2]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2916 VSS row_n[11] adc_array_wafflecap_8_8_0[10|5]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2917 adc_array_wafflecap_8_8_0[13|24]/adc_array_circuit_150n_0/vint1 col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2918 adc_array_wafflecap_8_8_0[11|12]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|12]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2919 adc_array_wafflecap_8_8_0[10|21]/adc_array_circuit_150n_0/vdrv row_n[11] adc_array_wafflecap_8_8_0[10|21]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2920 adc_array_wafflecap_8_8_0[7|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2921 adc_array_wafflecap_8_8_0[4|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2922 adc_array_wafflecap_8_8_0[0|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2923 adc_array_wafflecap_8_8_0[11|2]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|2]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2924 adc_array_wafflecap_8_8_0[5|28]/adc_array_circuit_150n_0/vint1 col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2925 adc_array_wafflecap_8_8_0[3|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2926 adc_array_wafflecap_8_8_0[6|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2927 adc_array_wafflecap_8_8_1[12]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[12]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2928 adc_array_wafflecap_8_8_0[13|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2929 adc_array_wafflecap_8_8_0[8|15]/adc_array_circuit_150n_0/vint1 col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2930 adc_array_wafflecap_8_8_0[8|5]/adc_array_circuit_150n_0/vint1 col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2931 adc_array_wafflecap_8_8_0[4|20]/adc_array_circuit_150n_0/vint2 col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2932 adc_array_wafflecap_8_8_0[0|21]/adc_array_circuit_150n_0/vint2 col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2933 adc_array_wafflecap_8_Dummy_4[4]/adc_array_circuit_150n_0/vint2 col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2934 adc_array_wafflecap_8_Dummy_4[14]/adc_array_circuit_150n_0/vint2 col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2935 VSS row_n[14] adc_array_wafflecap_8_8_0[13|17]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2936 VSS row_n[5] adc_array_wafflecap_8_8_0[4|30]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2937 adc_array_wafflecap_8_8_0[7|23]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|23]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2938 adc_array_wafflecap_8_8_0[6|11]/adc_array_circuit_150n_0/vint2 col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2939 vcm adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|22]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2940 adc_array_wafflecap_8_8_0[3|23]/adc_array_circuit_150n_0/vdrv row_n[4] adc_array_wafflecap_8_8_0[3|23]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2941 adc_array_wafflecap_8_Dummy_1[1]/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_1[1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2942 adc_array_wafflecap_8_8_0[2|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2943 adc_array_wafflecap_8_8_0[5|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2944 adc_array_wafflecap_8_8_0[3|24]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|24]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2945 adc_array_wafflecap_8_8_0[1|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2946 adc_array_wafflecap_8_8_0[14|9]/adc_array_circuit_150n_0/vdrv row_n[15] adc_array_wafflecap_8_8_0[14|9]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2947 VSS row_n[1] adc_array_wafflecap_8_8_0[0|6]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2948 adc_array_wafflecap_8_8_0[13|13]/adc_array_circuit_150n_0/vdrv row_n[14] adc_array_wafflecap_8_8_0[13|13]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2949 adc_array_wafflecap_8_Dummy_2[4]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_2[4]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2950 adc_array_wafflecap_8_8_0[14|26]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|26]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2951 adc_array_wafflecap_8_8_0[13|3]/adc_array_circuit_150n_0/vdrv row_n[14] adc_array_wafflecap_8_8_0[13|3]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2952 adc_array_wafflecap_8_8_0[12|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2953 adc_array_wafflecap_8_8_0[11|24]/adc_array_circuit_150n_0/vint2 rowon_n[12] adc_array_wafflecap_8_8_0[11|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2954 adc_array_wafflecap_8_8_0[10|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2955 adc_array_wafflecap_8_8_0[10|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2956 vcm adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|3]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2957 vcm adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|13]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2958 adc_array_wafflecap_8_8_0[2|25]/adc_array_circuit_150n_0/vint2 col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2959 adc_array_wafflecap_8_8_0[6|11]/adc_array_circuit_150n_0/vdrv row_n[7] adc_array_wafflecap_8_8_0[6|11]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2960 adc_array_wafflecap_8_8_0[5|3]/adc_array_circuit_150n_0/vint2 col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2961 adc_array_wafflecap_8_8_0[3|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2962 adc_array_wafflecap_8_8_0[1|4]/adc_array_circuit_150n_0/vint2 col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2963 adc_array_wafflecap_8_Dummy_8[4]/adc_array_circuit_150n_0/vint1 col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2964 adc_array_wafflecap_8_8_0[7|20]/adc_array_circuit_150n_0/vint2 col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2965 VSS VSS adc_array_wafflecap_8_Dummy_1[2]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2966 adc_array_wafflecap_8_8_0[0|25]/adc_array_circuit_150n_0/vdrv row_n[1] adc_array_wafflecap_8_8_0[0|25]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2967 adc_array_wafflecap_8_8_0[13|17]/adc_array_circuit_150n_0/vint2 rowon_n[14] adc_array_wafflecap_8_8_0[13|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2968 adc_array_wafflecap_8_8_0[5|27]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|27]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2969 adc_array_wafflecap_8_Dummy_8[0]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2970 adc_array_wafflecap_8_8_0[1|28]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|28]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2971 adc_array_wafflecap_8_8_0[9|19]/adc_array_circuit_150n_0/vint1 col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2972 adc_array_wafflecap_8_8_0[5|9]/adc_array_circuit_150n_0/vint2 rowon_n[6] adc_array_wafflecap_8_8_0[5|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2973 adc_array_wafflecap_8_8_0[2|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2974 adc_array_wafflecap_8_8_0[1|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2975 adc_array_wafflecap_8_8_0[1|4]/adc_array_circuit_150n_0/vdrv row_n[2] adc_array_wafflecap_8_8_0[1|4]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2976 VDD rowon_n[12] adc_array_wafflecap_8_8_0[11|3]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2977 VDD rowon_n[12] adc_array_wafflecap_8_8_0[11|13]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2978 VSS row_n[12] adc_array_wafflecap_8_8_0[11|13]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2979 adc_array_wafflecap_8_8_0[12|19]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|19]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2980 VSS row_n[12] adc_array_wafflecap_8_8_0[11|3]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2981 VDD rowon_n[5] adc_array_wafflecap_8_8_0[4|27]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2982 adc_array_wafflecap_8_8_0[8|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2983 VSS row_n[7] adc_array_wafflecap_8_8_0[6|21]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2984 adc_array_wafflecap_8_8_1[13]/adc_array_circuit_150n_0/vdrv row_n[0] adc_array_wafflecap_8_8_1[13]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2985 VSS row_n[15] adc_array_wafflecap_8_8_0[14|11]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2986 adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/vint2 rowon_n[7] adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2987 VSS row_n[15] adc_array_wafflecap_8_8_0[14|1]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2988 adc_array_wafflecap_8_8_0[0|2]/adc_array_circuit_150n_0/vint2 rowon_n[1] adc_array_wafflecap_8_8_0[0|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2989 adc_array_wafflecap_8_8_0[10|12]/adc_array_circuit_150n_0/vint2 col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2990 VSS row_n[9] adc_array_wafflecap_8_8_0[8|16]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2991 adc_array_wafflecap_8_8_0[4|1]/adc_array_circuit_150n_0/vint2 rowon_n[5] adc_array_wafflecap_8_8_0[4|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2992 adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2993 adc_array_wafflecap_8_8_0[3|14]/adc_array_circuit_150n_0/vint2 rowon_n[4] adc_array_wafflecap_8_8_0[3|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2994 VSS row_n[0] adc_array_wafflecap_8_8_1[19]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2995 adc_array_wafflecap_8_8_0[0|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2996 adc_array_wafflecap_8_8_0[10|2]/adc_array_circuit_150n_0/vint2 col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2997 VDD rowon_n[4] adc_array_wafflecap_8_8_0[3|4]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2998 adc_array_wafflecap_8_8_1[17]/adc_array_circuit_150n_0/vint2 col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2999 VSS row_n[6] adc_array_wafflecap_8_8_0[5|10]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3000 vcm adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|20]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3001 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.64e+07u l=1.6e+07u
X3002 vcm adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|20]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3003 adc_array_wafflecap_8_8_0[12|11]/adc_array_circuit_150n_0/vint1 col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3004 adc_array_wafflecap_8_8_0[9|8]/adc_array_circuit_150n_0/vdrv row_n[10] adc_array_wafflecap_8_8_0[9|8]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3005 adc_array_wafflecap_8_8_0[8|21]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|21]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3006 adc_array_wafflecap_8_8_0[7|19]/adc_array_circuit_150n_0/vint2 rowon_n[8] adc_array_wafflecap_8_8_0[7|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3007 adc_array_wafflecap_8_8_0[6|21]/adc_array_circuit_150n_0/vint1 col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3008 adc_array_wafflecap_8_8_0[3|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3009 adc_array_wafflecap_8_8_0[2|22]/adc_array_circuit_150n_0/vint1 col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3010 adc_array_wafflecap_8_8_0[2|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3011 VDD rowon_n[3] adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3012 adc_array_wafflecap_8_8_0[12|1]/adc_array_circuit_150n_0/vint1 col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3013 VDD rowon_n[7] adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3014 adc_array_wafflecap_8_8_0[5|0]/adc_array_circuit_150n_0/vint1 col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3015 VDD VSS adc_array_wafflecap_8_Dummy_8[0]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3016 adc_array_wafflecap_8_8_0[12|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3017 adc_array_wafflecap_8_8_0[9|25]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|25]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3018 adc_array_wafflecap_8_8_0[8|2]/adc_array_circuit_150n_0/vdrv row_n[9] adc_array_wafflecap_8_8_0[8|2]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3019 adc_array_wafflecap_8_8_0[8|12]/adc_array_circuit_150n_0/vdrv row_n[9] adc_array_wafflecap_8_8_0[8|12]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3020 adc_array_wafflecap_8_8_0[12|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3021 adc_array_wafflecap_8_8_0[2|6]/adc_array_circuit_150n_0/vint2 rowon_n[3] adc_array_wafflecap_8_8_0[2|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3022 adc_array_wafflecap_8_8_0[11|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3023 vcm adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|11]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3024 adc_array_wafflecap_8_Dummy_4[25]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[25]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3025 adc_array_wafflecap_8_8_0[13|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3026 adc_array_wafflecap_8_8_0[11|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3027 vcm adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|1]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3028 adc_array_wafflecap_8_8_0[3|29]/adc_array_circuit_150n_0/vint2 col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3029 vcm adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|9]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3030 VSS row_n[5] adc_array_wafflecap_8_8_0[4|2]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3031 VSS row_n[1] adc_array_wafflecap_8_8_0[0|3]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3032 VSS row_n[4] adc_array_wafflecap_8_8_0[3|15]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3033 vcm adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|25]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3034 adc_array_wafflecap_8_Dummy_4[21]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3035 adc_array_wafflecap_8_8_0[14|1]/adc_array_circuit_150n_0/vint2 rowon_n[15] adc_array_wafflecap_8_8_0[14|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3036 adc_array_wafflecap_8_8_0[14|11]/adc_array_circuit_150n_0/vint2 rowon_n[15] adc_array_wafflecap_8_8_0[14|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3037 VSS row_n[12] adc_array_wafflecap_8_8_0[11|21]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3038 adc_array_wafflecap_8_8_0[3|5]/adc_array_circuit_150n_0/vint1 col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3039 VDD rowon_n[1] adc_array_wafflecap_8_8_0[0|6]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3040 adc_array_wafflecap_8_8_0[13|15]/adc_array_circuit_150n_0/vint2 rowon_n[14] adc_array_wafflecap_8_8_0[13|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3041 adc_array_wafflecap_8_8_0[12|27]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|27]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3042 adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/vint2 col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3043 adc_array_wafflecap_8_8_1[23]/adc_array_circuit_150n_0/vint1 col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3044 adc_array_wafflecap_8_8_0[13|5]/adc_array_circuit_150n_0/vint2 rowon_n[14] adc_array_wafflecap_8_8_0[13|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3045 VDD sample adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3046 adc_array_wafflecap_8_Dummy_8[1]/adc_array_circuit_150n_0/vint1 col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3047 adc_array_wafflecap_8_8_0[0|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3048 VSS row_n[8] adc_array_wafflecap_8_8_0[7|8]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3049 VDD rowon_n[14] adc_array_wafflecap_8_8_0[13|20]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3050 adc_array_wafflecap_8_8_0[6|7]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|7]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3051 vcm adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|13]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3052 vcm adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|14]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3053 VDD rowon_n[13] adc_array_wafflecap_8_8_0[12|11]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3054 adc_array_wafflecap_8_8_0[9|30]/adc_array_circuit_150n_0/vint1 col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3055 adc_array_wafflecap_8_8_0[6|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3056 VDD rowon_n[13] adc_array_wafflecap_8_8_0[12|1]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3057 adc_array_wafflecap_8_8_0[1|21]/adc_array_circuit_150n_0/vint2 rowon_n[2] adc_array_wafflecap_8_8_0[1|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3058 adc_array_wafflecap_8_Dummy_4[33]/adc_array_circuit_150n_0/vint2 VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3059 adc_array_wafflecap_8_8_0[5|20]/adc_array_circuit_150n_0/vint2 rowon_n[6] adc_array_wafflecap_8_8_0[5|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3060 adc_array_wafflecap_8_Dummy_2[5]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_2[5]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3061 VSS VDD adc_array_wafflecap_8_Dummy_4[10]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3062 adc_array_wafflecap_8_8_0[12|6]/adc_array_circuit_150n_0/vint2 col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3063 adc_array_wafflecap_8_Dummy_6/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3064 VSS VDD adc_array_wafflecap_8_Dummy_4[0]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3065 adc_array_wafflecap_8_8_0[7|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3066 adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3067 vcm adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[5]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3068 adc_array_wafflecap_8_8_0[1|0]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|0]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3069 adc_array_wafflecap_8_8_0[14|28]/adc_array_circuit_150n_0/vdrv row_n[15] adc_array_wafflecap_8_8_0[14|28]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3070 adc_array_wafflecap_8_8_0[11|0]/adc_array_circuit_150n_0/vint2 col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3071 adc_array_wafflecap_8_8_0[11|10]/adc_array_circuit_150n_0/vint2 col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3072 adc_array_wafflecap_8_Dummy_2[3]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_2[3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3073 adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/vdrv row_n[14] adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3074 vcm adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3075 VDD rowon_n[2] adc_array_wafflecap_8_8_0[1|21]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3076 adc_array_wafflecap_8_8_0[2|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3077 adc_array_wafflecap_8_8_0[3|25]/adc_array_circuit_150n_0/vint2 rowon_n[4] adc_array_wafflecap_8_8_0[3|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3078 vcm VSS adc_array_wafflecap_8_Dummy_2[1]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3079 vcm adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|17]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3080 adc_array_wafflecap_8_8_0[14|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3081 adc_array_wafflecap_8_8_0[13|9]/adc_array_circuit_150n_0/vint1 col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3082 vcm adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3083 adc_array_wafflecap_8_8_0[10|6]/adc_array_circuit_150n_0/vdrv row_n[11] adc_array_wafflecap_8_8_0[10|6]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3084 adc_array_wafflecap_8_8_0[9|19]/adc_array_circuit_150n_0/vdrv row_n[10] adc_array_wafflecap_8_8_0[9|19]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3085 adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3086 adc_array_wafflecap_8_8_0[7|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3087 adc_array_wafflecap_8_8_0[13|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3088 adc_array_wafflecap_8_8_0[13|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3089 adc_array_wafflecap_8_8_0[10|23]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|23]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3090 adc_array_wafflecap_8_8_0[9|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3091 VSS row_n[3] adc_array_wafflecap_8_8_0[2|28]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3092 adc_array_wafflecap_8_8_0[9|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3093 adc_array_wafflecap_8_8_0[9|0]/adc_array_circuit_150n_0/vint2 rowon_n[10] adc_array_wafflecap_8_8_0[9|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3094 adc_array_wafflecap_8_8_0[9|10]/adc_array_circuit_150n_0/vint2 rowon_n[10] adc_array_wafflecap_8_8_0[9|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3095 adc_array_wafflecap_8_8_0[7|8]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|8]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3096 vcm adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|28]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3097 adc_array_wafflecap_8_8_0[5|20]/adc_array_circuit_150n_0/vdrv row_n[6] adc_array_wafflecap_8_8_0[5|20]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3098 adc_array_wafflecap_8_8_0[5|21]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|21]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3099 adc_array_wafflecap_8_8_0[0|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3100 vcm adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|7]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3101 adc_array_wafflecap_8_8_0[5|30]/adc_array_circuit_150n_0/vint1 col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3102 adc_array_wafflecap_8_8_0[3|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3103 adc_array_wafflecap_8_8_1[14]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[14]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3104 adc_array_wafflecap_8_Dummy_4[10]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3105 adc_array_wafflecap_8_Dummy_4[32]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[32]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3106 adc_array_wafflecap_8_8_0[14|24]/adc_array_circuit_150n_0/vint2 col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3107 VSS row_n[13] adc_array_wafflecap_8_8_0[12|28]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3108 adc_array_wafflecap_8_8_0[6|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3109 adc_array_wafflecap_8_Dummy_4[0]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3110 VSS row_n[12] adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3111 adc_array_wafflecap_8_8_0[8|29]/adc_array_circuit_150n_0/vint2 col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3112 adc_array_wafflecap_8_8_0[0|28]/adc_array_circuit_150n_0/vint1 col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3113 adc_array_wafflecap_8_8_0[14|11]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|11]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3114 adc_array_wafflecap_8_8_0[4|9]/adc_array_circuit_150n_0/vdrv row_n[5] adc_array_wafflecap_8_8_0[4|9]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3115 adc_array_wafflecap_8_8_0[4|22]/adc_array_circuit_150n_0/vint2 col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3116 adc_array_wafflecap_8_8_1[12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_1[12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3117 adc_array_wafflecap_8_8_0[0|23]/adc_array_circuit_150n_0/vint2 col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3118 adc_array_wafflecap_8_8_0[1|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3119 adc_array_wafflecap_8_8_0[14|1]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|1]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3120 VDD rowon_n[15] adc_array_wafflecap_8_8_0[14|27]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3121 VDD rowon_n[8] adc_array_wafflecap_8_8_0[7|0]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3122 VDD rowon_n[8] adc_array_wafflecap_8_8_0[7|10]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3123 VSS row_n[5] adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3124 adc_array_wafflecap_8_8_0[3|1]/adc_array_circuit_150n_0/vint2 col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3125 adc_array_wafflecap_8_8_0[13|15]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|15]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3126 VDD rowon_n[14] adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3127 adc_array_wafflecap_8_8_0[12|24]/adc_array_circuit_150n_0/vdrv row_n[13] adc_array_wafflecap_8_8_0[12|24]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3128 adc_array_wafflecap_8_8_0[10|28]/adc_array_circuit_150n_0/vint1 col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3129 adc_array_wafflecap_8_8_0[6|13]/adc_array_circuit_150n_0/vint2 col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3130 adc_array_wafflecap_8_8_0[13|5]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|5]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3131 VDD rowon_n[14] adc_array_wafflecap_8_8_0[13|9]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3132 adc_array_wafflecap_8_8_0[3|25]/adc_array_circuit_150n_0/vdrv row_n[4] adc_array_wafflecap_8_8_0[3|25]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3133 adc_array_wafflecap_8_8_0[3|26]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|26]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3134 adc_array_wafflecap_8_8_0[5|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3135 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X3136 adc_array_wafflecap_8_8_0[6|4]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|4]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3137 adc_array_wafflecap_8_Dummy_2[6]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_2[6]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3138 adc_array_wafflecap_8_8_0[3|7]/adc_array_circuit_150n_0/vint2 rowon_n[4] adc_array_wafflecap_8_8_0[3|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3139 adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3140 adc_array_wafflecap_8_8_0[9|27]/adc_array_circuit_150n_0/vdrv row_n[10] adc_array_wafflecap_8_8_0[9|27]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3141 adc_array_wafflecap_8_8_0[3|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3142 adc_array_wafflecap_8_8_0[2|14]/adc_array_circuit_150n_0/vdrv row_n[3] adc_array_wafflecap_8_8_0[2|14]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3143 adc_array_wafflecap_8_8_0[7|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3144 adc_array_wafflecap_8_8_0[6|13]/adc_array_circuit_150n_0/vdrv row_n[7] adc_array_wafflecap_8_8_0[6|13]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3145 adc_array_wafflecap_8_8_0[5|5]/adc_array_circuit_150n_0/vint2 col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3146 adc_array_wafflecap_8_Dummy_4[27]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[27]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3147 vcm adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|25]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3148 adc_array_wafflecap_8_8_0[12|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3149 adc_array_wafflecap_8_8_0[9|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3150 adc_array_wafflecap_8_Dummy_3[2]/adc_array_circuit_150n_0/vint2 col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3151 vcm adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|30]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3152 adc_array_wafflecap_8_8_0[8|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3153 adc_array_wafflecap_8_Dummy_4[21]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3154 vcm adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|6]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3155 vcm adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|16]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3156 adc_array_wafflecap_8_8_0[11|21]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|21]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3157 adc_array_wafflecap_8_8_0[5|11]/adc_array_circuit_150n_0/vint2 rowon_n[6] adc_array_wafflecap_8_8_0[5|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3158 adc_array_wafflecap_8_Dummy_8[2]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3159 adc_array_wafflecap_8_8_0[1|12]/adc_array_circuit_150n_0/vint2 rowon_n[2] adc_array_wafflecap_8_8_0[1|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3160 adc_array_wafflecap_8_8_0[1|30]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|30]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3161 adc_array_wafflecap_8_8_0[1|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3162 VDD rowon_n[6] adc_array_wafflecap_8_8_0[5|1]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3163 VSS row_n[4] adc_array_wafflecap_8_8_0[3|8]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3164 adc_array_wafflecap_8_8_0[4|19]/adc_array_circuit_150n_0/vint1 col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3165 adc_array_wafflecap_8_8_0[10|8]/adc_array_circuit_150n_0/vint2 rowon_n[11] adc_array_wafflecap_8_8_0[10|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3166 adc_array_wafflecap_8_8_0[10|30]/adc_array_circuit_150n_0/vint2 rowon_n[11] adc_array_wafflecap_8_8_0[10|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3167 adc_array_wafflecap_8_8_0[9|23]/adc_array_circuit_150n_0/vint2 col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3168 VSS row_n[8] adc_array_wafflecap_8_8_0[7|27]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3169 adc_array_wafflecap_8_8_0[5|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3170 adc_array_wafflecap_8_8_0[4|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3171 VDD rowon_n[5] adc_array_wafflecap_8_8_0[4|29]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3172 adc_array_wafflecap_8_8_0[1|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3173 adc_array_wafflecap_8_8_0[4|17]/adc_array_circuit_150n_0/vdrv row_n[5] adc_array_wafflecap_8_8_0[4|17]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3174 adc_array_wafflecap_8_8_0[4|18]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|18]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3175 adc_array_wafflecap_8_8_0[0|19]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|19]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3176 vcm adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|18]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3177 adc_array_wafflecap_8_8_0[7|19]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|19]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3178 VDD rowon_n[2] adc_array_wafflecap_8_8_0[1|12]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3179 adc_array_wafflecap_8_8_0[4|3]/adc_array_circuit_150n_0/vint2 rowon_n[5] adc_array_wafflecap_8_8_0[4|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3180 VDD rowon_n[0] adc_array_wafflecap_8_8_1[26]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3181 adc_array_wafflecap_8_8_0[0|4]/adc_array_circuit_150n_0/vint2 rowon_n[1] adc_array_wafflecap_8_8_0[0|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3182 VDD rowon_n[15] adc_array_wafflecap_8_8_0[14|25]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3183 adc_array_wafflecap_8_8_0[11|22]/adc_array_circuit_150n_0/vint1 col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3184 adc_array_wafflecap_8_8_0[9|0]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|0]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3185 adc_array_wafflecap_8_8_0[9|10]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|10]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3186 VDD rowon_n[10] adc_array_wafflecap_8_8_0[9|26]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3187 adc_array_wafflecap_8_8_0[3|16]/adc_array_circuit_150n_0/vint2 rowon_n[4] adc_array_wafflecap_8_8_0[3|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3188 VSS row_n[0] adc_array_wafflecap_8_8_1[21]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3189 adc_array_wafflecap_8_8_0[7|23]/adc_array_circuit_150n_0/vdrv row_n[8] adc_array_wafflecap_8_8_0[7|23]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3190 adc_array_wafflecap_8_8_0[5|26]/adc_array_circuit_150n_0/vint2 col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3191 adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/vint2 rowon_n[0] adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3192 VSS row_n[3] adc_array_wafflecap_8_8_0[2|0]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3193 adc_array_wafflecap_8_Dummy_4[10]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[10]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3194 VDD rowon_n[9] adc_array_wafflecap_8_8_0[8|8]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3195 VDD rowon_n[9] adc_array_wafflecap_8_8_0[8|30]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3196 VSS row_n[6] adc_array_wafflecap_8_8_0[5|12]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3197 VDD rowon_n[4] adc_array_wafflecap_8_8_0[3|6]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3198 VSS row_n[2] adc_array_wafflecap_8_8_0[1|13]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3199 adc_array_wafflecap_8_Dummy_4[0]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[0]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3200 vcm adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|22]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3201 adc_array_wafflecap_8_8_0[2|24]/adc_array_circuit_150n_0/vint1 col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3202 adc_array_wafflecap_8_8_0[10|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3203 vcm adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|0]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3204 adc_array_wafflecap_8_8_0[5|2]/adc_array_circuit_150n_0/vint1 col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3205 adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3206 adc_array_wafflecap_8_8_0[2|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3207 adc_array_wafflecap_8_8_0[5|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3208 VDD VSS adc_array_wafflecap_8_Dummy_8[2]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3209 adc_array_wafflecap_8_8_0[12|15]/adc_array_circuit_150n_0/vint2 col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3210 VSS row_n[12] adc_array_wafflecap_8_8_0[11|6]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3211 adc_array_wafflecap_8_8_0[7|16]/adc_array_circuit_150n_0/vint2 col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3212 VSS sample_n adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3213 adc_array_wafflecap_8_8_0[0|0]/adc_array_circuit_150n_0/vint1 col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3214 adc_array_wafflecap_8_8_0[12|5]/adc_array_circuit_150n_0/vint2 col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3215 VSS row_n[5] adc_array_wafflecap_8_8_0[4|4]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3216 adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/vint2 col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3217 VSS row_n[1] adc_array_wafflecap_8_8_0[0|5]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3218 adc_array_wafflecap_8_8_0[1|13]/adc_array_circuit_150n_0/vint1 col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3219 vcm adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|11]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3220 vcm VSS adc_array_wafflecap_8_Dummy_4[24]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3221 adc_array_wafflecap_8_8_0[14|14]/adc_array_circuit_150n_0/vint1 col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3222 adc_array_wafflecap_8_8_0[11|11]/adc_array_circuit_150n_0/vdrv row_n[12] adc_array_wafflecap_8_8_0[11|11]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3223 adc_array_wafflecap_8_8_0[9|22]/adc_array_circuit_150n_0/vint2 rowon_n[10] adc_array_wafflecap_8_8_0[9|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3224 adc_array_wafflecap_8_8_0[8|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3225 adc_array_wafflecap_8_8_0[14|4]/adc_array_circuit_150n_0/vint1 col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3226 adc_array_wafflecap_8_8_0[13|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3227 adc_array_wafflecap_8_8_0[11|1]/adc_array_circuit_150n_0/vdrv row_n[12] adc_array_wafflecap_8_8_0[11|1]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3228 adc_array_wafflecap_8_8_0[3|18]/adc_array_circuit_150n_0/vint2 rowon_n[4] adc_array_wafflecap_8_8_0[3|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3229 adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3230 adc_array_wafflecap_8_8_0[10|5]/adc_array_circuit_150n_0/vdrv row_n[11] adc_array_wafflecap_8_8_0[10|5]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3231 adc_array_wafflecap_8_8_0[10|15]/adc_array_circuit_150n_0/vdrv row_n[11] adc_array_wafflecap_8_8_0[10|15]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3232 adc_array_wafflecap_8_8_0[10|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3233 adc_array_wafflecap_8_8_0[14|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3234 adc_array_wafflecap_8_8_0[14|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3235 adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3236 VSS row_n[4] adc_array_wafflecap_8_8_0[3|16]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3237 adc_array_wafflecap_8_Dummy_4[18]/adc_array_circuit_150n_0/vint2 col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3238 vcm adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|14]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3239 adc_array_wafflecap_8_8_0[8|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3240 adc_array_wafflecap_8_Dummy_8[3]/adc_array_circuit_150n_0/vint1 col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3241 adc_array_wafflecap_8_8_0[0|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3242 vcm adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|4]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3243 adc_array_wafflecap_8_8_0[7|27]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|27]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3244 VDD sample adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3245 VDD rowon_n[8] adc_array_wafflecap_8_8_0[7|22]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3246 vcm adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|15]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3247 vcm adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|16]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3248 VSS row_n[15] adc_array_wafflecap_8_8_0[14|20]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3249 VSS row_n[14] adc_array_wafflecap_8_8_0[13|24]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3250 adc_array_wafflecap_8_8_0[10|21]/adc_array_circuit_150n_0/vint2 col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3251 adc_array_wafflecap_8_8_0[6|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3252 adc_array_wafflecap_8_8_1[17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3253 adc_array_wafflecap_8_8_1[7]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[7]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3254 adc_array_wafflecap_8_8_0[1|23]/adc_array_circuit_150n_0/vint2 rowon_n[2] adc_array_wafflecap_8_8_0[1|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3255 adc_array_wafflecap_8_8_0[14|30]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|30]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3256 adc_array_wafflecap_8_8_0[13|17]/adc_array_circuit_150n_0/vdrv row_n[14] adc_array_wafflecap_8_8_0[13|17]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3257 adc_array_wafflecap_8_8_0[11|28]/adc_array_circuit_150n_0/vint2 rowon_n[12] adc_array_wafflecap_8_8_0[11|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3258 vcm adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|17]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3259 adc_array_wafflecap_8_8_0[14|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3260 adc_array_wafflecap_8_8_0[1|2]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|2]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3261 VDD VDD adc_array_wafflecap_8_Dummy_4[24]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3262 adc_array_wafflecap_8_8_0[13|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3263 adc_array_wafflecap_8_8_0[12|20]/adc_array_circuit_150n_0/vint1 col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3264 adc_array_wafflecap_8_8_0[10|8]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|8]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3265 VSS row_n[9] adc_array_wafflecap_8_8_0[8|15]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3266 VDD rowon_n[15] adc_array_wafflecap_8_8_0[14|14]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3267 adc_array_wafflecap_8_8_0[13|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3268 VSS row_n[9] adc_array_wafflecap_8_8_0[8|5]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3269 adc_array_wafflecap_8_8_0[6|6]/adc_array_circuit_150n_0/vint2 col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3270 VDD rowon_n[15] adc_array_wafflecap_8_8_0[14|4]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3271 adc_array_wafflecap_8_8_0[8|21]/adc_array_circuit_150n_0/vdrv row_n[9] adc_array_wafflecap_8_8_0[8|21]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3272 adc_array_wafflecap_8_Dummy_2[5]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_2[5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3273 VDD rowon_n[2] adc_array_wafflecap_8_8_0[1|23]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3274 adc_array_wafflecap_8_8_0[2|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3275 adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3276 adc_array_wafflecap_8_8_0[3|28]/adc_array_circuit_150n_0/vint1 col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3277 adc_array_wafflecap_8_8_0[1|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3278 adc_array_wafflecap_8_8_0[11|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3279 VDD sample adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3280 adc_array_wafflecap_8_8_0[14|9]/adc_array_circuit_150n_0/vint2 col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3281 adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3282 adc_array_wafflecap_8_Dummy_2[4]/adc_array_circuit_150n_0/vint2 col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3283 adc_array_wafflecap_8_8_0[2|20]/adc_array_circuit_150n_0/vint2 col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3284 adc_array_wafflecap_8_8_0[14|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3285 adc_array_wafflecap_8_8_0[13|3]/adc_array_circuit_150n_0/vint2 col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3286 adc_array_wafflecap_8_8_0[13|13]/adc_array_circuit_150n_0/vint2 col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3287 VSS row_n[12] adc_array_wafflecap_8_8_0[11|17]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3288 adc_array_wafflecap_8_8_0[6|6]/adc_array_circuit_150n_0/vdrv row_n[7] adc_array_wafflecap_8_8_0[6|6]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3289 VSS row_n[3] adc_array_wafflecap_8_8_0[2|30]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3290 adc_array_wafflecap_8_8_0[8|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3291 vcm adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|22]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3292 adc_array_wafflecap_8_8_0[0|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3293 vcm adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|30]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3294 adc_array_wafflecap_8_8_0[5|22]/adc_array_circuit_150n_0/vdrv row_n[6] adc_array_wafflecap_8_8_0[5|22]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3295 adc_array_wafflecap_8_8_0[5|23]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|23]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3296 adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/vint1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3297 adc_array_wafflecap_8_8_0[3|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3298 adc_array_wafflecap_8_8_0[1|24]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|24]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3299 adc_array_wafflecap_8_Dummy_4[3]/adc_array_circuit_150n_0/vint1 col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3300 adc_array_wafflecap_8_Dummy_4[13]/adc_array_circuit_150n_0/vint1 col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3301 adc_array_wafflecap_8_8_0[12|9]/adc_array_circuit_150n_0/vdrv row_n[13] adc_array_wafflecap_8_8_0[12|9]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3302 adc_array_wafflecap_8_8_0[9|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3303 adc_array_wafflecap_8_8_0[9|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3304 VSS VSS adc_array_wafflecap_8_Dummy_8[4]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3305 adc_array_wafflecap_8_8_0[8|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3306 adc_array_wafflecap_8_8_0[6|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3307 adc_array_wafflecap_8_8_0[0|20]/adc_array_circuit_150n_0/vdrv row_n[1] adc_array_wafflecap_8_8_0[0|20]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3308 adc_array_wafflecap_8_8_0[12|26]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|26]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3309 adc_array_wafflecap_8_8_0[10|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3310 adc_array_wafflecap_8_8_0[8|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3311 vcm adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[28]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3312 adc_array_wafflecap_8_8_0[0|30]/adc_array_circuit_150n_0/vint1 col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3313 adc_array_wafflecap_8_8_0[0|25]/adc_array_circuit_150n_0/vint2 col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3314 adc_array_wafflecap_8_8_0[1|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3315 adc_array_wafflecap_8_8_0[4|11]/adc_array_circuit_150n_0/vdrv row_n[5] adc_array_wafflecap_8_8_0[4|11]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3316 adc_array_wafflecap_8_8_0[3|3]/adc_array_circuit_150n_0/vint2 col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3317 adc_array_wafflecap_8_8_1[14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_1[14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3318 VSS row_n[10] adc_array_wafflecap_8_8_0[9|19]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3319 vcm adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|19]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3320 adc_array_wafflecap_8_8_0[6|15]/adc_array_circuit_150n_0/vint2 col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3321 vcm adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|10]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3322 adc_array_wafflecap_8_8_1[8]/adc_array_circuit_150n_0/vdrv row_n[0] adc_array_wafflecap_8_8_1[8]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3323 vcm adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|0]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3324 adc_array_wafflecap_8_8_0[8|15]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|15]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3325 adc_array_wafflecap_8_8_0[6|6]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|6]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3326 adc_array_wafflecap_8_8_0[6|26]/adc_array_circuit_150n_0/vint2 rowon_n[7] adc_array_wafflecap_8_8_0[6|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3327 VDD rowon_n[12] adc_array_wafflecap_8_8_0[11|18]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3328 adc_array_wafflecap_8_8_0[8|5]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|5]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3329 adc_array_wafflecap_8_Dummy_3[0]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_3[0]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3330 adc_array_wafflecap_8_8_1[13]/adc_array_circuit_150n_0/vint2 col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3331 adc_array_wafflecap_8_Dummy_4[29]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[29]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3332 adc_array_wafflecap_8_8_0[11|17]/adc_array_circuit_150n_0/vint2 rowon_n[12] adc_array_wafflecap_8_8_0[11|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3333 adc_array_wafflecap_8_8_0[3|27]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|27]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3334 adc_array_wafflecap_8_8_0[3|9]/adc_array_circuit_150n_0/vint2 rowon_n[4] adc_array_wafflecap_8_8_0[3|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3335 adc_array_wafflecap_8_8_0[0|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3336 adc_array_wafflecap_8_8_0[7|19]/adc_array_circuit_150n_0/vint1 col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3337 adc_array_wafflecap_8_8_0[14|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3338 VDD rowon_n[10] adc_array_wafflecap_8_8_0[9|3]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3339 VDD rowon_n[10] adc_array_wafflecap_8_8_0[9|13]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3340 adc_array_wafflecap_8_8_0[6|15]/adc_array_circuit_150n_0/vdrv row_n[7] adc_array_wafflecap_8_8_0[6|15]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3341 VDD VDD adc_array_wafflecap_8_Dummy_4[13]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3342 adc_array_wafflecap_8_8_0[10|19]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|19]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3343 VDD rowon_n[3] adc_array_wafflecap_8_8_0[2|27]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3344 VDD VDD adc_array_wafflecap_8_Dummy_4[3]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3345 VDD rowon_n[7] adc_array_wafflecap_8_8_0[6|26]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3346 VSS row_n[13] adc_array_wafflecap_8_8_0[12|11]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3347 adc_array_wafflecap_8_8_0[9|8]/adc_array_circuit_150n_0/vint2 col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3348 VSS row_n[13] adc_array_wafflecap_8_8_0[12|1]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3349 adc_array_wafflecap_8_Dummy_8[0]/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_8[0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3350 adc_array_wafflecap_8_8_0[2|1]/adc_array_circuit_150n_0/vint2 rowon_n[3] adc_array_wafflecap_8_8_0[2|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3351 adc_array_wafflecap_8_8_0[8|12]/adc_array_circuit_150n_0/vint2 col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3352 adc_array_wafflecap_8_Dummy_8[4]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3353 adc_array_wafflecap_8_8_0[1|14]/adc_array_circuit_150n_0/vint2 rowon_n[2] adc_array_wafflecap_8_8_0[1|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3354 adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3355 adc_array_wafflecap_8_8_0[11|30]/adc_array_circuit_150n_0/vdrv row_n[12] adc_array_wafflecap_8_8_0[11|30]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3356 adc_array_wafflecap_8_8_0[8|2]/adc_array_circuit_150n_0/vint2 col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3357 adc_array_wafflecap_8_8_0[5|13]/adc_array_circuit_150n_0/vint2 rowon_n[6] adc_array_wafflecap_8_8_0[5|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3358 adc_array_wafflecap_8_Dummy_4[20]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3359 adc_array_wafflecap_8_8_0[11|7]/adc_array_circuit_150n_0/vint1 col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3360 adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3361 VDD rowon_n[6] adc_array_wafflecap_8_8_0[5|3]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3362 VSS row_n[4] adc_array_wafflecap_8_8_0[3|10]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3363 vcm adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|20]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3364 vcm adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|20]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3365 adc_array_wafflecap_8_8_0[10|11]/adc_array_circuit_150n_0/vint1 col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3366 adc_array_wafflecap_8_8_0[7|8]/adc_array_circuit_150n_0/vdrv row_n[8] adc_array_wafflecap_8_8_0[7|8]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3367 adc_array_wafflecap_8_8_0[5|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3368 adc_array_wafflecap_8_8_0[4|21]/adc_array_circuit_150n_0/vint1 col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3369 adc_array_wafflecap_8_8_0[4|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3370 adc_array_wafflecap_8_8_0[0|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3371 adc_array_wafflecap_8_8_0[1|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3372 adc_array_wafflecap_8_8_0[10|1]/adc_array_circuit_150n_0/vint1 col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3373 VDD rowon_n[5] adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3374 adc_array_wafflecap_8_8_0[3|0]/adc_array_circuit_150n_0/vint1 col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3375 VDD rowon_n[1] adc_array_wafflecap_8_8_0[0|1]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3376 adc_array_wafflecap_8_8_0[10|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3377 adc_array_wafflecap_8_8_0[6|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3378 adc_array_wafflecap_8_8_1[18]/adc_array_circuit_150n_0/vint1 col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3379 adc_array_wafflecap_8_8_0[10|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3380 VDD rowon_n[0] adc_array_wafflecap_8_8_1[28]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3381 adc_array_wafflecap_8_8_0[0|6]/adc_array_circuit_150n_0/vint2 rowon_n[1] adc_array_wafflecap_8_8_0[0|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3382 VDD rowon_n[2] adc_array_wafflecap_8_8_0[1|14]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3383 adc_array_wafflecap_8_8_0[4|5]/adc_array_circuit_150n_0/vint2 rowon_n[5] adc_array_wafflecap_8_8_0[4|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3384 adc_array_wafflecap_8_8_1[16]/adc_array_circuit_150n_0/vdrv row_n[0] adc_array_wafflecap_8_8_1[16]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3385 adc_array_wafflecap_8_8_0[13|24]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|24]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3386 adc_array_wafflecap_8_8_0[11|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3387 adc_array_wafflecap_8_8_0[5|28]/adc_array_circuit_150n_0/vint2 col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3388 vcm adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|8]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3389 VSS VSS adc_array_wafflecap_8_Dummy_8[1]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3390 VSS row_n[0] adc_array_wafflecap_8_8_1[23]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3391 vcm adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|9]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3392 adc_array_wafflecap_8_8_0[1|29]/adc_array_circuit_150n_0/vint2 col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3393 adc_array_wafflecap_8_8_0[4|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3394 VSS row_n[3] adc_array_wafflecap_8_8_0[2|2]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3395 VSS row_n[6] adc_array_wafflecap_8_8_0[5|14]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3396 VSS row_n[2] adc_array_wafflecap_8_8_0[1|15]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3397 adc_array_wafflecap_8_8_0[13|20]/adc_array_circuit_150n_0/vint2 rowon_n[14] adc_array_wafflecap_8_8_0[13|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3398 VSS row_n[10] adc_array_wafflecap_8_8_0[9|30]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3399 adc_array_wafflecap_8_8_0[12|1]/adc_array_circuit_150n_0/vint2 rowon_n[13] adc_array_wafflecap_8_8_0[12|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3400 adc_array_wafflecap_8_8_0[12|11]/adc_array_circuit_150n_0/vint2 rowon_n[13] adc_array_wafflecap_8_8_0[12|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3401 vcm adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|2]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3402 adc_array_wafflecap_8_8_0[5|4]/adc_array_circuit_150n_0/vint1 col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3403 adc_array_wafflecap_8_8_0[5|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3404 VDD VSS adc_array_wafflecap_8_Dummy_8[4]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3405 vcm VSS adc_array_wafflecap_8_Dummy_4[9]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3406 adc_array_wafflecap_8_8_0[11|15]/adc_array_circuit_150n_0/vint2 rowon_n[12] adc_array_wafflecap_8_8_0[11|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3407 adc_array_wafflecap_8_8_0[10|27]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|27]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3408 adc_array_wafflecap_8_8_0[11|5]/adc_array_circuit_150n_0/vint2 rowon_n[12] adc_array_wafflecap_8_8_0[11|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3409 VDD sample adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3410 adc_array_wafflecap_8_Dummy_3[2]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3411 adc_array_wafflecap_8_8_0[0|2]/adc_array_circuit_150n_0/vint1 col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3412 adc_array_wafflecap_8_8_0[14|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3413 adc_array_wafflecap_8_8_0[14|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3414 VDD rowon_n[12] adc_array_wafflecap_8_8_0[11|29]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3415 adc_array_wafflecap_8_8_0[9|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3416 vcm adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[0]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3417 adc_array_wafflecap_8_8_0[1|29]/adc_array_circuit_150n_0/vdrv row_n[2] adc_array_wafflecap_8_8_0[1|29]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3418 VDD rowon_n[12] adc_array_wafflecap_8_8_0[11|7]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3419 vcm VSS adc_array_wafflecap_8_Dummy_1[5]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3420 adc_array_wafflecap_8_8_0[1|15]/adc_array_circuit_150n_0/vint1 col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3421 vcm adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|13]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3422 VDD rowon_n[11] adc_array_wafflecap_8_8_0[10|11]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3423 adc_array_wafflecap_8_8_0[7|30]/adc_array_circuit_150n_0/vint1 col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3424 VDD rowon_n[11] adc_array_wafflecap_8_8_0[10|1]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3425 adc_array_wafflecap_8_8_0[14|28]/adc_array_circuit_150n_0/vint2 col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3426 adc_array_wafflecap_8_8_0[3|20]/adc_array_circuit_150n_0/vint2 rowon_n[4] adc_array_wafflecap_8_8_0[3|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3427 adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/vint2 VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3428 VSS row_n[14] adc_array_wafflecap_8_8_0[13|9]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3429 adc_array_wafflecap_8_8_0[10|6]/adc_array_circuit_150n_0/vint2 col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3430 adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3431 adc_array_wafflecap_8_8_0[9|19]/adc_array_circuit_150n_0/vint2 col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3432 vcm adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|24]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3433 adc_array_wafflecap_8_Dummy_4[32]/adc_array_circuit_150n_0/vint1 col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3434 adc_array_wafflecap_8_8_0[12|28]/adc_array_circuit_150n_0/vdrv row_n[13] adc_array_wafflecap_8_8_0[12|28]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3435 adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3436 adc_array_wafflecap_8_8_0[6|17]/adc_array_circuit_150n_0/vint2 rowon_n[7] adc_array_wafflecap_8_8_0[6|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3437 adc_array_wafflecap_8_8_0[11|18]/adc_array_circuit_150n_0/vint1 col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3438 adc_array_wafflecap_8_8_0[0|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3439 adc_array_wafflecap_8_Dummy_4[31]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3440 adc_array_wafflecap_8_8_1[9]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[9]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3441 vcm adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|17]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3442 adc_array_wafflecap_8_8_0[1|25]/adc_array_circuit_150n_0/vint2 rowon_n[2] adc_array_wafflecap_8_8_0[1|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3443 adc_array_wafflecap_8_8_0[12|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3444 vcm adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3445 adc_array_wafflecap_8_8_0[8|6]/adc_array_circuit_150n_0/vdrv row_n[9] adc_array_wafflecap_8_8_0[8|6]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3446 adc_array_wafflecap_8_8_0[7|19]/adc_array_circuit_150n_0/vdrv row_n[8] adc_array_wafflecap_8_8_0[7|19]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3447 adc_array_wafflecap_8_8_0[6|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3448 adc_array_wafflecap_8_8_0[11|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3449 adc_array_wafflecap_8_8_0[11|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3450 VDD rowon_n[7] adc_array_wafflecap_8_8_0[6|17]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3451 adc_array_wafflecap_8_8_1[7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_1[7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3452 VSS row_n[1] adc_array_wafflecap_8_8_0[0|28]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3453 VSS row_n[5] adc_array_wafflecap_8_8_0[4|27]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3454 adc_array_wafflecap_8_8_0[6|8]/adc_array_circuit_150n_0/vint2 col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3455 adc_array_wafflecap_8_8_0[14|27]/adc_array_circuit_150n_0/vint2 rowon_n[15] adc_array_wafflecap_8_8_0[14|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3456 adc_array_wafflecap_8_8_0[8|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3457 adc_array_wafflecap_8_8_0[7|0]/adc_array_circuit_150n_0/vint2 rowon_n[8] adc_array_wafflecap_8_8_0[7|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3458 adc_array_wafflecap_8_8_0[7|10]/adc_array_circuit_150n_0/vint2 rowon_n[8] adc_array_wafflecap_8_8_0[7|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3459 VSS row_n[7] adc_array_wafflecap_8_8_0[6|18]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3460 adc_array_wafflecap_8_8_0[3|20]/adc_array_circuit_150n_0/vdrv row_n[4] adc_array_wafflecap_8_8_0[3|20]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3461 adc_array_wafflecap_8_8_0[3|21]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|21]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3462 adc_array_wafflecap_8_1_0/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_1_0/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3463 VDD rowon_n[2] adc_array_wafflecap_8_8_0[1|25]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3464 vcm adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|7]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3465 adc_array_wafflecap_8_8_0[8|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3466 adc_array_wafflecap_8_8_0[5|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3467 adc_array_wafflecap_8_8_0[3|30]/adc_array_circuit_150n_0/vint1 col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3468 adc_array_wafflecap_8_8_0[1|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3469 adc_array_wafflecap_8_8_0[13|9]/adc_array_circuit_150n_0/vint2 rowon_n[14] adc_array_wafflecap_8_8_0[13|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3470 adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/vint2 rowon_n[14] adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3471 adc_array_wafflecap_8_8_0[12|24]/adc_array_circuit_150n_0/vint2 col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3472 VSS row_n[11] adc_array_wafflecap_8_8_0[10|28]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3473 VDD sample_n adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3474 adc_array_wafflecap_8_Dummy_3[3]/adc_array_circuit_150n_0/vint1 col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3475 vcm VSS adc_array_wafflecap_8_Dummy_4[20]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3476 adc_array_wafflecap_8_Dummy_4[15]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3477 adc_array_wafflecap_8_8_0[14|23]/adc_array_circuit_150n_0/vint1 col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3478 adc_array_wafflecap_8_8_0[12|11]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|11]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3479 adc_array_wafflecap_8_8_0[2|9]/adc_array_circuit_150n_0/vdrv row_n[3] adc_array_wafflecap_8_8_0[2|9]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3480 adc_array_wafflecap_8_Dummy_2[6]/adc_array_circuit_150n_0/vint2 col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3481 adc_array_wafflecap_8_8_0[2|22]/adc_array_circuit_150n_0/vint2 col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3482 adc_array_wafflecap_8_Dummy_4[5]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3483 adc_array_wafflecap_8_8_0[12|1]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|1]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3484 VDD rowon_n[13] adc_array_wafflecap_8_8_0[12|27]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3485 adc_array_wafflecap_8_8_0[6|8]/adc_array_circuit_150n_0/vdrv row_n[7] adc_array_wafflecap_8_8_0[6|8]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3486 adc_array_wafflecap_8_8_0[6|18]/adc_array_circuit_150n_0/vint1 col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3487 adc_array_wafflecap_8_8_0[5|0]/adc_array_circuit_150n_0/vint2 col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3488 adc_array_wafflecap_8_8_0[1|1]/adc_array_circuit_150n_0/vint2 col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3489 adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3490 VSS row_n[3] adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3491 adc_array_wafflecap_8_8_0[11|15]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|15]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3492 adc_array_wafflecap_8_8_0[10|24]/adc_array_circuit_150n_0/vdrv row_n[11] adc_array_wafflecap_8_8_0[10|24]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3493 adc_array_wafflecap_8_8_0[9|27]/adc_array_circuit_150n_0/vint2 col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3494 adc_array_wafflecap_8_8_0[8|28]/adc_array_circuit_150n_0/vint1 col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3495 adc_array_wafflecap_8_8_0[11|5]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|5]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3496 adc_array_wafflecap_8_8_0[1|26]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|26]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3497 adc_array_wafflecap_8_Dummy_4[27]/adc_array_circuit_150n_0/vint2 col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3498 vcm adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3499 adc_array_wafflecap_8_8_0[5|25]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|25]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3500 adc_array_wafflecap_8_8_0[3|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3501 adc_array_wafflecap_8_8_0[11|26]/adc_array_circuit_150n_0/vint1 col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3502 adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/vint1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3503 adc_array_wafflecap_8_8_0[0|22]/adc_array_circuit_150n_0/vdrv row_n[1] adc_array_wafflecap_8_8_0[0|22]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3504 vcm adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[30]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3505 adc_array_wafflecap_8_Dummy_0[0]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3506 adc_array_wafflecap_8_8_0[1|7]/adc_array_circuit_150n_0/vint2 rowon_n[2] adc_array_wafflecap_8_8_0[1|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3507 adc_array_wafflecap_8_8_0[1|1]/adc_array_circuit_150n_0/vdrv row_n[2] adc_array_wafflecap_8_8_0[1|1]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3508 adc_array_wafflecap_8_8_0[7|27]/adc_array_circuit_150n_0/vdrv row_n[8] adc_array_wafflecap_8_8_0[7|27]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3509 adc_array_wafflecap_8_8_0[5|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3510 adc_array_wafflecap_8_8_0[1|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3511 adc_array_wafflecap_8_8_0[7|26]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|26]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3512 adc_array_wafflecap_8_8_0[4|13]/adc_array_circuit_150n_0/vdrv row_n[5] adc_array_wafflecap_8_8_0[4|13]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3513 adc_array_wafflecap_8_8_0[4|14]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|14]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3514 adc_array_wafflecap_8_8_0[3|5]/adc_array_circuit_150n_0/vint2 col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3515 adc_array_wafflecap_8_8_0[13|26]/adc_array_circuit_150n_0/vdrv row_n[14] adc_array_wafflecap_8_8_0[13|26]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3516 vcm adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|25]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3517 adc_array_wafflecap_8_8_0[10|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3518 adc_array_wafflecap_8_8_1[10]/adc_array_circuit_150n_0/vdrv row_n[0] adc_array_wafflecap_8_8_1[10]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3519 adc_array_wafflecap_8_8_0[6|28]/adc_array_circuit_150n_0/vint2 rowon_n[7] adc_array_wafflecap_8_8_0[6|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3520 VDD rowon_n[2] adc_array_wafflecap_8_8_0[1|7]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3521 adc_array_wafflecap_8_8_0[13|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3522 vcm adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|6]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3523 vcm adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|16]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3524 adc_array_wafflecap_8_8_0[3|11]/adc_array_circuit_150n_0/vint2 rowon_n[4] adc_array_wafflecap_8_8_0[3|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3525 adc_array_wafflecap_8_8_1[26]/adc_array_circuit_150n_0/vint2 rowon_n[0] adc_array_wafflecap_8_8_1[26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3526 vcm VSS adc_array_wafflecap_8_Dummy_4[28]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3527 adc_array_wafflecap_8_8_0[14|25]/adc_array_circuit_150n_0/vint2 rowon_n[15] adc_array_wafflecap_8_8_0[14|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3528 adc_array_wafflecap_8_8_0[9|26]/adc_array_circuit_150n_0/vint2 rowon_n[10] adc_array_wafflecap_8_8_0[9|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3529 VSS row_n[6] adc_array_wafflecap_8_8_0[5|7]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3530 VDD rowon_n[4] adc_array_wafflecap_8_8_0[3|1]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3531 VSS row_n[2] adc_array_wafflecap_8_8_0[1|8]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3532 adc_array_wafflecap_8_8_0[2|19]/adc_array_circuit_150n_0/vint1 col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3533 adc_array_wafflecap_8_8_0[8|8]/adc_array_circuit_150n_0/vint2 rowon_n[9] adc_array_wafflecap_8_8_0[8|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3534 adc_array_wafflecap_8_8_0[8|30]/adc_array_circuit_150n_0/vint2 rowon_n[9] adc_array_wafflecap_8_8_0[8|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3535 adc_array_wafflecap_8_8_0[7|23]/adc_array_circuit_150n_0/vint2 col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3536 VDD rowon_n[7] adc_array_wafflecap_8_8_0[6|28]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3537 adc_array_wafflecap_8_8_0[3|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3538 adc_array_wafflecap_8_8_0[2|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3539 VDD rowon_n[3] adc_array_wafflecap_8_8_0[2|29]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3540 adc_array_wafflecap_8_8_0[14|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3541 adc_array_wafflecap_8_8_0[2|17]/adc_array_circuit_150n_0/vdrv row_n[3] adc_array_wafflecap_8_8_0[2|17]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3542 adc_array_wafflecap_8_8_0[2|18]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|18]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3543 VDD VSS adc_array_wafflecap_8_Dummy_0[0]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3544 adc_array_wafflecap_8_Dummy_2[2]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_2[2]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3545 vcm adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|18]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3546 adc_array_wafflecap_8_Dummy_8[2]/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_8[2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3547 adc_array_wafflecap_8_8_0[2|3]/adc_array_circuit_150n_0/vint2 rowon_n[3] adc_array_wafflecap_8_8_0[2|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3548 VDD rowon_n[13] adc_array_wafflecap_8_8_0[12|25]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3549 adc_array_wafflecap_8_8_0[9|22]/adc_array_circuit_150n_0/vint1 col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3550 VDD rowon_n[8] adc_array_wafflecap_8_8_0[7|26]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3551 adc_array_wafflecap_8_8_0[5|15]/adc_array_circuit_150n_0/vint2 rowon_n[6] adc_array_wafflecap_8_8_0[5|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3552 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X3553 adc_array_wafflecap_8_8_0[1|16]/adc_array_circuit_150n_0/vint2 rowon_n[2] adc_array_wafflecap_8_8_0[1|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3554 VDD rowon_n[12] adc_array_wafflecap_8_8_0[11|6]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3555 VDD rowon_n[12] adc_array_wafflecap_8_8_0[11|16]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3556 adc_array_wafflecap_8_8_0[3|26]/adc_array_circuit_150n_0/vint2 col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3557 VSS row_n[1] adc_array_wafflecap_8_8_0[0|0]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3558 adc_array_wafflecap_8_8_0[1|8]/adc_array_circuit_150n_0/vint1 col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3559 adc_array_wafflecap_8_8_0[13|9]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|9]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3560 VDD rowon_n[6] adc_array_wafflecap_8_8_0[5|5]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3561 VSS row_n[4] adc_array_wafflecap_8_8_0[3|12]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3562 VDD sample_n adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3563 vcm adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|22]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3564 adc_array_wafflecap_8_8_0[8|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3565 adc_array_wafflecap_8_8_0[6|29]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|29]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3566 adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3567 adc_array_wafflecap_8_8_0[4|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3568 adc_array_wafflecap_8_8_0[3|2]/adc_array_circuit_150n_0/vint1 col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3569 adc_array_wafflecap_8_8_0[0|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3570 adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3571 VSS row_n[15] adc_array_wafflecap_8_8_0[14|14]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3572 adc_array_wafflecap_8_8_0[3|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3573 VDD rowon_n[1] adc_array_wafflecap_8_8_0[0|3]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3574 VSS row_n[15] adc_array_wafflecap_8_8_0[14|4]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3575 adc_array_wafflecap_8_8_0[6|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3576 adc_array_wafflecap_8_8_1[20]/adc_array_circuit_150n_0/vint1 col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3577 adc_array_wafflecap_8_8_0[14|20]/adc_array_circuit_150n_0/vdrv row_n[15] adc_array_wafflecap_8_8_0[14|20]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3578 adc_array_wafflecap_8_8_0[10|15]/adc_array_circuit_150n_0/vint2 col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3579 adc_array_wafflecap_8_Dummy_0[1]/adc_array_circuit_150n_0/vint1 col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3580 VDD rowon_n[0] adc_array_wafflecap_8_8_1[30]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3581 VDD rowon_n[2] adc_array_wafflecap_8_8_0[1|16]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3582 adc_array_wafflecap_8_8_0[10|5]/adc_array_circuit_150n_0/vint2 col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3583 adc_array_wafflecap_8_8_0[5|30]/adc_array_circuit_150n_0/vint2 col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3584 vcm adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|10]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3585 VSS VSS adc_array_wafflecap_8_Dummy_8[3]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3586 vcm adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|11]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3587 adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/vint2 col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3588 VSS row_n[3] adc_array_wafflecap_8_8_0[2|4]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3589 vcm adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|23]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3590 adc_array_wafflecap_8_8_0[12|14]/adc_array_circuit_150n_0/vint1 col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3591 adc_array_wafflecap_8_8_0[9|11]/adc_array_circuit_150n_0/vdrv row_n[10] adc_array_wafflecap_8_8_0[9|11]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3592 adc_array_wafflecap_8_8_0[8|24]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|24]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3593 adc_array_wafflecap_8_8_0[7|22]/adc_array_circuit_150n_0/vint2 rowon_n[8] adc_array_wafflecap_8_8_0[7|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3594 adc_array_wafflecap_8_8_0[12|4]/adc_array_circuit_150n_0/vint1 col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3595 adc_array_wafflecap_8_8_0[11|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3596 adc_array_wafflecap_8_8_0[9|1]/adc_array_circuit_150n_0/vdrv row_n[10] adc_array_wafflecap_8_8_0[9|1]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3597 adc_array_wafflecap_8_8_0[1|18]/adc_array_circuit_150n_0/vint2 rowon_n[2] adc_array_wafflecap_8_8_0[1|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3598 adc_array_wafflecap_8_8_0[8|5]/adc_array_circuit_150n_0/vdrv row_n[9] adc_array_wafflecap_8_8_0[8|5]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3599 adc_array_wafflecap_8_8_0[8|15]/adc_array_circuit_150n_0/vdrv row_n[9] adc_array_wafflecap_8_8_0[8|15]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3600 VSS row_n[2] adc_array_wafflecap_8_8_0[1|16]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3601 adc_array_wafflecap_8_8_0[12|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3602 adc_array_wafflecap_8_8_0[12|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3603 adc_array_wafflecap_8_8_0[13|17]/adc_array_circuit_150n_0/vint2 col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3604 vcm adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|14]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3605 adc_array_wafflecap_8_8_0[4|19]/adc_array_circuit_150n_0/vint2 col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3606 adc_array_wafflecap_8_Dummy_3[4]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3607 adc_array_wafflecap_8_8_0[0|4]/adc_array_circuit_150n_0/vint1 col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3608 adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/vdrv row_n[2] adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3609 vcm adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|4]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3610 vcm VSS adc_array_wafflecap_8_2_0/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3611 vcm adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[2]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3612 vcm adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|15]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3613 VDD rowon_n[2] adc_array_wafflecap_8_8_0[1|18]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3614 adc_array_wafflecap_8_Dummy_4[17]/adc_array_circuit_150n_0/vint1 col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3615 adc_array_wafflecap_8_Dummy_4[24]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3616 VSS row_n[13] adc_array_wafflecap_8_8_0[12|20]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3617 adc_array_wafflecap_8_8_0[14|4]/adc_array_circuit_150n_0/vint2 rowon_n[15] adc_array_wafflecap_8_8_0[14|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3618 adc_array_wafflecap_8_8_0[14|14]/adc_array_circuit_150n_0/vint2 rowon_n[15] adc_array_wafflecap_8_8_0[14|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3619 VSS row_n[12] adc_array_wafflecap_8_8_0[11|24]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3620 adc_array_wafflecap_8_8_0[8|21]/adc_array_circuit_150n_0/vint2 col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3621 adc_array_wafflecap_8_8_0[1|16]/adc_array_circuit_150n_0/vint1 col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3622 adc_array_wafflecap_8_8_0[12|30]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|30]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3623 VDD rowon_n[15] adc_array_wafflecap_8_8_0[14|19]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3624 adc_array_wafflecap_8_8_0[12|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3625 VDD rowon_n[14] adc_array_wafflecap_8_8_0[13|23]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3626 adc_array_wafflecap_8_8_0[11|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3627 adc_array_wafflecap_8_8_0[10|20]/adc_array_circuit_150n_0/vint1 col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3628 vcm adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|26]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3629 VDD rowon_n[13] adc_array_wafflecap_8_8_0[12|14]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3630 adc_array_wafflecap_8_8_0[11|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3631 VDD rowon_n[13] adc_array_wafflecap_8_8_0[12|4]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3632 adc_array_wafflecap_8_8_0[0|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3633 adc_array_wafflecap_8_8_0[5|27]/adc_array_circuit_150n_0/vint1 col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3634 adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3635 adc_array_wafflecap_8_8_0[5|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3636 adc_array_wafflecap_8_8_1[11]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[11]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3637 VDD sample adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3638 adc_array_wafflecap_8_8_0[6|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3639 VSS VDD adc_array_wafflecap_8_Dummy_4[13]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3640 adc_array_wafflecap_8_8_0[12|9]/adc_array_circuit_150n_0/vint2 col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3641 VSS VDD adc_array_wafflecap_8_Dummy_4[3]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3642 adc_array_wafflecap_8_8_0[7|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3643 adc_array_wafflecap_8_8_0[0|20]/adc_array_circuit_150n_0/vint2 col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3644 adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/vdrv row_n[15] adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3645 adc_array_wafflecap_8_8_0[12|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3646 adc_array_wafflecap_8_8_0[11|3]/adc_array_circuit_150n_0/vint2 col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3647 adc_array_wafflecap_8_8_0[11|13]/adc_array_circuit_150n_0/vint2 col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3648 adc_array_wafflecap_8_8_0[4|6]/adc_array_circuit_150n_0/vdrv row_n[5] adc_array_wafflecap_8_8_0[4|6]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3649 VSS row_n[5] adc_array_wafflecap_8_8_0[4|29]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3650 adc_array_wafflecap_8_8_1[9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_1[9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3651 VSS row_n[1] adc_array_wafflecap_8_8_0[0|30]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3652 adc_array_wafflecap_8_8_0[6|22]/adc_array_circuit_150n_0/vint2 rowon_n[7] adc_array_wafflecap_8_8_0[6|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3653 adc_array_wafflecap_8_8_0[14|8]/adc_array_circuit_150n_0/vint1 col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3654 vcm adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|22]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3655 adc_array_wafflecap_8_8_0[6|10]/adc_array_circuit_150n_0/vint2 col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3656 adc_array_wafflecap_8_8_0[3|22]/adc_array_circuit_150n_0/vdrv row_n[4] adc_array_wafflecap_8_8_0[3|22]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3657 adc_array_wafflecap_8_Dummy_3[1]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_3[1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3658 adc_array_wafflecap_8_8_0[3|23]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|23]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3659 adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/vint1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3660 adc_array_wafflecap_8_8_0[1|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3661 adc_array_wafflecap_8_8_0[14|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3662 adc_array_wafflecap_8_8_0[13|2]/adc_array_circuit_150n_0/vint1 col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3663 adc_array_wafflecap_8_8_0[13|12]/adc_array_circuit_150n_0/vint1 col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3664 adc_array_wafflecap_8_8_0[10|9]/adc_array_circuit_150n_0/vdrv row_n[11] adc_array_wafflecap_8_8_0[10|9]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3665 adc_array_wafflecap_8_8_0[7|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3666 adc_array_wafflecap_8_8_0[7|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3667 adc_array_wafflecap_8_8_0[6|1]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|1]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3668 adc_array_wafflecap_8_Dummy_2[3]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_2[3]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3669 adc_array_wafflecap_8_8_1[8]/adc_array_circuit_150n_0/vint2 col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3670 adc_array_wafflecap_8_8_0[10|26]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|26]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3671 adc_array_wafflecap_8_Dummy_3[5]/adc_array_circuit_150n_0/vint1 col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3672 VDD rowon_n[7] adc_array_wafflecap_8_8_0[6|22]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3673 adc_array_wafflecap_8_Dummy_3[0]/adc_array_circuit_150n_0/vint2 col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3674 adc_array_wafflecap_8_8_0[6|10]/adc_array_circuit_150n_0/vdrv row_n[7] adc_array_wafflecap_8_8_0[6|10]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3675 adc_array_wafflecap_8_8_0[2|11]/adc_array_circuit_150n_0/vdrv row_n[3] adc_array_wafflecap_8_8_0[2|11]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3676 adc_array_wafflecap_8_8_0[1|3]/adc_array_circuit_150n_0/vint2 col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3677 VSS row_n[8] adc_array_wafflecap_8_8_0[7|19]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3678 adc_array_wafflecap_8_8_0[5|2]/adc_array_circuit_150n_0/vint2 col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3679 vcm adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|19]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3680 adc_array_wafflecap_8_8_0[9|3]/adc_array_circuit_150n_0/vint2 rowon_n[10] adc_array_wafflecap_8_8_0[9|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3681 adc_array_wafflecap_8_8_0[9|13]/adc_array_circuit_150n_0/vint2 rowon_n[10] adc_array_wafflecap_8_8_0[9|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3682 vcm adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|10]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3683 adc_array_wafflecap_8_8_0[7|1]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|1]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3684 adc_array_wafflecap_8_8_0[7|11]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|11]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3685 adc_array_wafflecap_8_Dummy_4[13]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3686 vcm adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|0]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3687 adc_array_wafflecap_8_Dummy_4[3]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3688 VDD rowon_n[10] adc_array_wafflecap_8_8_0[9|18]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3689 adc_array_wafflecap_8_8_0[13|28]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|28]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3690 adc_array_wafflecap_8_1_1/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3691 adc_array_wafflecap_8_8_0[1|9]/adc_array_circuit_150n_0/vint2 rowon_n[2] adc_array_wafflecap_8_8_0[1|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3692 adc_array_wafflecap_8_8_0[1|27]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|27]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3693 adc_array_wafflecap_8_8_0[5|8]/adc_array_circuit_150n_0/vint2 rowon_n[6] adc_array_wafflecap_8_8_0[5|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3694 adc_array_wafflecap_8_8_0[5|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3695 adc_array_wafflecap_8_8_0[1|3]/adc_array_circuit_150n_0/vdrv row_n[2] adc_array_wafflecap_8_8_0[1|3]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3696 adc_array_wafflecap_8_8_0[14|4]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|4]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3697 adc_array_wafflecap_8_8_0[14|14]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|14]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3698 adc_array_wafflecap_8_8_0[12|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3699 VDD rowon_n[8] adc_array_wafflecap_8_8_0[7|3]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3700 VDD rowon_n[8] adc_array_wafflecap_8_8_0[7|13]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3701 adc_array_wafflecap_8_8_0[4|15]/adc_array_circuit_150n_0/vdrv row_n[5] adc_array_wafflecap_8_8_0[4|15]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3702 adc_array_wafflecap_8_8_0[4|16]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|16]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3703 VDD rowon_n[14] adc_array_wafflecap_8_8_0[13|12]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3704 VDD rowon_n[14] adc_array_wafflecap_8_8_0[13|2]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3705 VDD rowon_n[5] adc_array_wafflecap_8_8_0[4|26]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3706 adc_array_wafflecap_8_8_1[12]/adc_array_circuit_150n_0/vdrv row_n[0] adc_array_wafflecap_8_8_1[12]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3707 VSS row_n[11] adc_array_wafflecap_8_8_0[10|11]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3708 adc_array_wafflecap_8_8_0[7|8]/adc_array_circuit_150n_0/vint2 col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3709 adc_array_wafflecap_8_8_0[6|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3710 adc_array_wafflecap_8_8_0[6|30]/adc_array_circuit_150n_0/vint2 rowon_n[7] adc_array_wafflecap_8_8_0[6|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3711 adc_array_wafflecap_8_8_0[5|24]/adc_array_circuit_150n_0/vint2 col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3712 VSS row_n[11] adc_array_wafflecap_8_8_0[10|1]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3713 adc_array_wafflecap_8_8_0[0|1]/adc_array_circuit_150n_0/vint2 rowon_n[1] adc_array_wafflecap_8_8_0[0|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3714 VDD rowon_n[2] adc_array_wafflecap_8_8_0[1|9]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3715 adc_array_wafflecap_8_8_0[4|0]/adc_array_circuit_150n_0/vint2 rowon_n[5] adc_array_wafflecap_8_8_0[4|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3716 adc_array_wafflecap_8_8_0[9|30]/adc_array_circuit_150n_0/vdrv row_n[10] adc_array_wafflecap_8_8_0[9|30]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3717 adc_array_wafflecap_8_8_0[3|13]/adc_array_circuit_150n_0/vint2 rowon_n[4] adc_array_wafflecap_8_8_0[3|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3718 adc_array_wafflecap_8_8_1[28]/adc_array_circuit_150n_0/vint2 rowon_n[0] adc_array_wafflecap_8_8_1[28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3719 VSS row_n[0] adc_array_wafflecap_8_8_1[18]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3720 adc_array_wafflecap_8_8_0[13|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3721 adc_array_wafflecap_8_8_0[9|7]/adc_array_circuit_150n_0/vint1 col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3722 adc_array_wafflecap_8_8_0[8|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3723 adc_array_wafflecap_8_8_1[16]/adc_array_circuit_150n_0/vint2 col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3724 adc_array_wafflecap_8_Dummy_4[30]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[30]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3725 adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3726 vcm adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|29]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3727 VSS row_n[6] adc_array_wafflecap_8_8_0[5|9]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3728 VDD rowon_n[4] adc_array_wafflecap_8_8_0[3|3]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3729 VSS row_n[2] adc_array_wafflecap_8_8_0[1|10]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3730 adc_array_wafflecap_8_8_0[9|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3731 adc_array_wafflecap_8_8_0[8|11]/adc_array_circuit_150n_0/vint1 col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3732 adc_array_wafflecap_8_8_0[3|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3733 adc_array_wafflecap_8_8_0[2|21]/adc_array_circuit_150n_0/vint1 col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3734 adc_array_wafflecap_8_8_0[2|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3735 adc_array_wafflecap_8_Dummy_2[6]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3736 adc_array_wafflecap_8_8_0[8|1]/adc_array_circuit_150n_0/vint1 col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3737 VDD rowon_n[7] adc_array_wafflecap_8_8_0[6|30]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3738 adc_array_wafflecap_8_8_0[5|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3739 VDD rowon_n[3] adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3740 VDD en_C0_n adc_array_wafflecap_8_1_1/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3741 adc_array_wafflecap_8_8_0[8|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3742 adc_array_wafflecap_8_Dummy_4[24]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3743 adc_array_wafflecap_8_8_0[8|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3744 adc_array_wafflecap_8_Dummy_8[4]/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_8[4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3745 adc_array_wafflecap_8_8_0[11|24]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|24]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3746 adc_array_wafflecap_8_8_0[2|5]/adc_array_circuit_150n_0/vint2 rowon_n[3] adc_array_wafflecap_8_8_0[2|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3747 adc_array_wafflecap_8_8_0[3|28]/adc_array_circuit_150n_0/vint2 col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3748 vcm VSS adc_array_wafflecap_8_Dummy_1[0]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3749 adc_array_wafflecap_8_8_0[1|10]/adc_array_circuit_150n_0/vint1 col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3750 vcm adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|8]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3751 VSS row_n[5] adc_array_wafflecap_8_8_0[4|1]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3752 VSS row_n[1] adc_array_wafflecap_8_8_0[0|2]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3753 adc_array_wafflecap_8_8_0[2|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3754 adc_array_wafflecap_8_8_0[11|20]/adc_array_circuit_150n_0/vint2 rowon_n[12] adc_array_wafflecap_8_8_0[11|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3755 VSS row_n[4] adc_array_wafflecap_8_8_0[3|14]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3756 adc_array_wafflecap_8_8_0[14|22]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|22]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3757 adc_array_wafflecap_8_8_0[10|11]/adc_array_circuit_150n_0/vint2 rowon_n[11] adc_array_wafflecap_8_8_0[10|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3758 VSS row_n[8] adc_array_wafflecap_8_8_0[7|30]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3759 adc_array_wafflecap_8_8_0[10|1]/adc_array_circuit_150n_0/vint2 rowon_n[11] adc_array_wafflecap_8_8_0[10|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3760 adc_array_wafflecap_8_8_0[8|9]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|9]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3761 adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3762 adc_array_wafflecap_8_8_0[4|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3763 adc_array_wafflecap_8_8_0[3|4]/adc_array_circuit_150n_0/vint1 col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3764 adc_array_wafflecap_8_8_0[3|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3765 VDD rowon_n[1] adc_array_wafflecap_8_8_0[0|5]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3766 vcm adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|8]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3767 VDD sample_n adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3768 adc_array_wafflecap_8_Dummy_8[0]/adc_array_circuit_150n_0/vint1 col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3769 adc_array_wafflecap_8_8_0[12|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3770 adc_array_wafflecap_8_8_0[12|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3771 adc_array_wafflecap_8_8_0[11|25]/adc_array_circuit_150n_0/vint1 col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3772 adc_array_wafflecap_8_8_0[9|3]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|3]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3773 adc_array_wafflecap_8_8_0[9|13]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|13]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3774 VDD rowon_n[10] adc_array_wafflecap_8_8_0[9|29]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3775 VDD rowon_n[10] adc_array_wafflecap_8_8_0[9|7]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3776 vcm adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|12]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3777 vcm adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|13]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3778 VDD rowon_n[9] adc_array_wafflecap_8_8_0[8|11]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3779 adc_array_wafflecap_8_8_0[5|19]/adc_array_circuit_150n_0/vdrv row_n[6] adc_array_wafflecap_8_8_0[5|19]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3780 adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/vint2 VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3781 VSS sample adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3782 VDD rowon_n[9] adc_array_wafflecap_8_8_0[8|1]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3783 VSS VDD adc_array_wafflecap_8_Dummy_4[32]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3784 adc_array_wafflecap_8_8_0[12|28]/adc_array_circuit_150n_0/vint2 col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3785 adc_array_wafflecap_8_8_0[1|20]/adc_array_circuit_150n_0/vint2 rowon_n[2] adc_array_wafflecap_8_8_0[1|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3786 adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/vint2 VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3787 VSS row_n[5] adc_array_wafflecap_8_8_0[4|23]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3788 VSS row_n[12] adc_array_wafflecap_8_8_0[11|9]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3789 adc_array_wafflecap_8_8_0[8|6]/adc_array_circuit_150n_0/vint2 col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3790 adc_array_wafflecap_8_8_0[7|19]/adc_array_circuit_150n_0/vint2 col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3791 adc_array_wafflecap_8_8_0[14|27]/adc_array_circuit_150n_0/vint1 col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3792 vcm adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[4]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3793 adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/vint1 col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3794 adc_array_wafflecap_8_8_0[10|28]/adc_array_circuit_150n_0/vdrv row_n[11] adc_array_wafflecap_8_8_0[10|28]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3795 adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3796 vcm VSS adc_array_wafflecap_8_Dummy_4[27]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3797 adc_array_wafflecap_8_8_0[11|14]/adc_array_circuit_150n_0/vdrv row_n[12] adc_array_wafflecap_8_8_0[11|14]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3798 adc_array_wafflecap_8_8_0[9|18]/adc_array_circuit_150n_0/vint1 col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3799 adc_array_wafflecap_8_Dummy_2[2]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_2[2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3800 VDD rowon_n[2] adc_array_wafflecap_8_8_0[1|20]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3801 adc_array_wafflecap_8_8_0[13|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3802 adc_array_wafflecap_8_8_0[11|4]/adc_array_circuit_150n_0/vdrv row_n[12] adc_array_wafflecap_8_8_0[11|4]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3803 vcm VSS adc_array_wafflecap_8_Dummy_2[0]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3804 adc_array_wafflecap_8_8_0[10|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3805 VDD rowon_n[5] adc_array_wafflecap_8_8_0[4|17]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3806 adc_array_wafflecap_8_8_0[7|30]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|30]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3807 VSS VSS adc_array_wafflecap_8_Dummy_3[3]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3808 VSS row_n[3] adc_array_wafflecap_8_8_0[2|27]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3809 adc_array_wafflecap_8_8_0[7|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3810 adc_array_wafflecap_8_8_0[14|16]/adc_array_circuit_150n_0/vdrv row_n[15] adc_array_wafflecap_8_8_0[14|16]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3811 VSS row_n[15] adc_array_wafflecap_8_8_0[14|23]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3812 adc_array_wafflecap_8_8_0[12|27]/adc_array_circuit_150n_0/vint2 rowon_n[13] adc_array_wafflecap_8_8_0[12|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3813 adc_array_wafflecap_8_8_0[1|21]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|21]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3814 adc_array_wafflecap_8_Dummy_4[21]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[21]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3815 adc_array_wafflecap_8_8_0[10|24]/adc_array_circuit_150n_0/vint2 col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3816 vcm adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|7]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3817 vcm adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|27]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3818 adc_array_wafflecap_8_8_0[5|20]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|20]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3819 adc_array_wafflecap_8_8_0[5|29]/adc_array_circuit_150n_0/vint1 col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3820 adc_array_wafflecap_8_8_0[5|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3821 adc_array_wafflecap_8_8_0[3|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3822 adc_array_wafflecap_8_8_0[11|9]/adc_array_circuit_150n_0/vint2 rowon_n[12] adc_array_wafflecap_8_8_0[11|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3823 adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/vint2 rowon_n[12] adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3824 VSS row_n[9] adc_array_wafflecap_8_8_0[8|28]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3825 adc_array_wafflecap_8_8_0[0|27]/adc_array_circuit_150n_0/vint1 col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3826 adc_array_wafflecap_8_8_0[14|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3827 adc_array_wafflecap_8_8_0[14|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3828 vcm adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|19]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3829 adc_array_wafflecap_8_8_0[13|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3830 adc_array_wafflecap_8_8_0[12|23]/adc_array_circuit_150n_0/vint1 col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3831 adc_array_wafflecap_8_8_0[10|11]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|11]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3832 adc_array_wafflecap_8_8_1[11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_1[11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3833 adc_array_wafflecap_8_8_0[0|22]/adc_array_circuit_150n_0/vint2 col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3834 adc_array_wafflecap_8_8_0[13|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3835 adc_array_wafflecap_8_8_0[10|1]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|1]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3836 VDD rowon_n[11] adc_array_wafflecap_8_8_0[10|27]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3837 adc_array_wafflecap_8_8_0[6|24]/adc_array_circuit_150n_0/vint2 rowon_n[7] adc_array_wafflecap_8_8_0[6|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3838 adc_array_wafflecap_8_8_0[4|8]/adc_array_circuit_150n_0/vdrv row_n[5] adc_array_wafflecap_8_8_0[4|8]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3839 adc_array_wafflecap_8_8_0[4|9]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|9]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3840 adc_array_wafflecap_8_8_0[4|18]/adc_array_circuit_150n_0/vint1 col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3841 VSS row_n[5] adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3842 adc_array_wafflecap_8_8_0[3|0]/adc_array_circuit_150n_0/vint2 col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3843 adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3844 VSS row_n[1] adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3845 adc_array_wafflecap_8_8_0[8|24]/adc_array_circuit_150n_0/vdrv row_n[9] adc_array_wafflecap_8_8_0[8|24]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3846 adc_array_wafflecap_8_8_0[7|27]/adc_array_circuit_150n_0/vint2 col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3847 adc_array_wafflecap_8_8_0[6|12]/adc_array_circuit_150n_0/vint2 col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3848 adc_array_wafflecap_8_8_1[5]/adc_array_circuit_150n_0/vdrv row_n[0] adc_array_wafflecap_8_8_1[5]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3849 adc_array_wafflecap_8_8_0[13|26]/adc_array_circuit_150n_0/vint2 col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3850 adc_array_wafflecap_8_8_0[3|25]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|25]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3851 adc_array_wafflecap_8_8_0[1|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3852 adc_array_wafflecap_8_8_0[6|3]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|3]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3853 adc_array_wafflecap_8_8_1[10]/adc_array_circuit_150n_0/vint2 col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3854 adc_array_wafflecap_8_8_0[11|22]/adc_array_circuit_150n_0/vdrv row_n[12] adc_array_wafflecap_8_8_0[11|22]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3855 adc_array_wafflecap_8_8_0[9|26]/adc_array_circuit_150n_0/vint1 col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3856 adc_array_wafflecap_8_Dummy_2[5]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_2[5]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3857 adc_array_wafflecap_8_Dummy_6/adc_array_circuit_150n_0/vint1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3858 adc_array_wafflecap_8_8_0[14|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3859 VDD rowon_n[7] adc_array_wafflecap_8_8_0[6|24]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3860 adc_array_wafflecap_8_8_0[3|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3861 adc_array_wafflecap_8_8_0[6|12]/adc_array_circuit_150n_0/vdrv row_n[7] adc_array_wafflecap_8_8_0[6|12]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3862 adc_array_wafflecap_8_8_0[2|13]/adc_array_circuit_150n_0/vdrv row_n[3] adc_array_wafflecap_8_8_0[2|13]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3863 adc_array_wafflecap_8_8_0[2|14]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|14]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3864 adc_array_wafflecap_8_8_0[1|5]/adc_array_circuit_150n_0/vint2 col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3865 vcm adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|25]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3866 adc_array_wafflecap_8_8_0[8|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3867 adc_array_wafflecap_8_Dummy_4[6]/adc_array_circuit_150n_0/vint1 col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3868 adc_array_wafflecap_8_Dummy_4[16]/adc_array_circuit_150n_0/vint1 col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3869 adc_array_wafflecap_8_8_0[9|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3870 adc_array_wafflecap_8_8_0[9|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3871 adc_array_wafflecap_8_8_0[11|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3872 adc_array_wafflecap_8_Dummy_0[0]/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_0[0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3873 adc_array_wafflecap_8_8_0[5|10]/adc_array_circuit_150n_0/vint2 rowon_n[6] adc_array_wafflecap_8_8_0[5|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3874 adc_array_wafflecap_8_8_0[1|11]/adc_array_circuit_150n_0/vint2 rowon_n[2] adc_array_wafflecap_8_8_0[1|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3875 adc_array_wafflecap_8_8_0[1|5]/adc_array_circuit_150n_0/vdrv row_n[2] adc_array_wafflecap_8_8_0[1|5]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3876 vcm adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|27]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3877 adc_array_wafflecap_8_8_0[12|25]/adc_array_circuit_150n_0/vint2 rowon_n[13] adc_array_wafflecap_8_8_0[12|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3878 VSS row_n[10] adc_array_wafflecap_8_8_0[9|22]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3879 adc_array_wafflecap_8_8_0[8|28]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|28]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3880 adc_array_wafflecap_8_8_0[7|26]/adc_array_circuit_150n_0/vint2 rowon_n[8] adc_array_wafflecap_8_8_0[7|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3881 VDD rowon_n[6] adc_array_wafflecap_8_8_0[5|0]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3882 VSS row_n[4] adc_array_wafflecap_8_8_0[3|7]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3883 VSS sample adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3884 vcm adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|13]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3885 adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3886 adc_array_wafflecap_8_8_0[7|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3887 adc_array_wafflecap_8_8_0[4|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3888 VDD rowon_n[5] adc_array_wafflecap_8_8_0[4|28]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3889 adc_array_wafflecap_8_8_1[14]/adc_array_circuit_150n_0/vdrv row_n[0] adc_array_wafflecap_8_8_1[14]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3890 adc_array_wafflecap_8_8_0[0|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3891 adc_array_wafflecap_8_8_0[1|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3892 vcm adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|3]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3893 adc_array_wafflecap_8_8_0[12|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3894 adc_array_wafflecap_8_8_0[0|18]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|18]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3895 VDD rowon_n[12] adc_array_wafflecap_8_8_0[11|21]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3896 adc_array_wafflecap_8_8_0[9|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3897 vcm adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|18]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3898 adc_array_wafflecap_8_8_0[6|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3899 adc_array_wafflecap_8_8_0[4|17]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|17]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3900 adc_array_wafflecap_8_Dummy_4[32]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[32]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3901 adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3902 VDD rowon_n[0] adc_array_wafflecap_8_8_1[25]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3903 adc_array_wafflecap_8_8_0[0|3]/adc_array_circuit_150n_0/vint2 rowon_n[1] adc_array_wafflecap_8_8_0[0|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3904 VDD rowon_n[2] adc_array_wafflecap_8_8_0[1|11]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3905 adc_array_wafflecap_8_Dummy_4[9]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3906 VDD rowon_n[11] adc_array_wafflecap_8_8_0[10|25]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3907 adc_array_wafflecap_8_8_0[7|22]/adc_array_circuit_150n_0/vint1 col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3908 adc_array_wafflecap_8_8_0[3|15]/adc_array_circuit_150n_0/vint2 rowon_n[4] adc_array_wafflecap_8_8_0[3|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3909 VSS row_n[0] adc_array_wafflecap_8_8_1[20]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3910 adc_array_wafflecap_8_8_0[14|20]/adc_array_circuit_150n_0/vint2 col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3911 VDD rowon_n[10] adc_array_wafflecap_8_8_0[9|6]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3912 VDD rowon_n[10] adc_array_wafflecap_8_8_0[9|16]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3913 adc_array_wafflecap_8_8_1[30]/adc_array_circuit_150n_0/vint2 rowon_n[0] adc_array_wafflecap_8_8_1[30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3914 VSS VSS adc_array_wafflecap_8_Dummy_0[1]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3915 adc_array_wafflecap_8_8_0[1|26]/adc_array_circuit_150n_0/vint2 col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3916 adc_array_wafflecap_8_8_0[11|9]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|9]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3917 VDD rowon_n[4] adc_array_wafflecap_8_8_0[3|5]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3918 VSS row_n[2] adc_array_wafflecap_8_8_0[1|12]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3919 VDD sample_n adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3920 VSS row_n[6] adc_array_wafflecap_8_8_0[5|11]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3921 adc_array_wafflecap_8_8_0[5|1]/adc_array_circuit_150n_0/vint1 col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3922 adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3923 adc_array_wafflecap_8_8_0[2|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3924 adc_array_wafflecap_8_Dummy_3[0]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3925 adc_array_wafflecap_8_8_0[14|7]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|7]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3926 VSS row_n[13] adc_array_wafflecap_8_8_0[12|14]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3927 adc_array_wafflecap_8_8_0[9|11]/adc_array_circuit_150n_0/vint2 col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3928 adc_array_wafflecap_8_8_0[5|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3929 VDD VSS adc_array_wafflecap_8_Dummy_8[1]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3930 adc_array_wafflecap_8_8_0[1|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3931 VSS row_n[13] adc_array_wafflecap_8_8_0[12|4]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3932 adc_array_wafflecap_8_8_0[9|1]/adc_array_circuit_150n_0/vint2 col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3933 adc_array_wafflecap_8_8_0[12|20]/adc_array_circuit_150n_0/vdrv row_n[13] adc_array_wafflecap_8_8_0[12|20]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3934 adc_array_wafflecap_8_8_0[8|15]/adc_array_circuit_150n_0/vint2 col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3935 adc_array_wafflecap_8_8_0[1|26]/adc_array_circuit_150n_0/vdrv row_n[2] adc_array_wafflecap_8_8_0[1|26]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3936 adc_array_wafflecap_8_8_0[8|5]/adc_array_circuit_150n_0/vint2 col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3937 vcm VSS adc_array_wafflecap_8_Dummy_1[2]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3938 adc_array_wafflecap_8_8_0[11|10]/adc_array_circuit_150n_0/vint1 col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3939 adc_array_wafflecap_8_8_0[3|30]/adc_array_circuit_150n_0/vint2 col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3940 VSS row_n[1] adc_array_wafflecap_8_8_0[0|4]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3941 adc_array_wafflecap_8_8_0[1|12]/adc_array_circuit_150n_0/vint1 col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3942 vcm adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|10]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3943 adc_array_wafflecap_8_Dummy_4[23]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3944 adc_array_wafflecap_8_8_0[11|0]/adc_array_circuit_150n_0/vint1 col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3945 vcm adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|23]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3946 adc_array_wafflecap_8_8_0[10|14]/adc_array_circuit_150n_0/vint1 col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3947 adc_array_wafflecap_8_8_0[7|11]/adc_array_circuit_150n_0/vdrv row_n[8] adc_array_wafflecap_8_8_0[7|11]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3948 adc_array_wafflecap_8_8_0[10|4]/adc_array_circuit_150n_0/vint1 col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3949 adc_array_wafflecap_8_8_0[7|1]/adc_array_circuit_150n_0/vdrv row_n[8] adc_array_wafflecap_8_8_0[7|1]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3950 VSS VDD adc_array_wafflecap_8_Dummy_4[17]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3951 adc_array_wafflecap_8_8_0[10|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3952 adc_array_wafflecap_8_8_0[10|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3953 adc_array_wafflecap_8_8_0[11|17]/adc_array_circuit_150n_0/vint2 col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3954 adc_array_wafflecap_8_Dummy_8[2]/adc_array_circuit_150n_0/vint1 col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3955 adc_array_wafflecap_8_8_0[2|19]/adc_array_circuit_150n_0/vint2 col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3956 vcm adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|21]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3957 adc_array_wafflecap_8_8_0[5|23]/adc_array_circuit_150n_0/vint1 col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3958 adc_array_wafflecap_8_8_0[14|19]/adc_array_circuit_150n_0/vint2 rowon_n[15] adc_array_wafflecap_8_8_0[14|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3959 vcm adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|15]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3960 adc_array_wafflecap_8_Dummy_4[13]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[13]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3961 adc_array_wafflecap_8_8_0[7|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3962 adc_array_wafflecap_8_8_0[7|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3963 adc_array_wafflecap_8_Dummy_4[3]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[3]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3964 adc_array_wafflecap_8_8_0[14|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3965 adc_array_wafflecap_8_8_0[13|16]/adc_array_circuit_150n_0/vint1 col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3966 adc_array_wafflecap_8_8_0[13|23]/adc_array_circuit_150n_0/vint2 rowon_n[14] adc_array_wafflecap_8_8_0[13|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3967 VSS row_n[11] adc_array_wafflecap_8_8_0[10|20]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3968 vcm adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|2]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3969 vcm adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|12]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3970 adc_array_wafflecap_8_8_0[12|4]/adc_array_circuit_150n_0/vint2 rowon_n[13] adc_array_wafflecap_8_8_0[12|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3971 adc_array_wafflecap_8_8_0[12|14]/adc_array_circuit_150n_0/vint2 rowon_n[13] adc_array_wafflecap_8_8_0[12|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3972 adc_array_wafflecap_8_8_1[6]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[6]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3973 adc_array_wafflecap_8_8_0[0|19]/adc_array_circuit_150n_0/vdrv row_n[1] adc_array_wafflecap_8_8_0[0|19]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3974 vcm VSS adc_array_wafflecap_8_Dummy_4[12]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3975 adc_array_wafflecap_8_8_0[10|30]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|30]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3976 VSS row_n[5] adc_array_wafflecap_8_8_0[4|25]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3977 adc_array_wafflecap_8_8_1[16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3978 vcm VSS adc_array_wafflecap_8_Dummy_4[2]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3979 VDD rowon_n[13] adc_array_wafflecap_8_8_0[12|19]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3980 VDD rowon_n[12] adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3981 adc_array_wafflecap_8_8_0[10|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3982 adc_array_wafflecap_8_8_0[8|20]/adc_array_circuit_150n_0/vint1 col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3983 VDD rowon_n[11] adc_array_wafflecap_8_8_0[10|14]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3984 VDD rowon_n[11] adc_array_wafflecap_8_8_0[10|4]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3985 adc_array_wafflecap_8_Dummy_2[4]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_2[4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3986 adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/vint2 col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3987 adc_array_wafflecap_8_8_0[3|27]/adc_array_circuit_150n_0/vint1 col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3988 adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3989 VSS row_n[15] adc_array_wafflecap_8_8_0[14|8]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3990 adc_array_wafflecap_8_8_0[3|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3991 VSS row_n[14] adc_array_wafflecap_8_8_0[13|12]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3992 adc_array_wafflecap_8_8_0[10|9]/adc_array_circuit_150n_0/vint2 col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3993 adc_array_wafflecap_8_8_0[14|18]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|18]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3994 VSS row_n[14] adc_array_wafflecap_8_8_0[13|2]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3995 adc_array_wafflecap_8_Dummy_2[3]/adc_array_circuit_150n_0/vint2 col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3996 adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/vdrv row_n[13] adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3997 adc_array_wafflecap_8_8_0[10|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3998 adc_array_wafflecap_8_8_0[2|6]/adc_array_circuit_150n_0/vdrv row_n[3] adc_array_wafflecap_8_8_0[2|6]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3999 VSS VSS adc_array_wafflecap_8_Dummy_3[5]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4000 VSS row_n[3] adc_array_wafflecap_8_8_0[2|29]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4001 VDD rowon_n[0] adc_array_wafflecap_8_8_1[16]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4002 adc_array_wafflecap_8_8_0[12|8]/adc_array_circuit_150n_0/vint1 col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4003 adc_array_wafflecap_8_8_0[5|22]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|22]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4004 adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/vint1 col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4005 adc_array_wafflecap_8_8_0[1|23]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|23]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4006 adc_array_wafflecap_8_8_0[12|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4007 adc_array_wafflecap_8_8_0[8|9]/adc_array_circuit_150n_0/vdrv row_n[9] adc_array_wafflecap_8_8_0[8|9]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4008 adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4009 vcm adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[27]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4010 adc_array_wafflecap_8_8_0[0|29]/adc_array_circuit_150n_0/vint1 col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4011 adc_array_wafflecap_8_8_0[11|7]/adc_array_circuit_150n_0/vdrv row_n[12] adc_array_wafflecap_8_8_0[11|7]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4012 adc_array_wafflecap_8_8_0[9|18]/adc_array_circuit_150n_0/vint2 rowon_n[10] adc_array_wafflecap_8_8_0[9|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4013 adc_array_wafflecap_8_8_0[5|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4014 VDD rowon_n[5] adc_array_wafflecap_8_8_0[4|22]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4015 vcm adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4016 adc_array_wafflecap_8_8_0[4|10]/adc_array_circuit_150n_0/vdrv row_n[5] adc_array_wafflecap_8_8_0[4|10]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4017 adc_array_wafflecap_8_8_1[13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_1[13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4018 adc_array_wafflecap_8_8_0[14|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4019 vcm adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|18]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4020 adc_array_wafflecap_8_8_0[4|11]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|11]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4021 adc_array_wafflecap_8_8_0[3|2]/adc_array_circuit_150n_0/vint2 col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4022 vcm adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|19]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4023 adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4024 adc_array_wafflecap_8_8_0[8|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4025 adc_array_wafflecap_8_8_0[7|3]/adc_array_circuit_150n_0/vint2 rowon_n[8] adc_array_wafflecap_8_8_0[7|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4026 adc_array_wafflecap_8_8_0[7|13]/adc_array_circuit_150n_0/vint2 rowon_n[8] adc_array_wafflecap_8_8_0[7|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4027 vcm adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|10]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4028 adc_array_wafflecap_8_8_0[8|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4029 adc_array_wafflecap_8_8_1[7]/adc_array_circuit_150n_0/vdrv row_n[0] adc_array_wafflecap_8_8_1[7]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4030 adc_array_wafflecap_8_Dummy_4[28]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4031 adc_array_wafflecap_8_8_0[13|12]/adc_array_circuit_150n_0/vint2 rowon_n[14] adc_array_wafflecap_8_8_0[13|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4032 vcm adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|0]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4033 adc_array_wafflecap_8_8_0[6|5]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|5]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4034 adc_array_wafflecap_8_8_1[17]/adc_array_circuit_150n_0/vint1 col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4035 adc_array_wafflecap_8_8_0[13|2]/adc_array_circuit_150n_0/vint2 rowon_n[14] adc_array_wafflecap_8_8_0[13|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4036 VDD rowon_n[8] adc_array_wafflecap_8_8_0[7|18]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4037 adc_array_wafflecap_8_8_1[12]/adc_array_circuit_150n_0/vint2 col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4038 adc_array_wafflecap_8_8_0[11|28]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|28]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4039 adc_array_wafflecap_8_8_0[12|14]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|14]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4040 adc_array_wafflecap_8_8_0[3|8]/adc_array_circuit_150n_0/vint2 rowon_n[4] adc_array_wafflecap_8_8_0[3|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4041 adc_array_wafflecap_8_8_0[3|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4042 adc_array_wafflecap_8_8_0[12|4]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|4]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4043 adc_array_wafflecap_8_8_0[10|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4044 adc_array_wafflecap_8_8_0[6|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4045 adc_array_wafflecap_8_8_0[2|15]/adc_array_circuit_150n_0/vdrv row_n[3] adc_array_wafflecap_8_8_0[2|15]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4046 adc_array_wafflecap_8_8_1[3]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[3]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4047 adc_array_wafflecap_8_8_0[9|30]/adc_array_circuit_150n_0/vint2 col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4048 adc_array_wafflecap_8_8_0[2|16]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|16]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4049 adc_array_wafflecap_8_Dummy_4[30]/adc_array_circuit_150n_0/vint2 col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4050 VSS row_n[10] adc_array_wafflecap_8_8_0[9|7]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X4051 VDD rowon_n[3] adc_array_wafflecap_8_8_0[2|26]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4052 VSS row_n[9] adc_array_wafflecap_8_8_0[8|11]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4053 adc_array_wafflecap_8_8_0[3|24]/adc_array_circuit_150n_0/vint2 col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4054 VDD rowon_n[15] adc_array_wafflecap_8_8_0[14|10]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4055 adc_array_wafflecap_8_8_0[11|29]/adc_array_circuit_150n_0/vint1 col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4056 adc_array_wafflecap_8_8_0[9|17]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|17]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4057 VSS row_n[9] adc_array_wafflecap_8_8_0[8|1]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4058 adc_array_wafflecap_8_1_1/adc_array_circuit_150n_0/vint2 en_C0_n adc_array_wafflecap_8_1_1/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4059 VDD rowon_n[15] adc_array_wafflecap_8_8_0[14|0]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4060 adc_array_wafflecap_8_8_0[2|0]/adc_array_circuit_150n_0/vint2 rowon_n[3] adc_array_wafflecap_8_8_0[2|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4061 adc_array_wafflecap_8_8_0[7|30]/adc_array_circuit_150n_0/vdrv row_n[8] adc_array_wafflecap_8_8_0[7|30]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4062 adc_array_wafflecap_8_8_0[1|13]/adc_array_circuit_150n_0/vint2 rowon_n[2] adc_array_wafflecap_8_8_0[1|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4063 adc_array_wafflecap_8_8_0[11|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4064 adc_array_wafflecap_8_8_0[7|7]/adc_array_circuit_150n_0/vint1 col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4065 adc_array_wafflecap_8_8_0[13|29]/adc_array_circuit_150n_0/vdrv row_n[14] adc_array_wafflecap_8_8_0[13|29]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4066 adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4067 vcm adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|29]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4068 VSS row_n[4] adc_array_wafflecap_8_8_0[3|9]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4069 adc_array_wafflecap_8_8_0[0|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4070 adc_array_wafflecap_8_8_0[1|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4071 adc_array_wafflecap_8_8_0[4|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4072 VDD rowon_n[5] adc_array_wafflecap_8_8_0[4|30]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4073 adc_array_wafflecap_8_8_0[3|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4074 VDD rowon_n[1] adc_array_wafflecap_8_8_0[0|0]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4075 adc_array_wafflecap_8_8_0[13|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4076 adc_array_wafflecap_8_8_0[6|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4077 VDD rowon_n[0] adc_array_wafflecap_8_8_1[27]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4078 VDD rowon_n[2] adc_array_wafflecap_8_8_0[1|13]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4079 adc_array_wafflecap_8_8_0[0|5]/adc_array_circuit_150n_0/vint2 rowon_n[1] adc_array_wafflecap_8_8_0[0|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4080 vcm adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|7]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4081 vcm adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|8]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4082 adc_array_wafflecap_8_8_0[1|28]/adc_array_circuit_150n_0/vint2 col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4083 vcm VSS adc_array_wafflecap_8_Dummy_4[31]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4084 adc_array_wafflecap_8_8_0[11|18]/adc_array_circuit_150n_0/vdrv row_n[12] adc_array_wafflecap_8_8_0[11|18]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4085 adc_array_wafflecap_8_8_0[9|29]/adc_array_circuit_150n_0/vint2 rowon_n[10] adc_array_wafflecap_8_8_0[9|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4086 adc_array_wafflecap_8_8_0[5|27]/adc_array_circuit_150n_0/vint2 col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4087 adc_array_wafflecap_8_8_0[4|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4088 VSS VSS adc_array_wafflecap_8_Dummy_8[0]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4089 adc_array_wafflecap_8_8_0[0|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4090 VSS row_n[3] adc_array_wafflecap_8_8_0[2|1]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4091 adc_array_wafflecap_8_8_0[9|7]/adc_array_circuit_150n_0/vint2 rowon_n[10] adc_array_wafflecap_8_8_0[9|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4092 VSS row_n[2] adc_array_wafflecap_8_8_0[1|14]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4093 adc_array_wafflecap_8_Dummy_4[8]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4094 adc_array_wafflecap_8_8_0[12|22]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|22]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4095 adc_array_wafflecap_8_8_0[8|11]/adc_array_circuit_150n_0/vint2 rowon_n[9] adc_array_wafflecap_8_8_0[8|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4096 adc_array_wafflecap_8_8_0[2|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4097 adc_array_wafflecap_8_8_0[8|1]/adc_array_circuit_150n_0/vint2 rowon_n[9] adc_array_wafflecap_8_8_0[8|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4098 VDD VSS adc_array_wafflecap_8_Dummy_8[3]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4099 adc_array_wafflecap_8_8_0[1|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4100 vcm adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|8]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4101 adc_array_wafflecap_8_8_0[5|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4102 adc_array_wafflecap_8_8_0[4|16]/adc_array_circuit_150n_0/vint2 col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4103 adc_array_wafflecap_8_8_0[10|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4104 adc_array_wafflecap_8_8_0[10|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4105 adc_array_wafflecap_8_8_0[9|25]/adc_array_circuit_150n_0/vint1 col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4106 VDD rowon_n[8] adc_array_wafflecap_8_8_0[7|7]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4107 VDD rowon_n[8] adc_array_wafflecap_8_8_0[7|29]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4108 vcm adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_7/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4109 adc_array_wafflecap_8_8_0[0|1]/adc_array_circuit_150n_0/vint1 col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4110 adc_array_wafflecap_8_8_0[1|28]/adc_array_circuit_150n_0/vdrv row_n[2] adc_array_wafflecap_8_8_0[1|28]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4111 vcm VSS adc_array_wafflecap_8_Dummy_1[4]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4112 vcm adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|12]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4113 VSS row_n[15] adc_array_wafflecap_8_8_0[14|27]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4114 adc_array_wafflecap_8_8_0[3|19]/adc_array_circuit_150n_0/vdrv row_n[4] adc_array_wafflecap_8_8_0[3|19]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4115 adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/vint2 VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4116 VSS sample adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4117 adc_array_wafflecap_8_8_0[1|14]/adc_array_circuit_150n_0/vint1 col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4118 VSS row_n[14] adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4119 adc_array_wafflecap_8_8_0[10|28]/adc_array_circuit_150n_0/vint2 col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4120 VSS row_n[10] adc_array_wafflecap_8_8_0[9|18]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4121 VSS row_n[3] adc_array_wafflecap_8_8_0[2|23]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4122 VDD VDD adc_array_wafflecap_8_Dummy_4[31]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4123 adc_array_wafflecap_8_8_0[14|23]/adc_array_circuit_150n_0/vdrv row_n[15] adc_array_wafflecap_8_8_0[14|23]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4124 adc_array_wafflecap_8_8_0[12|27]/adc_array_circuit_150n_0/vint1 col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4125 VDD VDD adc_array_wafflecap_8_Dummy_4[9]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4126 vcm adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|23]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4127 adc_array_wafflecap_8_8_0[8|28]/adc_array_circuit_150n_0/vdrv row_n[9] adc_array_wafflecap_8_8_0[8|28]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4128 adc_array_wafflecap_8_8_0[5|25]/adc_array_circuit_150n_0/vint1 col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4129 vcm adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|26]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4130 adc_array_wafflecap_8_8_0[9|14]/adc_array_circuit_150n_0/vdrv row_n[10] adc_array_wafflecap_8_8_0[9|14]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4131 adc_array_wafflecap_8_8_0[7|18]/adc_array_circuit_150n_0/vint1 col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4132 adc_array_wafflecap_8_8_0[0|23]/adc_array_circuit_150n_0/vint1 col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4133 adc_array_wafflecap_8_8_0[11|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4134 adc_array_wafflecap_8_8_0[9|4]/adc_array_circuit_150n_0/vdrv row_n[10] adc_array_wafflecap_8_8_0[9|4]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4135 adc_array_wafflecap_8_8_0[14|16]/adc_array_circuit_150n_0/vint2 col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4136 VDD rowon_n[3] adc_array_wafflecap_8_8_0[2|17]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4137 adc_array_wafflecap_8_8_1[6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_1[6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4138 adc_array_wafflecap_8_8_0[6|19]/adc_array_circuit_150n_0/vint2 rowon_n[7] adc_array_wafflecap_8_8_0[6|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4139 VSS row_n[5] adc_array_wafflecap_8_8_0[4|26]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4140 VSS row_n[1] adc_array_wafflecap_8_8_0[0|27]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4141 adc_array_wafflecap_8_8_0[6|7]/adc_array_circuit_150n_0/vint2 col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4142 adc_array_wafflecap_8_8_0[12|16]/adc_array_circuit_150n_0/vdrv row_n[13] adc_array_wafflecap_8_8_0[12|16]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4143 VSS row_n[13] adc_array_wafflecap_8_8_0[12|23]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4144 adc_array_wafflecap_8_8_0[10|27]/adc_array_circuit_150n_0/vint2 rowon_n[11] adc_array_wafflecap_8_8_0[10|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4145 VSS row_n[7] adc_array_wafflecap_8_8_0[6|17]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4146 adc_array_wafflecap_8_8_0[13|20]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|20]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4147 adc_array_wafflecap_8_8_0[8|24]/adc_array_circuit_150n_0/vint2 col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4148 adc_array_wafflecap_8_8_0[3|20]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|20]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4149 adc_array_wafflecap_8_8_0[3|29]/adc_array_circuit_150n_0/vint1 col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4150 adc_array_wafflecap_8_8_0[3|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4151 adc_array_wafflecap_8_8_0[1|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4152 adc_array_wafflecap_8_Dummy_4[19]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4153 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.64e+07u l=1.6e+07u
X4154 vcm adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|4]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4155 adc_array_wafflecap_8_8_1[5]/adc_array_circuit_150n_0/vint2 col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4156 adc_array_wafflecap_8_Dummy_3[2]/adc_array_circuit_150n_0/vint1 col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4157 VDD rowon_n[15] adc_array_wafflecap_8_8_0[14|22]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4158 adc_array_wafflecap_8_8_0[12|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4159 adc_array_wafflecap_8_8_0[12|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4160 vcm adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|19]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4161 adc_array_wafflecap_8_8_0[11|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4162 adc_array_wafflecap_8_8_0[10|23]/adc_array_circuit_150n_0/vint1 col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4163 VSS row_n[10] adc_array_wafflecap_8_8_0[9|26]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4164 VDD rowon_n[7] adc_array_wafflecap_8_8_0[6|19]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4165 adc_array_wafflecap_8_Dummy_2[5]/adc_array_circuit_150n_0/vint2 col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4166 adc_array_wafflecap_8_8_0[11|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4167 VDD rowon_n[9] adc_array_wafflecap_8_8_0[8|27]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4168 adc_array_wafflecap_8_8_0[6|7]/adc_array_circuit_150n_0/vdrv row_n[7] adc_array_wafflecap_8_8_0[6|7]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4169 adc_array_wafflecap_8_8_0[2|8]/adc_array_circuit_150n_0/vdrv row_n[3] adc_array_wafflecap_8_8_0[2|8]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4170 adc_array_wafflecap_8_8_0[2|9]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|9]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4171 adc_array_wafflecap_8_8_0[2|18]/adc_array_circuit_150n_0/vint1 col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4172 VSS VSS adc_array_wafflecap_8_Dummy_6/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4173 adc_array_wafflecap_8_8_0[1|0]/adc_array_circuit_150n_0/vint2 col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4174 VSS row_n[3] adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4175 vcm adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|17]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4176 adc_array_wafflecap_8_8_0[6|17]/adc_array_circuit_150n_0/vint1 col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4177 adc_array_wafflecap_8_8_0[11|26]/adc_array_circuit_150n_0/vint2 col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4178 adc_array_wafflecap_8_8_0[1|25]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|25]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4179 adc_array_wafflecap_8_8_0[9|22]/adc_array_circuit_150n_0/vdrv row_n[10] adc_array_wafflecap_8_8_0[9|22]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4180 VSS VDD adc_array_wafflecap_8_Dummy_4[16]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4181 adc_array_wafflecap_8_8_0[7|26]/adc_array_circuit_150n_0/vint1 col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4182 VSS VDD adc_array_wafflecap_8_Dummy_4[6]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4183 adc_array_wafflecap_8_8_0[7|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4184 vcm adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[29]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4185 adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/vint1 col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4186 adc_array_wafflecap_8_Dummy_4[22]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[22]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4187 adc_array_wafflecap_8_8_0[12|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4188 vcm adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|21]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4189 adc_array_wafflecap_8_8_0[5|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4190 VDD rowon_n[5] adc_array_wafflecap_8_8_0[4|24]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4191 adc_array_wafflecap_8_8_0[1|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4192 adc_array_wafflecap_8_8_0[1|0]/adc_array_circuit_150n_0/vdrv row_n[2] adc_array_wafflecap_8_8_0[1|0]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4193 adc_array_wafflecap_8_8_0[4|12]/adc_array_circuit_150n_0/vdrv row_n[5] adc_array_wafflecap_8_8_0[4|12]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4194 adc_array_wafflecap_8_8_0[4|13]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|13]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4195 adc_array_wafflecap_8_8_1[15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_1[15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4196 adc_array_wafflecap_8_8_0[0|14]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|14]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4197 vcm adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|25]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4198 VDD rowon_n[0] adc_array_wafflecap_8_8_1[21]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4199 adc_array_wafflecap_8_8_1[9]/adc_array_circuit_150n_0/vdrv row_n[0] adc_array_wafflecap_8_8_1[9]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4200 adc_array_wafflecap_8_8_0[13|5]/adc_array_circuit_150n_0/vint1 col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4201 adc_array_wafflecap_8_8_0[13|15]/adc_array_circuit_150n_0/vint1 col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4202 adc_array_wafflecap_8_8_0[7|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4203 adc_array_wafflecap_8_8_0[7|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4204 adc_array_wafflecap_8_8_0[5|21]/adc_array_circuit_150n_0/vint2 col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4205 adc_array_wafflecap_8_8_1[14]/adc_array_circuit_150n_0/vint2 col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4206 adc_array_wafflecap_8_8_0[3|10]/adc_array_circuit_150n_0/vint2 rowon_n[4] adc_array_wafflecap_8_8_0[3|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4207 adc_array_wafflecap_8_8_1[25]/adc_array_circuit_150n_0/vint2 rowon_n[0] adc_array_wafflecap_8_8_1[25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4208 adc_array_wafflecap_8_8_1[5]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[5]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4209 vcm adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|27]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4210 adc_array_wafflecap_8_8_0[10|25]/adc_array_circuit_150n_0/vint2 rowon_n[11] adc_array_wafflecap_8_8_0[10|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4211 VSS row_n[8] adc_array_wafflecap_8_8_0[7|22]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4212 adc_array_wafflecap_8_8_0[6|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4213 VDD rowon_n[4] adc_array_wafflecap_8_8_0[3|0]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4214 VSS row_n[2] adc_array_wafflecap_8_8_0[1|7]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4215 adc_array_wafflecap_8_8_0[9|16]/adc_array_circuit_150n_0/vint2 rowon_n[10] adc_array_wafflecap_8_8_0[9|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4216 VSS row_n[6] adc_array_wafflecap_8_8_0[5|6]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4217 adc_array_wafflecap_8_Dummy_4[17]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4218 vcm adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|13]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4219 adc_array_wafflecap_8_8_0[9|6]/adc_array_circuit_150n_0/vint2 rowon_n[10] adc_array_wafflecap_8_8_0[9|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4220 adc_array_wafflecap_8_8_0[7|4]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|4]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4221 adc_array_wafflecap_8_8_0[7|14]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|14]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4222 adc_array_wafflecap_8_8_0[2|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4223 VDD rowon_n[3] adc_array_wafflecap_8_8_0[2|28]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4224 adc_array_wafflecap_8_Dummy_2[3]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4225 adc_array_wafflecap_8_Dummy_4[7]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4226 vcm adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|3]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4227 adc_array_wafflecap_8_8_0[10|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4228 adc_array_wafflecap_8_Dummy_2[1]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_2[1]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4229 VDD rowon_n[10] adc_array_wafflecap_8_8_0[9|21]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4230 adc_array_wafflecap_8_8_0[2|17]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|17]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4231 adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4232 adc_array_wafflecap_8_8_0[6|4]/adc_array_circuit_150n_0/vint2 col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4233 adc_array_wafflecap_8_Dummy_8[1]/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_8[1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4234 adc_array_wafflecap_8_8_0[13|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4235 VDD rowon_n[9] adc_array_wafflecap_8_8_0[8|25]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4236 adc_array_wafflecap_8_8_0[1|15]/adc_array_circuit_150n_0/vint2 rowon_n[2] adc_array_wafflecap_8_8_0[1|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4237 adc_array_wafflecap_8_8_0[12|20]/adc_array_circuit_150n_0/vint2 col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4238 VDD rowon_n[8] adc_array_wafflecap_8_8_0[7|6]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4239 VDD rowon_n[8] adc_array_wafflecap_8_8_0[7|16]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4240 adc_array_wafflecap_8_8_0[1|7]/adc_array_circuit_150n_0/vint1 col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4241 VSS row_n[4] adc_array_wafflecap_8_8_0[3|11]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4242 adc_array_wafflecap_8_8_0[3|1]/adc_array_circuit_150n_0/vint1 col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4243 adc_array_wafflecap_8_8_0[0|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4244 adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4245 adc_array_wafflecap_8_8_0[14|19]/adc_array_circuit_150n_0/vint1 col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4246 adc_array_wafflecap_8_8_0[12|7]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|7]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4247 VSS row_n[11] adc_array_wafflecap_8_8_0[10|14]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4248 adc_array_wafflecap_8_8_0[7|11]/adc_array_circuit_150n_0/vint2 col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4249 adc_array_wafflecap_8_8_0[6|28]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|28]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4250 adc_array_wafflecap_8_8_0[3|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4251 VSS row_n[11] adc_array_wafflecap_8_8_0[10|4]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4252 adc_array_wafflecap_8_8_0[7|1]/adc_array_circuit_150n_0/vint2 col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4253 adc_array_wafflecap_8_8_0[6|4]/adc_array_circuit_150n_0/vdrv row_n[7] adc_array_wafflecap_8_8_0[6|4]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4254 adc_array_wafflecap_8_8_0[6|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4255 adc_array_wafflecap_8_8_0[10|20]/adc_array_circuit_150n_0/vdrv row_n[11] adc_array_wafflecap_8_8_0[10|20]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4256 adc_array_wafflecap_8_Dummy_0[0]/adc_array_circuit_150n_0/vint1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4257 VDD rowon_n[0] adc_array_wafflecap_8_8_1[29]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4258 VDD rowon_n[2] adc_array_wafflecap_8_8_0[1|15]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4259 adc_array_wafflecap_8_8_0[9|10]/adc_array_circuit_150n_0/vint1 col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4260 adc_array_wafflecap_8_8_0[8|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4261 VSS VSS adc_array_wafflecap_8_Dummy_8[2]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4262 adc_array_wafflecap_8_8_1[12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4263 vcm adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|10]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4264 adc_array_wafflecap_8_8_0[1|30]/adc_array_circuit_150n_0/vint2 col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4265 adc_array_wafflecap_8_8_0[13|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4266 adc_array_wafflecap_8_8_0[9|0]/adc_array_circuit_150n_0/vint1 col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4267 adc_array_wafflecap_8_8_0[5|16]/adc_array_circuit_150n_0/vdrv row_n[6] adc_array_wafflecap_8_8_0[5|16]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4268 adc_array_wafflecap_8_8_0[8|14]/adc_array_circuit_150n_0/vint1 col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4269 adc_array_wafflecap_8_8_0[8|4]/adc_array_circuit_150n_0/vint1 col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4270 adc_array_wafflecap_8_8_0[5|2]/adc_array_circuit_150n_0/vint2 rowon_n[6] adc_array_wafflecap_8_8_0[5|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4271 adc_array_wafflecap_8_Dummy_4[3]/adc_array_circuit_150n_0/vint2 col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4272 adc_array_wafflecap_8_Dummy_4[13]/adc_array_circuit_150n_0/vint2 col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4273 VSS row_n[14] adc_array_wafflecap_8_8_0[13|16]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4274 adc_array_wafflecap_8_8_0[8|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4275 adc_array_wafflecap_8_8_0[5|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4276 VSS row_n[5] adc_array_wafflecap_8_8_0[4|20]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4277 adc_array_wafflecap_8_8_0[8|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4278 adc_array_wafflecap_8_8_0[7|22]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|22]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4279 adc_array_wafflecap_8_8_0[4|18]/adc_array_circuit_150n_0/vint2 col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4280 adc_array_wafflecap_8_8_0[0|19]/adc_array_circuit_150n_0/vint2 col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4281 adc_array_wafflecap_8_8_0[3|23]/adc_array_circuit_150n_0/vint1 col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4282 vcm adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[1]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4283 adc_array_wafflecap_8_8_0[1|30]/adc_array_circuit_150n_0/vdrv row_n[2] adc_array_wafflecap_8_8_0[1|30]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4284 adc_array_wafflecap_8_8_0[14|8]/adc_array_circuit_150n_0/vdrv row_n[15] adc_array_wafflecap_8_8_0[14|8]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4285 adc_array_wafflecap_8_8_0[12|19]/adc_array_circuit_150n_0/vint2 rowon_n[13] adc_array_wafflecap_8_8_0[12|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4286 vcm VSS adc_array_wafflecap_8_Dummy_1[6]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4287 adc_array_wafflecap_8_8_0[13|12]/adc_array_circuit_150n_0/vdrv row_n[14] adc_array_wafflecap_8_8_0[13|12]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4288 adc_array_wafflecap_8_8_0[14|25]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|25]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4289 adc_array_wafflecap_8_8_0[13|2]/adc_array_circuit_150n_0/vdrv row_n[14] adc_array_wafflecap_8_8_0[13|2]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4290 adc_array_wafflecap_8_8_0[12|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4291 adc_array_wafflecap_8_8_0[11|23]/adc_array_circuit_150n_0/vint2 rowon_n[12] adc_array_wafflecap_8_8_0[11|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4292 VSS row_n[9] adc_array_wafflecap_8_8_0[8|20]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4293 vcm adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|2]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4294 vcm adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|12]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4295 adc_array_wafflecap_8_8_0[10|4]/adc_array_circuit_150n_0/vint2 rowon_n[11] adc_array_wafflecap_8_8_0[10|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4296 adc_array_wafflecap_8_8_0[10|14]/adc_array_circuit_150n_0/vint2 rowon_n[11] adc_array_wafflecap_8_8_0[10|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4297 adc_array_wafflecap_8_Dummy_2[2]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_2[2]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4298 vcm adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|1]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4299 vcm adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|11]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4300 VSS row_n[3] adc_array_wafflecap_8_8_0[2|25]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4301 VSS row_n[6] adc_array_wafflecap_8_8_0[5|3]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4302 VDD rowon_n[11] adc_array_wafflecap_8_8_0[10|19]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4303 adc_array_wafflecap_8_8_0[9|6]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|6]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4304 adc_array_wafflecap_8_8_0[9|16]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|16]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4305 VDD rowon_n[10] adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4306 vcm adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|25]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4307 VDD rowon_n[9] adc_array_wafflecap_8_8_0[8|14]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4308 VDD rowon_n[9] adc_array_wafflecap_8_8_0[8|4]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4309 adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/vint2 col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4310 adc_array_wafflecap_8_8_0[5|26]/adc_array_circuit_150n_0/vint1 col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4311 vcm adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[23]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4312 adc_array_wafflecap_8_8_0[0|25]/adc_array_circuit_150n_0/vint1 col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4313 VSS row_n[13] adc_array_wafflecap_8_8_0[12|8]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4314 adc_array_wafflecap_8_8_0[5|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4315 adc_array_wafflecap_8_8_1[16]/adc_array_circuit_150n_0/vint2 rowon_n[0] adc_array_wafflecap_8_8_1[16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4316 adc_array_wafflecap_8_8_0[1|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4317 VSS row_n[12] adc_array_wafflecap_8_8_0[11|12]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X4318 adc_array_wafflecap_8_8_0[8|9]/adc_array_circuit_150n_0/vint2 col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4319 vcm adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|14]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4320 adc_array_wafflecap_8_8_0[14|30]/adc_array_circuit_150n_0/vint1 col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4321 adc_array_wafflecap_8_8_0[12|18]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|18]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4322 VSS row_n[12] adc_array_wafflecap_8_8_0[11|2]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X4323 adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/vdrv row_n[11] adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4324 adc_array_wafflecap_8_8_0[8|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4325 adc_array_wafflecap_8_8_1[8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_1[8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4326 VSS row_n[1] adc_array_wafflecap_8_8_0[0|29]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4327 adc_array_wafflecap_8_8_0[6|21]/adc_array_circuit_150n_0/vint2 rowon_n[7] adc_array_wafflecap_8_8_0[6|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4328 adc_array_wafflecap_8_8_0[10|8]/adc_array_circuit_150n_0/vint1 col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4329 adc_array_wafflecap_8_8_0[3|22]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|22]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4330 adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/vint1 col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4331 adc_array_wafflecap_8_8_0[10|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4332 adc_array_wafflecap_8_8_0[6|0]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|0]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4333 adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4334 vcm adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|6]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4335 adc_array_wafflecap_8_8_1[7]/adc_array_circuit_150n_0/vint2 col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4336 adc_array_wafflecap_8_Dummy_3[4]/adc_array_circuit_150n_0/vint1 col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4337 VSS row_n[0] adc_array_wafflecap_8_8_1[17]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4338 adc_array_wafflecap_8_8_0[9|7]/adc_array_circuit_150n_0/vdrv row_n[10] adc_array_wafflecap_8_8_0[9|7]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4339 adc_array_wafflecap_8_8_0[8|20]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|20]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4340 adc_array_wafflecap_8_8_0[7|18]/adc_array_circuit_150n_0/vint2 rowon_n[8] adc_array_wafflecap_8_8_0[7|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4341 adc_array_wafflecap_8_8_0[3|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4342 VDD rowon_n[3] adc_array_wafflecap_8_8_0[2|22]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4343 VDD sample_n adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4344 vcm adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4345 VDD rowon_n[7] adc_array_wafflecap_8_8_0[6|21]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4346 adc_array_wafflecap_8_8_0[2|10]/adc_array_circuit_150n_0/vdrv row_n[3] adc_array_wafflecap_8_8_0[2|10]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4347 adc_array_wafflecap_8_Dummy_4[7]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[7]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4348 adc_array_wafflecap_8_8_0[12|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4349 adc_array_wafflecap_8_8_0[7|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4350 adc_array_wafflecap_8_8_0[7|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4351 vcm adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|18]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4352 adc_array_wafflecap_8_8_0[2|11]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|11]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4353 adc_array_wafflecap_8_8_0[1|2]/adc_array_circuit_150n_0/vint2 col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4354 adc_array_wafflecap_8_8_0[14|19]/adc_array_circuit_150n_0/vdrv row_n[15] adc_array_wafflecap_8_8_0[14|19]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4355 adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4356 vcm adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|10]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4357 adc_array_wafflecap_8_Dummy_4[24]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[24]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4358 adc_array_wafflecap_8_8_0[13|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4359 adc_array_wafflecap_8_8_0[11|12]/adc_array_circuit_150n_0/vint2 rowon_n[12] adc_array_wafflecap_8_8_0[11|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4360 vcm adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|0]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4361 adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4362 adc_array_wafflecap_8_8_0[11|2]/adc_array_circuit_150n_0/vint2 rowon_n[12] adc_array_wafflecap_8_8_0[11|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4363 adc_array_wafflecap_8_8_0[14|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4364 adc_array_wafflecap_8_8_0[14|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4365 adc_array_wafflecap_8_8_0[10|14]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|14]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4366 adc_array_wafflecap_8_8_0[5|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4367 vcm adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4368 adc_array_wafflecap_8_8_0[1|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4369 adc_array_wafflecap_8_8_0[1|8]/adc_array_circuit_150n_0/vint2 rowon_n[2] adc_array_wafflecap_8_8_0[1|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4370 adc_array_wafflecap_8_8_0[1|2]/adc_array_circuit_150n_0/vdrv row_n[2] adc_array_wafflecap_8_8_0[1|2]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4371 adc_array_wafflecap_8_8_0[14|0]/adc_array_circuit_150n_0/vint2 rowon_n[15] adc_array_wafflecap_8_8_0[14|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4372 adc_array_wafflecap_8_8_0[14|10]/adc_array_circuit_150n_0/vint2 rowon_n[15] adc_array_wafflecap_8_8_0[14|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4373 adc_array_wafflecap_8_8_0[10|4]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|4]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4374 adc_array_wafflecap_8_8_0[7|30]/adc_array_circuit_150n_0/vint2 col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4375 adc_array_wafflecap_8_8_0[4|15]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|15]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4376 adc_array_wafflecap_8_8_0[0|16]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|16]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4377 VSS row_n[8] adc_array_wafflecap_8_8_0[7|7]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X4378 VDD rowon_n[0] adc_array_wafflecap_8_8_1[23]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4379 adc_array_wafflecap_8_8_0[13|29]/adc_array_circuit_150n_0/vint2 col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4380 adc_array_wafflecap_8_8_1[11]/adc_array_circuit_150n_0/vdrv row_n[0] adc_array_wafflecap_8_8_1[11]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4381 adc_array_wafflecap_8_8_0[5|23]/adc_array_circuit_150n_0/vint2 col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4382 adc_array_wafflecap_8_8_0[1|24]/adc_array_circuit_150n_0/vint2 col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4383 VDD rowon_n[13] adc_array_wafflecap_8_8_0[12|10]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4384 adc_array_wafflecap_8_8_0[11|25]/adc_array_circuit_150n_0/vdrv row_n[12] adc_array_wafflecap_8_8_0[11|25]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4385 adc_array_wafflecap_8_8_0[9|29]/adc_array_circuit_150n_0/vint1 col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4386 adc_array_wafflecap_8_8_0[6|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4387 adc_array_wafflecap_8_8_0[4|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4388 VDD rowon_n[2] adc_array_wafflecap_8_8_0[1|8]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4389 VDD rowon_n[13] adc_array_wafflecap_8_8_0[12|0]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4390 adc_array_wafflecap_8_8_0[0|0]/adc_array_circuit_150n_0/vint2 rowon_n[1] adc_array_wafflecap_8_8_0[0|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4391 adc_array_wafflecap_8_Dummy_4[29]/adc_array_circuit_150n_0/vint1 col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4392 adc_array_wafflecap_8_8_0[9|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4393 adc_array_wafflecap_8_8_1[27]/adc_array_circuit_150n_0/vint2 rowon_n[0] adc_array_wafflecap_8_8_1[27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4394 adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4395 VSS row_n[2] adc_array_wafflecap_8_8_0[1|9]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4396 adc_array_wafflecap_8_8_0[2|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4397 adc_array_wafflecap_8_Dummy_2[5]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4398 VDD rowon_n[3] adc_array_wafflecap_8_8_0[2|30]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4399 VDD VSS adc_array_wafflecap_8_Dummy_0[1]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4400 adc_array_wafflecap_8_8_0[1|24]/adc_array_circuit_150n_0/vdrv row_n[2] adc_array_wafflecap_8_8_0[1|24]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4401 adc_array_wafflecap_8_8_0[1|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4402 adc_array_wafflecap_8_8_0[14|27]/adc_array_circuit_150n_0/vdrv row_n[15] adc_array_wafflecap_8_8_0[14|27]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4403 adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4404 adc_array_wafflecap_8_8_0[11|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4405 adc_array_wafflecap_8_Dummy_8[3]/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_8[3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4406 vcm VSS adc_array_wafflecap_8_4_0/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4407 vcm adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|7]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4408 adc_array_wafflecap_8_8_0[14|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4409 vcm adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|30]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4410 adc_array_wafflecap_8_8_0[9|18]/adc_array_circuit_150n_0/vdrv row_n[10] adc_array_wafflecap_8_8_0[9|18]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4411 VSS row_n[10] adc_array_wafflecap_8_8_0[9|25]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4412 adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4413 adc_array_wafflecap_8_8_0[7|29]/adc_array_circuit_150n_0/vint2 rowon_n[8] adc_array_wafflecap_8_8_0[7|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4414 adc_array_wafflecap_8_8_0[3|27]/adc_array_circuit_150n_0/vint2 col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4415 adc_array_wafflecap_8_Dummy_2[1]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_2[1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4416 VSS row_n[1] adc_array_wafflecap_8_8_0[0|1]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4417 adc_array_wafflecap_8_8_0[1|9]/adc_array_circuit_150n_0/vint1 col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4418 adc_array_wafflecap_8_8_0[2|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4419 adc_array_wafflecap_8_8_0[8|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4420 adc_array_wafflecap_8_8_0[7|7]/adc_array_circuit_150n_0/vint2 rowon_n[8] adc_array_wafflecap_8_8_0[7|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4421 vcm adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|16]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4422 adc_array_wafflecap_8_8_0[13|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4423 adc_array_wafflecap_8_8_0[10|22]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|22]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4424 adc_array_wafflecap_8_8_0[0|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4425 vcm adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|6]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4426 adc_array_wafflecap_8_8_0[6|30]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|30]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4427 VDD rowon_n[12] adc_array_wafflecap_8_8_0[11|24]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4428 adc_array_wafflecap_8_8_0[9|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4429 adc_array_wafflecap_8_8_0[6|12]/adc_array_circuit_150n_0/vint2 rowon_n[7] adc_array_wafflecap_8_8_0[6|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4430 adc_array_wafflecap_8_8_0[3|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4431 adc_array_wafflecap_8_8_0[9|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4432 adc_array_wafflecap_8_8_0[6|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4433 adc_array_wafflecap_8_8_0[2|16]/adc_array_circuit_150n_0/vint2 col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4434 adc_array_wafflecap_8_8_0[7|7]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|7]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4435 adc_array_wafflecap_8_8_0[7|25]/adc_array_circuit_150n_0/vint1 col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4436 adc_array_wafflecap_8_1_1/adc_array_circuit_150n_0/vint1 en_C0_n VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4437 adc_array_wafflecap_8_8_1[28]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[28]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4438 adc_array_wafflecap_8_8_0[6|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4439 adc_array_wafflecap_8_8_0[5|20]/adc_array_circuit_150n_0/vint1 col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4440 vcm adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|12]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4441 adc_array_wafflecap_8_Dummy_4[9]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4442 adc_array_wafflecap_8_Dummy_4[31]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4443 adc_array_wafflecap_8_8_0[14|23]/adc_array_circuit_150n_0/vint2 col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4444 VSS row_n[13] adc_array_wafflecap_8_8_0[12|27]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4445 adc_array_wafflecap_8_8_0[5|18]/adc_array_circuit_150n_0/vdrv row_n[6] adc_array_wafflecap_8_8_0[5|18]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4446 adc_array_wafflecap_8_8_1[14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4447 VSS sample adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4448 adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/vint2 VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4449 VSS row_n[12] adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4450 adc_array_wafflecap_8_8_0[8|28]/adc_array_circuit_150n_0/vint2 col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4451 adc_array_wafflecap_8_8_0[5|19]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|19]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4452 VDD rowon_n[7] adc_array_wafflecap_8_8_0[6|12]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4453 adc_array_wafflecap_8_8_0[14|10]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|10]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4454 adc_array_wafflecap_8_8_0[9|14]/adc_array_circuit_150n_0/vint2 col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4455 adc_array_wafflecap_8_8_0[5|4]/adc_array_circuit_150n_0/vint2 rowon_n[6] adc_array_wafflecap_8_8_0[5|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4456 VSS row_n[1] adc_array_wafflecap_8_8_0[0|23]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4457 adc_array_wafflecap_8_8_0[0|16]/adc_array_circuit_150n_0/vdrv row_n[1] adc_array_wafflecap_8_8_0[0|16]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4458 adc_array_wafflecap_8_8_0[14|0]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|0]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4459 VDD rowon_n[15] adc_array_wafflecap_8_8_0[14|26]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4460 adc_array_wafflecap_8_8_0[9|4]/adc_array_circuit_150n_0/vint2 col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4461 VSS row_n[8] adc_array_wafflecap_8_8_0[7|18]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4462 VSS row_n[5] adc_array_wafflecap_8_8_0[4|22]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4463 VDD rowon_n[14] adc_array_wafflecap_8_8_0[13|30]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4464 adc_array_wafflecap_8_8_0[12|23]/adc_array_circuit_150n_0/vdrv row_n[13] adc_array_wafflecap_8_8_0[12|23]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4465 adc_array_wafflecap_8_8_0[10|27]/adc_array_circuit_150n_0/vint1 col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4466 adc_array_wafflecap_8_8_0[9|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4467 adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/vint2 rowon_n[5] adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4468 VDD rowon_n[14] adc_array_wafflecap_8_8_0[13|8]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4469 VSS row_n[7] adc_array_wafflecap_8_8_0[6|13]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4470 adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/vdrv row_n[2] adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4471 adc_array_wafflecap_8_8_0[11|13]/adc_array_circuit_150n_0/vint1 col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4472 adc_array_wafflecap_8_8_0[3|25]/adc_array_circuit_150n_0/vint1 col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4473 adc_array_wafflecap_8_Dummy_4[26]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4474 adc_array_wafflecap_8_8_0[11|3]/adc_array_circuit_150n_0/vint1 col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4475 vcm adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|26]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4476 adc_array_wafflecap_8_8_0[7|14]/adc_array_circuit_150n_0/vdrv row_n[8] adc_array_wafflecap_8_8_0[7|14]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4477 adc_array_wafflecap_8_Dummy_2[6]/adc_array_circuit_150n_0/vint1 col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4478 adc_array_wafflecap_8_8_0[7|4]/adc_array_circuit_150n_0/vdrv row_n[8] adc_array_wafflecap_8_8_0[7|4]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4479 adc_array_wafflecap_8_8_0[12|16]/adc_array_circuit_150n_0/vint2 col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4480 VSS sample_n adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4481 adc_array_wafflecap_8_8_0[7|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4482 adc_array_wafflecap_8_8_0[6|13]/adc_array_circuit_150n_0/vint1 col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4483 VSS row_n[6] adc_array_wafflecap_8_8_0[5|5]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4484 adc_array_wafflecap_8_8_0[14|22]/adc_array_circuit_150n_0/vint2 rowon_n[15] adc_array_wafflecap_8_8_0[14|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4485 VSS VSS adc_array_wafflecap_8_Dummy_3[2]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4486 VSS row_n[3] adc_array_wafflecap_8_8_0[2|26]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4487 adc_array_wafflecap_8_Dummy_4[6]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[6]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4488 adc_array_wafflecap_8_Dummy_4[16]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[16]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4489 adc_array_wafflecap_8_Dummy_4[20]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4490 adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4491 adc_array_wafflecap_8_8_0[10|16]/adc_array_circuit_150n_0/vdrv row_n[11] adc_array_wafflecap_8_8_0[10|16]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4492 VSS row_n[11] adc_array_wafflecap_8_8_0[10|23]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4493 vcm adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|5]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4494 vcm adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|15]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4495 adc_array_wafflecap_8_8_0[8|27]/adc_array_circuit_150n_0/vint2 rowon_n[9] adc_array_wafflecap_8_8_0[8|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4496 adc_array_wafflecap_8_8_0[11|20]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|20]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4497 vcm adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[25]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4498 adc_array_wafflecap_8_8_0[1|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4499 adc_array_wafflecap_8_8_0[1|20]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|20]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4500 vcm VSS adc_array_wafflecap_8_Dummy_4[15]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4501 adc_array_wafflecap_8_8_0[13|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4502 adc_array_wafflecap_8_8_0[5|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4503 vcm adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|4]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4504 vcm VSS adc_array_wafflecap_8_Dummy_4[5]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4505 vcm adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|16]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4506 VDD rowon_n[13] adc_array_wafflecap_8_8_0[12|22]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4507 adc_array_wafflecap_8_8_0[10|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4508 adc_array_wafflecap_8_8_0[10|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4509 adc_array_wafflecap_8_8_0[0|26]/adc_array_circuit_150n_0/vint1 col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4510 adc_array_wafflecap_8_8_0[9|22]/adc_array_circuit_150n_0/vint2 col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4511 adc_array_wafflecap_8_8_0[8|23]/adc_array_circuit_150n_0/vint1 col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4512 VSS row_n[8] adc_array_wafflecap_8_8_0[7|26]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4513 VDD rowon_n[5] adc_array_wafflecap_8_8_0[4|19]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4514 adc_array_wafflecap_8_8_0[4|7]/adc_array_circuit_150n_0/vdrv row_n[5] adc_array_wafflecap_8_8_0[4|7]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4515 adc_array_wafflecap_8_8_0[4|8]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|8]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4516 adc_array_wafflecap_8_8_1[10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_1[10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4517 VSS row_n[1] adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4518 adc_array_wafflecap_8_8_0[0|9]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|9]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4519 adc_array_wafflecap_8_Dummy_4[22]/adc_array_circuit_150n_0/vint2 col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4520 vcm adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|17]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4521 adc_array_wafflecap_8_8_0[7|18]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|18]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4522 adc_array_wafflecap_8_8_0[6|23]/adc_array_circuit_150n_0/vint2 rowon_n[7] adc_array_wafflecap_8_8_0[6|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4523 adc_array_wafflecap_8_8_0[4|17]/adc_array_circuit_150n_0/vint1 col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4524 adc_array_wafflecap_8_8_0[4|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4525 adc_array_wafflecap_8_8_0[11|21]/adc_array_circuit_150n_0/vint1 col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4526 adc_array_wafflecap_8_8_0[7|22]/adc_array_circuit_150n_0/vdrv row_n[8] adc_array_wafflecap_8_8_0[7|22]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4527 adc_array_wafflecap_8_8_0[6|2]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|2]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4528 adc_array_wafflecap_8_8_1[21]/adc_array_circuit_150n_0/vint2 rowon_n[0] adc_array_wafflecap_8_8_1[21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4529 adc_array_wafflecap_8_Dummy_4[9]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[9]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4530 VSS row_n[14] adc_array_wafflecap_8_8_0[13|15]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4531 adc_array_wafflecap_8_8_1[9]/adc_array_circuit_150n_0/vint2 col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4532 VSS row_n[14] adc_array_wafflecap_8_8_0[13|5]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4533 adc_array_wafflecap_8_8_0[13|21]/adc_array_circuit_150n_0/vdrv row_n[14] adc_array_wafflecap_8_8_0[13|21]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4534 adc_array_wafflecap_8_8_0[10|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4535 vcm adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|21]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4536 VDD rowon_n[7] adc_array_wafflecap_8_8_0[6|23]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4537 adc_array_wafflecap_8_8_0[3|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4538 VDD rowon_n[3] adc_array_wafflecap_8_8_0[2|24]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4539 adc_array_wafflecap_8_8_1[0]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[0]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4540 adc_array_wafflecap_8_8_0[6|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4541 adc_array_wafflecap_8_8_0[2|12]/adc_array_circuit_150n_0/vdrv row_n[3] adc_array_wafflecap_8_8_0[2|12]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4542 adc_array_wafflecap_8_8_0[2|13]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|13]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4543 adc_array_wafflecap_8_Dummy_1[5]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_1[5]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4544 VDD sample adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4545 adc_array_wafflecap_8_8_0[3|21]/adc_array_circuit_150n_0/vint2 col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4546 vcm VSS adc_array_wafflecap_8_Dummy_4[23]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4547 adc_array_wafflecap_8_8_0[11|10]/adc_array_circuit_150n_0/vdrv row_n[12] adc_array_wafflecap_8_8_0[11|10]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4548 adc_array_wafflecap_8_8_0[9|21]/adc_array_circuit_150n_0/vint2 rowon_n[10] adc_array_wafflecap_8_8_0[9|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4549 adc_array_wafflecap_8_8_0[8|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4550 adc_array_wafflecap_8_8_0[1|10]/adc_array_circuit_150n_0/vint2 rowon_n[2] adc_array_wafflecap_8_8_0[1|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4551 adc_array_wafflecap_8_8_0[11|0]/adc_array_circuit_150n_0/vdrv row_n[12] adc_array_wafflecap_8_8_0[11|0]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4552 adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4553 adc_array_wafflecap_8_8_0[6|24]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|24]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4554 adc_array_wafflecap_8_8_0[5|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4555 adc_array_wafflecap_8_8_0[8|25]/adc_array_circuit_150n_0/vint2 rowon_n[9] adc_array_wafflecap_8_8_0[8|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4556 adc_array_wafflecap_8_8_0[14|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4557 adc_array_wafflecap_8_8_0[14|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4558 adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4559 adc_array_wafflecap_8_8_0[7|16]/adc_array_circuit_150n_0/vint2 rowon_n[8] adc_array_wafflecap_8_8_0[7|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4560 VSS row_n[4] adc_array_wafflecap_8_8_0[3|6]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4561 adc_array_wafflecap_8_8_0[13|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4562 vcm adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|13]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4563 adc_array_wafflecap_8_8_0[8|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4564 adc_array_wafflecap_8_8_0[7|6]/adc_array_circuit_150n_0/vint2 rowon_n[8] adc_array_wafflecap_8_8_0[7|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4565 adc_array_wafflecap_8_8_0[0|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4566 adc_array_wafflecap_8_Dummy_4[31]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4567 adc_array_wafflecap_8_8_0[13|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4568 vcm adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|3]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4569 vcm adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|29]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4570 adc_array_wafflecap_8_8_0[0|17]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|17]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4571 VDD rowon_n[8] adc_array_wafflecap_8_8_0[7|21]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4572 adc_array_wafflecap_8_8_0[6|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4573 adc_array_wafflecap_8_8_0[5|25]/adc_array_circuit_150n_0/vint2 col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4574 adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4575 adc_array_wafflecap_8_8_0[4|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4576 VDD rowon_n[2] adc_array_wafflecap_8_8_0[1|10]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4577 VSS row_n[15] adc_array_wafflecap_8_8_0[14|19]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4578 adc_array_wafflecap_8_8_0[11|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4579 adc_array_wafflecap_8_8_0[10|20]/adc_array_circuit_150n_0/vint2 col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4580 adc_array_wafflecap_8_8_1[29]/adc_array_circuit_150n_0/vint2 rowon_n[0] adc_array_wafflecap_8_8_1[29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4581 VSS VSS adc_array_wafflecap_8_Dummy_0[0]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4582 adc_array_wafflecap_8_8_1[7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4583 VSS row_n[2] adc_array_wafflecap_8_8_0[1|11]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4584 VSS row_n[10] adc_array_wafflecap_8_8_0[9|0]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4585 VSS row_n[10] adc_array_wafflecap_8_8_0[9|10]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4586 adc_array_wafflecap_8_8_0[4|14]/adc_array_circuit_150n_0/vint2 col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4587 adc_array_wafflecap_8_1_0/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4588 adc_array_wafflecap_8_8_0[12|19]/adc_array_circuit_150n_0/vint1 col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4589 adc_array_wafflecap_8_8_0[10|7]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|7]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4590 VSS row_n[9] adc_array_wafflecap_8_8_0[8|14]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4591 adc_array_wafflecap_8_8_0[5|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4592 adc_array_wafflecap_8_8_0[1|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4593 VDD rowon_n[15] adc_array_wafflecap_8_8_0[14|13]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4594 adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/vint1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4595 VSS row_n[9] adc_array_wafflecap_8_8_0[8|4]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4596 adc_array_wafflecap_8_8_0[4|4]/adc_array_circuit_150n_0/vdrv row_n[5] adc_array_wafflecap_8_8_0[4|4]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4597 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X4598 VDD rowon_n[15] adc_array_wafflecap_8_8_0[14|3]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4599 adc_array_wafflecap_8_8_0[8|20]/adc_array_circuit_150n_0/vdrv row_n[9] adc_array_wafflecap_8_8_0[8|20]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4600 adc_array_wafflecap_8_Dummy_4[20]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[20]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4601 adc_array_wafflecap_8_8_0[11|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4602 adc_array_wafflecap_8_8_0[7|10]/adc_array_circuit_150n_0/vint1 col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4603 vcm VSS adc_array_wafflecap_8_Dummy_1[1]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4604 adc_array_wafflecap_8_8_0[1|11]/adc_array_circuit_150n_0/vint1 col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4605 adc_array_wafflecap_8_8_0[7|0]/adc_array_circuit_150n_0/vint1 col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4606 adc_array_wafflecap_8_8_0[3|16]/adc_array_circuit_150n_0/vdrv row_n[4] adc_array_wafflecap_8_8_0[3|16]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4607 adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n sample VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4608 adc_array_wafflecap_8_8_0[14|8]/adc_array_circuit_150n_0/vint2 col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4609 adc_array_wafflecap_8_8_0[3|2]/adc_array_circuit_150n_0/vint2 rowon_n[4] adc_array_wafflecap_8_8_0[3|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4610 adc_array_wafflecap_8_8_0[13|2]/adc_array_circuit_150n_0/vint2 col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4611 adc_array_wafflecap_8_8_0[13|12]/adc_array_circuit_150n_0/vint2 col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4612 VSS row_n[12] adc_array_wafflecap_8_8_0[11|16]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4613 adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4614 adc_array_wafflecap_8_8_0[6|14]/adc_array_circuit_150n_0/vint2 rowon_n[7] adc_array_wafflecap_8_8_0[6|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4615 adc_array_wafflecap_8_8_0[3|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4616 VSS row_n[3] adc_array_wafflecap_8_8_0[2|20]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4617 adc_array_wafflecap_8_Dummy_2[2]/adc_array_circuit_150n_0/vint2 col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4618 adc_array_wafflecap_8_8_0[2|18]/adc_array_circuit_150n_0/vint2 col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4619 vcm adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|20]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4620 adc_array_wafflecap_8_8_0[5|22]/adc_array_circuit_150n_0/vint1 col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4621 adc_array_wafflecap_8_8_1[30]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[30]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4622 adc_array_wafflecap_8_Dummy_4[2]/adc_array_circuit_150n_0/vint1 col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4623 adc_array_wafflecap_8_Dummy_4[12]/adc_array_circuit_150n_0/vint1 col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4624 adc_array_wafflecap_8_8_0[12|8]/adc_array_circuit_150n_0/vdrv row_n[13] adc_array_wafflecap_8_8_0[12|8]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4625 adc_array_wafflecap_8_8_0[10|19]/adc_array_circuit_150n_0/vint2 rowon_n[11] adc_array_wafflecap_8_8_0[10|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4626 adc_array_wafflecap_8_8_0[9|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4627 adc_array_wafflecap_8_8_0[9|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4628 adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/vint2 rowon_n[10] adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4629 adc_array_wafflecap_8_8_0[6|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4630 adc_array_wafflecap_8_8_0[5|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4631 VDD rowon_n[6] adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4632 adc_array_wafflecap_8_Dummy_4[11]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4633 adc_array_wafflecap_8_8_0[12|25]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|25]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4634 adc_array_wafflecap_8_8_0[10|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4635 adc_array_wafflecap_8_8_0[0|20]/adc_array_circuit_150n_0/vint1 col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4636 adc_array_wafflecap_8_Dummy_4[1]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4637 adc_array_wafflecap_8_8_0[8|4]/adc_array_circuit_150n_0/vint2 rowon_n[9] adc_array_wafflecap_8_8_0[8|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4638 adc_array_wafflecap_8_8_0[8|14]/adc_array_circuit_150n_0/vint2 rowon_n[9] adc_array_wafflecap_8_8_0[8|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4639 VDD rowon_n[7] adc_array_wafflecap_8_8_0[6|14]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4640 adc_array_wafflecap_8_8_0[5|6]/adc_array_circuit_150n_0/vint2 rowon_n[6] adc_array_wafflecap_8_8_0[5|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4641 adc_array_wafflecap_8_8_0[0|18]/adc_array_circuit_150n_0/vdrv row_n[1] adc_array_wafflecap_8_8_0[0|18]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4642 vcm adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|1]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4643 vcm adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|11]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4644 VSS row_n[5] adc_array_wafflecap_8_8_0[4|24]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4645 ctop sw_n analog_in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4646 VSS row_n[1] adc_array_wafflecap_8_8_0[0|25]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4647 adc_array_wafflecap_8_8_0[6|29]/adc_array_circuit_150n_0/vint2 col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4648 vcm adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|9]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4649 VSS row_n[4] adc_array_wafflecap_8_8_0[3|3]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4650 VDD rowon_n[9] adc_array_wafflecap_8_8_0[8|19]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4651 VDD rowon_n[8] adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4652 VSS row_n[7] adc_array_wafflecap_8_8_0[6|15]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4653 VSS row_n[15] adc_array_wafflecap_8_8_0[14|30]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4654 adc_array_wafflecap_8_Dummy_4[28]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[28]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4655 adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/vint2 col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4656 adc_array_wafflecap_8_8_0[3|26]/adc_array_circuit_150n_0/vint1 col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4657 adc_array_wafflecap_8_Dummy_3[0]/adc_array_circuit_150n_0/vint1 col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4658 VSS row_n[11] adc_array_wafflecap_8_8_0[10|8]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4659 adc_array_wafflecap_8_8_0[3|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4660 adc_array_wafflecap_8_8_0[14|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4661 adc_array_wafflecap_8_8_0[6|29]/adc_array_circuit_150n_0/vdrv row_n[7] adc_array_wafflecap_8_8_0[6|29]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4662 vcm adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|1]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4663 adc_array_wafflecap_8_8_0[10|18]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|18]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4664 adc_array_wafflecap_8_8_0[6|15]/adc_array_circuit_150n_0/vint1 col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4665 vcm adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|14]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4666 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X4667 VDD VDD adc_array_wafflecap_8_Dummy_4[12]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4668 adc_array_wafflecap_8_8_0[12|30]/adc_array_circuit_150n_0/vint1 col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4669 VDD VDD adc_array_wafflecap_8_Dummy_4[2]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4670 adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/vdrv row_n[9] adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4671 VSS VSS adc_array_wafflecap_8_Dummy_3[4]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4672 adc_array_wafflecap_8_8_0[9|7]/adc_array_circuit_150n_0/vint2 col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4673 adc_array_wafflecap_8_8_0[8|8]/adc_array_circuit_150n_0/vint1 col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4674 adc_array_wafflecap_8_8_0[1|22]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|22]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4675 adc_array_wafflecap_8_Dummy_4[7]/adc_array_circuit_150n_0/vint2 col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4676 adc_array_wafflecap_8_8_0[14|19]/adc_array_circuit_150n_0/vint2 col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4677 adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4678 adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4679 adc_array_wafflecap_8_8_0[11|6]/adc_array_circuit_150n_0/vint1 col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4680 vcm adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|6]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4681 adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4682 adc_array_wafflecap_8_8_0[7|7]/adc_array_circuit_150n_0/vdrv row_n[8] adc_array_wafflecap_8_8_0[7|7]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4683 adc_array_wafflecap_8_8_0[5|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4684 vcm adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[26]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4685 adc_array_wafflecap_8_8_0[1|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4686 vcm adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4687 VDD rowon_n[5] adc_array_wafflecap_8_8_0[4|21]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4688 adc_array_wafflecap_8_8_0[13|6]/adc_array_circuit_150n_0/vdrv row_n[14] adc_array_wafflecap_8_8_0[13|6]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4689 adc_array_wafflecap_8_8_0[10|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4690 adc_array_wafflecap_8_8_0[6|25]/adc_array_circuit_150n_0/vint2 rowon_n[7] adc_array_wafflecap_8_8_0[6|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4691 vcm adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|17]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4692 adc_array_wafflecap_8_8_0[4|10]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|10]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4693 adc_array_wafflecap_8_8_0[0|11]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|11]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4694 vcm adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|18]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4695 adc_array_wafflecap_8_8_0[12|19]/adc_array_circuit_150n_0/vdrv row_n[13] adc_array_wafflecap_8_8_0[12|19]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4696 adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4697 VDD rowon_n[0] adc_array_wafflecap_8_8_1[18]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4698 adc_array_wafflecap_8_8_0[13|23]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|23]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4699 adc_array_wafflecap_8_8_1[6]/adc_array_circuit_150n_0/vdrv row_n[0] adc_array_wafflecap_8_8_1[6]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4700 adc_array_wafflecap_8_8_0[11|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4701 adc_array_wafflecap_8_8_1[23]/adc_array_circuit_150n_0/vint2 rowon_n[0] adc_array_wafflecap_8_8_1[23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4702 adc_array_wafflecap_8_8_1[16]/adc_array_circuit_150n_0/vint1 col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4703 VSS row_n[6] adc_array_wafflecap_8_8_0[5|28]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4704 adc_array_wafflecap_8_8_0[4|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4705 adc_array_wafflecap_8_8_1[11]/adc_array_circuit_150n_0/vint2 col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4706 adc_array_wafflecap_8_8_0[12|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4707 adc_array_wafflecap_8_8_0[12|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4708 adc_array_wafflecap_8_8_0[12|10]/adc_array_circuit_150n_0/vint2 rowon_n[13] adc_array_wafflecap_8_8_0[12|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4709 VSS row_n[10] adc_array_wafflecap_8_8_0[9|29]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4710 adc_array_wafflecap_8_8_0[3|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4711 adc_array_wafflecap_8_8_0[12|0]/adc_array_circuit_150n_0/vint2 rowon_n[13] adc_array_wafflecap_8_8_0[12|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4712 VDD rowon_n[7] adc_array_wafflecap_8_8_0[6|25]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4713 adc_array_wafflecap_8_8_0[6|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4714 adc_array_wafflecap_8_8_1[2]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[2]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4715 vcm VSS adc_array_wafflecap_8_Dummy_4[8]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4716 VSS VDD adc_array_wafflecap_8_Dummy_4[29]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4717 adc_array_wafflecap_8_8_0[2|15]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|15]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4718 adc_array_wafflecap_8_2_0/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_2_0/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4719 VDD rowon_n[12] adc_array_wafflecap_8_8_0[11|28]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4720 adc_array_wafflecap_8_8_0[11|29]/adc_array_circuit_150n_0/vint2 col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4721 adc_array_wafflecap_8_8_0[3|23]/adc_array_circuit_150n_0/vint2 col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4722 VDD rowon_n[11] adc_array_wafflecap_8_8_0[10|10]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4723 adc_array_wafflecap_8_8_0[9|25]/adc_array_circuit_150n_0/vdrv row_n[10] adc_array_wafflecap_8_8_0[9|25]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4724 adc_array_wafflecap_8_8_0[7|29]/adc_array_circuit_150n_0/vint1 col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4725 adc_array_wafflecap_8_8_0[2|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4726 VDD rowon_n[11] adc_array_wafflecap_8_8_0[10|0]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4727 adc_array_wafflecap_8_8_0[6|1]/adc_array_circuit_150n_0/vint2 col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4728 adc_array_wafflecap_8_Dummy_0[1]/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_0[1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4729 adc_array_wafflecap_8_Dummy_4[25]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[25]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4730 adc_array_wafflecap_8_8_0[14|27]/adc_array_circuit_150n_0/vint2 col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4731 adc_array_wafflecap_8_8_0[13|28]/adc_array_circuit_150n_0/vint1 col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4732 vcm adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|24]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4733 adc_array_wafflecap_8_8_0[7|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4734 adc_array_wafflecap_8_8_0[6|26]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|26]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4735 adc_array_wafflecap_8_8_0[9|18]/adc_array_circuit_150n_0/vint2 col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4736 adc_array_wafflecap_8_8_0[0|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4737 adc_array_wafflecap_8_8_0[12|27]/adc_array_circuit_150n_0/vdrv row_n[13] adc_array_wafflecap_8_8_0[12|27]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4738 adc_array_wafflecap_8_8_0[6|1]/adc_array_circuit_150n_0/vdrv row_n[7] adc_array_wafflecap_8_8_0[6|1]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4739 adc_array_wafflecap_8_8_0[6|7]/adc_array_circuit_150n_0/vint2 rowon_n[7] adc_array_wafflecap_8_8_0[6|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4740 vcm adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4741 adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4742 adc_array_wafflecap_8_8_0[6|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4743 adc_array_wafflecap_8_8_0[5|14]/adc_array_circuit_150n_0/vdrv row_n[6] adc_array_wafflecap_8_8_0[5|14]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4744 adc_array_wafflecap_8_8_0[11|17]/adc_array_circuit_150n_0/vint1 col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4745 adc_array_wafflecap_8_Dummy_4[30]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4746 vcm adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|7]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4747 adc_array_wafflecap_8_8_0[12|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4748 vcm adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|30]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4749 adc_array_wafflecap_8_8_0[7|18]/adc_array_circuit_150n_0/vdrv row_n[8] adc_array_wafflecap_8_8_0[7|18]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4750 VSS row_n[8] adc_array_wafflecap_8_8_0[7|25]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4751 VSS en_C0_n adc_array_wafflecap_8_1_1/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4752 adc_array_wafflecap_8_8_1[9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4753 adc_array_wafflecap_8_8_0[0|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4754 adc_array_wafflecap_8_8_0[1|27]/adc_array_circuit_150n_0/vint2 col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4755 vcm adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|16]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4756 adc_array_wafflecap_8_8_0[11|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4757 VDD rowon_n[7] adc_array_wafflecap_8_8_0[6|7]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4758 adc_array_wafflecap_8_Dummy_3[1]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4759 vcm adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|6]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4760 VDD rowon_n[10] adc_array_wafflecap_8_8_0[9|24]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4761 adc_array_wafflecap_8_8_0[1|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4762 adc_array_wafflecap_8_8_0[4|27]/adc_array_circuit_150n_0/vint2 rowon_n[5] adc_array_wafflecap_8_8_0[4|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4763 adc_array_wafflecap_8_8_0[0|16]/adc_array_circuit_150n_0/vint2 col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4764 adc_array_wafflecap_8_8_0[14|26]/adc_array_circuit_150n_0/vint2 rowon_n[15] adc_array_wafflecap_8_8_0[14|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4765 VSS row_n[7] adc_array_wafflecap_8_8_0[6|8]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4766 adc_array_wafflecap_8_8_0[1|27]/adc_array_circuit_150n_0/vdrv row_n[2] adc_array_wafflecap_8_8_0[1|27]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4767 adc_array_wafflecap_8_8_0[12|23]/adc_array_circuit_150n_0/vint2 col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4768 adc_array_wafflecap_8_8_0[3|20]/adc_array_circuit_150n_0/vint1 col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4769 vcm VSS adc_array_wafflecap_8_Dummy_1[3]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4770 adc_array_wafflecap_8_8_1[3]/adc_array_circuit_150n_0/vdrv row_n[0] adc_array_wafflecap_8_8_1[3]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4771 adc_array_wafflecap_8_8_0[13|8]/adc_array_circuit_150n_0/vint2 rowon_n[14] adc_array_wafflecap_8_8_0[13|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4772 adc_array_wafflecap_8_8_0[13|30]/adc_array_circuit_150n_0/vint2 rowon_n[14] adc_array_wafflecap_8_8_0[13|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4773 VSS row_n[11] adc_array_wafflecap_8_8_0[10|27]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4774 adc_array_wafflecap_8_8_0[3|18]/adc_array_circuit_150n_0/vdrv row_n[4] adc_array_wafflecap_8_8_0[3|18]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4775 adc_array_wafflecap_8_8_0[3|19]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|19]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4776 vcm VSS adc_array_wafflecap_8_Dummy_4[19]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4777 VDD rowon_n[5] adc_array_wafflecap_8_8_0[4|12]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4778 adc_array_wafflecap_8_8_0[14|22]/adc_array_circuit_150n_0/vint1 col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4779 adc_array_wafflecap_8_8_0[12|10]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|10]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4780 adc_array_wafflecap_8_8_0[7|14]/adc_array_circuit_150n_0/vint2 col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4781 adc_array_wafflecap_8_8_0[3|4]/adc_array_circuit_150n_0/vint2 rowon_n[4] adc_array_wafflecap_8_8_0[3|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4782 adc_array_wafflecap_8_2_0/adc_array_circuit_150n_0/vdrv en_n_bit[1] adc_array_wafflecap_8_2_0/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4783 VSS VSS adc_array_wafflecap_8_Dummy_2[6]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4784 adc_array_wafflecap_8_8_0[12|0]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|0]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4785 VDD rowon_n[13] adc_array_wafflecap_8_8_0[12|26]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4786 adc_array_wafflecap_8_8_0[7|4]/adc_array_circuit_150n_0/vint2 col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4787 adc_array_wafflecap_8_8_0[6|8]/adc_array_circuit_150n_0/vint1 col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4788 adc_array_wafflecap_8_8_0[6|16]/adc_array_circuit_150n_0/vint2 rowon_n[7] adc_array_wafflecap_8_8_0[6|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4789 adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/vint2 rowon_n[3] adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4790 VSS row_n[3] adc_array_wafflecap_8_8_0[2|22]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4791 VDD rowon_n[12] adc_array_wafflecap_8_8_0[11|17]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4792 adc_array_wafflecap_8_8_0[10|23]/adc_array_circuit_150n_0/vdrv row_n[11] adc_array_wafflecap_8_8_0[10|23]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4793 adc_array_wafflecap_8_8_0[8|27]/adc_array_circuit_150n_0/vint1 col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4794 adc_array_wafflecap_8_8_0[7|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4795 VSS row_n[6] adc_array_wafflecap_8_8_0[5|0]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4796 adc_array_wafflecap_8_8_0[9|13]/adc_array_circuit_150n_0/vint1 col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4797 vcm adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|22]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4798 adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4799 adc_array_wafflecap_8_8_0[5|24]/adc_array_circuit_150n_0/vint1 col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4800 adc_array_wafflecap_8_8_0[5|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4801 adc_array_wafflecap_8_8_0[13|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4802 adc_array_wafflecap_8_8_0[9|3]/adc_array_circuit_150n_0/vint1 col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4803 adc_array_wafflecap_8_8_0[0|22]/adc_array_circuit_150n_0/vint1 col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4804 VDD rowon_n[7] adc_array_wafflecap_8_8_0[6|16]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4805 vcm adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[20]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4806 VDD rowon_n[1] adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4807 adc_array_wafflecap_8_Dummy_4[6]/adc_array_circuit_150n_0/vint2 col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4808 adc_array_wafflecap_8_Dummy_4[16]/adc_array_circuit_150n_0/vint2 col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4809 adc_array_wafflecap_8_8_0[10|16]/adc_array_circuit_150n_0/vint2 col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4810 VSS sample_n adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4811 adc_array_wafflecap_8_8_0[7|25]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|25]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4812 vcm adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|11]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4813 adc_array_wafflecap_8_8_0[4|13]/adc_array_circuit_150n_0/vint1 col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4814 adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/vint2 col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4815 VSS row_n[4] adc_array_wafflecap_8_8_0[3|5]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4816 adc_array_wafflecap_8_8_0[14|1]/adc_array_circuit_150n_0/vdrv row_n[15] adc_array_wafflecap_8_8_0[14|1]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4817 adc_array_wafflecap_8_8_0[14|11]/adc_array_circuit_150n_0/vdrv row_n[15] adc_array_wafflecap_8_8_0[14|11]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4818 adc_array_wafflecap_8_8_0[12|22]/adc_array_circuit_150n_0/vint2 rowon_n[13] adc_array_wafflecap_8_8_0[12|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4819 VSS row_n[1] adc_array_wafflecap_8_8_0[0|26]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4820 adc_array_wafflecap_8_8_0[6|18]/adc_array_circuit_150n_0/vint2 rowon_n[7] adc_array_wafflecap_8_8_0[6|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4821 adc_array_wafflecap_8_8_0[13|5]/adc_array_circuit_150n_0/vdrv row_n[14] adc_array_wafflecap_8_8_0[13|5]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4822 adc_array_wafflecap_8_8_0[13|15]/adc_array_circuit_150n_0/vdrv row_n[14] adc_array_wafflecap_8_8_0[13|15]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4823 adc_array_wafflecap_8_8_0[13|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4824 adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4825 adc_array_wafflecap_8_8_0[9|29]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|29]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4826 adc_array_wafflecap_8_8_0[8|16]/adc_array_circuit_150n_0/vdrv row_n[9] adc_array_wafflecap_8_8_0[8|16]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4827 VSS row_n[9] adc_array_wafflecap_8_8_0[8|23]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4828 vcm adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|5]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4829 vcm adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|15]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4830 VSS row_n[7] adc_array_wafflecap_8_8_0[6|16]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4831 vcm adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|14]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4832 adc_array_wafflecap_8_8_0[11|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4833 adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/vdrv row_n[7] adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4834 vcm adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|3]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4835 adc_array_wafflecap_8_8_0[3|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4836 vcm adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|4]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4837 vcm adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|4]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4838 vcm adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|16]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4839 VDD rowon_n[11] adc_array_wafflecap_8_8_0[10|22]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4840 adc_array_wafflecap_8_Dummy_3[1]/adc_array_circuit_150n_0/vint1 col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4841 adc_array_wafflecap_8_8_0[7|22]/adc_array_circuit_150n_0/vint2 col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4842 VDD rowon_n[7] adc_array_wafflecap_8_8_0[6|18]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4843 VDD rowon_n[3] adc_array_wafflecap_8_8_0[2|19]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4844 adc_array_wafflecap_8_8_0[2|7]/adc_array_circuit_150n_0/vdrv row_n[3] adc_array_wafflecap_8_8_0[2|7]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4845 adc_array_wafflecap_8_8_0[2|8]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|8]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4846 adc_array_wafflecap_8_Dummy_1[0]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_1[0]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4847 adc_array_wafflecap_8_8_0[13|21]/adc_array_circuit_150n_0/vint2 col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4848 vcm adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|17]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4849 adc_array_wafflecap_8_8_0[6|16]/adc_array_circuit_150n_0/vint1 col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4850 adc_array_wafflecap_8_8_0[2|17]/adc_array_circuit_150n_0/vint1 col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4851 adc_array_wafflecap_8_8_0[2|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4852 adc_array_wafflecap_8_8_0[9|21]/adc_array_circuit_150n_0/vint1 col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4853 VDD rowon_n[12] adc_array_wafflecap_8_8_0[11|5]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4854 VDD rowon_n[12] adc_array_wafflecap_8_8_0[11|15]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4855 adc_array_wafflecap_8_Dummy_4[21]/adc_array_circuit_150n_0/vint1 col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4856 adc_array_wafflecap_8_8_0[13|8]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|8]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4857 VSS row_n[12] adc_array_wafflecap_8_8_0[11|15]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4858 adc_array_wafflecap_8_8_0[9|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4859 VSS row_n[12] adc_array_wafflecap_8_8_0[11|5]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4860 adc_array_wafflecap_8_8_0[8|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4861 adc_array_wafflecap_8_8_0[5|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4862 VDD rowon_n[5] adc_array_wafflecap_8_8_0[4|23]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4863 adc_array_wafflecap_8_8_0[1|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4864 adc_array_wafflecap_8_8_0[0|13]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|13]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4865 VDD sample adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4866 adc_array_wafflecap_8_8_0[4|12]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|12]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4867 VDD rowon_n[0] adc_array_wafflecap_8_8_1[20]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4868 adc_array_wafflecap_8_8_0[5|20]/adc_array_circuit_150n_0/vint2 col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4869 adc_array_wafflecap_8_8_0[1|21]/adc_array_circuit_150n_0/vint2 col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4870 VSS row_n[6] adc_array_wafflecap_8_8_0[5|30]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4871 adc_array_wafflecap_8_8_0[4|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4872 vcm adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|22]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4873 adc_array_wafflecap_8_8_0[9|10]/adc_array_circuit_150n_0/vdrv row_n[10] adc_array_wafflecap_8_8_0[9|10]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4874 adc_array_wafflecap_8_8_0[8|23]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|23]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4875 adc_array_wafflecap_8_8_0[7|21]/adc_array_circuit_150n_0/vint2 rowon_n[8] adc_array_wafflecap_8_8_0[7|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4876 adc_array_wafflecap_8_8_0[9|0]/adc_array_circuit_150n_0/vdrv row_n[10] adc_array_wafflecap_8_8_0[9|0]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4877 adc_array_wafflecap_8_8_0[3|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4878 adc_array_wafflecap_8_8_1[4]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[4]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4879 adc_array_wafflecap_8_Dummy_4[10]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[10]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4880 adc_array_wafflecap_8_8_0[12|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4881 adc_array_wafflecap_8_8_0[7|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4882 adc_array_wafflecap_8_8_0[7|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4883 adc_array_wafflecap_8_8_0[6|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4884 VSS row_n[2] adc_array_wafflecap_8_8_0[1|6]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4885 adc_array_wafflecap_8_Dummy_4[0]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[0]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4886 adc_array_wafflecap_8_8_0[12|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4887 VSS sample_n adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4888 vcm adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|9]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4889 adc_array_wafflecap_8_8_0[11|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4890 vcm adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|13]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4891 adc_array_wafflecap_8_8_0[4|9]/adc_array_circuit_150n_0/vint2 col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4892 adc_array_wafflecap_8_Dummy_2[2]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4893 adc_array_wafflecap_8_8_0[1|21]/adc_array_circuit_150n_0/vdrv row_n[2] adc_array_wafflecap_8_8_0[1|21]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4894 adc_array_wafflecap_8_Dummy_4[27]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[27]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4895 adc_array_wafflecap_8_8_0[13|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4896 adc_array_wafflecap_8_8_0[11|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4897 vcm adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|3]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4898 adc_array_wafflecap_8_Dummy_2[0]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_2[0]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4899 adc_array_wafflecap_8_8_1[2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_1[2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4900 vcm adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|29]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4901 adc_array_wafflecap_8_8_0[3|25]/adc_array_circuit_150n_0/vint2 col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4902 adc_array_wafflecap_8_8_0[6|3]/adc_array_circuit_150n_0/vint2 col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4903 adc_array_wafflecap_8_8_0[2|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4904 VSS row_n[13] adc_array_wafflecap_8_8_0[12|19]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4905 adc_array_wafflecap_8_8_0[14|3]/adc_array_circuit_150n_0/vint2 rowon_n[15] adc_array_wafflecap_8_8_0[14|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4906 adc_array_wafflecap_8_8_0[14|13]/adc_array_circuit_150n_0/vint2 rowon_n[15] adc_array_wafflecap_8_8_0[14|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4907 adc_array_wafflecap_8_8_0[8|20]/adc_array_circuit_150n_0/vint2 col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4908 adc_array_wafflecap_8_8_0[1|6]/adc_array_circuit_150n_0/vint1 col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4909 VDD rowon_n[15] adc_array_wafflecap_8_8_0[14|18]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4910 VSS row_n[8] adc_array_wafflecap_8_8_0[7|0]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4911 VSS row_n[8] adc_array_wafflecap_8_8_0[7|10]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4912 adc_array_wafflecap_8_8_0[2|14]/adc_array_circuit_150n_0/vint2 col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4913 adc_array_wafflecap_8_8_0[10|19]/adc_array_circuit_150n_0/vint1 col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4914 adc_array_wafflecap_8_8_0[6|27]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|27]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4915 adc_array_wafflecap_8_8_0[6|9]/adc_array_circuit_150n_0/vint2 rowon_n[7] adc_array_wafflecap_8_8_0[6|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4916 adc_array_wafflecap_8_8_0[3|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4917 adc_array_wafflecap_8_8_0[2|4]/adc_array_circuit_150n_0/vdrv row_n[3] adc_array_wafflecap_8_8_0[2|4]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4918 VDD rowon_n[13] adc_array_wafflecap_8_8_0[12|13]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4919 adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/vint1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4920 adc_array_wafflecap_8_8_0[6|3]/adc_array_circuit_150n_0/vdrv row_n[7] adc_array_wafflecap_8_8_0[6|3]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4921 VDD rowon_n[13] adc_array_wafflecap_8_8_0[12|3]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4922 adc_array_wafflecap_8_8_0[13|19]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|19]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4923 VDD rowon_n[6] adc_array_wafflecap_8_8_0[5|27]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4924 adc_array_wafflecap_8_8_0[0|14]/adc_array_circuit_150n_0/vdrv row_n[1] adc_array_wafflecap_8_8_0[0|14]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4925 adc_array_wafflecap_8_8_1[11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4926 adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n sample VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4927 VSS VDD adc_array_wafflecap_8_Dummy_4[12]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4928 adc_array_wafflecap_8_8_0[12|8]/adc_array_circuit_150n_0/vint2 col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4929 VSS VDD adc_array_wafflecap_8_Dummy_4[2]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4930 adc_array_wafflecap_8_8_0[7|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4931 VDD rowon_n[7] adc_array_wafflecap_8_8_0[6|9]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4932 adc_array_wafflecap_8_8_0[5|1]/adc_array_circuit_150n_0/vint2 rowon_n[6] adc_array_wafflecap_8_8_0[5|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4933 adc_array_wafflecap_8_8_0[1|2]/adc_array_circuit_150n_0/vint2 rowon_n[2] adc_array_wafflecap_8_8_0[1|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4934 adc_array_wafflecap_8_8_0[14|30]/adc_array_circuit_150n_0/vdrv row_n[15] adc_array_wafflecap_8_8_0[14|30]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4935 adc_array_wafflecap_8_8_0[11|2]/adc_array_circuit_150n_0/vint2 col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4936 adc_array_wafflecap_8_8_0[11|12]/adc_array_circuit_150n_0/vint2 col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4937 VSS row_n[5] adc_array_wafflecap_8_8_0[4|19]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4938 VSS row_n[1] adc_array_wafflecap_8_8_0[0|20]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4939 adc_array_wafflecap_8_8_0[1|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4940 adc_array_wafflecap_8_8_0[4|29]/adc_array_circuit_150n_0/vint2 rowon_n[5] adc_array_wafflecap_8_8_0[4|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4941 adc_array_wafflecap_8_8_0[14|7]/adc_array_circuit_150n_0/vint1 col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4942 VSS row_n[7] adc_array_wafflecap_8_8_0[6|10]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4943 adc_array_wafflecap_8_8_0[4|17]/adc_array_circuit_150n_0/vint2 col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4944 adc_array_wafflecap_8_8_0[0|18]/adc_array_circuit_150n_0/vint2 col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4945 vcm adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|29]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4946 adc_array_wafflecap_8_8_0[3|22]/adc_array_circuit_150n_0/vint1 col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4947 adc_array_wafflecap_8_8_0[14|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4948 adc_array_wafflecap_8_8_0[13|1]/adc_array_circuit_150n_0/vint1 col_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4949 adc_array_wafflecap_8_8_0[13|11]/adc_array_circuit_150n_0/vint1 col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4950 adc_array_wafflecap_8_8_0[10|8]/adc_array_circuit_150n_0/vdrv row_n[11] adc_array_wafflecap_8_8_0[10|8]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4951 adc_array_wafflecap_8_8_0[8|19]/adc_array_circuit_150n_0/vint2 rowon_n[9] adc_array_wafflecap_8_8_0[8|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4952 adc_array_wafflecap_8_8_0[7|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4953 adc_array_wafflecap_8_8_0[7|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4954 adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/vint2 rowon_n[8] adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4955 adc_array_wafflecap_8_8_0[3|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4956 VDD rowon_n[4] adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4957 adc_array_wafflecap_8_8_0[13|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4958 adc_array_wafflecap_8_8_0[10|25]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|25]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4959 adc_array_wafflecap_8_Dummy_2[3]/adc_array_circuit_150n_0/vint1 col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4960 VDD rowon_n[2] adc_array_wafflecap_8_8_0[1|2]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4961 adc_array_wafflecap_8_8_0[13|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4962 VDD rowon_n[5] adc_array_wafflecap_8_8_0[4|14]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4963 adc_array_wafflecap_8_8_0[3|6]/adc_array_circuit_150n_0/vint2 rowon_n[4] adc_array_wafflecap_8_8_0[3|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4964 adc_array_wafflecap_8_Dummy_2[1]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_2[1]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4965 adc_array_wafflecap_8_8_0[9|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4966 VSS VSS adc_array_wafflecap_8_Dummy_3[0]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4967 VSS row_n[3] adc_array_wafflecap_8_8_0[2|24]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4968 adc_array_wafflecap_8_8_0[9|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4969 adc_array_wafflecap_8_8_0[6|10]/adc_array_circuit_150n_0/vint1 col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4970 VSS row_n[6] adc_array_wafflecap_8_8_0[5|2]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4971 vcm adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|9]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4972 VDD rowon_n[0] adc_array_wafflecap_8_8_1[11]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4973 VSS row_n[2] adc_array_wafflecap_8_8_0[1|3]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4974 adc_array_wafflecap_8_8_0[7|0]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|0]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4975 adc_array_wafflecap_8_8_0[7|10]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|10]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4976 adc_array_wafflecap_8_Dummy_4[12]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4977 VSS row_n[13] adc_array_wafflecap_8_8_0[12|30]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4978 adc_array_wafflecap_8_Dummy_4[2]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4979 VDD sample adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4980 adc_array_wafflecap_8_8_0[13|27]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|27]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4981 adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/vint2 col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4982 vcm adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[22]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4983 adc_array_wafflecap_8_8_0[0|24]/adc_array_circuit_150n_0/vint1 col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4984 adc_array_wafflecap_8_8_0[14|13]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|13]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4985 VSS row_n[9] adc_array_wafflecap_8_8_0[8|8]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4986 adc_array_wafflecap_8_8_0[4|29]/adc_array_circuit_150n_0/vdrv row_n[5] adc_array_wafflecap_8_8_0[4|29]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4987 adc_array_wafflecap_8_8_0[1|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4988 adc_array_wafflecap_8_8_0[14|3]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|3]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4989 VDD rowon_n[15] adc_array_wafflecap_8_8_0[14|7]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4990 VDD rowon_n[15] adc_array_wafflecap_8_8_0[14|29]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4991 adc_array_wafflecap_8_8_0[12|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4992 adc_array_wafflecap_8_8_0[1|3]/adc_array_circuit_150n_0/vint1 col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4993 vcm adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|1]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4994 vcm adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|13]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4995 adc_array_wafflecap_8_8_0[4|15]/adc_array_circuit_150n_0/vint1 col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4996 vcm adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|14]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4997 VDD rowon_n[14] adc_array_wafflecap_8_8_0[13|11]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4998 adc_array_wafflecap_8_8_0[10|30]/adc_array_circuit_150n_0/vint1 col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4999 VDD rowon_n[14] adc_array_wafflecap_8_8_0[13|1]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5000 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.64e+07u l=1.6e+07u
X5001 adc_array_wafflecap_8_8_0[7|7]/adc_array_circuit_150n_0/vint2 col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5002 adc_array_wafflecap_8_8_0[6|20]/adc_array_circuit_150n_0/vint2 rowon_n[7] adc_array_wafflecap_8_8_0[6|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5003 adc_array_wafflecap_8_8_1[12]/adc_array_circuit_150n_0/vint1 col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5004 adc_array_wafflecap_8_8_0[13|6]/adc_array_circuit_150n_0/vint2 col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5005 adc_array_wafflecap_8_8_0[12|19]/adc_array_circuit_150n_0/vint2 col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5006 adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5007 adc_array_wafflecap_8_8_1[18]/adc_array_circuit_150n_0/vint2 rowon_n[0] adc_array_wafflecap_8_8_1[18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5008 adc_array_wafflecap_8_8_0[9|6]/adc_array_circuit_150n_0/vint1 col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5009 adc_array_wafflecap_8_8_0[8|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5010 adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5011 vcm adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|5]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5012 adc_array_wafflecap_8_8_1[6]/adc_array_circuit_150n_0/vint2 col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5013 vcm adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|6]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5014 adc_array_wafflecap_8_Dummy_4[29]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[29]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5015 adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5016 vcm adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|28]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5017 VSS row_n[0] adc_array_wafflecap_8_8_1[16]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5018 adc_array_wafflecap_8_8_0[3|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5019 adc_array_wafflecap_8_8_0[14|18]/adc_array_circuit_150n_0/vint1 col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5020 vcm adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5021 VDD rowon_n[7] adc_array_wafflecap_8_8_0[6|20]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5022 VDD rowon_n[3] adc_array_wafflecap_8_8_0[2|21]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5023 adc_array_wafflecap_8_8_0[8|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5024 vcm adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|17]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5025 adc_array_wafflecap_8_8_0[2|10]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|10]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5026 adc_array_wafflecap_8_Dummy_1[2]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_1[2]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5027 adc_array_wafflecap_8_Dummy_4[23]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5028 adc_array_wafflecap_8_8_0[10|19]/adc_array_circuit_150n_0/vdrv row_n[11] adc_array_wafflecap_8_8_0[10|19]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5029 adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5030 adc_array_wafflecap_8_8_0[11|23]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|23]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5031 VSS row_n[4] adc_array_wafflecap_8_8_0[3|28]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5032 adc_array_wafflecap_8_8_0[2|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5033 adc_array_wafflecap_8_8_0[10|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5034 adc_array_wafflecap_8_8_0[10|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5035 adc_array_wafflecap_8_8_0[10|10]/adc_array_circuit_150n_0/vint2 rowon_n[11] adc_array_wafflecap_8_8_0[10|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5036 adc_array_wafflecap_8_8_0[9|25]/adc_array_circuit_150n_0/vint2 col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5037 VSS row_n[8] adc_array_wafflecap_8_8_0[7|29]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5038 adc_array_wafflecap_8_8_0[1|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5039 adc_array_wafflecap_8_8_0[10|0]/adc_array_circuit_150n_0/vint2 rowon_n[11] adc_array_wafflecap_8_8_0[10|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5040 adc_array_wafflecap_8_8_0[8|8]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|8]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5041 adc_array_wafflecap_8_8_0[6|21]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|21]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5042 VDD rowon_n[5] adc_array_wafflecap_8_8_0[4|25]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5043 adc_array_wafflecap_8_Dummy_4[25]/adc_array_circuit_150n_0/vint2 col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5044 vcm adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|7]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5045 VSS row_n[14] adc_array_wafflecap_8_8_0[13|28]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5046 adc_array_wafflecap_8_8_0[0|15]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|15]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5047 VDD rowon_n[0] adc_array_wafflecap_8_8_1[22]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5048 adc_array_wafflecap_8_8_0[11|24]/adc_array_circuit_150n_0/vint1 col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5049 adc_array_wafflecap_8_8_0[9|2]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|2]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5050 adc_array_wafflecap_8_8_0[9|12]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|12]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5051 VDD rowon_n[10] adc_array_wafflecap_8_8_0[9|28]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5052 adc_array_wafflecap_8_8_0[1|23]/adc_array_circuit_150n_0/vint2 col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5053 adc_array_wafflecap_8_Dummy_4[12]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[12]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5054 VDD VDD adc_array_wafflecap_8_Dummy_4[28]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5055 VDD rowon_n[9] adc_array_wafflecap_8_8_0[8|10]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5056 adc_array_wafflecap_8_8_0[7|25]/adc_array_circuit_150n_0/vdrv row_n[8] adc_array_wafflecap_8_8_0[7|25]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5057 adc_array_wafflecap_8_8_0[5|9]/adc_array_circuit_150n_0/vdrv row_n[6] adc_array_wafflecap_8_8_0[5|9]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5058 adc_array_wafflecap_8_8_0[5|22]/adc_array_circuit_150n_0/vint2 col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5059 VSS row_n[6] adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5060 adc_array_wafflecap_8_8_0[4|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5061 adc_array_wafflecap_8_8_0[0|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5062 adc_array_wafflecap_8_Dummy_4[2]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[2]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5063 VDD rowon_n[9] adc_array_wafflecap_8_8_0[8|0]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5064 adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5065 adc_array_wafflecap_8_8_0[13|24]/adc_array_circuit_150n_0/vdrv row_n[14] adc_array_wafflecap_8_8_0[13|24]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5066 adc_array_wafflecap_8_8_0[12|27]/adc_array_circuit_150n_0/vint2 col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5067 vcm adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|24]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5068 adc_array_wafflecap_8_8_0[6|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5069 adc_array_wafflecap_8_8_0[14|26]/adc_array_circuit_150n_0/vint1 col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5070 adc_array_wafflecap_8_8_0[7|18]/adc_array_circuit_150n_0/vint2 col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5071 adc_array_wafflecap_8_8_0[4|11]/adc_array_circuit_150n_0/vint2 col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5072 adc_array_wafflecap_8_Dummy_2[4]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5073 adc_array_wafflecap_8_8_0[1|23]/adc_array_circuit_150n_0/vdrv row_n[2] adc_array_wafflecap_8_8_0[1|23]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5074 adc_array_wafflecap_8_8_0[10|27]/adc_array_circuit_150n_0/vdrv row_n[11] adc_array_wafflecap_8_8_0[10|27]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5075 adc_array_wafflecap_8_8_0[4|1]/adc_array_circuit_150n_0/vdrv row_n[5] adc_array_wafflecap_8_8_0[4|1]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5076 adc_array_wafflecap_8_8_1[4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_1[4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5077 adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5078 vcm adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5079 adc_array_wafflecap_8_8_0[3|14]/adc_array_circuit_150n_0/vdrv row_n[4] adc_array_wafflecap_8_8_0[3|14]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5080 vcm VSS adc_array_wafflecap_8_Dummy_4[26]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5081 adc_array_wafflecap_8_8_0[11|13]/adc_array_circuit_150n_0/vdrv row_n[12] adc_array_wafflecap_8_8_0[11|13]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5082 adc_array_wafflecap_8_8_0[9|17]/adc_array_circuit_150n_0/vint1 col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5083 adc_array_wafflecap_8_8_0[9|24]/adc_array_circuit_150n_0/vint2 rowon_n[10] adc_array_wafflecap_8_8_0[9|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5084 adc_array_wafflecap_8_8_0[8|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5085 adc_array_wafflecap_8_8_0[6|5]/adc_array_circuit_150n_0/vint2 col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5086 adc_array_wafflecap_8_8_0[13|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5087 adc_array_wafflecap_8_8_0[11|3]/adc_array_circuit_150n_0/vdrv row_n[12] adc_array_wafflecap_8_8_0[11|3]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5088 vcm VSS adc_array_wafflecap_8_Dummy_8[5]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5089 adc_array_wafflecap_8_8_0[10|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5090 adc_array_wafflecap_8_Dummy_2[0]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_2[0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5091 adc_array_wafflecap_8_8_0[14|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5092 adc_array_wafflecap_8_8_0[14|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5093 adc_array_wafflecap_8_8_1[3]/adc_array_circuit_150n_0/vint2 col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5094 vcm adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|16]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5095 VDD rowon_n[5] adc_array_wafflecap_8_8_0[4|7]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5096 vcm adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|6]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5097 VDD rowon_n[8] adc_array_wafflecap_8_8_0[7|24]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5098 adc_array_wafflecap_8_8_0[6|5]/adc_array_circuit_150n_0/vdrv row_n[7] adc_array_wafflecap_8_8_0[6|5]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5099 adc_array_wafflecap_8_8_0[6|11]/adc_array_circuit_150n_0/vint2 rowon_n[7] adc_array_wafflecap_8_8_0[6|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5100 adc_array_wafflecap_8_8_0[2|27]/adc_array_circuit_150n_0/vint2 rowon_n[3] adc_array_wafflecap_8_8_0[2|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5101 adc_array_wafflecap_8_2_0/adc_array_circuit_150n_0/vint2 en_n_bit[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5102 VSS row_n[15] adc_array_wafflecap_8_8_0[14|22]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5103 adc_array_wafflecap_8_8_0[12|26]/adc_array_circuit_150n_0/vint2 rowon_n[13] adc_array_wafflecap_8_8_0[12|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X5104 adc_array_wafflecap_8_8_0[10|23]/adc_array_circuit_150n_0/vint2 col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5105 adc_array_wafflecap_8_8_0[6|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5106 adc_array_wafflecap_8_8_0[5|19]/adc_array_circuit_150n_0/vint1 col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5107 adc_array_wafflecap_8_8_0[5|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5108 adc_array_wafflecap_8_8_1[27]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[27]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5109 adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5110 adc_array_wafflecap_8_8_0[11|8]/adc_array_circuit_150n_0/vint2 rowon_n[12] adc_array_wafflecap_8_8_0[11|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5111 adc_array_wafflecap_8_8_0[11|30]/adc_array_circuit_150n_0/vint2 rowon_n[12] adc_array_wafflecap_8_8_0[11|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5112 VSS row_n[9] adc_array_wafflecap_8_8_0[8|27]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5113 VDD rowon_n[6] adc_array_wafflecap_8_8_0[5|29]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5114 adc_array_wafflecap_8_8_1[13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5115 adc_array_wafflecap_8_8_0[8|19]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|19]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5116 adc_array_wafflecap_8_8_0[5|17]/adc_array_circuit_150n_0/vdrv row_n[6] adc_array_wafflecap_8_8_0[5|17]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X5117 adc_array_wafflecap_8_8_0[5|18]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|18]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5118 adc_array_wafflecap_8_8_0[1|19]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|19]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5119 adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5120 adc_array_wafflecap_8_8_0[14|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5121 vcm adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|18]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5122 VSS row_n[10] adc_array_wafflecap_8_8_0[9|3]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5123 VSS row_n[10] adc_array_wafflecap_8_8_0[9|13]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5124 VDD rowon_n[7] adc_array_wafflecap_8_8_0[6|11]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5125 VDD rowon_n[3] adc_array_wafflecap_8_8_0[2|12]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5126 VDD rowon_n[1] adc_array_wafflecap_8_8_0[0|27]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5127 adc_array_wafflecap_8_8_0[1|4]/adc_array_circuit_150n_0/vint2 rowon_n[2] adc_array_wafflecap_8_8_0[1|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5128 VDD VDD adc_array_wafflecap_8_Dummy_4[26]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5129 adc_array_wafflecap_8_8_0[12|22]/adc_array_circuit_150n_0/vint1 col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5130 adc_array_wafflecap_8_8_0[10|10]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|10]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5131 adc_array_wafflecap_8_8_0[5|3]/adc_array_circuit_150n_0/vint2 rowon_n[6] adc_array_wafflecap_8_8_0[5|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5132 VDD rowon_n[15] adc_array_wafflecap_8_8_0[14|16]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5133 adc_array_wafflecap_8_8_0[10|0]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|0]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5134 VDD rowon_n[11] adc_array_wafflecap_8_8_0[10|26]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5135 adc_array_wafflecap_8_8_0[6|26]/adc_array_circuit_150n_0/vint2 col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5136 adc_array_wafflecap_8_8_0[4|8]/adc_array_circuit_150n_0/vint1 col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5137 VSS row_n[5] adc_array_wafflecap_8_8_0[4|21]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5138 adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/vint2 rowon_n[1] adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5139 VSS row_n[1] adc_array_wafflecap_8_8_0[0|22]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5140 VDD rowon_n[15] adc_array_wafflecap_8_8_0[14|6]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5141 VDD rowon_n[10] adc_array_wafflecap_8_8_0[9|17]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5142 adc_array_wafflecap_8_8_0[8|23]/adc_array_circuit_150n_0/vdrv row_n[9] adc_array_wafflecap_8_8_0[8|23]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5143 adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/vint2 rowon_n[5] adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5144 VSS row_n[4] adc_array_wafflecap_8_8_0[3|0]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5145 VSS row_n[7] adc_array_wafflecap_8_8_0[6|12]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5146 adc_array_wafflecap_8_8_0[7|13]/adc_array_circuit_150n_0/vint1 col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5147 adc_array_wafflecap_8_8_0[3|24]/adc_array_circuit_150n_0/vint1 col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5148 adc_array_wafflecap_8_8_0[3|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5149 adc_array_wafflecap_8_8_0[11|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5150 adc_array_wafflecap_8_8_0[7|3]/adc_array_circuit_150n_0/vint1 col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5151 adc_array_wafflecap_8_8_0[6|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5152 adc_array_wafflecap_8_8_0[14|11]/adc_array_circuit_150n_0/vint2 col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5153 adc_array_wafflecap_8_Dummy_2[5]/adc_array_circuit_150n_0/vint1 col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5154 VDD rowon_n[2] adc_array_wafflecap_8_8_0[1|4]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5155 adc_array_wafflecap_8_8_0[14|1]/adc_array_circuit_150n_0/vint2 col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5156 VDD rowon_n[5] adc_array_wafflecap_8_8_0[4|16]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5157 VDD VSS adc_array_wafflecap_8_Dummy_6/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5158 adc_array_wafflecap_8_8_0[13|5]/adc_array_circuit_150n_0/vint2 col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5159 adc_array_wafflecap_8_8_0[13|15]/adc_array_circuit_150n_0/vint2 col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5160 adc_array_wafflecap_8_8_0[8|16]/adc_array_circuit_150n_0/vint2 col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5161 adc_array_wafflecap_8_8_0[6|26]/adc_array_circuit_150n_0/vdrv row_n[7] adc_array_wafflecap_8_8_0[6|26]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5162 VSS sample_n adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5163 vcm adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|11]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5164 adc_array_wafflecap_8_8_0[2|13]/adc_array_circuit_150n_0/vint1 col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5165 adc_array_wafflecap_8_8_0[6|12]/adc_array_circuit_150n_0/vint1 col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5166 VSS row_n[6] adc_array_wafflecap_8_8_0[5|4]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5167 VDD rowon_n[0] adc_array_wafflecap_8_8_1[13]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5168 VSS row_n[2] adc_array_wafflecap_8_8_0[1|5]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5169 adc_array_wafflecap_8_Dummy_4[5]/adc_array_circuit_150n_0/vint1 col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5170 adc_array_wafflecap_8_Dummy_4[15]/adc_array_circuit_150n_0/vint1 col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5171 adc_array_wafflecap_8_8_0[12|1]/adc_array_circuit_150n_0/vdrv row_n[13] adc_array_wafflecap_8_8_0[12|1]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5172 adc_array_wafflecap_8_8_0[12|11]/adc_array_circuit_150n_0/vdrv row_n[13] adc_array_wafflecap_8_8_0[12|11]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5173 adc_array_wafflecap_8_8_0[10|22]/adc_array_circuit_150n_0/vint2 rowon_n[11] adc_array_wafflecap_8_8_0[10|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5174 adc_array_wafflecap_8_8_0[9|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5175 adc_array_wafflecap_8_8_0[9|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5176 VSS VSS adc_array_wafflecap_8_Dummy_3[1]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5177 adc_array_wafflecap_8_Dummy_4[14]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5178 adc_array_wafflecap_8_8_0[11|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5179 adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5180 adc_array_wafflecap_8_Dummy_4[4]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5181 vcm adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[24]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5182 vcm adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|14]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5183 adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/vdrv row_n[5] adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5184 vcm VSS adc_array_wafflecap_8_Dummy_8[2]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5185 adc_array_wafflecap_8_8_0[1|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5186 adc_array_wafflecap_8_8_0[1|5]/adc_array_circuit_150n_0/vint1 col_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5187 vcm adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|3]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5188 vcm adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|4]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5189 VSS row_n[10] adc_array_wafflecap_8_8_0[9|21]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5190 adc_array_wafflecap_8_8_0[8|27]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|27]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5191 vcm adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|15]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5192 vcm adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|16]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5193 VDD sample adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5194 VDD rowon_n[9] adc_array_wafflecap_8_8_0[8|22]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5195 VSS VDD adc_array_wafflecap_8_Dummy_4[21]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5196 vcm adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|12]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5197 adc_array_wafflecap_8_8_0[7|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5198 VDD rowon_n[5] adc_array_wafflecap_8_8_0[4|18]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5199 adc_array_wafflecap_8_8_1[28]/adc_array_circuit_150n_0/vdrv row_n[0] adc_array_wafflecap_8_8_1[28]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5200 vcm adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|2]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5201 adc_array_wafflecap_8_8_1[14]/adc_array_circuit_150n_0/vint1 col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5202 adc_array_wafflecap_8_8_0[0|8]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|8]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5203 VDD rowon_n[12] adc_array_wafflecap_8_8_0[11|20]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5204 adc_array_wafflecap_8_8_0[11|21]/adc_array_circuit_150n_0/vint2 col_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5205 vcm adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|17]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5206 adc_array_wafflecap_8_8_0[4|7]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|7]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5207 adc_array_wafflecap_8_8_0[4|16]/adc_array_circuit_150n_0/vint1 col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5208 adc_array_wafflecap_8_8_0[4|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5209 adc_array_wafflecap_8_8_0[0|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5210 adc_array_wafflecap_8_Dummy_4[31]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[31]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5211 adc_array_wafflecap_8_Dummy_4[8]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5212 adc_array_wafflecap_8_8_0[7|21]/adc_array_circuit_150n_0/vint1 col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5213 VDD rowon_n[10] adc_array_wafflecap_8_8_0[9|5]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5214 VDD rowon_n[10] adc_array_wafflecap_8_8_0[9|15]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5215 adc_array_wafflecap_8_8_1[20]/adc_array_circuit_150n_0/vint2 rowon_n[0] adc_array_wafflecap_8_8_1[20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5216 adc_array_wafflecap_8_8_0[13|20]/adc_array_circuit_150n_0/vint1 col_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5217 adc_array_wafflecap_8_8_0[11|8]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|8]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5218 adc_array_wafflecap_8_8_0[7|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5219 VDD VDD adc_array_wafflecap_8_Dummy_4[15]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5220 VDD VDD adc_array_wafflecap_8_Dummy_4[5]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5221 adc_array_wafflecap_8_8_0[3|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5222 VDD rowon_n[3] adc_array_wafflecap_8_8_0[2|23]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5223 adc_array_wafflecap_8_Dummy_7/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_7/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5224 adc_array_wafflecap_8_8_0[9|10]/adc_array_circuit_150n_0/vint2 col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5225 adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5226 adc_array_wafflecap_8_Dummy_1[4]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_1[4]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5227 adc_array_wafflecap_8_8_0[9|0]/adc_array_circuit_150n_0/vint2 col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5228 VDD sample adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5229 adc_array_wafflecap_8_8_0[2|12]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|12]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5230 adc_array_wafflecap_8_Dummy_4[0]/adc_array_circuit_150n_0/vint2 VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5231 adc_array_wafflecap_8_Dummy_4[10]/adc_array_circuit_150n_0/vint2 col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5232 adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/vdrv row_n[12] adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5233 adc_array_wafflecap_8_8_0[11|9]/adc_array_circuit_150n_0/vint1 col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5234 adc_array_wafflecap_8_8_0[3|20]/adc_array_circuit_150n_0/vint2 col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5235 adc_array_wafflecap_8_8_0[2|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5236 adc_array_wafflecap_8_Dummy_4[22]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5237 VSS row_n[4] adc_array_wafflecap_8_8_0[3|30]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5238 vcm adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|22]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5239 adc_array_wafflecap_8_8_0[7|10]/adc_array_circuit_150n_0/vdrv row_n[8] adc_array_wafflecap_8_8_0[7|10]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5240 adc_array_wafflecap_8_8_0[7|0]/adc_array_circuit_150n_0/vdrv row_n[8] adc_array_wafflecap_8_8_0[7|0]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5241 adc_array_wafflecap_8_8_0[1|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5242 adc_array_wafflecap_8_8_0[13|9]/adc_array_circuit_150n_0/vdrv row_n[14] adc_array_wafflecap_8_8_0[13|9]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5243 adc_array_wafflecap_8_8_0[10|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5244 vcm adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|9]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5245 adc_array_wafflecap_8_8_0[6|23]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|23]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5246 adc_array_wafflecap_8_8_0[10|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5247 VSS sample_n adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5248 VDD rowon_n[0] adc_array_wafflecap_8_8_1[24]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5249 adc_array_wafflecap_8_8_0[2|9]/adc_array_circuit_150n_0/vint2 col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5250 adc_array_wafflecap_8_8_0[13|26]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|26]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5251 adc_array_wafflecap_8_8_0[11|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5252 vcm adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|28]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5253 vcm adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|29]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5254 adc_array_wafflecap_8_8_0[14|18]/adc_array_circuit_150n_0/vint2 rowon_n[15] adc_array_wafflecap_8_8_0[14|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5255 adc_array_wafflecap_8_8_0[0|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5256 adc_array_wafflecap_8_8_0[1|25]/adc_array_circuit_150n_0/vint2 col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5257 vcm adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|19]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5258 adc_array_wafflecap_8_8_0[5|11]/adc_array_circuit_150n_0/vdrv row_n[6] adc_array_wafflecap_8_8_0[5|11]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5259 adc_array_wafflecap_8_8_0[4|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5260 VSS row_n[11] adc_array_wafflecap_8_8_0[10|19]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5261 VSS row_n[10] adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5262 adc_array_wafflecap_8_8_0[12|3]/adc_array_circuit_150n_0/vint2 rowon_n[13] adc_array_wafflecap_8_8_0[12|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5263 adc_array_wafflecap_8_8_0[12|13]/adc_array_circuit_150n_0/vint2 rowon_n[13] adc_array_wafflecap_8_8_0[12|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5264 adc_array_wafflecap_8_8_0[0|9]/adc_array_circuit_150n_0/vdrv row_n[1] adc_array_wafflecap_8_8_0[0|9]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5265 vcm VSS adc_array_wafflecap_8_Dummy_4[1]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5266 vcm VSS adc_array_wafflecap_8_Dummy_4[11]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5267 adc_array_wafflecap_8_8_1[6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5268 VDD rowon_n[13] adc_array_wafflecap_8_8_0[12|18]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5269 VDD rowon_n[12] adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5270 adc_array_wafflecap_8_8_0[4|13]/adc_array_circuit_150n_0/vint2 col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5271 adc_array_wafflecap_8_8_0[0|14]/adc_array_circuit_150n_0/vint2 col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5272 VDD rowon_n[12] adc_array_wafflecap_8_8_0[11|9]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5273 adc_array_wafflecap_8_8_0[8|19]/adc_array_circuit_150n_0/vint1 col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5274 adc_array_wafflecap_8_8_0[1|25]/adc_array_circuit_150n_0/vdrv row_n[2] adc_array_wafflecap_8_8_0[1|25]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5275 adc_array_wafflecap_8_8_0[1|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5276 adc_array_wafflecap_8_Dummy_4[19]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5277 VDD rowon_n[11] adc_array_wafflecap_8_8_0[10|13]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5278 adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/vint1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5279 adc_array_wafflecap_8_8_0[4|3]/adc_array_circuit_150n_0/vdrv row_n[5] adc_array_wafflecap_8_8_0[4|3]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5280 adc_array_wafflecap_8_8_0[4|4]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|4]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5281 VDD rowon_n[11] adc_array_wafflecap_8_8_0[10|3]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5282 adc_array_wafflecap_8_8_0[14|30]/adc_array_circuit_150n_0/vint2 col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5283 adc_array_wafflecap_8_8_0[11|19]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|19]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5284 adc_array_wafflecap_8_8_1[0]/adc_array_circuit_150n_0/vdrv row_n[0] adc_array_wafflecap_8_8_1[0]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5285 VSS row_n[15] adc_array_wafflecap_8_8_0[14|7]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X5286 VDD rowon_n[4] adc_array_wafflecap_8_8_0[3|27]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5287 adc_array_wafflecap_8_Dummy_1[5]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_1[5]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5288 VSS row_n[14] adc_array_wafflecap_8_8_0[13|11]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5289 adc_array_wafflecap_8_8_0[10|8]/adc_array_circuit_150n_0/vint2 col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5290 adc_array_wafflecap_8_8_0[14|17]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|17]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5291 VSS row_n[14] adc_array_wafflecap_8_8_0[13|1]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5292 VDD rowon_n[5] adc_array_wafflecap_8_8_0[4|9]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5293 adc_array_wafflecap_8_8_0[3|1]/adc_array_circuit_150n_0/vint2 rowon_n[4] adc_array_wafflecap_8_8_0[3|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5294 adc_array_wafflecap_8_8_0[12|30]/adc_array_circuit_150n_0/vdrv row_n[13] adc_array_wafflecap_8_8_0[12|30]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5295 adc_array_wafflecap_8_8_0[6|13]/adc_array_circuit_150n_0/vint2 rowon_n[7] adc_array_wafflecap_8_8_0[6|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5296 VSS VSS adc_array_wafflecap_8_Dummy_2[3]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5297 VSS row_n[3] adc_array_wafflecap_8_8_0[2|19]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5298 VDD rowon_n[0] adc_array_wafflecap_8_8_1[6]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5299 adc_array_wafflecap_8_8_0[2|29]/adc_array_circuit_150n_0/vint2 rowon_n[3] adc_array_wafflecap_8_8_0[2|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5300 adc_array_wafflecap_8_8_0[12|7]/adc_array_circuit_150n_0/vint1 col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5301 adc_array_wafflecap_8_Dummy_2[1]/adc_array_circuit_150n_0/vint2 col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5302 adc_array_wafflecap_8_8_0[2|17]/adc_array_circuit_150n_0/vint2 col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5303 adc_array_wafflecap_8_Dummy_4[33]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[33]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5304 vcm adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|29]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5305 adc_array_wafflecap_8_8_0[5|21]/adc_array_circuit_150n_0/vint1 col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5306 adc_array_wafflecap_8_8_1[29]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[29]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5307 adc_array_wafflecap_8_8_0[12|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5308 adc_array_wafflecap_8_8_0[9|21]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|21]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5309 adc_array_wafflecap_8_8_0[8|8]/adc_array_circuit_150n_0/vdrv row_n[9] adc_array_wafflecap_8_8_0[8|8]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5310 adc_array_wafflecap_8_8_0[6|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5311 adc_array_wafflecap_8_8_0[5|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5312 VDD rowon_n[6] adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5313 adc_array_wafflecap_8_8_1[11]/adc_array_circuit_150n_0/vint2 rowon_n[0] adc_array_wafflecap_8_8_1[11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5314 adc_array_wafflecap_8_8_0[1|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5315 adc_array_wafflecap_8_8_1[15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5316 adc_array_wafflecap_8_8_0[11|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5317 adc_array_wafflecap_8_8_0[0|19]/adc_array_circuit_150n_0/vint1 col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5318 adc_array_wafflecap_8_8_0[11|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5319 VDD rowon_n[7] adc_array_wafflecap_8_8_0[6|13]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5320 adc_array_wafflecap_8_8_0[5|5]/adc_array_circuit_150n_0/vint2 rowon_n[6] adc_array_wafflecap_8_8_0[5|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5321 VDD rowon_n[3] adc_array_wafflecap_8_8_0[2|14]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5322 adc_array_wafflecap_8_8_1[27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_1[27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5323 VDD rowon_n[1] adc_array_wafflecap_8_8_0[0|29]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5324 adc_array_wafflecap_8_8_0[1|6]/adc_array_circuit_150n_0/vint2 rowon_n[2] adc_array_wafflecap_8_8_0[1|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5325 VSS row_n[1] adc_array_wafflecap_8_8_0[0|24]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5326 adc_array_wafflecap_8_8_0[0|17]/adc_array_circuit_150n_0/vdrv row_n[1] adc_array_wafflecap_8_8_0[0|17]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5327 adc_array_wafflecap_8_8_0[6|28]/adc_array_circuit_150n_0/vint2 col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5328 vcm adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|8]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5329 adc_array_wafflecap_8_8_0[4|10]/adc_array_circuit_150n_0/vint1 col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5330 VSS row_n[4] adc_array_wafflecap_8_8_0[3|2]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5331 vcm adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|9]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5332 adc_array_wafflecap_8_8_0[14|7]/adc_array_circuit_150n_0/vint2 rowon_n[15] adc_array_wafflecap_8_8_0[14|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5333 adc_array_wafflecap_8_8_0[14|29]/adc_array_circuit_150n_0/vint2 rowon_n[15] adc_array_wafflecap_8_8_0[14|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5334 adc_array_wafflecap_8_8_0[5|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5335 VSS row_n[7] adc_array_wafflecap_8_8_0[6|14]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5336 adc_array_wafflecap_8_8_0[13|11]/adc_array_circuit_150n_0/vint2 rowon_n[14] adc_array_wafflecap_8_8_0[13|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5337 VSS row_n[11] adc_array_wafflecap_8_8_0[10|30]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5338 adc_array_wafflecap_8_8_1[7]/adc_array_circuit_150n_0/vint1 col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5339 adc_array_wafflecap_8_8_0[13|1]/adc_array_circuit_150n_0/vint2 rowon_n[14] adc_array_wafflecap_8_8_0[13|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5340 adc_array_wafflecap_8_8_0[11|27]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|27]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5341 adc_array_wafflecap_8_8_0[6|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5342 adc_array_wafflecap_8_1_0/adc_array_circuit_150n_0/vint1 en_n_bit[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5343 VSS row_n[0] adc_array_wafflecap_8_8_1[12]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5344 VDD rowon_n[2] adc_array_wafflecap_8_8_0[1|6]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5345 adc_array_wafflecap_8_Dummy_4[17]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5346 adc_array_wafflecap_8_8_0[12|13]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|13]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5347 adc_array_wafflecap_8_8_0[2|29]/adc_array_circuit_150n_0/vdrv row_n[3] adc_array_wafflecap_8_8_0[2|29]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5348 adc_array_wafflecap_8_Dummy_4[7]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5349 adc_array_wafflecap_8_8_0[14|25]/adc_array_circuit_150n_0/vint1 col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5350 adc_array_wafflecap_8_8_0[12|3]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|3]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5351 VDD rowon_n[13] adc_array_wafflecap_8_8_0[12|7]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5352 VDD rowon_n[13] adc_array_wafflecap_8_8_0[12|29]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5353 adc_array_wafflecap_8_8_0[10|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5354 adc_array_wafflecap_8_8_0[6|28]/adc_array_circuit_150n_0/vdrv row_n[7] adc_array_wafflecap_8_8_0[6|28]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5355 vcm adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|0]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5356 vcm adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|1]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5357 adc_array_wafflecap_8_8_0[8|30]/adc_array_circuit_150n_0/vint1 col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5358 adc_array_wafflecap_8_8_0[6|14]/adc_array_circuit_150n_0/vint1 col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5359 vcm adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|13]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5360 adc_array_wafflecap_8_8_0[2|15]/adc_array_circuit_150n_0/vint1 col_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5361 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X5362 VSS row_n[10] adc_array_wafflecap_8_8_0[9|6]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5363 VDD rowon_n[0] adc_array_wafflecap_8_8_1[15]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5364 adc_array_wafflecap_8_Dummy_4[29]/adc_array_circuit_150n_0/vint2 col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5365 VSS row_n[15] adc_array_wafflecap_8_8_0[14|18]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5366 adc_array_wafflecap_8_8_0[11|6]/adc_array_circuit_150n_0/vint2 col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5367 adc_array_wafflecap_8_8_0[10|19]/adc_array_circuit_150n_0/vint2 col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5368 adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5369 adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5370 adc_array_wafflecap_8_8_0[7|6]/adc_array_circuit_150n_0/vint1 col_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5371 vcm VSS adc_array_wafflecap_8_Dummy_8[4]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5372 vcm adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|5]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5373 adc_array_wafflecap_8_8_0[13|28]/adc_array_circuit_150n_0/vdrv row_n[14] adc_array_wafflecap_8_8_0[13|28]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5374 adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5375 vcm adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|28]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5376 adc_array_wafflecap_8_8_1[30]/adc_array_circuit_150n_0/vdrv row_n[0] adc_array_wafflecap_8_8_1[30]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5377 adc_array_wafflecap_8_8_0[1|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5378 adc_array_wafflecap_8_8_0[14|14]/adc_array_circuit_150n_0/vdrv row_n[15] adc_array_wafflecap_8_8_0[14|14]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5379 adc_array_wafflecap_8_8_0[12|18]/adc_array_circuit_150n_0/vint1 col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5380 VDD rowon_n[5] adc_array_wafflecap_8_8_0[4|20]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5381 adc_array_wafflecap_8_8_0[14|4]/adc_array_circuit_150n_0/vdrv row_n[15] adc_array_wafflecap_8_8_0[14|4]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5382 adc_array_wafflecap_8_8_0[0|10]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|10]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5383 vcm adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|17]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5384 adc_array_wafflecap_8_8_0[13|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5385 adc_array_wafflecap_8_8_0[8|19]/adc_array_circuit_150n_0/vdrv row_n[9] adc_array_wafflecap_8_8_0[8|19]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5386 VDD rowon_n[0] adc_array_wafflecap_8_8_1[17]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5387 adc_array_wafflecap_8_8_1[15]/adc_array_circuit_150n_0/vint1 col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5388 adc_array_wafflecap_8_8_0[11|17]/adc_array_circuit_150n_0/vdrv row_n[12] adc_array_wafflecap_8_8_0[11|17]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5389 adc_array_wafflecap_8_8_0[9|28]/adc_array_circuit_150n_0/vint2 rowon_n[10] adc_array_wafflecap_8_8_0[9|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5390 VSS row_n[6] adc_array_wafflecap_8_8_0[5|27]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5391 adc_array_wafflecap_8_8_0[4|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5392 adc_array_wafflecap_8_8_1[22]/adc_array_circuit_150n_0/vint2 rowon_n[0] adc_array_wafflecap_8_8_1[22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5393 adc_array_wafflecap_8_8_0[0|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5394 VSS row_n[2] adc_array_wafflecap_8_8_0[1|28]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5395 adc_array_wafflecap_8_8_0[8|10]/adc_array_circuit_150n_0/vint2 rowon_n[9] adc_array_wafflecap_8_8_0[8|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5396 adc_array_wafflecap_8_8_0[7|25]/adc_array_circuit_150n_0/vint2 col_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5397 adc_array_wafflecap_8_Dummy_4[28]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5398 adc_array_wafflecap_8_8_0[8|0]/adc_array_circuit_150n_0/vint2 rowon_n[9] adc_array_wafflecap_8_8_0[8|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5399 VDD rowon_n[3] adc_array_wafflecap_8_8_0[2|25]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5400 adc_array_wafflecap_8_8_1[1]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[1]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5401 adc_array_wafflecap_8_8_0[13|24]/adc_array_circuit_150n_0/vint2 col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5402 vcm adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|7]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5403 VSS row_n[12] adc_array_wafflecap_8_8_0[11|28]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5404 adc_array_wafflecap_8_8_0[6|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5405 adc_array_wafflecap_8_Dummy_1[6]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_1[6]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5406 adc_array_wafflecap_8_8_0[4|6]/adc_array_circuit_150n_0/vint2 col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5407 adc_array_wafflecap_8_8_0[9|24]/adc_array_circuit_150n_0/vint1 col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5408 VDD rowon_n[8] adc_array_wafflecap_8_8_0[7|28]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5409 adc_array_wafflecap_8_Dummy_7/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_Dummy_7/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5410 adc_array_wafflecap_8_8_0[1|28]/adc_array_circuit_150n_0/vint1 col_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5411 adc_array_wafflecap_8_Dummy_4[24]/adc_array_circuit_150n_0/vint1 col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5412 VSS row_n[15] adc_array_wafflecap_8_8_0[14|26]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5413 adc_array_wafflecap_8_8_0[13|11]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|11]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5414 VDD rowon_n[14] adc_array_wafflecap_8_8_0[13|27]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5415 adc_array_wafflecap_8_8_0[9|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5416 adc_array_wafflecap_8_8_0[3|9]/adc_array_circuit_150n_0/vdrv row_n[4] adc_array_wafflecap_8_8_0[3|9]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5417 adc_array_wafflecap_8_8_0[3|22]/adc_array_circuit_150n_0/vint2 col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5418 VSS row_n[4] adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5419 adc_array_wafflecap_8_Dummy_1[4]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_1[4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5420 adc_array_wafflecap_8_8_0[2|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5421 adc_array_wafflecap_8_8_0[13|1]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|1]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5422 adc_array_wafflecap_8_8_0[10|27]/adc_array_circuit_150n_0/vint2 col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5423 adc_array_wafflecap_8_8_0[6|0]/adc_array_circuit_150n_0/vint2 col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5424 adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5425 adc_array_wafflecap_8_8_0[6|25]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|25]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5426 VSS row_n[10] adc_array_wafflecap_8_8_0[9|17]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X5427 adc_array_wafflecap_8_8_0[14|22]/adc_array_circuit_150n_0/vdrv row_n[15] adc_array_wafflecap_8_8_0[14|22]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5428 adc_array_wafflecap_8_8_0[12|26]/adc_array_circuit_150n_0/vint1 col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5429 adc_array_wafflecap_8_8_0[2|11]/adc_array_circuit_150n_0/vint2 col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5430 adc_array_wafflecap_8_8_1[23]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[23]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5431 adc_array_wafflecap_8_8_0[8|27]/adc_array_circuit_150n_0/vdrv row_n[9] adc_array_wafflecap_8_8_0[8|27]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5432 adc_array_wafflecap_8_8_0[6|0]/adc_array_circuit_150n_0/vdrv row_n[7] adc_array_wafflecap_8_8_0[6|0]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5433 adc_array_wafflecap_8_8_0[6|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5434 vcm adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|30]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5435 adc_array_wafflecap_8_8_0[2|1]/adc_array_circuit_150n_0/vdrv row_n[3] adc_array_wafflecap_8_8_0[2|1]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5436 vcm adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5437 vcm adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|21]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5438 adc_array_wafflecap_8_8_0[5|13]/adc_array_circuit_150n_0/vdrv row_n[6] adc_array_wafflecap_8_8_0[5|13]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5439 adc_array_wafflecap_8_8_0[4|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5440 vcm adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|25]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5441 adc_array_wafflecap_8_8_0[9|13]/adc_array_circuit_150n_0/vdrv row_n[10] adc_array_wafflecap_8_8_0[9|13]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5442 adc_array_wafflecap_8_8_0[8|26]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|26]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5443 adc_array_wafflecap_8_8_0[7|17]/adc_array_circuit_150n_0/vint1 col_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5444 adc_array_wafflecap_8_8_0[7|24]/adc_array_circuit_150n_0/vint2 rowon_n[8] adc_array_wafflecap_8_8_0[7|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5445 adc_array_wafflecap_8_8_0[5|14]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|14]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5446 adc_array_wafflecap_8_8_0[11|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5447 adc_array_wafflecap_8_8_0[9|3]/adc_array_circuit_150n_0/vdrv row_n[10] adc_array_wafflecap_8_8_0[9|3]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5448 adc_array_wafflecap_8_8_1[8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5449 adc_array_wafflecap_8_8_0[0|11]/adc_array_circuit_150n_0/vdrv row_n[1] adc_array_wafflecap_8_8_0[0|11]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5450 adc_array_wafflecap_8_8_0[12|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5451 adc_array_wafflecap_8_8_0[12|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5452 vcm adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|16]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5453 adc_array_wafflecap_8_8_0[4|15]/adc_array_circuit_150n_0/vint2 col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5454 VDD rowon_n[3] adc_array_wafflecap_8_8_0[2|7]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5455 vcm adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|6]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5456 adc_array_wafflecap_8_8_0[4|5]/adc_array_circuit_150n_0/vdrv row_n[5] adc_array_wafflecap_8_8_0[4|5]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5457 adc_array_wafflecap_8_8_0[0|27]/adc_array_circuit_150n_0/vint2 rowon_n[1] adc_array_wafflecap_8_8_0[0|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5458 adc_array_wafflecap_8_8_0[4|6]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|6]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5459 adc_array_wafflecap_8_8_0[4|26]/adc_array_circuit_150n_0/vint2 rowon_n[5] adc_array_wafflecap_8_8_0[4|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5460 adc_array_wafflecap_8_Dummy_4[26]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5461 VSS row_n[13] adc_array_wafflecap_8_8_0[12|22]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5462 adc_array_wafflecap_8_8_0[10|26]/adc_array_circuit_150n_0/vint2 rowon_n[11] adc_array_wafflecap_8_8_0[10|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5463 VSS row_n[7] adc_array_wafflecap_8_8_0[6|7]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5464 adc_array_wafflecap_8_8_0[14|6]/adc_array_circuit_150n_0/vint2 rowon_n[15] adc_array_wafflecap_8_8_0[14|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5465 adc_array_wafflecap_8_8_0[14|16]/adc_array_circuit_150n_0/vint2 rowon_n[15] adc_array_wafflecap_8_8_0[14|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5466 adc_array_wafflecap_8_8_0[9|17]/adc_array_circuit_150n_0/vint2 rowon_n[10] adc_array_wafflecap_8_8_0[9|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5467 adc_array_wafflecap_8_8_0[8|23]/adc_array_circuit_150n_0/vint2 col_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5468 adc_array_wafflecap_8_8_0[3|19]/adc_array_circuit_150n_0/vint1 col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5469 adc_array_wafflecap_8_8_0[3|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5470 adc_array_wafflecap_8_8_1[2]/adc_array_circuit_150n_0/vdrv row_n[0] adc_array_wafflecap_8_8_1[2]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5471 adc_array_wafflecap_8_Dummy_4[18]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5472 adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5473 adc_array_wafflecap_8_8_0[3|17]/adc_array_circuit_150n_0/vdrv row_n[4] adc_array_wafflecap_8_8_0[3|17]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5474 VDD rowon_n[4] adc_array_wafflecap_8_8_0[3|29]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5475 adc_array_wafflecap_8_8_0[3|18]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|18]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5476 VDD rowon_n[15] adc_array_wafflecap_8_8_0[14|21]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5477 adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5478 adc_array_wafflecap_8_8_0[12|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5479 vcm adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|18]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5480 VSS row_n[8] adc_array_wafflecap_8_8_0[7|3]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5481 VSS row_n[8] adc_array_wafflecap_8_8_0[7|13]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5482 VDD rowon_n[5] adc_array_wafflecap_8_8_0[4|11]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5483 VDD VSS adc_array_wafflecap_8_Dummy_3[2]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5484 VDD rowon_n[14] adc_array_wafflecap_8_8_0[13|25]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5485 adc_array_wafflecap_8_8_0[10|22]/adc_array_circuit_150n_0/vint1 col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5486 adc_array_wafflecap_8_8_0[3|3]/adc_array_circuit_150n_0/vint2 rowon_n[4] adc_array_wafflecap_8_8_0[3|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5487 VDD rowon_n[13] adc_array_wafflecap_8_8_0[12|16]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5488 VDD rowon_n[9] adc_array_wafflecap_8_8_0[8|26]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5489 adc_array_wafflecap_8_8_0[6|15]/adc_array_circuit_150n_0/vint2 rowon_n[7] adc_array_wafflecap_8_8_0[6|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5490 adc_array_wafflecap_8_8_0[2|8]/adc_array_circuit_150n_0/vint1 col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5491 adc_array_wafflecap_8_Dummy_6/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_6/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5492 VSS VSS adc_array_wafflecap_8_Dummy_2[5]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5493 VSS row_n[3] adc_array_wafflecap_8_8_0[2|21]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5494 VDD rowon_n[13] adc_array_wafflecap_8_8_0[12|6]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5495 VDD rowon_n[8] adc_array_wafflecap_8_8_0[7|17]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5496 adc_array_wafflecap_8_8_0[6|7]/adc_array_circuit_150n_0/vint1 col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5497 VDD rowon_n[0] adc_array_wafflecap_8_8_1[8]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5498 VSS row_n[2] adc_array_wafflecap_8_8_0[1|0]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5499 adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/vint2 rowon_n[3] adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5500 adc_array_wafflecap_8_8_1[13]/adc_array_circuit_150n_0/vint2 rowon_n[0] adc_array_wafflecap_8_8_1[13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5501 adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5502 adc_array_wafflecap_8_8_0[1|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5503 adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5504 adc_array_wafflecap_8_8_0[5|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5505 VSS VDD adc_array_wafflecap_8_Dummy_4[15]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5506 adc_array_wafflecap_8_8_0[12|11]/adc_array_circuit_150n_0/vint2 col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5507 VSS VDD adc_array_wafflecap_8_Dummy_4[5]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5508 adc_array_wafflecap_8_8_0[12|1]/adc_array_circuit_150n_0/vint2 col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5509 adc_array_wafflecap_8_8_0[7|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5510 VDD rowon_n[3] adc_array_wafflecap_8_8_0[2|16]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5511 vcm adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[19]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5512 VDD rowon_n[1] adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5513 adc_array_wafflecap_8_8_0[0|21]/adc_array_circuit_150n_0/vint1 col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5514 adc_array_wafflecap_8_Dummy_4[21]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[21]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5515 adc_array_wafflecap_8_8_0[11|5]/adc_array_circuit_150n_0/vint2 col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5516 adc_array_wafflecap_8_8_0[11|15]/adc_array_circuit_150n_0/vint2 col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5517 vcm adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|20]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5518 VDD rowon_n[7] adc_array_wafflecap_8_8_0[6|15]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5519 adc_array_wafflecap_8_8_0[4|26]/adc_array_circuit_150n_0/vdrv row_n[5] adc_array_wafflecap_8_8_0[4|26]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5520 adc_array_wafflecap_8_8_1[29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_1[29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5521 vcm VSS adc_array_wafflecap_8_Dummy_0[0]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5522 adc_array_wafflecap_8_8_0[1|0]/adc_array_circuit_150n_0/vint1 col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5523 vcm adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|10]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5524 vcm adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|11]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5525 adc_array_wafflecap_8_8_0[14|10]/adc_array_circuit_150n_0/vint1 col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5526 adc_array_wafflecap_8_8_0[6|30]/adc_array_circuit_150n_0/vint2 col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5527 adc_array_wafflecap_8_8_0[4|12]/adc_array_circuit_150n_0/vint1 col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5528 adc_array_wafflecap_8_8_0[4|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5529 VSS row_n[4] adc_array_wafflecap_8_8_0[3|4]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5530 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.64e+07u l=1.6e+07u
X5531 adc_array_wafflecap_8_8_0[14|0]/adc_array_circuit_150n_0/vint1 col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5532 adc_array_wafflecap_8_8_0[13|4]/adc_array_circuit_150n_0/vint1 col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5533 adc_array_wafflecap_8_8_0[13|14]/adc_array_circuit_150n_0/vint1 col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5534 adc_array_wafflecap_8_8_0[10|1]/adc_array_circuit_150n_0/vdrv row_n[11] adc_array_wafflecap_8_8_0[10|1]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5535 adc_array_wafflecap_8_8_0[10|11]/adc_array_circuit_150n_0/vdrv row_n[11] adc_array_wafflecap_8_8_0[10|11]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5536 adc_array_wafflecap_8_8_0[9|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5537 adc_array_wafflecap_8_8_0[8|22]/adc_array_circuit_150n_0/vint2 rowon_n[9] adc_array_wafflecap_8_8_0[8|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5538 adc_array_wafflecap_8_8_0[7|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5539 adc_array_wafflecap_8_8_0[7|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5540 adc_array_wafflecap_8_8_1[9]/adc_array_circuit_150n_0/vint1 col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5541 adc_array_wafflecap_8_8_1[28]/adc_array_circuit_150n_0/vint2 col_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5542 adc_array_wafflecap_8_8_0[13|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5543 VSS row_n[0] adc_array_wafflecap_8_8_1[14]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5544 adc_array_wafflecap_8_8_0[13|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5545 adc_array_wafflecap_8_8_0[5|19]/adc_array_circuit_150n_0/vint2 col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5546 adc_array_wafflecap_8_8_0[6|30]/adc_array_circuit_150n_0/vdrv row_n[7] adc_array_wafflecap_8_8_0[6|30]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5547 vcm adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|2]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5548 vcm adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|3]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5549 adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/vdrv row_n[3] adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5550 VSS row_n[8] adc_array_wafflecap_8_8_0[7|21]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5551 vcm adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|15]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5552 adc_array_wafflecap_8_8_0[9|15]/adc_array_circuit_150n_0/vint2 rowon_n[10] adc_array_wafflecap_8_8_0[9|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5553 VSS row_n[14] adc_array_wafflecap_8_8_0[13|20]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5554 vcm adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|12]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5555 adc_array_wafflecap_8_8_0[9|5]/adc_array_circuit_150n_0/vint2 rowon_n[10] adc_array_wafflecap_8_8_0[9|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5556 adc_array_wafflecap_8_8_0[7|3]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|3]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5557 adc_array_wafflecap_8_8_0[7|13]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|13]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5558 VDD rowon_n[3] adc_array_wafflecap_8_8_0[2|18]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5559 adc_array_wafflecap_8_Dummy_4[15]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5560 vcm adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|2]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5561 adc_array_wafflecap_8_4_0/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_4_0/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5562 adc_array_wafflecap_8_Dummy_4[5]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5563 VDD rowon_n[10] adc_array_wafflecap_8_8_0[9|20]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5564 adc_array_wafflecap_8_8_0[2|7]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|7]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5565 adc_array_wafflecap_8_8_0[2|16]/adc_array_circuit_150n_0/vint1 col_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5566 adc_array_wafflecap_8_8_0[2|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5567 adc_array_wafflecap_8_Dummy_2[1]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5568 adc_array_wafflecap_8_8_0[13|30]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|30]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5569 VDD VDD adc_array_wafflecap_8_Dummy_4[20]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5570 adc_array_wafflecap_8_8_0[13|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5571 adc_array_wafflecap_8_8_0[14|6]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|6]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5572 adc_array_wafflecap_8_8_0[14|16]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|16]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5573 VDD rowon_n[15] adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5574 VDD rowon_n[8] adc_array_wafflecap_8_8_0[7|5]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5575 VDD rowon_n[8] adc_array_wafflecap_8_8_0[7|15]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5576 VDD rowon_n[14] adc_array_wafflecap_8_8_0[13|14]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5577 VDD rowon_n[14] adc_array_wafflecap_8_8_0[13|4]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5578 adc_array_wafflecap_8_8_0[1|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5579 adc_array_wafflecap_8_8_0[7|10]/adc_array_circuit_150n_0/vint2 col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5580 adc_array_wafflecap_8_8_0[6|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5581 adc_array_wafflecap_8_8_0[4|17]/adc_array_circuit_150n_0/vint2 rowon_n[5] adc_array_wafflecap_8_8_0[4|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5582 vcm adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|24]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5583 adc_array_wafflecap_8_8_0[0|12]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|12]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5584 adc_array_wafflecap_8_8_0[7|0]/adc_array_circuit_150n_0/vint2 col_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5585 VDD sample adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5586 VDD rowon_n[0] adc_array_wafflecap_8_8_1[19]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5587 adc_array_wafflecap_8_8_0[13|9]/adc_array_circuit_150n_0/vint2 col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5588 adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/vdrv row_n[10] adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5589 adc_array_wafflecap_8_8_0[13|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5590 adc_array_wafflecap_8_8_0[9|9]/adc_array_circuit_150n_0/vint1 col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5591 adc_array_wafflecap_8_8_0[8|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5592 adc_array_wafflecap_8_8_1[24]/adc_array_circuit_150n_0/vint2 rowon_n[0] adc_array_wafflecap_8_8_1[24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5593 adc_array_wafflecap_8_8_0[0|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5594 adc_array_wafflecap_8_8_0[1|20]/adc_array_circuit_150n_0/vint2 col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5595 adc_array_wafflecap_8_Dummy_4[32]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[32]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5596 vcm adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5597 adc_array_wafflecap_8_8_0[5|6]/adc_array_circuit_150n_0/vdrv row_n[6] adc_array_wafflecap_8_8_0[5|6]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5598 VSS row_n[6] adc_array_wafflecap_8_8_0[5|29]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5599 adc_array_wafflecap_8_8_0[4|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5600 VSS row_n[2] adc_array_wafflecap_8_8_0[1|30]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5601 adc_array_wafflecap_8_8_0[9|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5602 adc_array_wafflecap_8_Dummy_4[9]/adc_array_circuit_150n_0/vint1 col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5603 adc_array_wafflecap_8_8_0[9|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5604 adc_array_wafflecap_8_8_0[8|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5605 adc_array_wafflecap_8_Dummy_4[26]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5606 adc_array_wafflecap_8_8_0[8|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5607 adc_array_wafflecap_8_8_0[4|8]/adc_array_circuit_150n_0/vint2 col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5608 adc_array_wafflecap_8_8_0[0|9]/adc_array_circuit_150n_0/vint2 col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5609 adc_array_wafflecap_8_8_0[11|26]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|26]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5610 VSS row_n[5] adc_array_wafflecap_8_8_0[4|18]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5611 vcm VSS adc_array_wafflecap_8_Dummy_3[4]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5612 adc_array_wafflecap_8_8_1[1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_1[1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5613 adc_array_wafflecap_8_8_0[1|30]/adc_array_circuit_150n_0/vint1 col_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5614 adc_array_wafflecap_8_8_0[1|20]/adc_array_circuit_150n_0/vdrv row_n[2] adc_array_wafflecap_8_8_0[1|20]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5615 vcm adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|28]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5616 adc_array_wafflecap_8_8_0[14|7]/adc_array_circuit_150n_0/vdrv row_n[15] adc_array_wafflecap_8_8_0[14|7]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5617 adc_array_wafflecap_8_8_0[12|18]/adc_array_circuit_150n_0/vint2 rowon_n[13] adc_array_wafflecap_8_8_0[12|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5618 VDD sample_n adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5619 adc_array_wafflecap_8_Dummy_1[6]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_1[6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5620 adc_array_wafflecap_8_8_0[6|2]/adc_array_circuit_150n_0/vint2 col_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5621 adc_array_wafflecap_8_8_0[3|11]/adc_array_circuit_150n_0/vdrv row_n[4] adc_array_wafflecap_8_8_0[3|11]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5622 adc_array_wafflecap_8_8_0[2|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5623 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.64e+07u l=1.6e+07u
X5624 VSS row_n[9] adc_array_wafflecap_8_8_0[8|19]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5625 VSS row_n[8] adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5626 adc_array_wafflecap_8_8_0[10|3]/adc_array_circuit_150n_0/vint2 rowon_n[11] adc_array_wafflecap_8_8_0[10|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5627 adc_array_wafflecap_8_8_0[10|13]/adc_array_circuit_150n_0/vint2 rowon_n[11] adc_array_wafflecap_8_8_0[10|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5628 adc_array_wafflecap_8_8_0[8|11]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|11]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5629 adc_array_wafflecap_8_Dummy_1[0]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_1[0]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5630 vcm adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|0]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5631 vcm adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|10]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5632 adc_array_wafflecap_8_8_0[8|1]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|1]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5633 adc_array_wafflecap_8_Dummy_1[5]/adc_array_circuit_150n_0/vint2 col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5634 adc_array_wafflecap_8_8_1[0]/adc_array_circuit_150n_0/vint2 col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5635 VDD rowon_n[11] adc_array_wafflecap_8_8_0[10|18]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5636 adc_array_wafflecap_8_8_0[9|5]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|5]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5637 adc_array_wafflecap_8_8_0[9|15]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|15]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5638 VDD rowon_n[10] adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5639 adc_array_wafflecap_8_8_0[2|13]/adc_array_circuit_150n_0/vint2 col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5640 VDD rowon_n[10] adc_array_wafflecap_8_8_0[9|9]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5641 adc_array_wafflecap_8_8_0[6|8]/adc_array_circuit_150n_0/vint2 rowon_n[7] adc_array_wafflecap_8_8_0[6|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5642 vcm adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5643 adc_array_wafflecap_8_8_1[25]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[25]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5644 adc_array_wafflecap_8_Dummy_4[15]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[15]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5645 adc_array_wafflecap_8_8_0[13|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5646 VDD rowon_n[9] adc_array_wafflecap_8_8_0[8|13]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5647 adc_array_wafflecap_8_8_0[6|2]/adc_array_circuit_150n_0/vdrv row_n[7] adc_array_wafflecap_8_8_0[6|2]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5648 adc_array_wafflecap_8_8_0[6|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5649 adc_array_wafflecap_8_8_0[2|3]/adc_array_circuit_150n_0/vdrv row_n[3] adc_array_wafflecap_8_8_0[2|3]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5650 adc_array_wafflecap_8_8_0[2|4]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|4]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5651 adc_array_wafflecap_8_Dummy_4[5]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[5]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5652 VDD rowon_n[9] adc_array_wafflecap_8_8_0[8|3]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5653 adc_array_wafflecap_8_8_0[5|15]/adc_array_circuit_150n_0/vdrv row_n[6] adc_array_wafflecap_8_8_0[5|15]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5654 adc_array_wafflecap_8_8_0[5|16]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|16]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5655 adc_array_wafflecap_8_8_0[12|30]/adc_array_circuit_150n_0/vint2 col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5656 VSS row_n[13] adc_array_wafflecap_8_8_0[12|7]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5657 VDD rowon_n[6] adc_array_wafflecap_8_8_0[5|26]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5658 adc_array_wafflecap_8_8_1[6]/adc_array_circuit_150n_0/vint2 rowon_n[0] adc_array_wafflecap_8_8_1[6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5659 adc_array_wafflecap_8_8_0[0|13]/adc_array_circuit_150n_0/vdrv row_n[1] adc_array_wafflecap_8_8_0[0|13]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5660 adc_array_wafflecap_8_8_1[10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5661 adc_array_wafflecap_8_8_0[12|17]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|17]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5662 VSS row_n[12] adc_array_wafflecap_8_8_0[11|1]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5663 VSS row_n[12] adc_array_wafflecap_8_8_0[11|11]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5664 adc_array_wafflecap_8_8_0[8|8]/adc_array_circuit_150n_0/vint2 col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5665 adc_array_wafflecap_8_8_0[6|24]/adc_array_circuit_150n_0/vint2 col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5666 adc_array_wafflecap_8_8_0[14|29]/adc_array_circuit_150n_0/vint1 col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5667 adc_array_wafflecap_8_8_0[11|26]/adc_array_circuit_150n_0/vdrv row_n[12] adc_array_wafflecap_8_8_0[11|26]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5668 VDD rowon_n[7] adc_array_wafflecap_8_8_0[6|8]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5669 adc_array_wafflecap_8_8_0[5|0]/adc_array_circuit_150n_0/vint2 rowon_n[6] adc_array_wafflecap_8_8_0[5|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5670 VDD rowon_n[3] adc_array_wafflecap_8_8_0[2|9]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5671 adc_array_wafflecap_8_8_0[1|1]/adc_array_circuit_150n_0/vint2 rowon_n[2] adc_array_wafflecap_8_8_0[1|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5672 adc_array_wafflecap_8_8_0[10|30]/adc_array_circuit_150n_0/vdrv row_n[11] adc_array_wafflecap_8_8_0[10|30]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5673 VSS row_n[1] adc_array_wafflecap_8_8_0[0|19]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5674 adc_array_wafflecap_8_8_0[14|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5675 adc_array_wafflecap_8_8_0[4|28]/adc_array_circuit_150n_0/vint2 rowon_n[5] adc_array_wafflecap_8_8_0[4|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5676 adc_array_wafflecap_8_8_0[0|29]/adc_array_circuit_150n_0/vint2 rowon_n[1] adc_array_wafflecap_8_8_0[0|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5677 adc_array_wafflecap_8_8_0[10|7]/adc_array_circuit_150n_0/vint1 col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5678 adc_array_wafflecap_8_8_0[0|17]/adc_array_circuit_150n_0/vint2 col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5679 adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5680 vcm adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|29]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5681 VSS row_n[7] adc_array_wafflecap_8_8_0[6|9]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5682 adc_array_wafflecap_8_8_0[3|21]/adc_array_circuit_150n_0/vint1 col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5683 adc_array_wafflecap_8_8_1[4]/adc_array_circuit_150n_0/vdrv row_n[0] adc_array_wafflecap_8_8_1[4]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5684 adc_array_wafflecap_8_8_0[10|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5685 adc_array_wafflecap_8_8_0[3|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5686 VDD rowon_n[4] adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5687 adc_array_wafflecap_8_8_0[6|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5688 adc_array_wafflecap_8_8_0[6|24]/adc_array_circuit_150n_0/vdrv row_n[7] adc_array_wafflecap_8_8_0[6|24]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5689 adc_array_wafflecap_8_Dummy_2[2]/adc_array_circuit_150n_0/vint1 col_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5690 VSS row_n[0] adc_array_wafflecap_8_8_1[7]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5691 VDD rowon_n[2] adc_array_wafflecap_8_8_0[1|1]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5692 adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5693 VDD rowon_n[5] adc_array_wafflecap_8_8_0[4|13]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5694 adc_array_wafflecap_8_8_0[3|5]/adc_array_circuit_150n_0/vint2 rowon_n[4] adc_array_wafflecap_8_8_0[3|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5695 VDD VSS adc_array_wafflecap_8_Dummy_3[4]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5696 adc_array_wafflecap_8_Dummy_2[0]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_2[0]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5697 VSS en_n_bit[0] adc_array_wafflecap_8_1_0/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5698 adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5699 adc_array_wafflecap_8_8_0[7|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5700 adc_array_wafflecap_8_8_0[6|9]/adc_array_circuit_150n_0/vint1 col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5701 vcm adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|8]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5702 adc_array_wafflecap_8_8_0[2|10]/adc_array_circuit_150n_0/vint1 col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5703 VDD rowon_n[0] adc_array_wafflecap_8_8_1[10]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5704 VSS row_n[2] adc_array_wafflecap_8_8_0[1|2]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5705 adc_array_wafflecap_8_8_0[14|18]/adc_array_circuit_150n_0/vdrv row_n[15] adc_array_wafflecap_8_8_0[14|18]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5706 VSS row_n[15] adc_array_wafflecap_8_8_0[14|25]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5707 adc_array_wafflecap_8_8_0[12|7]/adc_array_circuit_150n_0/vint2 rowon_n[13] adc_array_wafflecap_8_8_0[12|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5708 adc_array_wafflecap_8_8_0[12|29]/adc_array_circuit_150n_0/vint2 rowon_n[13] adc_array_wafflecap_8_8_0[12|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5709 VSS row_n[6] adc_array_wafflecap_8_8_0[5|1]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5710 adc_array_wafflecap_8_8_0[3|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5711 adc_array_wafflecap_8_Dummy_4[23]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[23]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5712 adc_array_wafflecap_8_8_0[11|11]/adc_array_circuit_150n_0/vint2 rowon_n[12] adc_array_wafflecap_8_8_0[11|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5713 VSS row_n[9] adc_array_wafflecap_8_8_0[8|30]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5714 adc_array_wafflecap_8_8_0[5|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5715 adc_array_wafflecap_8_8_1[15]/adc_array_circuit_150n_0/vint2 rowon_n[0] adc_array_wafflecap_8_8_1[15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5716 adc_array_wafflecap_8_8_0[11|1]/adc_array_circuit_150n_0/vint2 rowon_n[12] adc_array_wafflecap_8_8_0[11|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5717 adc_array_wafflecap_8_8_0[14|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5718 adc_array_wafflecap_8_8_0[14|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5719 adc_array_wafflecap_8_8_0[13|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5720 adc_array_wafflecap_8_8_0[12|25]/adc_array_circuit_150n_0/vint1 col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5721 adc_array_wafflecap_8_8_0[10|13]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|13]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5722 adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5723 vcm adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[21]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5724 adc_array_wafflecap_8_8_0[13|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5725 adc_array_wafflecap_8_8_0[10|3]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|3]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5726 VDD rowon_n[11] adc_array_wafflecap_8_8_0[10|7]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5727 VDD rowon_n[11] adc_array_wafflecap_8_8_0[10|29]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5728 adc_array_wafflecap_8_8_0[4|28]/adc_array_circuit_150n_0/vdrv row_n[5] adc_array_wafflecap_8_8_0[4|28]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5729 adc_array_wafflecap_8_8_0[4|29]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|29]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5730 vcm VSS adc_array_wafflecap_8_1_1/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5731 adc_array_wafflecap_8_8_0[1|2]/adc_array_circuit_150n_0/vint1 col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5732 vcm adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|0]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5733 adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/vint2 VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5734 vcm adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|12]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5735 adc_array_wafflecap_8_8_0[4|14]/adc_array_circuit_150n_0/vint1 col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5736 vcm adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|13]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5737 VSS row_n[8] adc_array_wafflecap_8_8_0[7|6]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5738 VSS sample adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5739 adc_array_wafflecap_8_8_0[4|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5740 adc_array_wafflecap_8_8_1[25]/adc_array_circuit_150n_0/vdrv row_n[0] adc_array_wafflecap_8_8_1[25]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5741 adc_array_wafflecap_8_8_0[13|28]/adc_array_circuit_150n_0/vint2 col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5742 adc_array_wafflecap_8_8_1[11]/adc_array_circuit_150n_0/vint1 col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5743 adc_array_wafflecap_8_8_0[14|14]/adc_array_circuit_150n_0/vint2 col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5744 VSS row_n[13] adc_array_wafflecap_8_8_0[12|18]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5745 VSS row_n[6] adc_array_wafflecap_8_8_0[5|23]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5746 adc_array_wafflecap_8_8_1[30]/adc_array_circuit_150n_0/vint2 col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5747 adc_array_wafflecap_8_8_0[14|4]/adc_array_circuit_150n_0/vint2 col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5748 adc_array_wafflecap_8_Dummy_4[28]/adc_array_circuit_150n_0/vint1 col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5749 adc_array_wafflecap_8_8_0[14|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5750 adc_array_wafflecap_8_8_0[9|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5751 adc_array_wafflecap_8_8_0[8|19]/adc_array_circuit_150n_0/vint2 col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5752 adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5753 adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/vdrv row_n[7] adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5754 adc_array_wafflecap_8_8_1[17]/adc_array_circuit_150n_0/vint2 rowon_n[0] adc_array_wafflecap_8_8_1[17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5755 vcm adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|5]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5756 adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5757 VSS row_n[0] adc_array_wafflecap_8_8_1[15]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5758 adc_array_wafflecap_8_8_0[12|4]/adc_array_circuit_150n_0/vdrv row_n[13] adc_array_wafflecap_8_8_0[12|4]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5759 adc_array_wafflecap_8_8_0[12|14]/adc_array_circuit_150n_0/vdrv row_n[13] adc_array_wafflecap_8_8_0[12|14]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5760 adc_array_wafflecap_8_8_0[10|18]/adc_array_circuit_150n_0/vint1 col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5761 VDD rowon_n[3] adc_array_wafflecap_8_8_0[2|20]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5762 adc_array_wafflecap_8_Dummy_1[1]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_1[1]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5763 adc_array_wafflecap_8_8_0[11|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5764 VDD rowon_n[6] adc_array_wafflecap_8_8_0[5|17]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5765 adc_array_wafflecap_8_8_0[9|17]/adc_array_circuit_150n_0/vdrv row_n[10] adc_array_wafflecap_8_8_0[9|17]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5766 VSS row_n[10] adc_array_wafflecap_8_8_0[9|24]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5767 adc_array_wafflecap_8_8_0[8|30]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|30]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5768 adc_array_wafflecap_8_8_0[7|28]/adc_array_circuit_150n_0/vint2 rowon_n[8] adc_array_wafflecap_8_8_0[7|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5769 VSS row_n[4] adc_array_wafflecap_8_8_0[3|27]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5770 adc_array_wafflecap_8_4_0/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_4_0/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5771 adc_array_wafflecap_8_8_0[2|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5772 adc_array_wafflecap_8_8_0[8|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5773 VSS VDD adc_array_wafflecap_8_Dummy_4[24]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5774 vcm adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|15]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5775 adc_array_wafflecap_8_Dummy_4[17]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[17]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5776 vcm adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|5]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5777 adc_array_wafflecap_8_8_0[13|27]/adc_array_circuit_150n_0/vint2 rowon_n[14] adc_array_wafflecap_8_8_0[13|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5778 adc_array_wafflecap_8_8_0[6|20]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|20]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5779 VDD rowon_n[12] adc_array_wafflecap_8_8_0[11|23]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5780 adc_array_wafflecap_8_8_0[11|24]/adc_array_circuit_150n_0/vint2 col_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5781 adc_array_wafflecap_8_8_0[9|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5782 adc_array_wafflecap_8_8_0[6|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5783 vcm adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|26]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5784 adc_array_wafflecap_8_8_0[9|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5785 adc_array_wafflecap_8_8_0[2|6]/adc_array_circuit_150n_0/vint2 col_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5786 adc_array_wafflecap_8_Dummy_4[11]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5787 adc_array_wafflecap_8_8_0[7|24]/adc_array_circuit_150n_0/vint1 col_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5788 adc_array_wafflecap_8_Dummy_4[1]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5789 adc_array_wafflecap_8_8_0[14|22]/adc_array_circuit_150n_0/vint2 col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5790 adc_array_wafflecap_8_8_0[13|23]/adc_array_circuit_150n_0/vint1 col_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5791 VSS row_n[13] adc_array_wafflecap_8_8_0[12|26]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5792 adc_array_wafflecap_8_8_0[11|11]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|11]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5793 adc_array_wafflecap_8_8_0[7|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5794 adc_array_wafflecap_8_8_0[5|8]/adc_array_circuit_150n_0/vdrv row_n[6] adc_array_wafflecap_8_8_0[5|8]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5795 adc_array_wafflecap_8_8_0[4|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5796 adc_array_wafflecap_8_8_0[0|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5797 VSS row_n[2] adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5798 adc_array_wafflecap_8_8_0[1|22]/adc_array_circuit_150n_0/vint2 col_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5799 adc_array_wafflecap_8_8_0[11|1]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|1]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5800 adc_array_wafflecap_8_8_0[8|27]/adc_array_circuit_150n_0/vint2 col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5801 adc_array_wafflecap_8_8_0[5|9]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|9]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5802 adc_array_wafflecap_8_8_0[5|18]/adc_array_circuit_150n_0/vint1 col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5803 VSS row_n[6] adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5804 adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5805 adc_array_wafflecap_8_8_0[9|13]/adc_array_circuit_150n_0/vint2 col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5806 adc_array_wafflecap_8_8_0[0|6]/adc_array_circuit_150n_0/vdrv row_n[1] adc_array_wafflecap_8_8_0[0|6]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5807 adc_array_wafflecap_8_8_0[9|3]/adc_array_circuit_150n_0/vint2 col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5808 VSS row_n[8] adc_array_wafflecap_8_8_0[7|17]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5809 adc_array_wafflecap_8_8_0[4|22]/adc_array_circuit_150n_0/vint2 rowon_n[5] adc_array_wafflecap_8_8_0[4|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5810 adc_array_wafflecap_8_8_0[12|22]/adc_array_circuit_150n_0/vdrv row_n[13] adc_array_wafflecap_8_8_0[12|22]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5811 adc_array_wafflecap_8_8_0[10|26]/adc_array_circuit_150n_0/vint1 col_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5812 adc_array_wafflecap_8_8_0[4|10]/adc_array_circuit_150n_0/vint2 col_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5813 adc_array_wafflecap_8_8_0[0|11]/adc_array_circuit_150n_0/vint2 col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5814 adc_array_wafflecap_8_8_0[1|22]/adc_array_circuit_150n_0/vdrv row_n[2] adc_array_wafflecap_8_8_0[1|22]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5815 adc_array_wafflecap_8_8_0[11|12]/adc_array_circuit_150n_0/vint1 col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5816 adc_array_wafflecap_8_8_0[4|0]/adc_array_circuit_150n_0/vdrv row_n[5] adc_array_wafflecap_8_8_0[4|0]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5817 adc_array_wafflecap_8_8_1[3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_1[3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5818 adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/vint1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5819 vcm adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|30]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5820 adc_array_wafflecap_8_Dummy_4[25]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5821 vcm adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|21]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5822 adc_array_wafflecap_8_8_0[11|2]/adc_array_circuit_150n_0/vint1 col_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5823 adc_array_wafflecap_8_8_0[4|1]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|1]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5824 adc_array_wafflecap_8_8_0[3|13]/adc_array_circuit_150n_0/vdrv row_n[4] adc_array_wafflecap_8_8_0[3|13]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5825 adc_array_wafflecap_8_8_0[2|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5826 vcm adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|25]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5827 adc_array_wafflecap_8_8_0[7|13]/adc_array_circuit_150n_0/vdrv row_n[8] adc_array_wafflecap_8_8_0[7|13]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5828 adc_array_wafflecap_8_8_0[3|14]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|14]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5829 adc_array_wafflecap_8_8_0[7|3]/adc_array_circuit_150n_0/vdrv row_n[8] adc_array_wafflecap_8_8_0[7|3]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5830 adc_array_wafflecap_8_Dummy_1[2]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_1[2]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5831 adc_array_wafflecap_8_8_0[10|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5832 adc_array_wafflecap_8_8_0[10|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5833 adc_array_wafflecap_8_8_1[2]/adc_array_circuit_150n_0/vint2 col_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5834 adc_array_wafflecap_8_8_0[2|15]/adc_array_circuit_150n_0/vint2 col_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5835 adc_array_wafflecap_8_8_0[14|21]/adc_array_circuit_150n_0/vint2 rowon_n[15] adc_array_wafflecap_8_8_0[14|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5836 adc_array_wafflecap_8_8_0[6|10]/adc_array_circuit_150n_0/vint2 rowon_n[7] adc_array_wafflecap_8_8_0[6|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5837 adc_array_wafflecap_8_8_0[2|5]/adc_array_circuit_150n_0/vdrv row_n[3] adc_array_wafflecap_8_8_0[2|5]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5838 adc_array_wafflecap_8_Dummy_3[2]/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_3[2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5839 adc_array_wafflecap_8_8_0[2|6]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|6]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5840 analog_in sw ctop VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=500000u
X5841 adc_array_wafflecap_8_8_0[2|26]/adc_array_circuit_150n_0/vint2 rowon_n[3] adc_array_wafflecap_8_8_0[2|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5842 adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5843 adc_array_wafflecap_8_8_0[13|25]/adc_array_circuit_150n_0/vint2 rowon_n[14] adc_array_wafflecap_8_8_0[13|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5844 VSS row_n[11] adc_array_wafflecap_8_8_0[10|22]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5845 adc_array_wafflecap_8_8_0[8|26]/adc_array_circuit_150n_0/vint2 rowon_n[9] adc_array_wafflecap_8_8_0[8|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5846 adc_array_wafflecap_8_8_0[12|6]/adc_array_circuit_150n_0/vint2 rowon_n[13] adc_array_wafflecap_8_8_0[12|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5847 adc_array_wafflecap_8_8_0[12|16]/adc_array_circuit_150n_0/vint2 rowon_n[13] adc_array_wafflecap_8_8_0[12|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5848 adc_array_wafflecap_8_8_0[7|17]/adc_array_circuit_150n_0/vint2 rowon_n[8] adc_array_wafflecap_8_8_0[7|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5849 adc_array_wafflecap_8_8_1[8]/adc_array_circuit_150n_0/vint2 rowon_n[0] adc_array_wafflecap_8_8_1[8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5850 adc_array_wafflecap_8_8_1[26]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[26]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5851 adc_array_wafflecap_8_8_0[1|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5852 vcm VSS adc_array_wafflecap_8_Dummy_4[14]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5853 adc_array_wafflecap_8_8_0[13|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5854 adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5855 adc_array_wafflecap_8_8_0[8|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5856 adc_array_wafflecap_8_8_0[5|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5857 VDD rowon_n[6] adc_array_wafflecap_8_8_0[5|28]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5858 adc_array_wafflecap_8_8_0[0|15]/adc_array_circuit_150n_0/vdrv row_n[1] adc_array_wafflecap_8_8_0[0|15]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5859 vcm VSS adc_array_wafflecap_8_Dummy_4[4]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5860 adc_array_wafflecap_8_8_0[5|17]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|17]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5861 adc_array_wafflecap_8_8_0[1|18]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|18]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5862 VDD rowon_n[13] adc_array_wafflecap_8_8_0[12|21]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5863 adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5864 adc_array_wafflecap_8_8_0[10|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5865 VDD rowon_n[3] adc_array_wafflecap_8_8_0[2|11]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5866 VDD rowon_n[1] adc_array_wafflecap_8_8_0[0|26]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5867 VDD rowon_n[12] adc_array_wafflecap_8_8_0[11|2]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5868 VDD rowon_n[12] adc_array_wafflecap_8_8_0[11|12]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5869 adc_array_wafflecap_8_8_0[8|22]/adc_array_circuit_150n_0/vint1 col_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5870 VDD rowon_n[7] adc_array_wafflecap_8_8_0[6|10]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5871 adc_array_wafflecap_8_8_0[1|3]/adc_array_circuit_150n_0/vint2 rowon_n[2] adc_array_wafflecap_8_8_0[1|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5872 VDD rowon_n[11] adc_array_wafflecap_8_8_0[10|16]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5873 VSS row_n[1] adc_array_wafflecap_8_8_0[0|21]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5874 adc_array_wafflecap_8_Dummy_4[21]/adc_array_circuit_150n_0/vint2 col_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5875 VDD rowon_n[11] adc_array_wafflecap_8_8_0[10|6]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5876 adc_array_wafflecap_8_8_0[7|17]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|17]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5877 adc_array_wafflecap_8_8_0[4|7]/adc_array_circuit_150n_0/vint1 col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5878 adc_array_wafflecap_8_8_0[4|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5879 adc_array_wafflecap_8_8_0[4|30]/adc_array_circuit_150n_0/vint2 rowon_n[5] adc_array_wafflecap_8_8_0[4|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5880 adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/vint2 rowon_n[1] adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5881 VSS row_n[7] adc_array_wafflecap_8_8_0[6|11]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5882 VSS row_n[15] adc_array_wafflecap_8_8_0[14|10]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5883 VSS row_n[15] adc_array_wafflecap_8_8_0[14|0]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5884 adc_array_wafflecap_8_8_0[3|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5885 adc_array_wafflecap_8_Dummy_4[8]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[8]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5886 VSS row_n[14] adc_array_wafflecap_8_8_0[13|14]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5887 adc_array_wafflecap_8_8_0[10|11]/adc_array_circuit_150n_0/vint2 col_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5888 adc_array_wafflecap_8_8_0[6|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5889 VSS row_n[0] adc_array_wafflecap_8_8_1[9]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5890 VDD rowon_n[2] adc_array_wafflecap_8_8_0[1|3]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5891 VSS row_n[14] adc_array_wafflecap_8_8_0[13|4]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5892 adc_array_wafflecap_8_8_0[10|1]/adc_array_circuit_150n_0/vint2 col_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5893 adc_array_wafflecap_8_Dummy_2[4]/adc_array_circuit_150n_0/vint1 col_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5894 adc_array_wafflecap_8_8_0[13|20]/adc_array_circuit_150n_0/vdrv row_n[14] adc_array_wafflecap_8_8_0[13|20]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5895 vcm adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|20]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5896 VDD rowon_n[5] adc_array_wafflecap_8_8_0[4|15]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5897 adc_array_wafflecap_8_8_0[2|26]/adc_array_circuit_150n_0/vdrv row_n[3] adc_array_wafflecap_8_8_0[2|26]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5898 vcm adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|10]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5899 adc_array_wafflecap_8_8_0[12|10]/adc_array_circuit_150n_0/vint1 col_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5900 adc_array_wafflecap_8_8_0[6|11]/adc_array_circuit_150n_0/vint1 col_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5901 adc_array_wafflecap_8_8_0[2|12]/adc_array_circuit_150n_0/vint1 col_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5902 adc_array_wafflecap_8_8_0[2|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5903 VDD rowon_n[0] adc_array_wafflecap_8_8_1[12]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5904 VSS row_n[2] adc_array_wafflecap_8_8_0[1|4]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5905 adc_array_wafflecap_8_8_0[12|0]/adc_array_circuit_150n_0/vint1 col_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5906 adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n sample VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5907 adc_array_wafflecap_8_8_0[9|24]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|24]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5908 adc_array_wafflecap_8_8_0[8|1]/adc_array_circuit_150n_0/vdrv row_n[9] adc_array_wafflecap_8_8_0[8|1]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5909 adc_array_wafflecap_8_8_0[8|11]/adc_array_circuit_150n_0/vdrv row_n[9] adc_array_wafflecap_8_8_0[8|11]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5910 adc_array_wafflecap_8_8_0[11|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5911 adc_array_wafflecap_8_8_0[11|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5912 adc_array_wafflecap_8_8_0[9|20]/adc_array_circuit_150n_0/vint2 rowon_n[10] adc_array_wafflecap_8_8_0[9|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5913 adc_array_wafflecap_8_8_0[3|19]/adc_array_circuit_150n_0/vint2 col_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5914 adc_array_wafflecap_8_8_0[4|30]/adc_array_circuit_150n_0/vdrv row_n[5] adc_array_wafflecap_8_8_0[4|30]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5915 vcm VSS adc_array_wafflecap_8_Dummy_8[1]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5916 vcm adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|2]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5917 adc_array_wafflecap_8_8_0[14|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5918 adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5919 vcm adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|15]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5920 adc_array_wafflecap_8_8_0[1|4]/adc_array_circuit_150n_0/vint1 col_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5921 adc_array_wafflecap_8_Dummy_4[20]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5922 adc_array_wafflecap_8_8_0[14|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5923 adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/vint2 rowon_n[15] adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5924 adc_array_wafflecap_8_8_0[7|5]/adc_array_circuit_150n_0/vint2 rowon_n[8] adc_array_wafflecap_8_8_0[7|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5925 adc_array_wafflecap_8_8_0[7|15]/adc_array_circuit_150n_0/vint2 rowon_n[8] adc_array_wafflecap_8_8_0[7|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5926 VSS row_n[12] adc_array_wafflecap_8_8_0[11|20]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5927 vcm adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|12]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5928 adc_array_wafflecap_8_8_0[8|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5929 adc_array_wafflecap_8_8_0[8|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5930 adc_array_wafflecap_8_8_1[27]/adc_array_circuit_150n_0/vdrv row_n[0] adc_array_wafflecap_8_8_1[27]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5931 adc_array_wafflecap_8_Dummy_4[30]/adc_array_circuit_150n_0/cbot VDD vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5932 adc_array_wafflecap_8_8_0[13|14]/adc_array_circuit_150n_0/vint2 rowon_n[14] adc_array_wafflecap_8_8_0[13|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5933 vcm adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|2]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5934 adc_array_wafflecap_8_8_1[13]/adc_array_circuit_150n_0/vint1 col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5935 adc_array_wafflecap_8_8_0[0|7]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|7]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5936 adc_array_wafflecap_8_8_0[13|4]/adc_array_circuit_150n_0/vint2 rowon_n[14] adc_array_wafflecap_8_8_0[13|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5937 VDD rowon_n[8] adc_array_wafflecap_8_8_0[7|20]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5938 adc_array_wafflecap_8_8_0[0|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5939 adc_array_wafflecap_8_8_0[11|30]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|30]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5940 VSS row_n[6] adc_array_wafflecap_8_8_0[5|25]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5941 VDD rowon_n[14] adc_array_wafflecap_8_8_0[13|19]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5942 adc_array_wafflecap_8_8_0[11|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5943 adc_array_wafflecap_8_8_0[12|6]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|6]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5944 adc_array_wafflecap_8_8_0[12|16]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|16]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5945 VDD rowon_n[13] adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5946 adc_array_wafflecap_8_8_1[19]/adc_array_circuit_150n_0/vint2 rowon_n[0] adc_array_wafflecap_8_8_1[19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5947 adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/vint2 VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5948 adc_array_wafflecap_8_Dummy_4[32]/adc_array_circuit_150n_0/vint2 col_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5949 VSS row_n[10] adc_array_wafflecap_8_8_0[9|9]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5950 adc_array_wafflecap_8_Dummy_1[3]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_1[3]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5951 vcm adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|24]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5952 adc_array_wafflecap_8_8_0[2|17]/adc_array_circuit_150n_0/vint2 rowon_n[3] adc_array_wafflecap_8_8_0[2|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5953 VSS VDD adc_array_wafflecap_8_Dummy_4[9]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5954 adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/vint1 col_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5955 adc_array_wafflecap_8_Dummy_4[19]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[19]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5956 adc_array_wafflecap_8_8_0[11|9]/adc_array_circuit_150n_0/vint2 col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5957 adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/vdrv row_n[8] adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5958 adc_array_wafflecap_8_8_0[11|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5959 adc_array_wafflecap_8_8_0[7|9]/adc_array_circuit_150n_0/vint1 col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5960 adc_array_wafflecap_8_Dummy_1[1]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_1[1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5961 adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/vdrv row_n[14] adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5962 vcm adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5963 adc_array_wafflecap_8_8_0[3|6]/adc_array_circuit_150n_0/vdrv row_n[4] adc_array_wafflecap_8_8_0[3|6]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5964 VSS row_n[4] adc_array_wafflecap_8_8_0[3|29]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5965 adc_array_wafflecap_8_8_0[2|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5966 adc_array_wafflecap_8_8_0[14|7]/adc_array_circuit_150n_0/vint2 col_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5967 VDD rowon_n[1] adc_array_wafflecap_8_8_0[0|17]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5968 adc_array_wafflecap_8_8_0[13|8]/adc_array_circuit_150n_0/vint1 col_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5969 adc_array_wafflecap_8_8_0[7|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5970 adc_array_wafflecap_8_8_0[6|22]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|22]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5971 adc_array_wafflecap_8_8_0[13|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5972 adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5973 adc_array_wafflecap_8_Dummy_1[0]/adc_array_circuit_150n_0/vint2 col_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5974 adc_array_wafflecap_8_8_0[2|8]/adc_array_circuit_150n_0/vint2 col_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5975 vcm adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|27]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5976 adc_array_wafflecap_8_8_1[20]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_1[20]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5977 vcm adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|28]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5978 VSS row_n[3] adc_array_wafflecap_8_8_0[2|18]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5979 vcm VSS adc_array_wafflecap_8_Dummy_4[33]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5980 adc_array_wafflecap_8_8_0[12|7]/adc_array_circuit_150n_0/vdrv row_n[13] adc_array_wafflecap_8_8_0[12|7]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5981 adc_array_wafflecap_8_8_0[10|18]/adc_array_circuit_150n_0/vint2 rowon_n[11] adc_array_wafflecap_8_8_0[10|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5982 adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/vint2 rowon_n[10] adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5983 adc_array_wafflecap_8_8_0[6|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5984 VDD rowon_n[6] adc_array_wafflecap_8_8_0[5|22]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5985 VDD sample_n adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5986 adc_array_wafflecap_8_8_0[9|9]/adc_array_circuit_150n_0/vint2 rowon_n[10] adc_array_wafflecap_8_8_0[9|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5987 vcm adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|18]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5988 adc_array_wafflecap_8_8_0[5|10]/adc_array_circuit_150n_0/vdrv row_n[6] adc_array_wafflecap_8_8_0[5|10]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5989 adc_array_wafflecap_8_8_0[5|11]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|11]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5990 adc_array_wafflecap_8_8_0[0|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5991 adc_array_wafflecap_8_Dummy_4[10]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5992 adc_array_wafflecap_8_8_0[8|13]/adc_array_circuit_150n_0/vint2 rowon_n[9] adc_array_wafflecap_8_8_0[8|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5993 adc_array_wafflecap_8_Dummy_4[0]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5994 adc_array_wafflecap_8_8_0[8|3]/adc_array_circuit_150n_0/vint2 rowon_n[9] adc_array_wafflecap_8_8_0[8|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5995 adc_array_wafflecap_8_8_0[0|8]/adc_array_circuit_150n_0/vdrv row_n[1] adc_array_wafflecap_8_8_0[0|8]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5996 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.64e+07u l=1.6e+07u
X5997 vcm adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|0]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5998 vcm adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|10]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5999 adc_array_wafflecap_8_8_0[0|18]/adc_array_circuit_150n_0/vint1 col_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6000 VDD rowon_n[9] adc_array_wafflecap_8_8_0[8|18]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6001 adc_array_wafflecap_8_8_0[4|24]/adc_array_circuit_150n_0/vint2 rowon_n[5] adc_array_wafflecap_8_8_0[4|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6002 VDD rowon_n[8] adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6003 adc_array_wafflecap_8_8_0[4|12]/adc_array_circuit_150n_0/vint2 col_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6004 adc_array_wafflecap_8_8_0[0|13]/adc_array_circuit_150n_0/vint2 col_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6005 VDD rowon_n[8] adc_array_wafflecap_8_8_0[7|9]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6006 vcm adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6007 VSS row_n[15] adc_array_wafflecap_8_8_0[14|29]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6008 adc_array_wafflecap_8_8_0[13|14]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|14]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6009 adc_array_wafflecap_8_8_0[11|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6010 adc_array_wafflecap_8_8_0[4|2]/adc_array_circuit_150n_0/vdrv row_n[5] adc_array_wafflecap_8_8_0[4|2]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6011 adc_array_wafflecap_8_8_0[4|3]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|3]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6012 adc_array_wafflecap_8_8_1[5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_1[5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6013 adc_array_wafflecap_8_8_0[0|4]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|4]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6014 adc_array_wafflecap_8_8_0[13|4]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|4]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6015 adc_array_wafflecap_8_8_0[3|15]/adc_array_circuit_150n_0/vdrv row_n[4] adc_array_wafflecap_8_8_0[3|15]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6016 adc_array_wafflecap_8_8_0[3|16]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|16]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6017 adc_array_wafflecap_8_8_0[10|30]/adc_array_circuit_150n_0/vint2 col_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6018 adc_array_wafflecap_8_Dummy_7/adc_array_circuit_150n_0/vdrv row_n[0] adc_array_wafflecap_8_Dummy_7/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6019 VSS row_n[11] adc_array_wafflecap_8_8_0[10|7]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6020 VDD rowon_n[4] adc_array_wafflecap_8_8_0[3|26]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6021 adc_array_wafflecap_8_Dummy_1[4]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_1[4]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6022 adc_array_wafflecap_8_8_0[14|25]/adc_array_circuit_150n_0/vdrv row_n[15] adc_array_wafflecap_8_8_0[14|25]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6023 adc_array_wafflecap_8_8_0[10|17]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|17]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6024 adc_array_wafflecap_8_8_1[4]/adc_array_circuit_150n_0/vint2 col_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6025 VDD VDD adc_array_wafflecap_8_Dummy_4[11]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6026 adc_array_wafflecap_8_8_0[12|29]/adc_array_circuit_150n_0/vint1 col_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6027 adc_array_wafflecap_8_8_0[9|26]/adc_array_circuit_150n_0/vdrv row_n[10] adc_array_wafflecap_8_8_0[9|26]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6028 VDD rowon_n[5] adc_array_wafflecap_8_8_0[4|8]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6029 adc_array_wafflecap_8_8_0[3|0]/adc_array_circuit_150n_0/vint2 rowon_n[4] adc_array_wafflecap_8_8_0[3|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6030 VDD VDD adc_array_wafflecap_8_Dummy_4[1]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6031 adc_array_wafflecap_8_8_0[8|30]/adc_array_circuit_150n_0/vdrv row_n[9] adc_array_wafflecap_8_8_0[8|30]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6032 VSS VSS adc_array_wafflecap_8_Dummy_2[2]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6033 vcm adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|24]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6034 adc_array_wafflecap_8_8_0[12|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6035 adc_array_wafflecap_8_Dummy_3[4]/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_3[4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6036 adc_array_wafflecap_8_8_0[2|28]/adc_array_circuit_150n_0/vint2 rowon_n[3] adc_array_wafflecap_8_8_0[2|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6037 adc_array_wafflecap_8_8_0[9|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6038 adc_array_wafflecap_8_8_0[8|7]/adc_array_circuit_150n_0/vint1 col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6039 adc_array_wafflecap_8_Dummy_2[0]/adc_array_circuit_150n_0/vint2 col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6040 adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6041 vcm adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|29]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6042 adc_array_wafflecap_8_8_0[14|18]/adc_array_circuit_150n_0/vint2 col_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6043 adc_array_wafflecap_8_8_0[5|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6044 VDD rowon_n[6] adc_array_wafflecap_8_8_0[5|30]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6045 adc_array_wafflecap_8_8_0[4|24]/adc_array_circuit_150n_0/vdrv row_n[5] adc_array_wafflecap_8_8_0[4|24]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6046 adc_array_wafflecap_8_8_1[10]/adc_array_circuit_150n_0/vint2 rowon_n[0] adc_array_wafflecap_8_8_1[10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6047 adc_array_wafflecap_8_8_0[1|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6048 VSS sample adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6049 VDD rowon_n[3] adc_array_wafflecap_8_8_0[2|13]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6050 adc_array_wafflecap_8_8_1[26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_1[26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6051 VDD rowon_n[1] adc_array_wafflecap_8_8_0[0|28]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6052 adc_array_wafflecap_8_8_0[1|5]/adc_array_circuit_150n_0/vint2 rowon_n[2] adc_array_wafflecap_8_8_0[1|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6053 adc_array_wafflecap_8_8_0[6|27]/adc_array_circuit_150n_0/vint2 col_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6054 vcm adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|7]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6055 adc_array_wafflecap_8_8_0[4|9]/adc_array_circuit_150n_0/vint1 col_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6056 vcm adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|8]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6057 adc_array_wafflecap_8_8_0[12|18]/adc_array_circuit_150n_0/vdrv row_n[13] adc_array_wafflecap_8_8_0[12|18]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6058 VSS row_n[13] adc_array_wafflecap_8_8_0[12|25]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6059 adc_array_wafflecap_8_8_0[10|7]/adc_array_circuit_150n_0/vint2 rowon_n[11] adc_array_wafflecap_8_8_0[10|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6060 adc_array_wafflecap_8_8_0[10|29]/adc_array_circuit_150n_0/vint2 rowon_n[11] adc_array_wafflecap_8_8_0[10|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6061 adc_array_wafflecap_8_8_0[5|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6062 adc_array_wafflecap_8_8_0[4|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6063 VSS row_n[4] adc_array_wafflecap_8_8_0[3|1]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6064 adc_array_wafflecap_8_8_0[1|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6065 adc_array_wafflecap_8_8_0[13|22]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|22]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6066 adc_array_wafflecap_8_8_0[3|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6067 adc_array_wafflecap_8_8_1[25]/adc_array_circuit_150n_0/vint2 col_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6068 adc_array_wafflecap_8_8_1[6]/adc_array_circuit_150n_0/vint1 col_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6069 adc_array_wafflecap_8_8_0[6|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6070 VDD rowon_n[15] adc_array_wafflecap_8_8_0[14|24]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6071 adc_array_wafflecap_8_8_0[12|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6072 adc_array_wafflecap_8_8_0[12|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6073 VDD sample_n adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6074 adc_array_wafflecap_8_8_0[9|9]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|9]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6075 VSS row_n[0] adc_array_wafflecap_8_8_1[11]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6076 VDD rowon_n[2] adc_array_wafflecap_8_8_0[1|5]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6077 adc_array_wafflecap_8_8_0[11|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6078 adc_array_wafflecap_8_8_0[10|25]/adc_array_circuit_150n_0/vint1 col_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6079 adc_array_wafflecap_8_8_0[5|16]/adc_array_circuit_150n_0/vint2 col_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6080 adc_array_wafflecap_8_8_0[11|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6081 VDD rowon_n[9] adc_array_wafflecap_8_8_0[8|7]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6082 VDD rowon_n[9] adc_array_wafflecap_8_8_0[8|29]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6083 adc_array_wafflecap_8_8_0[6|27]/adc_array_circuit_150n_0/vdrv row_n[7] adc_array_wafflecap_8_8_0[6|27]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6084 adc_array_wafflecap_8_8_0[2|28]/adc_array_circuit_150n_0/vdrv row_n[3] adc_array_wafflecap_8_8_0[2|28]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6085 adc_array_wafflecap_8_8_0[2|29]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|29]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6086 adc_array_wafflecap_8_8_1[2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6087 vcm adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|0]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6088 VSS VDD adc_array_wafflecap_8_Dummy_4[28]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6089 vcm adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|12]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6090 adc_array_wafflecap_8_8_0[2|14]/adc_array_circuit_150n_0/vint1 col_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6091 VSS sample adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/sample_n VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6092 adc_array_wafflecap_8_8_0[2|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/sample_n vcm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6093 VDD rowon_n[0] adc_array_wafflecap_8_8_1[14]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6094 adc_array_wafflecap_8_8_0[11|28]/adc_array_circuit_150n_0/vint2 col_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6095 adc_array_wafflecap_8_8_0[12|14]/adc_array_circuit_150n_0/vint2 col_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6096 VSS row_n[11] adc_array_wafflecap_8_8_0[10|18]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6097 VSS row_n[4] adc_array_wafflecap_8_8_0[3|23]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6098 adc_array_wafflecap_8_8_0[12|4]/adc_array_circuit_150n_0/vint2 col_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6099 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.64e+07u l=1.6e+07u
X6100 adc_array_wafflecap_8_Dummy_4[24]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[24]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6101 adc_array_wafflecap_8_8_0[13|27]/adc_array_circuit_150n_0/vint1 col_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6102 adc_array_wafflecap_8_8_0[12|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6103 vcm adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|23]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6104 adc_array_wafflecap_8_8_0[7|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6105 adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/sample_n sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6106 adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/vdrv row_n[5] adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6107 vcm VSS adc_array_wafflecap_8_Dummy_8[3]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6108 adc_array_wafflecap_8_8_0[14|13]/adc_array_circuit_150n_0/vint1 col_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6109 adc_array_wafflecap_8_8_0[14|3]/adc_array_circuit_150n_0/vint1 col_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6110 adc_array_wafflecap_8_8_0[9|17]/adc_array_circuit_150n_0/vint2 col_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6111 adc_array_wafflecap_8_8_1[29]/adc_array_circuit_150n_0/vdrv row_n[0] adc_array_wafflecap_8_8_1[29]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
.ends

