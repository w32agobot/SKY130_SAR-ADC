magic
tech sky130A
magscale 1 2
timestamp 1659713046
<< error_p >>
rect 342 1238 1144 1266
rect 342 1206 364 1238
rect 364 1026 370 1032
rect 402 1026 424 1206
rect 1122 1032 1144 1238
rect 1116 1026 1144 1032
rect 358 1024 365 1026
rect 342 964 365 1024
rect 358 962 365 964
rect 396 962 428 1026
rect 1121 962 1154 1026
rect 364 956 370 962
rect 364 786 370 792
rect 402 786 424 962
rect 1116 956 1144 962
rect 1122 792 1144 956
rect 1116 786 1144 792
rect 358 784 365 786
rect 342 724 365 784
rect 358 722 365 724
rect 396 722 428 786
rect 1121 722 1154 786
rect 364 716 370 722
rect 364 546 370 552
rect 402 546 424 722
rect 1116 716 1144 722
rect 1122 552 1144 716
rect 1116 546 1144 552
rect 358 544 365 546
rect 342 484 365 544
rect 358 482 365 484
rect 396 482 428 546
rect 1121 482 1154 546
rect 364 476 370 482
rect 364 306 370 312
rect 402 306 424 482
rect 1116 476 1144 482
rect 1122 312 1144 476
rect 1116 306 1144 312
rect 358 304 365 306
rect 342 244 365 304
rect 358 242 365 244
rect 396 242 428 306
rect 1121 242 1154 306
rect 364 236 370 242
rect 402 92 424 242
rect 1116 236 1144 242
rect 402 64 1084 92
rect 1122 64 1144 236
rect 432 58 486 64
rect 582 58 636 64
rect 848 58 902 64
rect 998 58 1052 64
<< metal1 >>
rect 364 1212 432 1238
rect 486 1212 582 1238
rect 636 1212 848 1238
rect 902 1212 998 1238
rect 1052 1212 1084 1238
rect 364 1208 1084 1212
rect 364 58 1084 64
rect 364 32 432 58
rect 486 32 582 58
rect 636 32 848 58
rect 902 32 998 58
rect 1052 32 1084 58
<< via1 >>
rect 432 1212 486 1238
rect 582 1212 636 1238
rect 848 1212 902 1238
rect 998 1212 1052 1238
rect 432 32 486 58
rect 582 32 636 58
rect 848 32 902 58
rect 998 32 1052 58
<< metal2 >>
rect 364 1212 432 1238
rect 486 1212 582 1238
rect 636 1212 848 1238
rect 902 1212 998 1238
rect 1052 1212 1122 1238
rect 364 1206 1122 1212
rect 364 1184 686 1206
rect 798 1184 1122 1206
rect 364 1048 656 1184
rect 714 1154 770 1178
rect 686 1148 798 1154
rect 686 1086 696 1148
rect 788 1086 798 1148
rect 686 1078 798 1086
rect 364 942 686 1048
rect 364 806 656 942
rect 714 912 770 1078
rect 828 1048 1122 1184
rect 798 942 1122 1048
rect 686 906 798 912
rect 686 844 696 906
rect 788 844 798 906
rect 686 836 798 844
rect 364 702 686 806
rect 364 566 656 702
rect 714 672 770 836
rect 828 806 1122 942
rect 798 702 1122 806
rect 686 666 798 672
rect 686 604 696 666
rect 788 604 798 666
rect 686 596 798 604
rect 364 462 686 566
rect 364 326 656 462
rect 714 432 770 596
rect 828 566 1122 702
rect 798 462 1122 566
rect 686 426 798 432
rect 686 364 696 426
rect 788 364 798 426
rect 686 356 798 364
rect 364 222 686 326
rect 364 88 656 222
rect 714 192 770 356
rect 828 326 1122 462
rect 798 222 1122 326
rect 686 186 798 192
rect 686 124 696 186
rect 788 124 798 186
rect 686 116 798 124
rect 714 92 770 116
rect 828 88 1122 222
rect 364 64 686 88
rect 798 64 1122 88
rect 364 58 1122 64
rect 364 32 432 58
rect 486 32 582 58
rect 636 32 848 58
rect 902 32 998 58
rect 1052 32 1122 58
<< via2 >>
rect 696 1086 788 1148
rect 696 844 788 906
rect 696 604 788 666
rect 696 364 788 426
rect 696 124 788 186
<< metal3 >>
rect 686 1148 798 1154
rect 686 1146 696 1148
rect 470 1086 696 1146
rect 788 1146 798 1148
rect 788 1086 1016 1146
rect 686 1078 798 1086
rect 396 1024 402 1026
rect 1084 1024 1090 1026
rect 396 964 656 1024
rect 828 964 1090 1024
rect 396 962 402 964
rect 1084 962 1090 964
rect 686 906 798 912
rect 686 904 696 906
rect 470 844 696 904
rect 788 904 798 906
rect 788 844 1016 904
rect 686 836 798 844
rect 396 784 402 786
rect 1084 784 1090 786
rect 396 724 656 784
rect 828 724 1090 784
rect 396 722 402 724
rect 1084 722 1090 724
rect 686 666 798 672
rect 686 664 696 666
rect 470 604 696 664
rect 788 664 798 666
rect 788 604 1016 664
rect 686 596 798 604
rect 396 544 402 546
rect 1084 544 1090 546
rect 396 484 656 544
rect 828 484 1090 544
rect 396 482 402 484
rect 1084 482 1090 484
rect 686 426 798 432
rect 686 424 696 426
rect 470 364 696 424
rect 788 424 798 426
rect 788 364 1016 424
rect 686 356 798 364
rect 396 304 402 306
rect 1084 304 1090 306
rect 396 244 656 304
rect 828 244 1090 304
rect 396 242 402 244
rect 1084 242 1090 244
rect 686 186 798 192
rect 686 184 696 186
rect 470 124 696 184
rect 788 184 798 186
rect 788 124 1016 184
rect 686 116 798 124
<< via3 >>
rect 364 962 396 1026
rect 1090 962 1122 1026
rect 364 722 396 786
rect 1090 722 1122 786
rect 364 482 396 546
rect 1090 482 1122 546
rect 364 242 396 306
rect 1090 242 1122 306
<< metal4 >>
rect 364 1206 1122 1238
rect 364 1026 402 1206
rect 396 962 402 1026
rect 364 786 402 962
rect 396 722 402 786
rect 364 546 402 722
rect 396 482 402 546
rect 364 306 402 482
rect 396 242 402 306
rect 364 64 402 242
rect 1084 1026 1122 1206
rect 1084 962 1090 1026
rect 1084 786 1122 962
rect 1084 722 1090 786
rect 1084 546 1122 722
rect 1084 482 1090 546
rect 1084 306 1122 482
rect 1084 242 1090 306
rect 1084 64 1122 242
rect 364 32 1122 64
<< end >>
