* NGSPICE file created from adc_array_matrix_12bit.ext - technology: sky130A

.subckt adc_array_wafflecap_dummy sample_n colon_n col_n sample vcom row_n ctop VDD
+ VSS
X0 VDD colon_n a_170_252# VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1 a_662_574# row_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2 a_170_252# col_n a_662_574# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3 a_566_252# colon_n a_170_252# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4 VSS col_n a_566_252# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5 a_566_252# row_n VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_262_252# sample_n a_170_252# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X7 vcom sample a_262_252# VSS sky130_fd_pr__nfet_01v8 ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X8 a_262_252# sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=2.48e+11p ps=2.22e+06u w=800000u l=150000u
X9 a_170_252# sample a_262_252# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
.ends

.subckt adc_array_wafflecap_drv ctop colon_n col_n vcom row_n sample_i sample_n_i
+ sample_n_o sample_o VDD VSS
X0 VSS sample_i sample_n_o VSS sky130_fd_pr__nfet_01v8 ad=5.208e+11p pd=5.84e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1 sample_n_o sample_i VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VDD sample_i sample_n_o VDD sky130_fd_pr__pfet_01v8 ad=9.92e+11p pd=8.88e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3 sample_n_o sample_i VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4 sample_o sample_n_i VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5 VSS sample_n_i sample_o VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 sample_o sample_n_i VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7 VDD sample_n_i sample_o VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
.ends

.subckt adc_array_wafflecap_1 sample_n colon_n col_n sample vcom row_n en_n ctop VDD
+ VSS
X0 VDD en_n a_170_252# VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1 a_662_574# en_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2 a_170_252# en_n a_662_574# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3 a_566_252# en_n a_170_252# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4 VSS en_n a_566_252# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5 a_566_252# en_n VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_262_252# sample_n a_170_252# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X7 vcom sample a_262_252# VSS sky130_fd_pr__nfet_01v8 ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X8 a_262_252# sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=2.48e+11p ps=2.22e+06u w=800000u l=150000u
X9 a_170_252# sample a_262_252# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
.ends

.subckt adc_array_wafflecap_8 sample_n colon_n col_n sample vcom row_n ctop VDD VSS
X0 VDD colon_n a_170_252# VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1 a_662_574# row_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2 a_170_252# col_n a_662_574# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3 a_566_252# colon_n a_170_252# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4 VSS col_n a_566_252# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5 a_566_252# row_n VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_262_252# sample_n a_170_252# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X7 vcom sample a_262_252# VSS sky130_fd_pr__nfet_01v8 ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X8 a_262_252# sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=2.48e+11p ps=2.22e+06u w=800000u l=150000u
X9 a_170_252# sample a_262_252# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
.ends

.subckt adc_noise_decoup_cell1 nmoscap_top nmoscap_bot mimcap_top mimcap_bot pwell
X0 mimcap_top mimcap_bot sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X1 nmoscap_bot nmoscap_top nmoscap_bot pwell sky130_fd_pr__nfet_01v8 ad=2.296e+13p pd=6.84e+07u as=0p ps=0u w=1.64e+07u l=1.6e+07u
.ends

.subckt adc_array_wafflecap_4 sample_n colon_n col_n sample vcom row_n en_n ctop VDD
+ VSS
X0 VDD en_n a_170_252# VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1 a_662_574# en_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2 a_170_252# en_n a_662_574# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3 a_566_252# en_n a_170_252# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4 VSS en_n a_566_252# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5 a_566_252# en_n VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_262_252# sample_n a_170_252# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X7 vcom sample a_262_252# VSS sky130_fd_pr__nfet_01v8 ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X8 a_262_252# sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=2.48e+11p ps=2.22e+06u w=800000u l=150000u
X9 a_170_252# sample a_262_252# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
.ends

.subckt adc_array_wafflecap_2 sample_n colon_n col_n sample vcom row_n en_n ctop VDD
+ VSS
X0 VDD en_n a_170_252# VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1 a_662_574# en_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2 a_170_252# en_n a_662_574# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3 a_566_252# en_n a_170_252# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4 VSS en_n a_566_252# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5 a_566_252# en_n VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_262_252# sample_n a_170_252# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X7 vcom sample a_262_252# VSS sky130_fd_pr__nfet_01v8 ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
X8 a_262_252# sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=2.48e+11p ps=2.22e+06u w=800000u l=150000u
X9 a_170_252# sample a_262_252# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
.ends

.subckt adc_array_wafflecap_gate sample_n colon_n col_n sample vcom row_n sw_n in
+ sw ctop VDD VSS
X0 ctop sw in VSS sky130_fd_pr__nfet_01v8 ad=1.45e+11p pd=1.58e+06u as=2.9e+11p ps=3.16e+06u w=500000u l=500000u
X1 in sw ctop VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=500000u
X2 ctop sw_n in VDD sky130_fd_pr__pfet_01v8 ad=1.45e+11p pd=1.58e+06u as=2.9e+11p ps=3.16e+06u w=500000u l=500000u
X3 in sw_n ctop VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=500000u
.ends

.subckt adc_array_matrix_12bit VDD VSS vcm sample sample_n row_n[15] row_n[14] row_n[13]
+ row_n[12] row_n[11] row_n[10] row_n[9] row_n[8] row_n[7] row_n[6] row_n[5] row_n[4]
+ row_n[3] row_n[2] row_n[1] row_n[0] rowon_n[15] rowon_n[14] rowon_n[13] rowon_n[12]
+ rowon_n[11] rowon_n[10] rowon_n[9] rowon_n[8] rowon_n[7] rowon_n[6] rowon_n[5] rowon_n[4]
+ rowon_n[3] rowon_n[2] rowon_n[1] rowon_n[0] col_n[31] col_n[30] col_n[29] col_n[28]
+ col_n[27] col_n[26] col_n[25] col_n[24] col_n[23] col_n[22] col_n[21] col_n[20]
+ col_n[19] col_n[18] col_n[17] col_n[16] col_n[15] col_n[14] col_n[13] col_n[12]
+ col_n[11] col_n[10] col_n[9] col_n[8] col_n[7] col_n[6] col_n[5] col_n[4] col_n[3]
+ col_n[2] col_n[1] col_n[0] en_bit_n[2] en_bit_n[1] en_bit_n[0] en_C0_n sw sw_n analog_in
+ ctop
Xadc_array_wafflecap_dummy_5[0] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm VDD adc_array_wafflecap_dummy_5[0]/ctop VDD
+ VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_5[1] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm VDD adc_array_wafflecap_dummy_5[1]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_5[2] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm VDD adc_array_wafflecap_dummy_5[2]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_5[3] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm VDD adc_array_wafflecap_dummy_5[3]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_5[4] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm VDD adc_array_wafflecap_dummy_5[4]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_5[5] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm VDD adc_array_wafflecap_dummy_5[5]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_5[6] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm VDD adc_array_wafflecap_dummy_5[6]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_5[7] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm VDD adc_array_wafflecap_dummy_5[7]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_5[8] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm VDD adc_array_wafflecap_dummy_5[8]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_5[9] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm VDD adc_array_wafflecap_dummy_5[9]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_5[10] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10]
+ row_n[10] adc_array_wafflecap_8_0[9|9]/sample vcm VDD adc_array_wafflecap_dummy_5[10]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_5[11] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm VDD adc_array_wafflecap_dummy_5[11]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_5[12] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm VDD adc_array_wafflecap_dummy_5[12]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_5[13] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm VDD adc_array_wafflecap_dummy_5[13]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_5[14] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm VDD adc_array_wafflecap_dummy_5[14]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_5[15] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm VDD adc_array_wafflecap_dummy_5[15]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_7 adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[0] adc_array_wafflecap_dummy_7/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_6 VDD VSS VSS VSS vcm VDD adc_array_wafflecap_dummy_6/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_8[0] VDD VSS VSS VSS vcm col_n[2] adc_array_wafflecap_dummy_8[0]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_8[1] VDD VSS VSS VSS vcm col_n[3] adc_array_wafflecap_dummy_8[1]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_8[2] VDD VSS VSS VSS vcm col_n[4] adc_array_wafflecap_dummy_8[2]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_8[3] VDD VSS VSS VSS vcm col_n[5] adc_array_wafflecap_dummy_8[3]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_8[4] VDD VSS VSS VSS vcm col_n[6] adc_array_wafflecap_dummy_8[4]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_8[5] VDD VSS VSS VSS vcm col_n[7] adc_array_wafflecap_dummy_8[5]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_drv_0[0] adc_array_wafflecap_drv_0[0]/ctop rowon_n[0] row_n[0]
+ vcm VDD sample sample_n adc_array_wafflecap_8_1[9]/sample_n adc_array_wafflecap_8_1[9]/sample
+ VDD VSS adc_array_wafflecap_drv
Xadc_array_wafflecap_drv_0[1] adc_array_wafflecap_drv_0[1]/ctop rowon_n[1] row_n[1]
+ vcm VDD sample sample_n adc_array_wafflecap_8_0[0|9]/sample_n adc_array_wafflecap_8_0[0|9]/sample
+ VDD VSS adc_array_wafflecap_drv
Xadc_array_wafflecap_drv_0[2] adc_array_wafflecap_drv_0[2]/ctop rowon_n[2] row_n[2]
+ vcm VDD sample sample_n adc_array_wafflecap_8_0[1|9]/sample_n adc_array_wafflecap_8_0[1|9]/sample
+ VDD VSS adc_array_wafflecap_drv
Xadc_array_wafflecap_drv_0[3] adc_array_wafflecap_drv_0[3]/ctop rowon_n[3] row_n[3]
+ vcm VDD sample sample_n adc_array_wafflecap_8_0[2|9]/sample_n adc_array_wafflecap_8_0[2|9]/sample
+ VDD VSS adc_array_wafflecap_drv
Xadc_array_wafflecap_drv_0[4] adc_array_wafflecap_drv_0[4]/ctop rowon_n[4] row_n[4]
+ vcm VDD sample sample_n adc_array_wafflecap_8_0[3|9]/sample_n adc_array_wafflecap_8_0[3|9]/sample
+ VDD VSS adc_array_wafflecap_drv
Xadc_array_wafflecap_drv_0[5] adc_array_wafflecap_drv_0[5]/ctop rowon_n[5] row_n[5]
+ vcm VDD sample sample_n adc_array_wafflecap_8_0[4|9]/sample_n adc_array_wafflecap_8_0[4|9]/sample
+ VDD VSS adc_array_wafflecap_drv
Xadc_array_wafflecap_drv_0[6] adc_array_wafflecap_drv_0[6]/ctop rowon_n[6] row_n[6]
+ vcm VDD sample sample_n adc_array_wafflecap_8_0[5|9]/sample_n adc_array_wafflecap_8_0[5|9]/sample
+ VDD VSS adc_array_wafflecap_drv
Xadc_array_wafflecap_drv_0[7] adc_array_wafflecap_drv_0[7]/ctop rowon_n[7] row_n[7]
+ vcm VDD sample sample_n adc_array_wafflecap_8_0[6|9]/sample_n adc_array_wafflecap_8_0[6|9]/sample
+ VDD VSS adc_array_wafflecap_drv
Xadc_array_wafflecap_drv_0[8] adc_array_wafflecap_drv_0[8]/ctop rowon_n[8] row_n[8]
+ vcm VDD sample sample_n adc_array_wafflecap_8_0[7|9]/sample_n adc_array_wafflecap_8_0[7|9]/sample
+ VDD VSS adc_array_wafflecap_drv
Xadc_array_wafflecap_drv_0[9] adc_array_wafflecap_drv_0[9]/ctop rowon_n[9] row_n[9]
+ vcm VDD sample sample_n adc_array_wafflecap_8_0[8|9]/sample_n adc_array_wafflecap_8_0[8|9]/sample
+ VDD VSS adc_array_wafflecap_drv
Xadc_array_wafflecap_drv_0[10] adc_array_wafflecap_drv_0[10]/ctop rowon_n[10] row_n[10]
+ vcm VDD sample sample_n adc_array_wafflecap_8_0[9|9]/sample_n adc_array_wafflecap_8_0[9|9]/sample
+ VDD VSS adc_array_wafflecap_drv
Xadc_array_wafflecap_drv_0[11] adc_array_wafflecap_drv_0[11]/ctop rowon_n[11] row_n[11]
+ vcm VDD sample sample_n adc_array_wafflecap_8_0[10|9]/sample_n adc_array_wafflecap_8_0[10|9]/sample
+ VDD VSS adc_array_wafflecap_drv
Xadc_array_wafflecap_drv_0[12] adc_array_wafflecap_drv_0[12]/ctop rowon_n[12] row_n[12]
+ vcm VDD sample sample_n adc_array_wafflecap_8_0[11|9]/sample_n adc_array_wafflecap_8_0[11|9]/sample
+ VDD VSS adc_array_wafflecap_drv
Xadc_array_wafflecap_drv_0[13] adc_array_wafflecap_drv_0[13]/ctop rowon_n[13] row_n[13]
+ vcm VDD sample sample_n adc_array_wafflecap_8_0[12|9]/sample_n adc_array_wafflecap_8_0[12|9]/sample
+ VDD VSS adc_array_wafflecap_drv
Xadc_array_wafflecap_drv_0[14] adc_array_wafflecap_drv_0[14]/ctop rowon_n[14] row_n[14]
+ vcm VDD sample sample_n adc_array_wafflecap_8_0[13|9]/sample_n adc_array_wafflecap_8_0[13|9]/sample
+ VDD VSS adc_array_wafflecap_drv
Xadc_array_wafflecap_drv_0[15] adc_array_wafflecap_drv_0[15]/ctop rowon_n[15] row_n[15]
+ vcm VDD sample sample_n adc_array_wafflecap_8_0[14|9]/sample_n adc_array_wafflecap_8_0[14|9]/sample
+ VDD VSS adc_array_wafflecap_drv
Xadc_array_wafflecap_1_0 VDD VSS VSS VSS vcm col_n[24] en_bit_n[0] ctop VDD VSS adc_array_wafflecap_1
Xadc_array_wafflecap_1_1 VDD VSS VSS VSS vcm col_n[1] en_C0_n ctop VDD VSS adc_array_wafflecap_1
Xadc_array_wafflecap_8_0[0|0] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[0] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|0] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[0] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|0] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[0] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|0] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[0] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|0] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[0] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|0] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[0] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|0] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[0] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|0] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[0] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|0] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[0] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|0] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[0] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|0] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[0] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|0] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[0] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|0] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[0] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|0] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[0] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|0] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[0] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|1] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[1] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|1] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[1] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|1] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[1] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|1] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[1] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|1] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[1] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|1] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[1] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|1] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[1] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|1] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[1] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|1] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[1] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|1] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[1] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|1] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[1] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|1] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[1] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|1] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[1] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|1] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[1] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|1] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[1] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|2] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[2] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|2] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[2] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|2] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[2] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|2] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[2] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|2] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[2] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|2] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[2] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|2] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[2] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|2] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[2] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|2] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[2] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|2] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[2] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|2] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[2] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|2] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[2] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|2] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[2] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|2] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[2] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|2] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[2] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|3] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[3] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|3] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[3] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|3] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[3] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|3] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[3] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|3] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[3] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|3] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[3] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|3] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[3] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|3] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[3] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|3] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[3] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|3] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[3] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|3] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[3] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|3] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[3] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|3] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[3] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|3] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[3] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|3] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[3] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|4] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[4] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|4] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[4] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|4] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[4] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|4] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[4] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|4] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[4] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|4] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[4] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|4] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[4] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|4] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[4] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|4] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[4] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|4] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[4] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|4] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[4] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|4] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[4] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|4] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[4] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|4] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[4] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|4] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[4] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|5] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[5] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|5] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[5] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|5] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[5] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|5] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[5] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|5] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[5] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|5] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[5] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|5] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[5] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|5] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[5] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|5] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[5] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|5] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[5] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|5] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[5] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|5] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[5] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|5] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[5] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|5] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[5] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|5] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[5] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|6] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[6] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|6] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[6] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|6] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[6] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|6] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[6] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|6] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[6] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|6] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[6] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|6] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[6] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|6] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[6] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|6] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[6] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|6] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[6] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|6] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[6] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|6] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[6] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|6] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[6] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|6] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[6] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|6] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[6] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|7] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[7] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|7] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[7] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|7] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[7] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|7] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[7] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|7] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[7] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|7] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[7] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|7] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[7] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|7] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[7] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|7] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[7] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|7] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[7] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|7] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[7] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|7] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[7] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|7] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[7] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|7] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[7] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|7] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[7] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|8] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[8] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|8] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[8] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|8] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[8] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|8] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[8] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|8] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[8] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|8] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[8] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|8] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[8] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|8] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[8] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|8] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[8] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|8] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[8] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|8] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[8] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|8] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[8] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|8] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[8] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|8] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[8] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|8] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[8] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|9] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[9] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|9] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[9] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|9] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[9] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|9] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[9] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|9] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[9] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|9] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[9] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|9] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[9] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|9] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[9] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|9] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[9] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|9] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[9] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|9] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[9] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|9] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[9] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|9] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[9] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|9] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[9] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|9] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[9] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|10] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[10] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|10] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[10] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|10] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[10] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|10] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[10] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|10] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[10] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|10] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[10] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|10] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[10] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|10] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[10] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|10] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[10] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|10] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[10] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|10] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[10] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|10] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[10] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|10] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[10] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|10] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[10] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|10] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[10] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|11] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[11] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|11] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[11] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|11] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[11] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|11] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[11] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|11] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[11] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|11] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[11] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|11] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[11] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|11] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[11] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|11] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[11] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|11] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[11] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|11] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[11] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|11] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[11] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|11] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[11] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|11] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[11] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|11] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[11] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|12] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[12] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|12] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[12] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|12] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[12] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|12] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[12] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|12] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[12] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|12] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[12] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|12] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[12] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|12] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[12] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|12] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[12] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|12] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[12] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|12] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[12] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|12] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[12] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|12] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[12] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|12] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[12] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|12] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[12] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|13] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[13] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|13] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[13] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|13] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[13] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|13] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[13] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|13] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[13] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|13] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[13] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|13] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[13] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|13] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[13] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|13] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[13] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|13] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[13] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|13] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[13] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|13] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[13] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|13] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[13] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|13] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[13] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|13] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[13] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|14] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[14] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|14] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[14] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|14] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[14] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|14] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[14] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|14] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[14] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|14] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[14] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|14] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[14] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|14] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[14] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|14] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[14] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|14] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[14] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|14] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[14] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|14] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[14] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|14] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[14] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|14] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[14] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|14] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[14] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|15] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[15] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|15] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[15] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|15] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[15] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|15] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[15] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|15] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[15] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|15] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[15] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|15] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[15] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|15] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[15] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|15] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[15] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|15] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[15] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|15] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[15] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|15] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[15] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|15] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[15] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|15] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[15] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|15] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[15] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|16] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[16] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|16] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[16] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|16] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[16] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|16] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[16] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|16] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[16] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|16] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[16] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|16] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[16] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|16] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[16] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|16] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[16] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|16] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[16] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|16] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[16] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|16] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[16] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|16] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[16] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|16] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[16] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|16] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[16] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|17] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[17] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|17] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[17] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|17] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[17] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|17] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[17] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|17] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[17] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|17] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[17] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|17] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[17] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|17] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[17] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|17] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[17] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|17] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[17] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|17] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[17] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|17] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[17] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|17] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[17] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|17] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[17] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|17] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[17] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|18] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[18] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|18] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[18] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|18] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[18] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|18] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[18] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|18] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[18] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|18] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[18] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|18] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[18] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|18] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[18] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|18] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[18] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|18] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[18] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|18] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[18] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|18] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[18] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|18] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[18] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|18] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[18] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|18] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[18] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|19] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[19] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|19] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[19] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|19] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[19] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|19] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[19] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|19] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[19] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|19] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[19] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|19] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[19] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|19] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[19] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|19] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[19] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|19] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[19] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|19] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[19] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|19] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[19] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|19] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[19] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|19] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[19] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|19] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[19] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|20] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[20] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|20] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[20] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|20] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[20] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|20] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[20] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|20] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[20] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|20] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[20] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|20] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[20] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|20] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[20] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|20] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[20] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|20] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[20] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|20] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[20] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|20] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[20] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|20] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[20] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|20] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[20] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|20] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[20] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|21] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[21] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|21] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[21] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|21] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[21] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|21] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[21] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|21] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[21] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|21] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[21] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|21] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[21] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|21] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[21] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|21] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[21] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|21] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[21] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|21] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[21] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|21] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[21] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|21] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[21] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|21] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[21] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|21] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[21] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|22] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[22] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|22] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[22] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|22] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[22] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|22] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[22] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|22] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[22] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|22] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[22] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|22] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[22] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|22] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[22] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|22] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[22] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|22] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[22] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|22] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[22] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|22] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[22] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|22] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[22] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|22] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[22] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|22] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[22] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|23] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[23] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|23] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[23] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|23] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[23] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|23] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[23] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|23] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[23] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|23] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[23] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|23] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[23] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|23] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[23] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|23] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[23] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|23] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[23] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|23] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[23] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|23] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[23] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|23] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[23] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|23] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[23] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|23] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[23] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|24] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[24] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|24] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[24] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|24] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[24] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|24] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[24] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|24] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[24] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|24] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[24] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|24] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[24] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|24] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[24] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|24] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[24] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|24] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[24] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|24] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[24] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|24] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[24] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|24] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[24] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|24] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[24] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|24] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[24] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|25] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[25] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|25] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[25] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|25] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[25] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|25] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[25] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|25] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[25] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|25] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[25] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|25] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[25] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|25] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[25] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|25] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[25] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|25] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[25] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|25] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[25] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|25] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[25] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|25] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[25] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|25] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[25] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|25] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[25] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|26] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[26] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|26] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[26] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|26] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[26] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|26] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[26] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|26] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[26] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|26] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[26] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|26] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[26] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|26] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[26] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|26] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[26] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|26] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[26] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|26] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[26] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|26] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[26] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|26] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[26] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|26] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[26] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|26] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[26] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|27] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[27] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|27] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[27] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|27] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[27] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|27] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[27] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|27] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[27] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|27] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[27] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|27] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[27] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|27] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[27] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|27] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[27] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|27] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[27] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|27] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[27] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|27] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[27] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|27] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[27] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|27] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[27] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|27] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[27] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|28] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[28] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|28] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[28] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|28] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[28] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|28] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[28] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|28] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[28] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|28] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[28] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|28] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[28] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|28] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[28] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|28] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[28] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|28] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[28] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|28] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[28] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|28] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[28] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|28] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[28] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|28] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[28] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|28] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[28] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|29] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[29] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|29] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[29] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|29] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[29] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|29] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[29] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|29] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[29] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|29] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[29] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|29] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[29] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|29] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[29] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|29] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[29] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|29] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[29] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|29] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[29] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|29] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[29] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|29] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[29] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|29] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[29] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|29] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[29] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|30] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[30] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|30] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[30] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|30] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[30] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|30] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[30] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|30] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[30] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|30] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[30] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|30] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[30] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|30] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[30] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|30] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[30] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|30] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[30] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|30] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[30] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|30] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[30] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|30] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[30] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|30] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[30] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|30] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[30] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|31] adc_array_wafflecap_8_0[0|9]/sample_n rowon_n[1] row_n[1]
+ adc_array_wafflecap_8_0[0|9]/sample vcm col_n[31] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|31] adc_array_wafflecap_8_0[1|9]/sample_n rowon_n[2] row_n[2]
+ adc_array_wafflecap_8_0[1|9]/sample vcm col_n[31] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|31] adc_array_wafflecap_8_0[2|9]/sample_n rowon_n[3] row_n[3]
+ adc_array_wafflecap_8_0[2|9]/sample vcm col_n[31] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|31] adc_array_wafflecap_8_0[3|9]/sample_n rowon_n[4] row_n[4]
+ adc_array_wafflecap_8_0[3|9]/sample vcm col_n[31] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|31] adc_array_wafflecap_8_0[4|9]/sample_n rowon_n[5] row_n[5]
+ adc_array_wafflecap_8_0[4|9]/sample vcm col_n[31] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|31] adc_array_wafflecap_8_0[5|9]/sample_n rowon_n[6] row_n[6]
+ adc_array_wafflecap_8_0[5|9]/sample vcm col_n[31] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|31] adc_array_wafflecap_8_0[6|9]/sample_n rowon_n[7] row_n[7]
+ adc_array_wafflecap_8_0[6|9]/sample vcm col_n[31] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|31] adc_array_wafflecap_8_0[7|9]/sample_n rowon_n[8] row_n[8]
+ adc_array_wafflecap_8_0[7|9]/sample vcm col_n[31] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|31] adc_array_wafflecap_8_0[8|9]/sample_n rowon_n[9] row_n[9]
+ adc_array_wafflecap_8_0[8|9]/sample vcm col_n[31] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|31] adc_array_wafflecap_8_0[9|9]/sample_n rowon_n[10] row_n[10]
+ adc_array_wafflecap_8_0[9|9]/sample vcm col_n[31] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|31] adc_array_wafflecap_8_0[10|9]/sample_n rowon_n[11]
+ row_n[11] adc_array_wafflecap_8_0[10|9]/sample vcm col_n[31] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|31] adc_array_wafflecap_8_0[11|9]/sample_n rowon_n[12]
+ row_n[12] adc_array_wafflecap_8_0[11|9]/sample vcm col_n[31] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|31] adc_array_wafflecap_8_0[12|9]/sample_n rowon_n[13]
+ row_n[13] adc_array_wafflecap_8_0[12|9]/sample vcm col_n[31] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|31] adc_array_wafflecap_8_0[13|9]/sample_n rowon_n[14]
+ row_n[14] adc_array_wafflecap_8_0[13|9]/sample vcm col_n[31] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|31] adc_array_wafflecap_8_0[14|9]/sample_n rowon_n[15]
+ row_n[15] adc_array_wafflecap_8_0[14|9]/sample vcm col_n[31] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[0] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[1] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[1] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[2] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[2] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[3] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[3] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[4] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[4] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[5] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[5] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[6] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[6] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[7] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[7] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[8] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[8] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[9] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[9] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[10] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[10] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[11] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[11] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[12] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[12] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[13] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[13] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[14] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[14] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[15] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[15] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[16] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[16] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[17] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[17] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[18] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[18] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[19] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[19] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[20] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[20] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[21] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[21] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[22] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[22] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[23] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[23] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[24] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[24] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[25] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[25] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[26] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[26] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[27] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[27] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[28] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[28] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[29] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[29] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[30] ctop VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[30] adc_array_wafflecap_8_1[9]/sample_n rowon_n[0] row_n[0]
+ adc_array_wafflecap_8_1[9]/sample vcm col_n[31] ctop VDD VSS adc_array_wafflecap_8
Xadc_noise_decoup_cell1_0[0] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[1] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[2] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[3] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[4] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[5] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[0] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[1] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[2] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[3] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[4] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[5] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[6] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[7] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[8] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_array_wafflecap_4_0 VDD VSS VSS VSS vcm col_n[8] en_bit_n[2] ctop VDD VSS adc_array_wafflecap_4
Xadc_array_wafflecap_2_0 VDD VSS VSS VSS vcm col_n[16] en_bit_n[1] ctop VDD VSS adc_array_wafflecap_2
Xadc_array_wafflecap_dummy_0[0] VDD VSS VSS VSS vcm VDD adc_array_wafflecap_dummy_0[0]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_0[1] VDD VSS VSS VSS vcm col_n[0] adc_array_wafflecap_dummy_0[1]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_1[0] VDD VSS VSS VSS vcm col_n[9] adc_array_wafflecap_dummy_1[0]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_1[1] VDD VSS VSS VSS vcm col_n[10] adc_array_wafflecap_dummy_1[1]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_1[2] VDD VSS VSS VSS vcm col_n[11] adc_array_wafflecap_dummy_1[2]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_1[3] VDD VSS VSS VSS vcm col_n[12] ctop VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_1[4] VDD VSS VSS VSS vcm col_n[13] adc_array_wafflecap_dummy_1[4]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_1[5] VDD VSS VSS VSS vcm col_n[14] adc_array_wafflecap_dummy_1[5]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_1[6] VDD VSS VSS VSS vcm col_n[15] adc_array_wafflecap_dummy_1[6]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_2[0] VDD VSS VSS VSS vcm col_n[17] adc_array_wafflecap_dummy_2[0]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_2[1] VDD VSS VSS VSS vcm col_n[18] adc_array_wafflecap_dummy_2[1]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_2[2] VDD VSS VSS VSS vcm col_n[19] adc_array_wafflecap_dummy_2[2]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_2[3] VDD VSS VSS VSS vcm col_n[20] adc_array_wafflecap_dummy_2[3]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_2[4] VDD VSS VSS VSS vcm col_n[21] adc_array_wafflecap_dummy_2[4]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_2[5] VDD VSS VSS VSS vcm col_n[22] adc_array_wafflecap_dummy_2[5]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_2[6] VDD VSS VSS VSS vcm col_n[23] adc_array_wafflecap_dummy_2[6]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_3[0] VDD VSS VSS VSS vcm col_n[25] adc_array_wafflecap_dummy_3[0]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_3[1] VDD VSS VSS VSS vcm col_n[26] adc_array_wafflecap_dummy_3[1]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_3[2] VDD VSS VSS VSS vcm col_n[27] adc_array_wafflecap_dummy_3[2]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_3[3] VDD VSS VSS VSS vcm col_n[28] adc_array_wafflecap_dummy_3[3]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_3[4] VDD VSS VSS VSS vcm col_n[29] adc_array_wafflecap_dummy_3[4]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_3[5] VDD VSS VSS VSS vcm col_n[30] adc_array_wafflecap_dummy_3[5]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[0] VDD VDD VDD VSS vcm VDD adc_array_wafflecap_dummy_4[0]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[1] VDD VDD VDD VSS vcm col_n[0] adc_array_wafflecap_dummy_4[1]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[2] VDD VDD VDD VSS vcm col_n[1] adc_array_wafflecap_dummy_4[2]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[3] VDD VDD VDD VSS vcm col_n[2] adc_array_wafflecap_dummy_4[3]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[4] VDD VDD VDD VSS vcm col_n[3] adc_array_wafflecap_dummy_4[4]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[5] VDD VDD VDD VSS vcm col_n[4] adc_array_wafflecap_dummy_4[5]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[6] VDD VDD VDD VSS vcm col_n[5] adc_array_wafflecap_dummy_4[6]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[7] VDD VDD VDD VSS vcm col_n[6] adc_array_wafflecap_dummy_4[7]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[8] VDD VDD VDD VSS vcm col_n[7] adc_array_wafflecap_dummy_4[8]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[9] VDD VDD VDD VSS vcm col_n[8] adc_array_wafflecap_dummy_4[9]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[10] VDD VDD VDD VSS vcm col_n[9] adc_array_wafflecap_dummy_4[10]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[11] VDD VDD VDD VSS vcm col_n[10] adc_array_wafflecap_dummy_4[11]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[12] VDD VDD VDD VSS vcm col_n[11] adc_array_wafflecap_dummy_4[12]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[13] VDD VDD VDD VSS vcm col_n[12] adc_array_wafflecap_dummy_4[13]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[14] VDD VDD VDD VSS vcm col_n[13] adc_array_wafflecap_dummy_4[14]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[15] VDD VDD VDD VSS vcm col_n[14] adc_array_wafflecap_dummy_4[15]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[16] VDD VDD VDD VSS vcm col_n[15] adc_array_wafflecap_dummy_4[16]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[17] VDD VDD VDD VSS vcm col_n[16] adc_array_wafflecap_dummy_4[17]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[18] VDD VDD VDD VSS vcm col_n[17] adc_array_wafflecap_dummy_4[18]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[19] VDD VDD VDD VSS vcm col_n[18] adc_array_wafflecap_dummy_4[19]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[20] VDD VDD VDD VSS vcm col_n[19] adc_array_wafflecap_dummy_4[20]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[21] VDD VDD VDD VSS vcm col_n[20] adc_array_wafflecap_dummy_4[21]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[22] VDD VDD VDD VSS vcm col_n[21] adc_array_wafflecap_dummy_4[22]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[23] VDD VDD VDD VSS vcm col_n[22] adc_array_wafflecap_dummy_4[23]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[24] VDD VDD VDD VSS vcm col_n[23] adc_array_wafflecap_dummy_4[24]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[25] VDD VDD VDD VSS vcm col_n[24] adc_array_wafflecap_dummy_4[25]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[26] VDD VDD VDD VSS vcm col_n[25] adc_array_wafflecap_dummy_4[26]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[27] VDD VDD VDD VSS vcm col_n[26] adc_array_wafflecap_dummy_4[27]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[28] VDD VDD VDD VSS vcm col_n[27] adc_array_wafflecap_dummy_4[28]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[29] VDD VDD VDD VSS vcm col_n[28] adc_array_wafflecap_dummy_4[29]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[30] VDD VDD VDD VSS vcm col_n[29] adc_array_wafflecap_dummy_4[30]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[31] VDD VDD VDD VSS vcm col_n[30] adc_array_wafflecap_dummy_4[31]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[32] VDD VDD VDD VSS vcm col_n[31] adc_array_wafflecap_dummy_4[32]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[33] VDD VDD VDD VSS vcm VDD adc_array_wafflecap_dummy_4[33]/ctop
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_gate_0 VDD VSS VSS VSS vcm col_n[31] sw_n analog_in sw ctop VDD
+ VSS adc_array_wafflecap_gate
.ends

