* NGSPICE file created from sky130_mm_sc_hd_dlyxnsB.ext - technology: sky130A

.subckt sky130_mm_sc_hd_dlyxnsB in out VPWR VGND VNB VPB
X0 a_1184_80# out VPWR VNB sky130_fd_pr__nfet_01v8 ad=3.99e+11p pd=4.42e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1 VPWR out a_1184_80# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND out a_1162_296# VPB sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=7.52e+11p ps=6.68e+06u w=800000u l=150000u
X3 a_1162_296# out VGND VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4 cap_top in VGND VNB sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=2.478e+11p ps=2.86e+06u w=420000u l=3.995e+06u
X5 a_1162_296# cap_top VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.72e+11p ps=4.38e+06u w=800000u l=150000u
X6 out cap_top a_1162_296# VPB sky130_fd_pr__pfet_01v8 ad=2.4e+11p pd=2.2e+06u as=0p ps=0u w=800000u l=150000u
X7 cap_top in VPWR VPB sky130_fd_pr__pfet_01v8_lvt ad=2.32e+11p pd=2.18e+06u as=0p ps=0u w=800000u l=3.995e+06u
X8 out cap_top a_1184_80# VNB sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=0p ps=0u w=420000u l=150000u
X9 a_1184_80# cap_top VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
C0 in out 0.03fF
C1 VGND a_1184_80# 1.07fF
C2 VPB out 0.07fF
C3 VPWR a_1184_80# 0.10fF
C4 VPB in 0.22fF
C5 cap_top out 0.05fF
C6 cap_top in 0.07fF
C7 cap_top VPB 0.06fF
C8 out a_1184_80# 0.35fF
C9 in a_1184_80# 0.02fF
C10 VPB a_1184_80# 0.00fF
C11 cap_top a_1184_80# 0.01fF
C12 VGND a_1162_296# 0.16fF
C13 VPWR a_1162_296# 1.12fF
C14 out a_1162_296# 0.41fF
C15 in a_1162_296# 0.03fF
C16 VPB a_1162_296# 0.03fF
C17 cap_top a_1162_296# 0.01fF
C18 a_1184_80# a_1162_296# 0.02fF
C19 VPWR VGND 0.32fF
C20 VGND out 0.14fF
C21 VPWR out 0.15fF
C22 VGND in 0.14fF
C23 VPWR in 0.17fF
C24 VGND VPB 0.09fF
C25 VPWR VPB 0.27fF
C26 VGND cap_top 0.12fF
C27 VPWR cap_top 0.15fF
.ends

