VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO adc_comp_latch
  CLASS BLOCK ;
  FOREIGN adc_comp_latch ;
  ORIGIN 0.000 0.000 ;
  SIZE 30.050 BY 27.980 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 18.380 18.020 26.290 18.040 ;
        RECT 6.590 16.000 26.290 18.020 ;
        RECT 6.590 15.910 18.050 16.000 ;
        RECT 9.220 15.900 10.430 15.910 ;
        RECT 12.260 14.160 18.050 15.910 ;
        RECT 21.240 15.760 26.290 16.000 ;
        RECT 4.230 12.070 6.440 14.060 ;
        RECT 22.040 12.300 24.610 12.560 ;
        RECT 18.560 10.280 24.610 12.300 ;
      LAYER li1 ;
        RECT 18.390 17.650 21.130 18.140 ;
        RECT 21.680 17.690 25.910 17.860 ;
        RECT 5.700 17.190 11.060 17.430 ;
        RECT 13.280 17.240 16.900 17.480 ;
        RECT 5.700 14.060 6.130 17.190 ;
        RECT 6.840 17.100 10.850 17.190 ;
        RECT 6.840 16.390 7.010 17.100 ;
        RECT 7.800 16.390 7.970 17.100 ;
        RECT 8.760 16.390 8.930 17.100 ;
        RECT 9.720 16.390 9.890 17.100 ;
        RECT 10.680 16.390 10.850 17.100 ;
        RECT 14.960 17.070 15.410 17.240 ;
        RECT 14.110 16.900 16.200 17.070 ;
        RECT 14.110 14.640 14.280 16.900 ;
        RECT 15.070 14.640 15.240 16.900 ;
        RECT 16.030 14.640 16.200 16.900 ;
        RECT 19.280 16.290 19.450 17.650 ;
        RECT 20.240 16.290 20.410 17.650 ;
        RECT 4.100 13.860 6.130 14.060 ;
        RECT 4.100 12.940 4.280 13.860 ;
        RECT 4.540 13.700 4.960 13.860 ;
        RECT 5.230 12.940 5.450 13.860 ;
        RECT 5.710 13.700 6.130 13.860 ;
        RECT 4.100 12.750 4.980 12.940 ;
        RECT 5.230 12.750 6.150 12.940 ;
        RECT 19.280 10.650 19.450 12.010 ;
        RECT 20.240 10.650 20.410 12.010 ;
        RECT 20.850 10.650 21.130 17.650 ;
        RECT 22.440 16.250 22.610 17.690 ;
        RECT 24.920 16.250 25.090 17.690 ;
        RECT 18.400 10.630 21.130 10.650 ;
        RECT 23.240 10.630 23.410 12.070 ;
        RECT 18.400 10.460 24.230 10.630 ;
      LAYER mcon ;
        RECT 18.860 17.860 19.040 18.040 ;
        RECT 19.240 17.860 19.420 18.040 ;
        RECT 19.620 17.860 19.800 18.040 ;
        RECT 20.000 17.860 20.180 18.040 ;
        RECT 20.380 17.860 20.560 18.040 ;
        RECT 20.760 17.860 20.940 18.040 ;
        RECT 5.760 17.220 5.930 17.400 ;
        RECT 6.150 17.220 6.320 17.400 ;
        RECT 6.510 17.220 6.680 17.400 ;
        RECT 6.930 17.220 7.100 17.390 ;
        RECT 7.350 17.220 7.520 17.390 ;
        RECT 7.770 17.220 7.940 17.390 ;
        RECT 8.190 17.220 8.360 17.390 ;
        RECT 8.610 17.220 8.780 17.390 ;
        RECT 9.030 17.220 9.200 17.390 ;
        RECT 9.450 17.220 9.620 17.390 ;
        RECT 9.870 17.220 10.040 17.390 ;
        RECT 10.290 17.220 10.460 17.390 ;
        RECT 10.740 17.220 10.910 17.390 ;
        RECT 13.470 17.270 13.640 17.440 ;
        RECT 13.890 17.270 14.060 17.440 ;
        RECT 14.310 17.270 14.480 17.440 ;
        RECT 14.730 17.270 14.900 17.440 ;
        RECT 15.150 17.270 15.320 17.440 ;
        RECT 15.570 17.270 15.740 17.440 ;
        RECT 15.990 17.270 16.160 17.440 ;
        RECT 16.410 17.270 16.580 17.440 ;
        RECT 4.660 13.890 4.840 14.060 ;
        RECT 5.830 13.890 6.010 14.060 ;
      LAYER met1 ;
        RECT 0.000 17.700 29.920 18.850 ;
        RECT 5.700 17.190 11.060 17.700 ;
        RECT 13.280 17.240 16.900 17.700 ;
        RECT 4.500 13.860 4.990 14.090 ;
        RECT 5.670 13.860 6.160 14.090 ;
      LAYER via ;
        RECT 0.320 17.790 1.120 18.740 ;
        RECT 29.020 17.790 29.820 18.740 ;
      LAYER met2 ;
        RECT 0.230 17.700 1.230 18.850 ;
        RECT 28.920 17.700 29.920 18.850 ;
      LAYER via2 ;
        RECT 0.320 17.790 1.120 18.740 ;
        RECT 29.020 17.790 29.820 18.740 ;
      LAYER met3 ;
        RECT 0.230 17.700 1.230 18.850 ;
        RECT 28.920 17.700 29.920 18.850 ;
      LAYER via3 ;
        RECT 0.320 17.790 1.120 18.740 ;
        RECT 29.020 17.790 29.820 18.740 ;
      LAYER met4 ;
        RECT 0.230 0.000 1.230 27.980 ;
        RECT 28.920 0.000 29.920 27.980 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER pwell ;
        RECT 7.320 25.990 9.720 26.890 ;
        RECT 20.220 25.990 22.620 26.890 ;
        RECT 5.020 25.590 11.270 25.990 ;
        RECT 14.520 25.590 15.420 25.990 ;
        RECT 18.670 25.590 24.920 25.990 ;
        RECT 5.020 20.290 24.920 25.590 ;
        RECT 5.020 19.890 11.270 20.290 ;
        RECT 14.520 19.890 15.420 20.290 ;
        RECT 18.670 19.890 24.920 20.290 ;
        RECT 7.320 18.990 9.720 19.890 ;
        RECT 20.220 18.990 22.620 19.890 ;
        RECT 7.320 8.040 9.720 8.940 ;
        RECT 20.220 8.040 22.620 8.940 ;
        RECT 5.020 7.640 11.270 8.040 ;
        RECT 14.520 7.640 15.420 8.040 ;
        RECT 18.670 7.640 24.920 8.040 ;
        RECT 5.020 2.340 24.920 7.640 ;
        RECT 5.020 1.940 11.270 2.340 ;
        RECT 14.520 1.940 15.420 2.340 ;
        RECT 18.670 1.940 24.920 2.340 ;
        RECT 7.320 1.040 9.720 1.940 ;
        RECT 20.220 1.040 22.620 1.940 ;
      LAYER li1 ;
        RECT 2.940 26.990 27.330 27.980 ;
        RECT 2.940 24.540 4.120 26.990 ;
        RECT 7.370 26.490 9.670 26.990 ;
        RECT 20.270 26.490 22.570 26.990 ;
        RECT 4.520 26.090 25.420 26.490 ;
        RECT 2.940 0.990 3.930 24.540 ;
        RECT 4.520 19.790 4.920 26.090 ;
        RECT 7.370 26.040 9.670 26.090 ;
        RECT 20.270 26.040 22.570 26.090 ;
        RECT 5.720 24.890 24.220 25.490 ;
        RECT 8.320 24.290 8.670 24.890 ;
        RECT 6.070 24.090 8.670 24.290 ;
        RECT 8.320 23.490 8.670 24.090 ;
        RECT 6.070 23.290 8.670 23.490 ;
        RECT 9.270 23.390 9.470 24.890 ;
        RECT 10.070 23.390 10.270 24.890 ;
        RECT 10.870 23.390 11.070 24.890 ;
        RECT 11.670 23.390 11.870 24.890 ;
        RECT 12.470 23.390 12.670 24.890 ;
        RECT 13.270 23.390 13.470 24.890 ;
        RECT 14.070 23.390 14.270 24.890 ;
        RECT 14.870 23.390 15.070 24.890 ;
        RECT 15.670 23.390 15.870 24.890 ;
        RECT 16.470 23.390 16.670 24.890 ;
        RECT 17.270 23.390 17.470 24.890 ;
        RECT 18.070 23.390 18.270 24.890 ;
        RECT 18.870 23.390 19.070 24.890 ;
        RECT 19.670 23.390 19.870 24.890 ;
        RECT 20.470 23.390 20.670 24.890 ;
        RECT 21.270 24.290 21.620 24.890 ;
        RECT 21.270 24.090 23.870 24.290 ;
        RECT 21.270 23.490 21.620 24.090 ;
        RECT 21.270 23.290 23.820 23.490 ;
        RECT 6.070 22.390 8.670 22.590 ;
        RECT 8.320 21.790 8.670 22.390 ;
        RECT 6.070 21.590 8.670 21.790 ;
        RECT 8.320 20.990 8.670 21.590 ;
        RECT 9.270 20.990 9.470 22.490 ;
        RECT 10.070 20.990 10.270 22.490 ;
        RECT 10.870 20.990 11.070 22.490 ;
        RECT 11.670 20.990 11.870 22.490 ;
        RECT 12.470 20.990 12.670 22.490 ;
        RECT 13.270 20.990 13.470 22.490 ;
        RECT 14.070 20.990 14.270 22.490 ;
        RECT 14.870 20.990 15.070 22.490 ;
        RECT 15.670 20.990 15.870 22.490 ;
        RECT 16.470 20.990 16.670 22.490 ;
        RECT 17.270 20.990 17.470 22.490 ;
        RECT 18.070 20.990 18.270 22.490 ;
        RECT 18.870 20.990 19.070 22.490 ;
        RECT 19.670 20.990 19.870 22.490 ;
        RECT 20.470 20.990 20.670 22.490 ;
        RECT 21.270 22.390 23.820 22.590 ;
        RECT 21.270 21.790 21.620 22.390 ;
        RECT 21.270 21.590 23.870 21.790 ;
        RECT 21.270 20.990 21.620 21.590 ;
        RECT 5.720 20.390 24.220 20.990 ;
        RECT 7.370 19.790 9.670 19.840 ;
        RECT 20.270 19.790 22.570 19.840 ;
        RECT 25.020 19.790 25.420 26.090 ;
        RECT 4.520 19.390 25.420 19.790 ;
        RECT 7.370 18.990 9.670 19.390 ;
        RECT 20.270 18.990 22.570 19.390 ;
        RECT 19.280 14.410 19.450 15.200 ;
        RECT 20.240 14.410 20.410 15.200 ;
        RECT 21.960 14.740 22.130 15.440 ;
        RECT 24.440 14.740 24.610 15.440 ;
        RECT 26.340 14.740 27.330 26.990 ;
        RECT 21.830 14.480 27.330 14.740 ;
        RECT 18.740 14.320 20.520 14.410 ;
        RECT 18.060 13.980 20.520 14.320 ;
        RECT 4.520 11.060 4.980 11.230 ;
        RECT 5.690 11.060 6.150 11.230 ;
        RECT 4.540 10.530 4.960 11.060 ;
        RECT 5.710 10.530 6.130 11.060 ;
        RECT 7.320 10.310 7.490 11.570 ;
        RECT 8.280 10.310 8.450 11.560 ;
        RECT 9.240 10.310 9.410 11.560 ;
        RECT 10.200 10.310 10.370 11.560 ;
        RECT 14.110 10.450 14.280 13.030 ;
        RECT 15.070 10.450 15.240 13.030 ;
        RECT 16.030 10.450 16.200 13.030 ;
        RECT 18.060 12.350 18.400 13.980 ;
        RECT 18.740 13.890 20.520 13.980 ;
        RECT 19.280 13.100 19.450 13.890 ;
        RECT 20.240 13.100 20.410 13.890 ;
        RECT 22.640 13.590 23.070 14.480 ;
        RECT 22.760 12.880 22.930 13.590 ;
        RECT 17.710 12.010 18.400 12.350 ;
        RECT 7.320 10.240 10.370 10.310 ;
        RECT 14.080 10.260 16.340 10.450 ;
        RECT 17.710 10.260 18.110 12.010 ;
        RECT 6.750 10.030 10.840 10.240 ;
        RECT 7.370 8.540 9.670 10.030 ;
        RECT 17.710 9.910 22.570 10.260 ;
        RECT 20.270 8.540 22.570 9.910 ;
        RECT 4.520 8.140 25.420 8.540 ;
        RECT 4.520 1.840 4.920 8.140 ;
        RECT 7.370 8.090 9.670 8.140 ;
        RECT 20.270 8.090 22.570 8.140 ;
        RECT 5.720 6.940 24.220 7.540 ;
        RECT 8.320 6.340 8.670 6.940 ;
        RECT 6.070 6.140 8.670 6.340 ;
        RECT 8.320 5.540 8.670 6.140 ;
        RECT 6.070 5.340 8.670 5.540 ;
        RECT 9.270 5.440 9.470 6.940 ;
        RECT 10.070 5.440 10.270 6.940 ;
        RECT 10.870 5.440 11.070 6.940 ;
        RECT 11.670 5.440 11.870 6.940 ;
        RECT 12.470 5.440 12.670 6.940 ;
        RECT 13.270 5.440 13.470 6.940 ;
        RECT 14.070 5.440 14.270 6.940 ;
        RECT 14.870 5.440 15.070 6.940 ;
        RECT 15.670 5.440 15.870 6.940 ;
        RECT 16.470 5.440 16.670 6.940 ;
        RECT 17.270 5.440 17.470 6.940 ;
        RECT 18.070 5.440 18.270 6.940 ;
        RECT 18.870 5.440 19.070 6.940 ;
        RECT 19.670 5.440 19.870 6.940 ;
        RECT 20.470 5.440 20.670 6.940 ;
        RECT 21.270 6.340 21.620 6.940 ;
        RECT 21.270 6.140 23.870 6.340 ;
        RECT 21.270 5.540 21.620 6.140 ;
        RECT 21.270 5.340 23.820 5.540 ;
        RECT 6.070 4.440 8.670 4.640 ;
        RECT 8.320 3.840 8.670 4.440 ;
        RECT 6.070 3.640 8.670 3.840 ;
        RECT 8.320 3.040 8.670 3.640 ;
        RECT 9.270 3.040 9.470 4.540 ;
        RECT 10.070 3.040 10.270 4.540 ;
        RECT 10.870 3.040 11.070 4.540 ;
        RECT 11.670 3.040 11.870 4.540 ;
        RECT 12.470 3.040 12.670 4.540 ;
        RECT 13.270 3.040 13.470 4.540 ;
        RECT 14.070 3.040 14.270 4.540 ;
        RECT 14.870 3.040 15.070 4.540 ;
        RECT 15.670 3.040 15.870 4.540 ;
        RECT 16.470 3.040 16.670 4.540 ;
        RECT 17.270 3.040 17.470 4.540 ;
        RECT 18.070 3.040 18.270 4.540 ;
        RECT 18.870 3.040 19.070 4.540 ;
        RECT 19.670 3.040 19.870 4.540 ;
        RECT 20.470 3.040 20.670 4.540 ;
        RECT 21.270 4.440 23.820 4.640 ;
        RECT 21.270 3.840 21.620 4.440 ;
        RECT 21.270 3.640 23.870 3.840 ;
        RECT 21.270 3.040 21.620 3.640 ;
        RECT 5.720 2.440 24.220 3.040 ;
        RECT 7.370 1.840 9.670 1.890 ;
        RECT 20.270 1.840 22.570 1.890 ;
        RECT 25.020 1.840 25.420 8.140 ;
        RECT 4.520 1.440 25.420 1.840 ;
        RECT 7.370 0.990 9.670 1.440 ;
        RECT 20.270 0.990 22.570 1.440 ;
        RECT 26.340 0.990 27.330 14.480 ;
        RECT 2.940 0.000 27.330 0.990 ;
      LAYER mcon ;
        RECT 3.120 24.740 3.770 26.740 ;
        RECT 3.040 21.840 3.720 24.040 ;
        RECT 3.040 19.090 3.820 21.240 ;
        RECT 5.820 24.990 6.420 25.490 ;
        RECT 6.620 24.990 7.220 25.490 ;
        RECT 7.420 24.990 8.020 25.490 ;
        RECT 8.220 24.990 8.820 25.490 ;
        RECT 21.120 24.990 21.720 25.490 ;
        RECT 21.920 24.990 22.520 25.490 ;
        RECT 22.720 24.990 23.320 25.490 ;
        RECT 23.520 24.990 24.120 25.490 ;
        RECT 5.820 20.390 6.420 20.890 ;
        RECT 6.620 20.390 7.220 20.890 ;
        RECT 7.420 20.390 8.020 20.890 ;
        RECT 8.220 20.390 8.820 20.890 ;
        RECT 21.120 20.390 21.720 20.890 ;
        RECT 21.920 20.390 22.520 20.890 ;
        RECT 22.720 20.390 23.320 20.890 ;
        RECT 23.520 20.390 24.120 20.890 ;
        RECT 3.020 10.610 3.190 10.780 ;
        RECT 3.380 10.610 3.550 10.780 ;
        RECT 3.740 10.610 3.910 10.780 ;
        RECT 4.660 10.560 4.840 10.730 ;
        RECT 5.830 10.560 6.010 10.730 ;
        RECT 3.020 10.250 3.190 10.420 ;
        RECT 3.380 10.250 3.550 10.420 ;
        RECT 3.740 10.250 3.910 10.420 ;
        RECT 14.200 10.270 14.380 10.450 ;
        RECT 14.660 10.270 14.840 10.450 ;
        RECT 15.120 10.270 15.300 10.450 ;
        RECT 15.580 10.270 15.760 10.450 ;
        RECT 16.040 10.270 16.220 10.450 ;
        RECT 26.410 10.610 26.580 10.780 ;
        RECT 26.770 10.610 26.940 10.780 ;
        RECT 27.130 10.610 27.300 10.780 ;
        RECT 3.020 9.890 3.190 10.060 ;
        RECT 3.380 9.890 3.550 10.060 ;
        RECT 3.740 9.890 3.910 10.060 ;
        RECT 6.870 10.050 7.050 10.230 ;
        RECT 7.460 10.050 7.640 10.230 ;
        RECT 8.050 10.050 8.230 10.230 ;
        RECT 8.640 10.050 8.820 10.230 ;
        RECT 9.230 10.050 9.410 10.230 ;
        RECT 9.820 10.050 10.000 10.230 ;
        RECT 10.410 10.050 10.590 10.230 ;
        RECT 3.020 9.530 3.190 9.700 ;
        RECT 3.380 9.530 3.550 9.700 ;
        RECT 3.740 9.530 3.910 9.700 ;
        RECT 3.010 9.170 3.180 9.340 ;
        RECT 3.370 9.170 3.540 9.340 ;
        RECT 3.730 9.170 3.900 9.340 ;
        RECT 3.030 6.690 3.820 8.840 ;
        RECT 17.750 9.980 17.930 10.160 ;
        RECT 18.120 9.990 18.300 10.170 ;
        RECT 18.520 9.990 18.700 10.170 ;
        RECT 18.920 9.990 19.100 10.170 ;
        RECT 19.320 9.990 19.500 10.170 ;
        RECT 26.410 10.250 26.580 10.420 ;
        RECT 26.770 10.250 26.940 10.420 ;
        RECT 27.130 10.250 27.300 10.420 ;
        RECT 26.410 9.890 26.580 10.060 ;
        RECT 26.770 9.890 26.940 10.060 ;
        RECT 27.130 9.890 27.300 10.060 ;
        RECT 26.410 9.530 26.580 9.700 ;
        RECT 26.770 9.530 26.940 9.700 ;
        RECT 27.130 9.530 27.300 9.700 ;
        RECT 26.410 9.170 26.580 9.340 ;
        RECT 26.770 9.170 26.940 9.340 ;
        RECT 27.130 9.170 27.300 9.340 ;
        RECT 3.070 3.890 3.720 6.090 ;
        RECT 3.070 1.190 3.870 3.240 ;
        RECT 5.820 7.040 6.420 7.540 ;
        RECT 6.620 7.040 7.220 7.540 ;
        RECT 7.420 7.040 8.020 7.540 ;
        RECT 8.220 7.040 8.820 7.540 ;
        RECT 21.120 7.040 21.720 7.540 ;
        RECT 21.920 7.040 22.520 7.540 ;
        RECT 22.720 7.040 23.320 7.540 ;
        RECT 23.520 7.040 24.120 7.540 ;
        RECT 5.820 2.440 6.420 2.940 ;
        RECT 6.620 2.440 7.220 2.940 ;
        RECT 7.420 2.440 8.020 2.940 ;
        RECT 8.220 2.440 8.820 2.940 ;
        RECT 21.120 2.440 21.720 2.940 ;
        RECT 21.920 2.440 22.520 2.940 ;
        RECT 22.720 2.440 23.320 2.940 ;
        RECT 23.520 2.440 24.120 2.940 ;
      LAYER met1 ;
        RECT 2.940 25.690 7.320 26.890 ;
        RECT 22.620 25.690 25.820 26.890 ;
        RECT 2.940 25.540 6.420 25.690 ;
        RECT 23.520 25.540 25.820 25.690 ;
        RECT 2.940 25.390 14.520 25.540 ;
        RECT 15.420 25.390 25.820 25.540 ;
        RECT 2.940 24.940 8.920 25.390 ;
        RECT 21.020 24.940 25.820 25.390 ;
        RECT 2.940 24.540 5.320 24.940 ;
        RECT 5.770 24.890 14.520 24.940 ;
        RECT 2.940 21.740 3.820 24.140 ;
        RECT 4.120 24.040 5.320 24.540 ;
        RECT 5.920 23.540 6.070 24.890 ;
        RECT 6.520 23.540 6.670 24.890 ;
        RECT 7.120 23.540 7.270 24.890 ;
        RECT 7.720 23.540 7.870 24.890 ;
        RECT 8.320 24.790 14.520 24.890 ;
        RECT 15.420 24.890 24.170 24.940 ;
        RECT 15.420 24.790 21.620 24.890 ;
        RECT 8.320 24.340 8.920 24.790 ;
        RECT 21.020 24.340 21.620 24.790 ;
        RECT 8.320 24.190 14.520 24.340 ;
        RECT 15.420 24.190 21.620 24.340 ;
        RECT 8.320 23.740 8.920 24.190 ;
        RECT 21.020 23.740 21.620 24.190 ;
        RECT 8.320 23.590 14.520 23.740 ;
        RECT 15.420 23.590 21.620 23.740 ;
        RECT 8.320 23.390 8.920 23.590 ;
        RECT 21.020 23.390 21.620 23.590 ;
        RECT 22.070 23.540 22.220 24.890 ;
        RECT 22.670 23.540 22.820 24.890 ;
        RECT 23.270 23.540 23.420 24.890 ;
        RECT 23.870 23.540 24.020 24.890 ;
        RECT 24.620 24.040 25.820 24.940 ;
        RECT 4.120 21.340 5.320 21.840 ;
        RECT 2.940 20.940 5.320 21.340 ;
        RECT 5.920 20.990 6.070 22.290 ;
        RECT 6.520 20.990 6.670 22.290 ;
        RECT 7.120 20.990 7.270 22.290 ;
        RECT 7.720 20.990 7.870 22.290 ;
        RECT 8.320 22.140 14.520 22.290 ;
        RECT 15.420 22.140 21.620 22.290 ;
        RECT 8.320 21.690 8.920 22.140 ;
        RECT 21.020 21.690 21.620 22.140 ;
        RECT 8.320 21.540 14.520 21.690 ;
        RECT 15.420 21.540 21.620 21.690 ;
        RECT 8.320 21.090 8.920 21.540 ;
        RECT 21.020 21.090 21.620 21.540 ;
        RECT 8.320 20.990 14.520 21.090 ;
        RECT 5.770 20.940 14.520 20.990 ;
        RECT 15.420 20.990 21.620 21.090 ;
        RECT 22.070 20.990 22.220 22.290 ;
        RECT 22.670 20.990 22.820 22.290 ;
        RECT 23.270 20.990 23.420 22.290 ;
        RECT 23.870 20.990 24.020 22.290 ;
        RECT 15.420 20.940 24.170 20.990 ;
        RECT 24.620 20.940 25.820 21.840 ;
        RECT 2.940 20.490 8.920 20.940 ;
        RECT 21.020 20.490 25.820 20.940 ;
        RECT 2.940 20.340 14.520 20.490 ;
        RECT 15.420 20.340 25.820 20.490 ;
        RECT 2.940 20.190 6.420 20.340 ;
        RECT 23.520 20.190 25.820 20.340 ;
        RECT 2.940 18.990 7.320 20.190 ;
        RECT 22.620 18.990 25.820 20.190 ;
        RECT 2.940 10.780 3.940 10.880 ;
        RECT 2.940 10.260 6.210 10.780 ;
        RECT 14.080 10.260 16.340 10.480 ;
        RECT 26.340 10.260 27.330 10.880 ;
        RECT 0.000 9.100 28.570 10.260 ;
        RECT 2.930 7.740 7.320 8.940 ;
        RECT 22.620 7.740 25.820 8.940 ;
        RECT 2.930 7.590 6.420 7.740 ;
        RECT 23.520 7.590 25.820 7.740 ;
        RECT 2.930 7.440 14.520 7.590 ;
        RECT 15.420 7.440 25.820 7.590 ;
        RECT 2.930 6.990 8.920 7.440 ;
        RECT 21.020 6.990 25.820 7.440 ;
        RECT 2.930 6.590 5.320 6.990 ;
        RECT 5.770 6.940 14.520 6.990 ;
        RECT 2.940 3.790 3.820 6.190 ;
        RECT 4.120 6.090 5.320 6.590 ;
        RECT 5.920 5.590 6.070 6.940 ;
        RECT 6.520 5.590 6.670 6.940 ;
        RECT 7.120 5.590 7.270 6.940 ;
        RECT 7.720 5.590 7.870 6.940 ;
        RECT 8.320 6.840 14.520 6.940 ;
        RECT 15.420 6.940 24.170 6.990 ;
        RECT 15.420 6.840 21.620 6.940 ;
        RECT 8.320 6.390 8.920 6.840 ;
        RECT 21.020 6.390 21.620 6.840 ;
        RECT 8.320 6.240 14.520 6.390 ;
        RECT 15.420 6.240 21.620 6.390 ;
        RECT 8.320 5.790 8.920 6.240 ;
        RECT 21.020 5.790 21.620 6.240 ;
        RECT 8.320 5.640 14.520 5.790 ;
        RECT 15.420 5.640 21.620 5.790 ;
        RECT 8.320 5.440 8.920 5.640 ;
        RECT 21.020 5.440 21.620 5.640 ;
        RECT 22.070 5.590 22.220 6.940 ;
        RECT 22.670 5.590 22.820 6.940 ;
        RECT 23.270 5.590 23.420 6.940 ;
        RECT 23.870 5.590 24.020 6.940 ;
        RECT 24.620 6.090 25.820 6.990 ;
        RECT 4.120 3.390 5.320 3.890 ;
        RECT 2.940 2.990 5.320 3.390 ;
        RECT 5.920 3.040 6.070 4.340 ;
        RECT 6.520 3.040 6.670 4.340 ;
        RECT 7.120 3.040 7.270 4.340 ;
        RECT 7.720 3.040 7.870 4.340 ;
        RECT 8.320 4.190 14.520 4.340 ;
        RECT 15.420 4.190 21.620 4.340 ;
        RECT 8.320 3.740 8.920 4.190 ;
        RECT 21.020 3.740 21.620 4.190 ;
        RECT 8.320 3.590 14.520 3.740 ;
        RECT 15.420 3.590 21.620 3.740 ;
        RECT 8.320 3.140 8.920 3.590 ;
        RECT 21.020 3.140 21.620 3.590 ;
        RECT 8.320 3.040 14.520 3.140 ;
        RECT 5.770 2.990 14.520 3.040 ;
        RECT 15.420 3.040 21.620 3.140 ;
        RECT 22.070 3.040 22.220 4.340 ;
        RECT 22.670 3.040 22.820 4.340 ;
        RECT 23.270 3.040 23.420 4.340 ;
        RECT 23.870 3.040 24.020 4.340 ;
        RECT 15.420 2.990 24.170 3.040 ;
        RECT 24.620 2.990 25.820 3.890 ;
        RECT 2.940 2.540 8.920 2.990 ;
        RECT 21.020 2.540 25.820 2.990 ;
        RECT 2.940 2.390 14.520 2.540 ;
        RECT 15.420 2.390 25.820 2.540 ;
        RECT 2.940 2.240 6.420 2.390 ;
        RECT 23.520 2.240 25.820 2.390 ;
        RECT 2.940 1.040 7.320 2.240 ;
        RECT 22.620 1.040 25.820 2.240 ;
      LAYER via ;
        RECT 3.120 24.740 3.770 26.740 ;
        RECT 4.220 25.790 5.220 26.790 ;
        RECT 6.220 25.790 7.220 26.790 ;
        RECT 22.720 25.790 23.720 26.790 ;
        RECT 24.720 25.790 25.720 26.790 ;
        RECT 4.220 24.190 5.220 25.190 ;
        RECT 3.040 21.840 3.720 24.040 ;
        RECT 24.720 24.190 25.720 25.190 ;
        RECT 4.220 20.690 5.220 21.690 ;
        RECT 24.720 20.690 25.720 21.690 ;
        RECT 4.220 19.090 5.220 20.090 ;
        RECT 6.220 19.090 7.220 20.090 ;
        RECT 22.720 19.090 23.720 20.090 ;
        RECT 24.720 19.090 25.720 20.090 ;
        RECT 1.720 9.190 2.520 10.140 ;
        RECT 4.220 9.290 7.000 10.120 ;
        RECT 27.670 9.190 28.470 10.140 ;
        RECT 4.220 7.840 5.220 8.840 ;
        RECT 6.220 7.840 7.220 8.840 ;
        RECT 22.720 7.840 23.720 8.840 ;
        RECT 24.720 7.840 25.720 8.840 ;
        RECT 4.220 6.240 5.220 7.240 ;
        RECT 3.070 3.890 3.720 6.090 ;
        RECT 24.720 6.240 25.720 7.240 ;
        RECT 3.070 1.190 3.730 3.240 ;
        RECT 4.220 2.740 5.220 3.740 ;
        RECT 24.720 2.740 25.720 3.740 ;
        RECT 4.220 1.140 5.220 2.140 ;
        RECT 6.220 1.140 7.220 2.140 ;
        RECT 22.720 1.140 23.720 2.140 ;
        RECT 24.720 1.140 25.720 2.140 ;
      LAYER met2 ;
        RECT 2.940 25.690 7.320 26.890 ;
        RECT 22.620 25.690 25.820 26.890 ;
        RECT 2.940 24.740 6.070 25.690 ;
        RECT 23.870 24.740 25.820 25.690 ;
        RECT 2.940 24.590 8.070 24.740 ;
        RECT 2.940 24.540 6.070 24.590 ;
        RECT 4.120 24.140 6.070 24.540 ;
        RECT 2.940 21.740 3.820 24.140 ;
        RECT 4.120 24.040 8.070 24.140 ;
        RECT 5.520 23.990 8.070 24.040 ;
        RECT 5.520 23.390 6.070 23.990 ;
        RECT 5.520 23.090 8.070 23.390 ;
        RECT 8.670 23.090 8.820 24.740 ;
        RECT 9.270 23.090 9.420 24.740 ;
        RECT 9.870 23.090 10.020 24.740 ;
        RECT 10.470 23.090 10.620 24.740 ;
        RECT 11.070 23.090 11.220 24.740 ;
        RECT 11.670 23.090 11.820 24.740 ;
        RECT 12.270 23.090 12.420 24.740 ;
        RECT 12.870 23.090 13.020 24.740 ;
        RECT 13.470 23.090 13.620 24.740 ;
        RECT 14.070 23.090 14.220 24.740 ;
        RECT 14.670 23.090 15.270 24.740 ;
        RECT 15.720 23.090 15.870 24.740 ;
        RECT 16.320 23.090 16.470 24.740 ;
        RECT 16.920 23.090 17.070 24.740 ;
        RECT 17.520 23.090 17.670 24.740 ;
        RECT 18.120 23.090 18.270 24.740 ;
        RECT 18.720 23.090 18.870 24.740 ;
        RECT 19.320 23.090 19.470 24.740 ;
        RECT 19.920 23.090 20.070 24.740 ;
        RECT 20.520 23.090 20.670 24.740 ;
        RECT 21.120 23.090 21.270 24.740 ;
        RECT 21.870 24.590 25.820 24.740 ;
        RECT 23.870 24.140 25.820 24.590 ;
        RECT 21.870 24.040 25.820 24.140 ;
        RECT 21.870 23.990 24.420 24.040 ;
        RECT 23.870 23.390 24.420 23.990 ;
        RECT 21.870 23.090 24.420 23.390 ;
        RECT 5.520 22.790 24.420 23.090 ;
        RECT 5.520 22.340 8.070 22.790 ;
        RECT 5.520 21.890 6.070 22.340 ;
        RECT 5.520 21.840 8.070 21.890 ;
        RECT 4.120 21.740 8.070 21.840 ;
        RECT 4.120 21.290 6.070 21.740 ;
        RECT 4.120 21.140 8.070 21.290 ;
        RECT 8.670 21.140 8.820 22.790 ;
        RECT 9.270 21.140 9.420 22.790 ;
        RECT 9.870 21.140 10.020 22.790 ;
        RECT 10.470 21.140 10.620 22.790 ;
        RECT 11.070 21.140 11.220 22.790 ;
        RECT 11.670 21.140 11.820 22.790 ;
        RECT 12.270 21.140 12.420 22.790 ;
        RECT 12.870 21.140 13.020 22.790 ;
        RECT 13.470 21.140 13.620 22.790 ;
        RECT 14.070 21.140 14.220 22.790 ;
        RECT 14.670 21.140 15.270 22.790 ;
        RECT 15.720 21.140 15.870 22.790 ;
        RECT 16.320 21.140 16.470 22.790 ;
        RECT 16.920 21.140 17.070 22.790 ;
        RECT 17.520 21.140 17.670 22.790 ;
        RECT 18.120 21.140 18.270 22.790 ;
        RECT 18.720 21.140 18.870 22.790 ;
        RECT 19.320 21.140 19.470 22.790 ;
        RECT 19.920 21.140 20.070 22.790 ;
        RECT 20.520 21.140 20.670 22.790 ;
        RECT 21.120 21.140 21.270 22.790 ;
        RECT 21.870 22.340 24.420 22.790 ;
        RECT 23.870 21.890 24.420 22.340 ;
        RECT 21.870 21.840 24.420 21.890 ;
        RECT 21.870 21.740 25.820 21.840 ;
        RECT 23.870 21.290 25.820 21.740 ;
        RECT 21.870 21.140 25.820 21.290 ;
        RECT 4.120 20.190 6.070 21.140 ;
        RECT 23.870 20.190 25.820 21.140 ;
        RECT 4.120 18.990 7.320 20.190 ;
        RECT 22.620 18.990 25.820 20.190 ;
        RECT 1.610 9.100 2.610 10.260 ;
        RECT 4.080 9.260 7.230 10.260 ;
        RECT 4.120 8.940 7.270 9.260 ;
        RECT 27.570 9.100 28.570 10.260 ;
        RECT 4.120 7.740 7.320 8.940 ;
        RECT 22.620 7.740 25.820 8.940 ;
        RECT 4.120 6.790 6.070 7.740 ;
        RECT 23.870 6.790 25.820 7.740 ;
        RECT 4.120 6.640 8.070 6.790 ;
        RECT 4.120 6.190 6.070 6.640 ;
        RECT 2.940 3.790 3.820 6.190 ;
        RECT 4.120 6.090 8.070 6.190 ;
        RECT 5.520 6.040 8.070 6.090 ;
        RECT 5.520 5.440 6.070 6.040 ;
        RECT 5.520 5.140 8.070 5.440 ;
        RECT 8.670 5.140 8.820 6.790 ;
        RECT 9.270 5.140 9.420 6.790 ;
        RECT 9.870 5.140 10.020 6.790 ;
        RECT 10.470 5.140 10.620 6.790 ;
        RECT 11.070 5.140 11.220 6.790 ;
        RECT 11.670 5.140 11.820 6.790 ;
        RECT 12.270 5.140 12.420 6.790 ;
        RECT 12.870 5.140 13.020 6.790 ;
        RECT 13.470 5.140 13.620 6.790 ;
        RECT 14.070 5.140 14.220 6.790 ;
        RECT 14.670 5.140 15.270 6.790 ;
        RECT 15.720 5.140 15.870 6.790 ;
        RECT 16.320 5.140 16.470 6.790 ;
        RECT 16.920 5.140 17.070 6.790 ;
        RECT 17.520 5.140 17.670 6.790 ;
        RECT 18.120 5.140 18.270 6.790 ;
        RECT 18.720 5.140 18.870 6.790 ;
        RECT 19.320 5.140 19.470 6.790 ;
        RECT 19.920 5.140 20.070 6.790 ;
        RECT 20.520 5.140 20.670 6.790 ;
        RECT 21.120 5.140 21.270 6.790 ;
        RECT 21.870 6.640 25.820 6.790 ;
        RECT 23.870 6.190 25.820 6.640 ;
        RECT 21.870 6.090 25.820 6.190 ;
        RECT 21.870 6.040 24.420 6.090 ;
        RECT 23.870 5.440 24.420 6.040 ;
        RECT 21.870 5.140 24.420 5.440 ;
        RECT 5.520 4.840 24.420 5.140 ;
        RECT 5.520 4.390 8.070 4.840 ;
        RECT 5.520 3.940 6.070 4.390 ;
        RECT 5.520 3.890 8.070 3.940 ;
        RECT 4.120 3.790 8.070 3.890 ;
        RECT 4.120 3.390 6.070 3.790 ;
        RECT 2.940 3.340 6.070 3.390 ;
        RECT 2.940 3.190 8.070 3.340 ;
        RECT 8.670 3.190 8.820 4.840 ;
        RECT 9.270 3.190 9.420 4.840 ;
        RECT 9.870 3.190 10.020 4.840 ;
        RECT 10.470 3.190 10.620 4.840 ;
        RECT 11.070 3.190 11.220 4.840 ;
        RECT 11.670 3.190 11.820 4.840 ;
        RECT 12.270 3.190 12.420 4.840 ;
        RECT 12.870 3.190 13.020 4.840 ;
        RECT 13.470 3.190 13.620 4.840 ;
        RECT 14.070 3.190 14.220 4.840 ;
        RECT 14.670 3.190 15.270 4.840 ;
        RECT 15.720 3.190 15.870 4.840 ;
        RECT 16.320 3.190 16.470 4.840 ;
        RECT 16.920 3.190 17.070 4.840 ;
        RECT 17.520 3.190 17.670 4.840 ;
        RECT 18.120 3.190 18.270 4.840 ;
        RECT 18.720 3.190 18.870 4.840 ;
        RECT 19.320 3.190 19.470 4.840 ;
        RECT 19.920 3.190 20.070 4.840 ;
        RECT 20.520 3.190 20.670 4.840 ;
        RECT 21.120 3.190 21.270 4.840 ;
        RECT 21.870 4.390 24.420 4.840 ;
        RECT 23.870 3.940 24.420 4.390 ;
        RECT 21.870 3.890 24.420 3.940 ;
        RECT 21.870 3.790 25.820 3.890 ;
        RECT 23.870 3.340 25.820 3.790 ;
        RECT 21.870 3.190 25.820 3.340 ;
        RECT 2.940 2.240 6.070 3.190 ;
        RECT 23.870 2.240 25.820 3.190 ;
        RECT 2.940 1.040 7.320 2.240 ;
        RECT 22.620 1.040 25.820 2.240 ;
      LAYER via2 ;
        RECT 3.120 24.740 3.770 26.740 ;
        RECT 3.040 21.840 3.720 24.040 ;
        RECT 1.720 9.190 2.520 10.140 ;
        RECT 4.220 9.290 7.000 10.120 ;
        RECT 27.670 9.190 28.470 10.140 ;
        RECT 3.070 3.890 3.720 6.090 ;
        RECT 3.070 1.190 3.730 3.240 ;
      LAYER met3 ;
        RECT 2.940 24.540 3.810 26.890 ;
        RECT 4.120 25.640 7.320 26.890 ;
        RECT 9.720 26.040 20.220 26.890 ;
        RECT 22.620 25.640 25.820 26.890 ;
        RECT 4.120 24.490 25.820 25.640 ;
        RECT 2.940 21.740 3.820 24.140 ;
        RECT 4.120 21.740 4.970 24.140 ;
        RECT 5.370 21.390 24.570 24.490 ;
        RECT 24.970 21.740 25.820 24.140 ;
        RECT 4.120 20.240 25.820 21.390 ;
        RECT 4.120 18.990 7.320 20.240 ;
        RECT 9.720 18.990 20.220 19.840 ;
        RECT 22.620 18.990 25.820 20.240 ;
        RECT 1.610 9.100 2.610 10.260 ;
        RECT 4.080 9.260 7.230 10.260 ;
        RECT 27.570 9.100 28.570 10.260 ;
        RECT 4.120 7.690 7.320 8.940 ;
        RECT 9.720 8.090 20.220 8.940 ;
        RECT 22.620 7.690 25.820 8.940 ;
        RECT 4.120 6.540 25.820 7.690 ;
        RECT 2.940 3.790 3.820 6.190 ;
        RECT 4.120 3.790 4.970 6.190 ;
        RECT 5.370 3.440 24.570 6.540 ;
        RECT 24.970 3.790 25.820 6.190 ;
        RECT 2.940 1.040 3.800 3.390 ;
        RECT 4.120 2.290 25.820 3.440 ;
        RECT 4.120 1.040 7.320 2.290 ;
        RECT 9.720 1.040 20.220 1.890 ;
        RECT 22.620 1.040 25.820 2.290 ;
      LAYER via3 ;
        RECT 3.120 24.740 3.770 26.740 ;
        RECT 4.220 25.940 5.070 26.790 ;
        RECT 6.320 25.940 7.170 26.790 ;
        RECT 9.820 26.140 10.470 26.790 ;
        RECT 10.620 26.140 11.270 26.790 ;
        RECT 18.670 26.140 19.320 26.790 ;
        RECT 19.470 26.140 20.120 26.790 ;
        RECT 22.770 25.940 23.620 26.790 ;
        RECT 24.870 25.940 25.720 26.790 ;
        RECT 4.220 24.640 5.070 25.490 ;
        RECT 24.870 24.640 25.720 25.490 ;
        RECT 3.040 21.840 3.720 24.040 ;
        RECT 4.220 23.040 4.870 24.040 ;
        RECT 4.220 21.840 4.870 22.840 ;
        RECT 25.070 23.040 25.720 24.040 ;
        RECT 25.070 21.840 25.720 22.840 ;
        RECT 4.220 20.390 5.070 21.240 ;
        RECT 24.870 20.390 25.720 21.240 ;
        RECT 4.220 19.090 5.070 19.940 ;
        RECT 6.320 19.090 7.170 19.940 ;
        RECT 9.820 19.090 10.470 19.740 ;
        RECT 10.620 19.090 11.270 19.740 ;
        RECT 18.670 19.090 19.320 19.740 ;
        RECT 19.470 19.090 20.120 19.740 ;
        RECT 22.770 19.090 23.620 19.940 ;
        RECT 24.870 19.090 25.720 19.940 ;
        RECT 1.720 9.190 2.520 10.140 ;
        RECT 27.670 9.190 28.470 10.140 ;
        RECT 4.220 7.990 5.070 8.840 ;
        RECT 6.320 7.990 7.170 8.840 ;
        RECT 9.820 8.190 10.470 8.840 ;
        RECT 10.620 8.190 11.270 8.840 ;
        RECT 18.670 8.190 19.320 8.840 ;
        RECT 19.470 8.190 20.120 8.840 ;
        RECT 22.770 7.990 23.620 8.840 ;
        RECT 24.870 7.990 25.720 8.840 ;
        RECT 4.220 6.690 5.070 7.540 ;
        RECT 24.870 6.690 25.720 7.540 ;
        RECT 3.070 3.890 3.720 6.090 ;
        RECT 4.220 5.090 4.870 6.090 ;
        RECT 4.220 3.890 4.870 4.890 ;
        RECT 25.070 5.090 25.720 6.090 ;
        RECT 25.070 3.890 25.720 4.890 ;
        RECT 3.070 1.190 3.730 3.240 ;
        RECT 4.220 2.440 5.070 3.290 ;
        RECT 24.870 2.440 25.720 3.290 ;
        RECT 4.220 1.140 5.070 1.990 ;
        RECT 6.320 1.140 7.170 1.990 ;
        RECT 9.820 1.140 10.470 1.790 ;
        RECT 10.620 1.140 11.270 1.790 ;
        RECT 18.670 1.140 19.320 1.790 ;
        RECT 19.470 1.140 20.120 1.790 ;
        RECT 22.770 1.140 23.620 1.990 ;
        RECT 24.870 1.140 25.720 1.990 ;
      LAYER met4 ;
        RECT 1.610 0.000 2.610 27.980 ;
        RECT 2.940 25.840 7.270 26.890 ;
        RECT 2.940 24.540 5.170 25.840 ;
        RECT 9.720 25.440 20.220 26.890 ;
        RECT 22.670 25.840 25.820 26.890 ;
        RECT 5.570 24.140 24.370 25.440 ;
        RECT 24.770 24.540 25.820 25.840 ;
        RECT 2.940 21.740 25.820 24.140 ;
        RECT 4.120 20.040 5.170 21.340 ;
        RECT 5.570 20.440 24.370 21.740 ;
        RECT 4.120 18.990 7.270 20.040 ;
        RECT 9.720 18.990 20.220 20.440 ;
        RECT 24.770 20.040 25.820 21.340 ;
        RECT 22.670 18.990 25.820 20.040 ;
        RECT 4.120 7.890 7.270 8.940 ;
        RECT 4.120 6.590 5.170 7.890 ;
        RECT 9.720 7.490 20.220 8.940 ;
        RECT 22.670 7.890 25.820 8.940 ;
        RECT 5.570 6.190 24.370 7.490 ;
        RECT 24.770 6.590 25.820 7.890 ;
        RECT 2.940 3.790 25.820 6.190 ;
        RECT 2.940 2.090 5.170 3.390 ;
        RECT 5.570 2.490 24.370 3.790 ;
        RECT 2.940 1.040 7.270 2.090 ;
        RECT 9.720 1.040 20.220 2.490 ;
        RECT 24.770 2.090 25.820 3.390 ;
        RECT 22.670 1.040 25.820 2.090 ;
        RECT 27.570 0.000 28.570 27.980 ;
    END
  END VSS
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.189000 ;
    PORT
      LAYER li1 ;
        RECT 4.100 11.790 4.370 12.120 ;
      LAYER mcon ;
        RECT 4.180 11.870 4.350 12.040 ;
      LAYER met1 ;
        RECT 4.070 12.030 4.380 12.120 ;
        RECT 0.000 11.890 4.380 12.030 ;
        RECT 4.070 11.790 4.380 11.890 ;
    END
  END clk
  PIN inp
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.200000 ;
    PORT
      LAYER li1 ;
        RECT 9.630 15.220 9.990 15.520 ;
      LAYER mcon ;
        RECT 9.710 15.270 9.910 15.470 ;
      LAYER met1 ;
        RECT 0.000 15.410 9.990 15.550 ;
        RECT 9.630 15.220 9.990 15.410 ;
    END
  END inp
  PIN inn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.200000 ;
    PORT
      LAYER li1 ;
        RECT 7.670 14.970 8.030 15.270 ;
      LAYER mcon ;
        RECT 7.750 15.020 7.950 15.220 ;
      LAYER met1 ;
        RECT 0.000 15.130 8.030 15.270 ;
        RECT 7.670 14.970 8.030 15.130 ;
    END
  END inn
  PIN comp_trig
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.756400 ;
    PORT
      LAYER li1 ;
        RECT 22.280 11.230 22.450 13.340 ;
        RECT 23.240 12.880 23.510 13.340 ;
        RECT 23.340 12.780 23.510 12.880 ;
        RECT 23.340 12.590 25.370 12.780 ;
        RECT 24.200 11.230 24.370 12.590 ;
        RECT 24.690 12.540 25.370 12.590 ;
      LAYER mcon ;
        RECT 22.280 12.960 22.450 13.260 ;
        RECT 23.240 12.960 23.410 13.260 ;
        RECT 24.750 12.570 24.930 12.750 ;
        RECT 25.130 12.570 25.310 12.750 ;
      LAYER met1 ;
        RECT 22.250 13.180 22.480 13.320 ;
        RECT 23.210 13.180 23.440 13.320 ;
        RECT 22.250 13.040 23.440 13.180 ;
        RECT 22.250 12.900 22.480 13.040 ;
        RECT 23.210 12.900 23.440 13.040 ;
        RECT 24.690 12.730 25.370 12.780 ;
        RECT 24.690 12.590 30.050 12.730 ;
        RECT 24.690 12.540 25.370 12.590 ;
    END
  END comp_trig
  PIN latch_qn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.303000 ;
    ANTENNADIFFAREA 0.756400 ;
    PORT
      LAYER li1 ;
        RECT 22.060 15.810 22.390 16.070 ;
        RECT 23.960 14.980 24.130 17.090 ;
        RECT 25.880 15.730 26.050 17.090 ;
        RECT 25.020 15.540 26.170 15.730 ;
        RECT 25.020 15.440 25.190 15.540 ;
        RECT 25.500 15.490 26.170 15.540 ;
        RECT 24.920 14.980 25.190 15.440 ;
      LAYER mcon ;
        RECT 22.140 15.860 22.310 16.030 ;
        RECT 25.560 15.520 25.740 15.700 ;
        RECT 25.930 15.520 26.110 15.700 ;
        RECT 23.960 15.060 24.130 15.360 ;
        RECT 24.920 15.060 25.090 15.360 ;
      LAYER met1 ;
        RECT 22.060 16.050 22.390 16.070 ;
        RECT 21.400 15.870 23.190 16.050 ;
        RECT 22.060 15.810 22.390 15.870 ;
        RECT 23.010 15.310 23.190 15.870 ;
        RECT 25.500 15.680 26.170 15.730 ;
        RECT 25.500 15.540 30.050 15.680 ;
        RECT 25.500 15.490 26.170 15.540 ;
        RECT 23.930 15.310 24.160 15.420 ;
        RECT 23.010 15.280 24.160 15.310 ;
        RECT 24.890 15.280 25.120 15.420 ;
        RECT 23.010 15.140 25.120 15.280 ;
        RECT 23.010 15.130 24.160 15.140 ;
        RECT 23.930 15.000 24.160 15.130 ;
        RECT 24.890 15.000 25.120 15.140 ;
    END
  END latch_qn
  PIN latch_q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.303000 ;
    ANTENNADIFFAREA 0.756400 ;
    PORT
      LAYER li1 ;
        RECT 21.480 14.980 21.650 17.090 ;
        RECT 23.400 15.780 23.570 17.090 ;
        RECT 24.540 15.810 24.870 16.070 ;
        RECT 23.400 15.730 23.640 15.780 ;
        RECT 22.540 15.540 23.640 15.730 ;
        RECT 22.540 15.440 22.710 15.540 ;
        RECT 22.440 14.980 22.710 15.440 ;
      LAYER mcon ;
        RECT 24.620 15.860 24.790 16.030 ;
        RECT 23.440 15.580 23.610 15.750 ;
        RECT 21.480 15.060 21.650 15.360 ;
        RECT 22.440 15.060 22.610 15.360 ;
      LAYER met1 ;
        RECT 24.540 16.060 24.870 16.070 ;
        RECT 24.480 16.050 26.070 16.060 ;
        RECT 23.460 16.020 26.070 16.050 ;
        RECT 23.460 15.880 30.050 16.020 ;
        RECT 23.460 15.870 24.870 15.880 ;
        RECT 23.460 15.810 23.640 15.870 ;
        RECT 24.540 15.810 24.870 15.870 ;
        RECT 23.400 15.520 23.640 15.810 ;
        RECT 21.450 15.280 21.680 15.420 ;
        RECT 22.410 15.280 22.640 15.420 ;
        RECT 21.450 15.140 22.640 15.280 ;
        RECT 21.450 15.000 21.680 15.140 ;
        RECT 22.410 15.000 22.640 15.140 ;
    END
  END latch_q
  OBS
      LAYER li1 ;
        RECT 5.320 24.490 8.120 24.690 ;
        RECT 5.320 23.890 5.870 24.490 ;
        RECT 5.320 23.690 8.120 23.890 ;
        RECT 5.320 23.090 5.870 23.690 ;
        RECT 8.870 23.140 9.070 24.690 ;
        RECT 9.670 23.140 9.870 24.690 ;
        RECT 10.470 23.140 10.670 24.690 ;
        RECT 11.270 23.140 11.470 24.690 ;
        RECT 12.070 23.140 12.270 24.690 ;
        RECT 12.870 23.140 13.070 24.690 ;
        RECT 13.670 23.140 13.870 24.690 ;
        RECT 14.470 23.140 14.670 24.690 ;
        RECT 15.270 23.140 15.470 24.690 ;
        RECT 16.070 23.140 16.270 24.690 ;
        RECT 16.870 23.140 17.070 24.690 ;
        RECT 17.670 23.140 17.870 24.690 ;
        RECT 18.470 23.140 18.670 24.690 ;
        RECT 19.270 23.140 19.470 24.690 ;
        RECT 20.070 23.140 20.270 24.690 ;
        RECT 20.870 23.140 21.070 24.690 ;
        RECT 21.820 24.490 24.620 24.690 ;
        RECT 24.070 23.890 24.620 24.490 ;
        RECT 21.820 23.690 24.620 23.890 ;
        RECT 8.870 23.090 21.070 23.140 ;
        RECT 24.070 23.090 24.620 23.690 ;
        RECT 5.320 22.790 24.620 23.090 ;
        RECT 5.320 22.190 5.870 22.790 ;
        RECT 8.870 22.740 21.070 22.790 ;
        RECT 5.320 21.990 8.120 22.190 ;
        RECT 5.320 21.390 5.870 21.990 ;
        RECT 5.320 21.190 8.120 21.390 ;
        RECT 8.870 21.190 9.070 22.740 ;
        RECT 9.670 21.190 9.870 22.740 ;
        RECT 10.470 21.190 10.670 22.740 ;
        RECT 11.270 21.190 11.470 22.740 ;
        RECT 12.070 21.190 12.270 22.740 ;
        RECT 12.870 21.190 13.070 22.740 ;
        RECT 13.670 21.190 13.870 22.740 ;
        RECT 14.470 21.240 14.670 22.740 ;
        RECT 15.270 21.240 15.470 22.740 ;
        RECT 16.070 21.190 16.270 22.740 ;
        RECT 16.870 21.190 17.070 22.740 ;
        RECT 17.670 21.190 17.870 22.740 ;
        RECT 18.470 21.190 18.670 22.740 ;
        RECT 19.270 21.190 19.470 22.740 ;
        RECT 20.070 21.190 20.270 22.740 ;
        RECT 20.870 21.190 21.070 22.740 ;
        RECT 24.070 22.190 24.620 22.790 ;
        RECT 21.820 21.990 24.620 22.190 ;
        RECT 24.070 21.390 24.620 21.990 ;
        RECT 21.820 21.190 24.620 21.390 ;
        RECT 7.320 16.090 7.490 16.930 ;
        RECT 8.280 16.090 8.450 16.930 ;
        RECT 7.320 15.920 8.450 16.090 ;
        RECT 9.240 16.090 9.410 16.930 ;
        RECT 10.200 16.090 10.370 16.930 ;
        RECT 11.320 16.290 12.270 17.240 ;
        RECT 12.500 16.850 13.630 17.020 ;
        RECT 9.240 15.920 10.370 16.090 ;
        RECT 6.300 15.620 6.630 15.910 ;
        RECT 4.540 13.400 4.960 13.430 ;
        RECT 5.710 13.400 6.130 13.430 ;
        RECT 4.520 13.210 4.980 13.400 ;
        RECT 5.690 13.210 6.150 13.400 ;
        RECT 4.520 12.310 4.980 12.480 ;
        RECT 5.690 12.310 6.150 12.480 ;
        RECT 4.540 12.070 4.960 12.310 ;
        RECT 5.270 12.070 5.540 12.120 ;
        RECT 4.540 11.840 5.540 12.070 ;
        RECT 4.540 11.670 4.960 11.840 ;
        RECT 5.270 11.790 5.540 11.840 ;
        RECT 5.710 12.070 6.130 12.310 ;
        RECT 6.400 12.070 6.630 15.620 ;
        RECT 7.320 14.800 7.490 15.920 ;
        RECT 8.210 14.800 8.450 15.100 ;
        RECT 7.320 14.630 8.450 14.800 ;
        RECT 5.710 11.920 6.630 12.070 ;
        RECT 6.840 12.150 7.010 14.360 ;
        RECT 7.320 12.320 7.490 14.630 ;
        RECT 7.800 12.150 7.970 14.360 ;
        RECT 8.280 12.320 8.450 14.630 ;
        RECT 9.240 14.810 9.410 15.920 ;
        RECT 9.240 14.640 11.620 14.810 ;
        RECT 8.760 12.150 8.930 14.360 ;
        RECT 9.240 12.320 9.410 14.640 ;
        RECT 9.720 12.150 9.890 14.360 ;
        RECT 10.200 12.320 10.370 14.640 ;
        RECT 10.680 12.150 10.850 14.360 ;
        RECT 11.240 14.190 11.620 14.640 ;
        RECT 11.850 14.360 12.230 16.290 ;
        RECT 11.240 13.130 12.230 14.190 ;
        RECT 12.500 14.050 12.670 16.850 ;
        RECT 12.980 14.390 13.150 16.680 ;
        RECT 13.460 14.640 13.630 16.850 ;
        RECT 16.680 16.850 17.810 17.020 ;
        RECT 14.590 14.390 14.760 16.680 ;
        RECT 12.980 14.220 14.760 14.390 ;
        RECT 15.550 14.390 15.720 16.680 ;
        RECT 16.680 14.640 16.850 16.850 ;
        RECT 17.160 14.390 17.330 16.680 ;
        RECT 15.550 14.220 17.330 14.390 ;
        RECT 17.640 15.950 17.810 16.850 ;
        RECT 17.640 15.260 18.630 15.950 ;
        RECT 18.800 15.900 18.970 17.330 ;
        RECT 18.800 15.560 19.590 15.900 ;
        RECT 19.760 15.720 19.930 17.330 ;
        RECT 21.480 17.260 21.810 17.520 ;
        RECT 23.960 17.260 24.290 17.520 ;
        RECT 21.960 16.250 22.130 17.090 ;
        RECT 22.920 16.250 23.090 17.090 ;
        RECT 24.440 16.250 24.610 17.090 ;
        RECT 25.400 16.250 25.570 17.090 ;
        RECT 20.300 15.720 20.600 15.770 ;
        RECT 17.640 14.050 17.810 15.260 ;
        RECT 18.800 14.660 18.970 15.560 ;
        RECT 19.760 15.530 20.670 15.720 ;
        RECT 19.760 14.660 19.930 15.530 ;
        RECT 20.300 15.470 20.600 15.530 ;
        RECT 12.420 13.880 14.480 14.050 ;
        RECT 14.660 13.880 17.870 14.050 ;
        RECT 14.310 13.710 14.480 13.880 ;
        RECT 14.310 13.540 15.660 13.710 ;
        RECT 6.840 11.970 10.850 12.150 ;
        RECT 5.710 11.840 6.670 11.920 ;
        RECT 5.710 11.670 6.130 11.840 ;
        RECT 4.520 11.500 4.980 11.670 ;
        RECT 5.690 11.500 6.150 11.670 ;
        RECT 6.340 11.650 6.670 11.840 ;
        RECT 4.540 11.470 4.960 11.500 ;
        RECT 5.710 11.470 6.130 11.500 ;
        RECT 6.840 11.020 7.010 11.970 ;
        RECT 7.800 11.020 7.970 11.970 ;
        RECT 8.760 11.020 8.930 11.970 ;
        RECT 9.720 11.020 9.890 11.970 ;
        RECT 10.680 11.020 10.850 11.970 ;
        RECT 11.850 11.840 12.230 13.130 ;
        RECT 11.820 10.890 12.770 11.840 ;
        RECT 14.590 10.990 14.760 13.540 ;
        RECT 15.880 13.370 16.050 13.880 ;
        RECT 15.550 13.200 16.050 13.370 ;
        RECT 16.930 13.210 17.540 13.550 ;
        RECT 15.550 10.990 15.720 13.200 ;
        RECT 18.800 12.740 18.970 13.640 ;
        RECT 19.760 12.770 19.930 13.640 ;
        RECT 20.320 12.770 20.620 12.820 ;
        RECT 18.800 12.400 19.590 12.740 ;
        RECT 19.760 12.580 20.680 12.770 ;
        RECT 18.800 10.970 18.970 12.400 ;
        RECT 19.760 10.970 19.930 12.580 ;
        RECT 20.320 12.520 20.620 12.580 ;
        RECT 21.300 11.060 21.540 14.730 ;
        RECT 21.710 12.280 21.950 14.260 ;
        RECT 22.860 12.250 23.190 12.510 ;
        RECT 22.760 11.230 22.930 12.070 ;
        RECT 23.720 11.230 23.890 12.070 ;
        RECT 21.300 10.800 22.610 11.060 ;
        RECT 13.180 10.400 13.900 10.670 ;
        RECT 5.320 6.540 8.120 6.740 ;
        RECT 5.320 5.940 5.870 6.540 ;
        RECT 5.320 5.740 8.120 5.940 ;
        RECT 5.320 5.140 5.870 5.740 ;
        RECT 8.870 5.190 9.070 6.740 ;
        RECT 9.670 5.190 9.870 6.740 ;
        RECT 10.470 5.190 10.670 6.740 ;
        RECT 11.270 5.190 11.470 6.740 ;
        RECT 12.070 5.190 12.270 6.740 ;
        RECT 12.870 5.190 13.070 6.740 ;
        RECT 13.670 5.190 13.870 6.740 ;
        RECT 14.470 5.190 14.670 6.740 ;
        RECT 15.270 5.190 15.470 6.740 ;
        RECT 16.070 5.190 16.270 6.740 ;
        RECT 16.870 5.190 17.070 6.740 ;
        RECT 17.670 5.190 17.870 6.740 ;
        RECT 18.470 5.190 18.670 6.740 ;
        RECT 19.270 5.190 19.470 6.740 ;
        RECT 20.070 5.190 20.270 6.740 ;
        RECT 20.870 5.190 21.070 6.740 ;
        RECT 21.820 6.540 24.620 6.740 ;
        RECT 24.070 5.940 24.620 6.540 ;
        RECT 21.820 5.740 24.620 5.940 ;
        RECT 8.870 5.140 21.070 5.190 ;
        RECT 24.070 5.140 24.620 5.740 ;
        RECT 5.320 4.840 24.620 5.140 ;
        RECT 5.320 4.240 5.870 4.840 ;
        RECT 8.870 4.790 21.070 4.840 ;
        RECT 5.320 4.040 8.120 4.240 ;
        RECT 5.320 3.440 5.870 4.040 ;
        RECT 5.320 3.240 8.120 3.440 ;
        RECT 8.870 3.240 9.070 4.790 ;
        RECT 9.670 3.240 9.870 4.790 ;
        RECT 10.470 3.240 10.670 4.790 ;
        RECT 11.270 3.240 11.470 4.790 ;
        RECT 12.070 3.240 12.270 4.790 ;
        RECT 12.870 3.240 13.070 4.790 ;
        RECT 13.670 3.240 13.870 4.790 ;
        RECT 14.470 3.290 14.670 4.790 ;
        RECT 15.270 3.290 15.470 4.790 ;
        RECT 16.070 3.240 16.270 4.790 ;
        RECT 16.870 3.240 17.070 4.790 ;
        RECT 17.670 3.240 17.870 4.790 ;
        RECT 18.470 3.240 18.670 4.790 ;
        RECT 19.270 3.240 19.470 4.790 ;
        RECT 20.070 3.240 20.270 4.790 ;
        RECT 20.870 3.240 21.070 4.790 ;
        RECT 24.070 4.240 24.620 4.840 ;
        RECT 21.820 4.040 24.620 4.240 ;
        RECT 24.070 3.440 24.620 4.040 ;
        RECT 21.820 3.240 24.620 3.440 ;
      LAYER mcon ;
        RECT 5.420 23.540 5.670 23.790 ;
        RECT 5.420 23.090 5.670 23.340 ;
        RECT 24.270 23.490 24.520 23.740 ;
        RECT 24.270 23.040 24.520 23.290 ;
        RECT 5.420 22.590 5.670 22.840 ;
        RECT 5.420 22.140 5.670 22.390 ;
        RECT 24.270 22.540 24.520 22.790 ;
        RECT 24.270 22.090 24.520 22.340 ;
        RECT 11.420 16.390 12.170 17.140 ;
        RECT 4.600 13.220 4.900 13.390 ;
        RECT 5.770 13.220 6.070 13.390 ;
        RECT 4.600 12.310 4.900 12.480 ;
        RECT 5.770 12.310 6.070 12.480 ;
        RECT 5.350 11.870 5.520 12.040 ;
        RECT 8.240 14.890 8.420 15.070 ;
        RECT 11.950 15.240 12.130 15.420 ;
        RECT 11.950 14.870 12.130 15.050 ;
        RECT 11.950 14.500 12.130 14.680 ;
        RECT 11.950 13.950 12.130 14.130 ;
        RECT 18.420 15.700 18.600 15.870 ;
        RECT 18.420 15.340 18.600 15.510 ;
        RECT 24.040 17.320 24.210 17.490 ;
        RECT 20.330 15.530 20.510 15.710 ;
        RECT 11.950 13.570 12.130 13.750 ;
        RECT 11.950 13.200 12.130 13.380 ;
        RECT 11.920 10.990 12.670 11.740 ;
        RECT 16.960 13.290 17.140 13.470 ;
        RECT 17.330 13.290 17.510 13.470 ;
        RECT 20.360 12.580 20.530 12.760 ;
        RECT 21.330 12.640 21.510 12.820 ;
        RECT 21.740 14.020 21.920 14.200 ;
        RECT 21.740 12.340 21.920 12.520 ;
        RECT 22.940 12.290 23.110 12.460 ;
        RECT 13.260 10.450 13.430 10.620 ;
        RECT 13.650 10.450 13.820 10.620 ;
        RECT 5.420 5.590 5.670 5.840 ;
        RECT 5.420 5.140 5.670 5.390 ;
        RECT 24.270 5.540 24.520 5.790 ;
        RECT 24.270 5.090 24.520 5.340 ;
        RECT 5.420 4.640 5.670 4.890 ;
        RECT 5.420 4.190 5.670 4.440 ;
        RECT 24.270 4.590 24.520 4.840 ;
        RECT 24.270 4.140 24.520 4.390 ;
      LAYER met1 ;
        RECT 9.720 25.690 20.220 26.890 ;
        RECT 14.670 25.240 15.270 25.690 ;
        RECT 9.070 25.090 20.870 25.240 ;
        RECT 4.120 23.240 5.770 23.890 ;
        RECT 6.220 23.240 6.370 24.740 ;
        RECT 6.820 23.240 6.970 24.740 ;
        RECT 7.420 23.240 7.570 24.740 ;
        RECT 8.020 23.240 8.170 24.740 ;
        RECT 14.670 24.640 15.270 25.090 ;
        RECT 9.070 24.490 20.870 24.640 ;
        RECT 14.670 24.040 15.270 24.490 ;
        RECT 9.070 23.890 20.870 24.040 ;
        RECT 14.670 23.440 15.270 23.890 ;
        RECT 9.070 23.290 20.870 23.440 ;
        RECT 4.120 23.140 8.170 23.240 ;
        RECT 14.670 23.140 15.270 23.290 ;
        RECT 21.770 23.240 21.920 24.740 ;
        RECT 22.370 23.240 22.520 24.740 ;
        RECT 22.970 23.240 23.120 24.740 ;
        RECT 23.570 23.240 23.720 24.740 ;
        RECT 24.170 23.240 25.820 23.840 ;
        RECT 21.770 23.140 25.820 23.240 ;
        RECT 4.120 22.440 25.820 23.140 ;
        RECT 4.120 22.040 5.770 22.440 ;
        RECT 6.220 21.140 6.370 22.440 ;
        RECT 6.820 21.140 6.970 22.440 ;
        RECT 7.420 21.140 7.570 22.440 ;
        RECT 8.020 21.140 8.170 22.440 ;
        RECT 14.670 21.990 15.270 22.440 ;
        RECT 9.070 21.840 20.870 21.990 ;
        RECT 14.670 21.390 15.270 21.840 ;
        RECT 9.070 21.240 20.870 21.390 ;
        RECT 14.670 20.790 15.270 21.240 ;
        RECT 21.770 21.140 21.920 22.440 ;
        RECT 22.370 21.140 22.520 22.440 ;
        RECT 22.970 21.140 23.120 22.440 ;
        RECT 23.570 21.140 23.720 22.440 ;
        RECT 24.170 21.990 25.820 22.440 ;
        RECT 9.070 20.640 20.870 20.790 ;
        RECT 14.670 20.190 15.270 20.640 ;
        RECT 9.720 18.990 20.220 20.190 ;
        RECT 20.600 17.520 21.820 17.550 ;
        RECT 20.600 17.380 24.270 17.520 ;
        RECT 11.320 16.290 12.270 17.240 ;
        RECT 8.180 15.080 8.450 15.100 ;
        RECT 11.890 15.080 12.190 15.470 ;
        RECT 18.350 15.250 18.630 15.950 ;
        RECT 20.600 15.770 20.780 17.380 ;
        RECT 23.960 17.290 24.270 17.380 ;
        RECT 20.300 15.470 20.780 15.770 ;
        RECT 8.180 15.010 12.190 15.080 ;
        RECT 8.170 14.820 12.190 15.010 ;
        RECT 11.890 14.470 12.190 14.820 ;
        RECT 20.600 14.260 20.780 15.470 ;
        RECT 4.560 12.250 4.950 13.460 ;
        RECT 5.730 12.250 6.120 13.460 ;
        RECT 11.890 13.390 12.190 14.160 ;
        RECT 20.600 14.070 21.950 14.260 ;
        RECT 21.710 13.960 21.950 14.070 ;
        RECT 16.910 13.390 17.560 13.550 ;
        RECT 11.890 13.210 17.560 13.390 ;
        RECT 11.890 13.170 12.190 13.210 ;
        RECT 20.320 12.770 20.620 12.820 ;
        RECT 21.300 12.770 21.540 12.880 ;
        RECT 20.320 12.580 21.540 12.770 ;
        RECT 20.320 12.520 20.620 12.580 ;
        RECT 21.710 12.450 21.950 12.580 ;
        RECT 22.860 12.450 23.190 12.510 ;
        RECT 21.710 12.270 23.190 12.450 ;
        RECT 21.710 12.260 22.200 12.270 ;
        RECT 22.860 12.250 23.190 12.270 ;
        RECT 5.270 11.950 5.550 12.120 ;
        RECT 5.270 11.790 6.570 11.950 ;
        RECT 6.360 10.670 6.570 11.790 ;
        RECT 11.820 10.890 12.770 11.840 ;
        RECT 6.360 10.400 13.900 10.670 ;
        RECT 9.720 7.740 20.220 8.940 ;
        RECT 14.670 7.290 15.270 7.740 ;
        RECT 9.070 7.140 20.870 7.290 ;
        RECT 4.120 5.290 5.770 5.940 ;
        RECT 6.220 5.290 6.370 6.790 ;
        RECT 6.820 5.290 6.970 6.790 ;
        RECT 7.420 5.290 7.570 6.790 ;
        RECT 8.020 5.290 8.170 6.790 ;
        RECT 14.670 6.690 15.270 7.140 ;
        RECT 9.070 6.540 20.870 6.690 ;
        RECT 14.670 6.090 15.270 6.540 ;
        RECT 9.070 5.940 20.870 6.090 ;
        RECT 14.670 5.490 15.270 5.940 ;
        RECT 9.070 5.340 20.870 5.490 ;
        RECT 4.120 5.190 8.170 5.290 ;
        RECT 14.670 5.190 15.270 5.340 ;
        RECT 21.770 5.290 21.920 6.790 ;
        RECT 22.370 5.290 22.520 6.790 ;
        RECT 22.970 5.290 23.120 6.790 ;
        RECT 23.570 5.290 23.720 6.790 ;
        RECT 24.170 5.290 25.820 5.890 ;
        RECT 21.770 5.190 25.820 5.290 ;
        RECT 4.120 4.490 25.820 5.190 ;
        RECT 4.120 4.090 5.770 4.490 ;
        RECT 6.220 3.190 6.370 4.490 ;
        RECT 6.820 3.190 6.970 4.490 ;
        RECT 7.420 3.190 7.570 4.490 ;
        RECT 8.020 3.190 8.170 4.490 ;
        RECT 14.670 4.040 15.270 4.490 ;
        RECT 9.070 3.890 20.870 4.040 ;
        RECT 14.670 3.440 15.270 3.890 ;
        RECT 9.070 3.290 20.870 3.440 ;
        RECT 14.670 2.840 15.270 3.290 ;
        RECT 21.770 3.190 21.920 4.490 ;
        RECT 22.370 3.190 22.520 4.490 ;
        RECT 22.970 3.190 23.120 4.490 ;
        RECT 23.570 3.190 23.720 4.490 ;
        RECT 24.170 4.040 25.820 4.490 ;
        RECT 9.070 2.690 20.870 2.840 ;
        RECT 14.670 2.240 15.270 2.690 ;
        RECT 9.720 1.040 20.220 2.240 ;
      LAYER via ;
        RECT 9.820 25.790 10.820 26.790 ;
        RECT 10.920 25.790 11.920 26.790 ;
        RECT 14.520 25.790 15.420 26.790 ;
        RECT 18.020 25.790 19.020 26.790 ;
        RECT 19.120 25.790 20.120 26.790 ;
        RECT 4.220 23.190 5.220 23.740 ;
        RECT 24.720 23.190 25.720 23.740 ;
        RECT 4.220 22.140 5.220 22.690 ;
        RECT 24.720 22.140 25.720 22.690 ;
        RECT 9.820 19.090 10.820 20.090 ;
        RECT 10.920 19.090 11.920 20.090 ;
        RECT 14.520 19.090 15.420 20.090 ;
        RECT 18.020 19.090 19.020 20.090 ;
        RECT 19.120 19.090 20.120 20.090 ;
        RECT 11.420 16.390 12.170 17.140 ;
        RECT 11.920 10.990 12.670 11.740 ;
        RECT 9.820 7.840 10.820 8.840 ;
        RECT 10.920 7.840 11.920 8.840 ;
        RECT 14.520 7.840 15.420 8.840 ;
        RECT 18.020 7.840 19.020 8.840 ;
        RECT 19.120 7.840 20.120 8.840 ;
        RECT 4.220 5.240 5.220 5.790 ;
        RECT 24.720 5.240 25.720 5.790 ;
        RECT 4.220 4.190 5.220 4.740 ;
        RECT 24.720 4.190 25.720 4.740 ;
        RECT 9.820 1.140 10.820 2.140 ;
        RECT 10.920 1.140 11.920 2.140 ;
        RECT 14.520 1.140 15.420 2.140 ;
        RECT 18.020 1.140 19.020 2.140 ;
        RECT 19.120 1.140 20.120 2.140 ;
      LAYER met2 ;
        RECT 9.720 25.490 20.220 26.890 ;
        RECT 6.220 24.890 23.720 25.490 ;
        RECT 8.220 24.440 8.520 24.890 ;
        RECT 6.220 24.290 8.520 24.440 ;
        RECT 8.220 23.840 8.520 24.290 ;
        RECT 4.120 22.040 5.320 23.840 ;
        RECT 6.220 23.690 8.520 23.840 ;
        RECT 8.220 23.240 8.520 23.690 ;
        RECT 8.970 23.240 9.120 24.890 ;
        RECT 9.570 23.240 9.720 24.890 ;
        RECT 10.170 23.240 10.320 24.890 ;
        RECT 10.770 23.240 10.920 24.890 ;
        RECT 11.370 23.240 11.520 24.890 ;
        RECT 11.970 23.240 12.120 24.890 ;
        RECT 12.570 23.240 12.720 24.890 ;
        RECT 13.170 23.240 13.320 24.890 ;
        RECT 13.770 23.240 13.920 24.890 ;
        RECT 14.370 23.240 14.520 24.890 ;
        RECT 15.420 23.240 15.570 24.890 ;
        RECT 16.020 23.240 16.170 24.890 ;
        RECT 16.620 23.240 16.770 24.890 ;
        RECT 17.220 23.240 17.370 24.890 ;
        RECT 17.820 23.240 17.970 24.890 ;
        RECT 18.420 23.240 18.570 24.890 ;
        RECT 19.020 23.240 19.170 24.890 ;
        RECT 19.620 23.240 19.770 24.890 ;
        RECT 20.220 23.240 20.370 24.890 ;
        RECT 20.820 23.240 20.970 24.890 ;
        RECT 21.420 24.440 21.720 24.890 ;
        RECT 21.420 24.290 23.720 24.440 ;
        RECT 21.420 23.840 21.720 24.290 ;
        RECT 21.420 23.690 23.720 23.840 ;
        RECT 21.420 23.240 21.720 23.690 ;
        RECT 8.220 22.190 8.520 22.640 ;
        RECT 6.220 22.040 8.520 22.190 ;
        RECT 8.220 21.590 8.520 22.040 ;
        RECT 6.220 21.440 8.520 21.590 ;
        RECT 8.220 20.990 8.520 21.440 ;
        RECT 8.970 20.990 9.120 22.640 ;
        RECT 9.570 20.990 9.720 22.640 ;
        RECT 10.170 20.990 10.320 22.640 ;
        RECT 10.770 20.990 10.920 22.640 ;
        RECT 11.370 20.990 11.520 22.640 ;
        RECT 11.970 20.990 12.120 22.640 ;
        RECT 12.570 20.990 12.720 22.640 ;
        RECT 13.170 20.990 13.320 22.640 ;
        RECT 13.770 20.990 13.920 22.640 ;
        RECT 14.370 20.990 14.520 22.640 ;
        RECT 15.420 20.990 15.570 22.640 ;
        RECT 16.020 20.990 16.170 22.640 ;
        RECT 16.620 20.990 16.770 22.640 ;
        RECT 17.220 20.990 17.370 22.640 ;
        RECT 17.820 20.990 17.970 22.640 ;
        RECT 18.420 20.990 18.570 22.640 ;
        RECT 19.020 20.990 19.170 22.640 ;
        RECT 19.620 20.990 19.770 22.640 ;
        RECT 20.220 20.990 20.370 22.640 ;
        RECT 20.820 20.990 20.970 22.640 ;
        RECT 21.420 22.190 21.720 22.640 ;
        RECT 21.420 22.040 23.720 22.190 ;
        RECT 24.620 22.040 25.820 23.840 ;
        RECT 21.420 21.590 21.720 22.040 ;
        RECT 21.420 21.440 23.720 21.590 ;
        RECT 21.420 20.990 21.720 21.440 ;
        RECT 6.220 20.390 23.720 20.990 ;
        RECT 9.720 18.990 20.220 20.390 ;
        RECT 11.320 16.290 12.270 18.990 ;
        RECT 11.820 8.940 12.770 11.840 ;
        RECT 9.720 7.540 20.220 8.940 ;
        RECT 6.220 6.940 23.720 7.540 ;
        RECT 8.220 6.490 8.520 6.940 ;
        RECT 6.220 6.340 8.520 6.490 ;
        RECT 8.220 5.890 8.520 6.340 ;
        RECT 4.120 4.090 5.320 5.890 ;
        RECT 6.220 5.740 8.520 5.890 ;
        RECT 8.220 5.290 8.520 5.740 ;
        RECT 8.970 5.290 9.120 6.940 ;
        RECT 9.570 5.290 9.720 6.940 ;
        RECT 10.170 5.290 10.320 6.940 ;
        RECT 10.770 5.290 10.920 6.940 ;
        RECT 11.370 5.290 11.520 6.940 ;
        RECT 11.970 5.290 12.120 6.940 ;
        RECT 12.570 5.290 12.720 6.940 ;
        RECT 13.170 5.290 13.320 6.940 ;
        RECT 13.770 5.290 13.920 6.940 ;
        RECT 14.370 5.290 14.520 6.940 ;
        RECT 15.420 5.290 15.570 6.940 ;
        RECT 16.020 5.290 16.170 6.940 ;
        RECT 16.620 5.290 16.770 6.940 ;
        RECT 17.220 5.290 17.370 6.940 ;
        RECT 17.820 5.290 17.970 6.940 ;
        RECT 18.420 5.290 18.570 6.940 ;
        RECT 19.020 5.290 19.170 6.940 ;
        RECT 19.620 5.290 19.770 6.940 ;
        RECT 20.220 5.290 20.370 6.940 ;
        RECT 20.820 5.290 20.970 6.940 ;
        RECT 21.420 6.490 21.720 6.940 ;
        RECT 21.420 6.340 23.720 6.490 ;
        RECT 21.420 5.890 21.720 6.340 ;
        RECT 21.420 5.740 23.720 5.890 ;
        RECT 21.420 5.290 21.720 5.740 ;
        RECT 8.220 4.240 8.520 4.690 ;
        RECT 6.220 4.090 8.520 4.240 ;
        RECT 8.220 3.640 8.520 4.090 ;
        RECT 6.220 3.490 8.520 3.640 ;
        RECT 8.220 3.040 8.520 3.490 ;
        RECT 8.970 3.040 9.120 4.690 ;
        RECT 9.570 3.040 9.720 4.690 ;
        RECT 10.170 3.040 10.320 4.690 ;
        RECT 10.770 3.040 10.920 4.690 ;
        RECT 11.370 3.040 11.520 4.690 ;
        RECT 11.970 3.040 12.120 4.690 ;
        RECT 12.570 3.040 12.720 4.690 ;
        RECT 13.170 3.040 13.320 4.690 ;
        RECT 13.770 3.040 13.920 4.690 ;
        RECT 14.370 3.040 14.520 4.690 ;
        RECT 15.420 3.040 15.570 4.690 ;
        RECT 16.020 3.040 16.170 4.690 ;
        RECT 16.620 3.040 16.770 4.690 ;
        RECT 17.220 3.040 17.370 4.690 ;
        RECT 17.820 3.040 17.970 4.690 ;
        RECT 18.420 3.040 18.570 4.690 ;
        RECT 19.020 3.040 19.170 4.690 ;
        RECT 19.620 3.040 19.770 4.690 ;
        RECT 20.220 3.040 20.370 4.690 ;
        RECT 20.820 3.040 20.970 4.690 ;
        RECT 21.420 4.240 21.720 4.690 ;
        RECT 21.420 4.090 23.720 4.240 ;
        RECT 24.620 4.090 25.820 5.890 ;
        RECT 21.420 3.640 21.720 4.090 ;
        RECT 21.420 3.490 23.720 3.640 ;
        RECT 21.420 3.040 21.720 3.490 ;
        RECT 6.220 2.440 23.720 3.040 ;
        RECT 9.720 1.040 20.220 2.440 ;
  END
END adc_comp_latch
END LIBRARY

