magic
tech sky130A
timestamp 1686123651
<< nwell >>
rect 100 605 2064 678
rect 90 185 2075 605
rect 100 112 2064 185
<< pwell >>
rect 0 678 2170 790
rect 0 605 100 678
rect 2064 605 2170 678
rect 0 185 90 605
rect 2075 185 2170 605
rect 0 112 100 185
rect 2064 112 2170 185
rect 0 0 2170 112
<< varactor >>
rect 165 200 2005 590
<< psubdiff >>
rect 325 740 555 750
rect 325 715 340 740
rect 540 715 555 740
rect 325 705 555 715
rect 1615 740 1845 750
rect 1615 715 1630 740
rect 1830 715 1845 740
rect 1615 705 1845 715
rect 325 75 555 85
rect 325 50 340 75
rect 540 50 555 75
rect 325 40 555 50
rect 1615 75 1845 85
rect 1615 50 1630 75
rect 1830 50 1845 75
rect 1615 40 1845 50
<< nsubdiff >>
rect 165 650 2005 660
rect 165 615 250 650
rect 1920 615 2005 650
rect 165 590 2005 615
rect 165 175 2005 200
rect 165 140 250 175
rect 1920 140 2005 175
rect 165 130 2005 140
<< psubdiffcont >>
rect 340 715 540 740
rect 1630 715 1830 740
rect 340 50 540 75
rect 1630 50 1830 75
<< nsubdiffcont >>
rect 250 615 1920 650
rect 250 140 1920 175
<< poly >>
rect 105 525 165 590
rect 105 500 120 525
rect 145 500 165 525
rect 105 480 165 500
rect 105 455 120 480
rect 145 455 165 480
rect 105 435 165 455
rect 105 410 120 435
rect 145 410 165 435
rect 105 385 165 410
rect 105 360 120 385
rect 145 360 165 385
rect 105 340 165 360
rect 105 315 120 340
rect 145 315 165 340
rect 105 295 165 315
rect 105 270 120 295
rect 145 270 165 295
rect 105 200 165 270
rect 2005 520 2060 590
rect 2005 495 2025 520
rect 2050 495 2060 520
rect 2005 475 2060 495
rect 2005 450 2025 475
rect 2050 450 2060 475
rect 2005 430 2060 450
rect 2005 405 2025 430
rect 2050 405 2060 430
rect 2005 380 2060 405
rect 2005 355 2025 380
rect 2050 355 2060 380
rect 2005 335 2060 355
rect 2005 310 2025 335
rect 2050 310 2060 335
rect 2005 290 2060 310
rect 2005 265 2025 290
rect 2050 265 2060 290
rect 2005 200 2060 265
<< polycont >>
rect 120 500 145 525
rect 120 455 145 480
rect 120 410 145 435
rect 120 360 145 385
rect 120 315 145 340
rect 120 270 145 295
rect 2025 495 2050 520
rect 2025 450 2050 475
rect 2025 405 2050 430
rect 2025 355 2050 380
rect 2025 310 2050 335
rect 2025 265 2050 290
<< locali >>
rect 325 750 555 790
rect 1615 750 1845 790
rect 40 740 2130 750
rect 40 715 340 740
rect 540 715 1630 740
rect 1830 715 2130 740
rect 40 710 2130 715
rect 40 80 80 710
rect 325 705 555 710
rect 1615 705 1845 710
rect 160 600 170 650
rect 230 600 250 650
rect 310 600 330 615
rect 390 600 410 615
rect 470 600 1700 615
rect 1760 600 1780 615
rect 1840 600 1860 615
rect 1920 600 1940 650
rect 2000 600 2010 650
rect 160 590 2010 600
rect 120 550 400 570
rect 120 525 175 550
rect 420 530 455 590
rect 145 500 175 525
rect 195 510 455 530
rect 120 490 175 500
rect 120 480 400 490
rect 155 470 400 480
rect 155 455 175 470
rect 120 435 175 455
rect 420 450 455 510
rect 155 410 175 435
rect 195 430 455 450
rect 475 415 495 570
rect 515 440 535 590
rect 555 415 575 570
rect 595 440 615 590
rect 635 415 655 570
rect 675 440 695 590
rect 715 415 735 570
rect 755 440 775 590
rect 795 415 815 570
rect 835 440 855 590
rect 875 415 895 570
rect 915 440 935 590
rect 955 415 975 570
rect 995 440 1015 590
rect 1035 415 1055 570
rect 1075 440 1095 590
rect 1115 415 1135 570
rect 1155 440 1175 590
rect 1195 415 1215 570
rect 1235 440 1255 590
rect 1275 415 1295 570
rect 1315 440 1335 590
rect 1355 415 1375 570
rect 1395 440 1415 590
rect 1435 415 1455 570
rect 1475 440 1495 590
rect 1515 415 1535 570
rect 1555 440 1575 590
rect 1595 415 1615 570
rect 1635 440 1655 590
rect 1675 415 1695 570
rect 1715 530 1750 590
rect 1770 550 2050 570
rect 1715 510 1975 530
rect 1995 520 2050 550
rect 1715 450 1750 510
rect 1995 495 2025 520
rect 1995 490 2050 495
rect 1770 475 2050 490
rect 1770 470 2015 475
rect 1995 450 2015 470
rect 1715 430 1970 450
rect 1995 430 2050 450
rect 475 410 1695 415
rect 1995 410 2015 430
rect 120 405 2015 410
rect 120 385 2050 405
rect 155 380 2050 385
rect 155 360 175 380
rect 475 375 1695 380
rect 120 340 175 360
rect 195 340 455 360
rect 155 320 175 340
rect 155 315 400 320
rect 120 300 400 315
rect 120 295 175 300
rect 145 270 175 295
rect 420 280 455 340
rect 120 240 175 270
rect 195 260 455 280
rect 120 220 400 240
rect 420 200 455 260
rect 475 220 495 375
rect 515 200 535 350
rect 555 220 575 375
rect 595 200 615 350
rect 635 220 655 375
rect 675 200 695 350
rect 715 220 735 375
rect 755 200 775 350
rect 795 220 815 375
rect 835 200 855 350
rect 875 220 895 375
rect 915 200 935 350
rect 955 220 975 375
rect 995 200 1015 350
rect 1035 225 1055 375
rect 1075 200 1095 350
rect 1115 225 1135 375
rect 1155 200 1175 350
rect 1195 220 1215 375
rect 1235 200 1255 350
rect 1275 220 1295 375
rect 1315 200 1335 350
rect 1355 220 1375 375
rect 1395 200 1415 350
rect 1435 220 1455 375
rect 1475 200 1495 350
rect 1515 220 1535 375
rect 1555 200 1575 350
rect 1595 220 1615 375
rect 1635 200 1655 350
rect 1675 220 1695 375
rect 1715 340 1970 360
rect 1995 355 2015 380
rect 1715 280 1750 340
rect 1995 335 2050 355
rect 1995 320 2015 335
rect 1770 310 2015 320
rect 1770 300 2050 310
rect 1995 290 2050 300
rect 1715 260 1975 280
rect 1995 265 2025 290
rect 1715 200 1750 260
rect 1995 240 2050 265
rect 1770 220 2050 240
rect 160 190 2010 200
rect 160 140 170 190
rect 230 140 250 190
rect 310 175 330 190
rect 390 175 410 190
rect 470 175 1700 190
rect 1760 175 1780 190
rect 1840 175 1860 190
rect 1920 140 1940 190
rect 2000 140 2010 190
rect 325 80 555 85
rect 1615 80 1845 85
rect 2090 80 2130 710
rect 40 75 2130 80
rect 40 50 340 75
rect 540 50 1630 75
rect 1830 50 2130 75
rect 40 40 2130 50
rect 325 0 555 40
rect 1615 0 1845 40
<< viali >>
rect 170 600 230 650
rect 250 615 310 650
rect 330 615 390 650
rect 410 615 470 650
rect 1700 615 1760 650
rect 1780 615 1840 650
rect 1860 615 1920 650
rect 250 600 310 615
rect 330 600 390 615
rect 410 600 470 615
rect 1700 600 1760 615
rect 1780 600 1840 615
rect 1860 600 1920 615
rect 1940 600 2000 650
rect 130 455 145 480
rect 145 455 155 480
rect 130 410 145 435
rect 145 410 155 435
rect 2015 450 2025 475
rect 2025 450 2040 475
rect 2015 405 2025 430
rect 2025 405 2040 430
rect 130 360 145 385
rect 145 360 155 385
rect 130 315 145 340
rect 145 315 155 340
rect 2015 355 2025 380
rect 2025 355 2040 380
rect 2015 310 2025 335
rect 2025 310 2040 335
rect 170 140 230 190
rect 250 175 310 190
rect 330 175 390 190
rect 410 175 470 190
rect 1700 175 1760 190
rect 1780 175 1840 190
rect 1860 175 1920 190
rect 250 140 310 175
rect 330 140 390 175
rect 410 140 470 175
rect 1700 140 1760 175
rect 1780 140 1840 175
rect 1860 140 1920 175
rect 1940 140 2000 190
<< metal1 >>
rect 0 780 320 790
rect 0 680 10 780
rect 110 680 210 780
rect 310 680 320 780
rect 0 670 320 680
rect 560 780 1610 790
rect 560 680 570 780
rect 670 680 680 780
rect 780 680 1040 780
rect 1130 680 1390 780
rect 1490 680 1500 780
rect 1600 680 1610 780
rect 560 670 1610 680
rect 1850 780 2170 790
rect 1850 680 1860 780
rect 1960 680 2060 780
rect 2160 680 2170 780
rect 1850 670 2170 680
rect 0 655 230 670
rect 0 650 1040 655
rect 0 620 170 650
rect 0 520 10 620
rect 110 600 170 620
rect 230 600 250 650
rect 310 600 330 650
rect 390 600 410 650
rect 470 640 1040 650
rect 470 600 480 640
rect 1055 625 1115 670
rect 1940 655 2170 670
rect 1130 650 2170 655
rect 1130 640 1700 650
rect 495 610 1675 625
rect 110 595 480 600
rect 110 520 120 595
rect 165 590 1040 595
rect 0 505 120 520
rect 0 480 165 490
rect 0 475 130 480
rect 0 420 10 475
rect 110 455 130 475
rect 155 455 165 480
rect 180 455 195 590
rect 110 435 165 455
rect 110 420 130 435
rect 0 410 130 420
rect 155 425 165 435
rect 210 425 225 575
rect 240 455 255 590
rect 270 425 285 575
rect 300 455 315 590
rect 330 425 345 575
rect 360 455 375 590
rect 420 580 1040 590
rect 390 425 405 575
rect 420 535 480 580
rect 1055 565 1115 610
rect 1690 600 1700 640
rect 1760 600 1780 650
rect 1840 600 1860 650
rect 1920 600 1940 650
rect 2000 620 2170 650
rect 2000 600 2060 620
rect 1690 595 2060 600
rect 1130 590 2005 595
rect 1130 580 1750 590
rect 495 550 1675 565
rect 420 520 1040 535
rect 420 475 480 520
rect 1055 505 1115 550
rect 1690 535 1750 580
rect 1130 520 1750 535
rect 495 490 1675 505
rect 420 460 1040 475
rect 420 440 480 460
rect 1055 445 1115 490
rect 1690 475 1750 520
rect 1130 460 1750 475
rect 495 430 1675 445
rect 1690 440 1750 460
rect 155 415 405 425
rect 1055 415 1115 430
rect 1765 425 1780 575
rect 1795 455 1810 590
rect 1825 425 1840 575
rect 1855 455 1870 590
rect 1885 425 1900 575
rect 1915 455 1930 590
rect 1945 425 1960 575
rect 1975 455 1990 590
rect 2050 520 2060 595
rect 2160 520 2170 620
rect 2050 505 2170 520
rect 2005 475 2170 485
rect 2005 450 2015 475
rect 2040 450 2060 475
rect 2005 430 2060 450
rect 2005 425 2015 430
rect 1765 415 2015 425
rect 155 410 2015 415
rect 0 405 2015 410
rect 2040 420 2060 430
rect 2160 420 2170 475
rect 2040 405 2170 420
rect 0 385 2170 405
rect 0 370 130 385
rect 0 315 10 370
rect 110 360 130 370
rect 155 380 2170 385
rect 155 360 2015 380
rect 110 355 2015 360
rect 2040 370 2170 380
rect 2040 355 2060 370
rect 110 345 2060 355
rect 110 340 165 345
rect 110 315 130 340
rect 155 315 165 340
rect 0 305 165 315
rect 0 270 120 285
rect 0 170 10 270
rect 110 195 120 270
rect 180 200 195 330
rect 210 215 225 345
rect 240 200 255 330
rect 270 215 285 345
rect 300 200 315 330
rect 330 215 345 345
rect 360 200 375 330
rect 390 215 405 345
rect 420 315 1040 330
rect 420 270 480 315
rect 1055 300 1115 345
rect 1130 315 1750 330
rect 495 285 1675 300
rect 420 255 1040 270
rect 420 210 480 255
rect 1055 240 1115 285
rect 1690 270 1750 315
rect 1130 255 1750 270
rect 495 225 1675 240
rect 420 200 1040 210
rect 165 195 1040 200
rect 110 190 480 195
rect 110 170 170 190
rect 0 140 170 170
rect 230 140 250 190
rect 310 140 330 190
rect 390 140 410 190
rect 470 150 480 190
rect 1055 180 1115 225
rect 1690 210 1750 255
rect 1765 215 1780 345
rect 1130 200 1750 210
rect 1795 200 1810 330
rect 1825 215 1840 345
rect 1855 200 1870 330
rect 1885 215 1900 345
rect 1915 200 1930 330
rect 1945 215 1960 345
rect 2005 335 2060 345
rect 1975 200 1990 330
rect 2005 310 2015 335
rect 2040 315 2060 335
rect 2160 315 2170 370
rect 2040 310 2170 315
rect 2005 300 2170 310
rect 2050 270 2170 285
rect 1130 195 2005 200
rect 2050 195 2060 270
rect 1690 190 2060 195
rect 495 165 1675 180
rect 470 140 1040 150
rect 0 135 1040 140
rect 0 120 230 135
rect 1055 120 1115 165
rect 1690 150 1700 190
rect 1130 140 1700 150
rect 1760 140 1780 190
rect 1840 140 1860 190
rect 1920 140 1940 190
rect 2000 170 2060 190
rect 2160 170 2170 270
rect 2000 140 2170 170
rect 1130 135 2170 140
rect 1940 120 2170 135
rect 0 110 320 120
rect 0 10 10 110
rect 110 10 210 110
rect 310 10 320 110
rect 0 0 320 10
rect 560 110 1610 120
rect 560 10 570 110
rect 670 10 680 110
rect 780 10 1040 110
rect 1130 10 1390 110
rect 1490 10 1500 110
rect 1600 10 1610 110
rect 560 0 1610 10
rect 1850 110 2170 120
rect 1850 10 1860 110
rect 1960 10 2060 110
rect 2160 10 2170 110
rect 1850 0 2170 10
<< via1 >>
rect 10 680 110 780
rect 210 680 310 780
rect 570 680 670 780
rect 680 680 780 780
rect 1040 680 1130 780
rect 1390 680 1490 780
rect 1500 680 1600 780
rect 1860 680 1960 780
rect 2060 680 2160 780
rect 10 520 110 620
rect 10 420 110 475
rect 2060 520 2160 620
rect 2060 420 2160 475
rect 10 315 110 370
rect 10 170 110 270
rect 2060 315 2160 370
rect 2060 170 2160 270
rect 10 10 110 110
rect 210 10 310 110
rect 570 10 670 110
rect 680 10 780 110
rect 1040 10 1130 110
rect 1390 10 1490 110
rect 1500 10 1600 110
rect 1860 10 1960 110
rect 2060 10 2160 110
<< metal2 >>
rect 0 780 320 790
rect 0 680 10 780
rect 110 680 210 780
rect 310 680 320 780
rect 0 670 320 680
rect 560 780 1610 790
rect 560 680 570 780
rect 670 680 680 780
rect 780 680 1040 780
rect 1130 680 1390 780
rect 1490 680 1500 780
rect 1600 680 1610 780
rect 0 620 195 670
rect 560 650 1610 680
rect 1850 780 2170 790
rect 1850 680 1860 780
rect 1960 680 2060 780
rect 2160 680 2170 780
rect 1850 670 2170 680
rect 0 520 10 620
rect 110 575 195 620
rect 210 590 1960 650
rect 1975 620 2170 670
rect 110 560 395 575
rect 110 520 195 560
rect 410 545 440 590
rect 210 530 440 545
rect 0 515 195 520
rect 0 505 395 515
rect 140 500 395 505
rect 0 475 120 485
rect 0 420 10 475
rect 110 420 120 475
rect 0 370 120 420
rect 0 315 10 370
rect 110 315 120 370
rect 0 305 120 315
rect 140 440 195 500
rect 410 485 440 530
rect 210 470 440 485
rect 140 410 395 440
rect 410 425 440 470
rect 455 410 470 575
rect 485 425 500 590
rect 515 410 530 575
rect 545 425 560 590
rect 575 410 590 575
rect 605 425 620 590
rect 635 410 650 575
rect 665 425 680 590
rect 695 410 710 575
rect 725 425 740 590
rect 755 410 770 575
rect 785 425 800 590
rect 815 410 830 575
rect 845 425 860 590
rect 875 410 890 575
rect 905 425 920 590
rect 935 410 950 575
rect 965 425 980 590
rect 995 410 1010 575
rect 1025 425 1040 590
rect 1055 410 1115 575
rect 1130 425 1145 590
rect 1160 410 1175 575
rect 1190 425 1205 590
rect 1220 410 1235 575
rect 1250 425 1265 590
rect 1280 410 1295 575
rect 1310 425 1325 590
rect 1340 410 1355 575
rect 1370 425 1385 590
rect 1400 410 1415 575
rect 1430 425 1445 590
rect 1460 410 1475 575
rect 1490 425 1505 590
rect 1520 410 1535 575
rect 1550 425 1565 590
rect 1580 410 1595 575
rect 1610 425 1625 590
rect 1640 410 1655 575
rect 1670 425 1685 590
rect 1700 410 1715 575
rect 1730 545 1760 590
rect 1975 575 2060 620
rect 1775 560 2060 575
rect 1730 530 1960 545
rect 1730 485 1760 530
rect 1975 520 2060 560
rect 2160 520 2170 620
rect 1975 515 2170 520
rect 1775 505 2170 515
rect 1775 500 2030 505
rect 1730 470 1960 485
rect 1730 425 1760 470
rect 1975 440 2030 500
rect 1775 410 2030 440
rect 140 380 2030 410
rect 140 335 395 380
rect 140 290 195 335
rect 410 320 440 365
rect 210 305 440 320
rect 140 285 395 290
rect 0 275 395 285
rect 0 270 195 275
rect 0 170 10 270
rect 110 230 195 270
rect 410 260 440 305
rect 210 245 440 260
rect 110 215 395 230
rect 110 170 195 215
rect 410 200 440 245
rect 455 215 470 380
rect 485 200 500 365
rect 515 215 530 380
rect 545 200 560 365
rect 575 215 590 380
rect 605 200 620 365
rect 635 215 650 380
rect 665 200 680 365
rect 695 215 710 380
rect 725 200 740 365
rect 755 215 770 380
rect 785 200 800 365
rect 815 215 830 380
rect 845 200 860 365
rect 875 215 890 380
rect 905 200 920 365
rect 935 215 950 380
rect 965 200 980 365
rect 995 215 1010 380
rect 1025 200 1040 365
rect 1055 215 1115 380
rect 1130 200 1145 365
rect 1160 215 1175 380
rect 1190 200 1205 365
rect 1220 215 1235 380
rect 1250 200 1265 365
rect 1280 215 1295 380
rect 1310 200 1325 365
rect 1340 215 1355 380
rect 1370 200 1385 365
rect 1400 215 1415 380
rect 1430 200 1445 365
rect 1460 215 1475 380
rect 1490 200 1505 365
rect 1520 215 1535 380
rect 1550 200 1565 365
rect 1580 215 1595 380
rect 1610 200 1625 365
rect 1640 215 1655 380
rect 1670 200 1685 365
rect 1700 215 1715 380
rect 1730 320 1760 365
rect 1775 335 2030 380
rect 1730 305 1960 320
rect 1730 260 1760 305
rect 1975 290 2030 335
rect 2050 475 2170 485
rect 2050 420 2060 475
rect 2160 420 2170 475
rect 2050 370 2170 420
rect 2050 315 2060 370
rect 2160 315 2170 370
rect 2050 305 2170 315
rect 1775 285 2030 290
rect 1775 275 2170 285
rect 1975 270 2170 275
rect 1730 245 1960 260
rect 1730 200 1760 245
rect 1975 230 2060 270
rect 1775 215 2060 230
rect 0 120 195 170
rect 210 140 1960 200
rect 1975 170 2060 215
rect 2160 170 2170 270
rect 0 110 320 120
rect 0 10 10 110
rect 110 10 210 110
rect 310 10 320 110
rect 0 0 320 10
rect 560 110 1610 140
rect 1975 120 2170 170
rect 560 10 570 110
rect 670 10 680 110
rect 780 10 1040 110
rect 1130 10 1390 110
rect 1490 10 1500 110
rect 1600 10 1610 110
rect 560 0 1610 10
rect 1850 110 2170 120
rect 1850 10 1860 110
rect 1960 10 2060 110
rect 2160 10 2170 110
rect 1850 0 2170 10
<< metal3 >>
rect 0 780 320 790
rect 0 695 10 780
rect 95 695 220 780
rect 305 695 320 780
rect 560 780 1610 790
rect 560 715 570 780
rect 635 715 650 780
rect 715 715 1455 780
rect 1520 715 1535 780
rect 1600 715 1610 780
rect 560 705 1610 715
rect 1850 780 2170 790
rect 0 665 320 695
rect 1850 695 1865 780
rect 1950 695 2075 780
rect 2160 695 2170 780
rect 1850 665 2170 695
rect 0 650 2170 665
rect 0 565 10 650
rect 95 565 2075 650
rect 2160 565 2170 650
rect 0 550 2170 565
rect 0 505 85 515
rect 0 405 10 505
rect 75 405 85 505
rect 0 385 85 405
rect 0 285 10 385
rect 75 285 85 385
rect 0 275 85 285
rect 125 240 2045 550
rect 2085 505 2170 515
rect 2085 405 2095 505
rect 2160 405 2170 505
rect 2085 385 2170 405
rect 2085 285 2095 385
rect 2160 285 2170 385
rect 2085 275 2170 285
rect 0 225 2170 240
rect 0 140 10 225
rect 95 140 2075 225
rect 2160 140 2170 225
rect 0 125 2170 140
rect 0 95 320 125
rect 0 10 10 95
rect 95 10 220 95
rect 305 10 320 95
rect 1850 95 2170 125
rect 0 0 320 10
rect 560 75 1610 85
rect 560 10 570 75
rect 635 10 650 75
rect 715 10 1455 75
rect 1520 10 1535 75
rect 1600 10 1610 75
rect 560 0 1610 10
rect 1850 10 1865 95
rect 1950 10 2075 95
rect 2160 10 2170 95
rect 1850 0 2170 10
<< via3 >>
rect 10 695 95 780
rect 220 695 305 780
rect 570 715 635 780
rect 650 715 715 780
rect 1455 715 1520 780
rect 1535 715 1600 780
rect 1865 695 1950 780
rect 2075 695 2160 780
rect 10 565 95 650
rect 2075 565 2160 650
rect 10 405 75 505
rect 10 285 75 385
rect 2095 405 2160 505
rect 2095 285 2160 385
rect 10 140 95 225
rect 2075 140 2160 225
rect 10 10 95 95
rect 220 10 305 95
rect 570 10 635 75
rect 650 10 715 75
rect 1455 10 1520 75
rect 1535 10 1600 75
rect 1865 10 1950 95
rect 2075 10 2160 95
<< mimcap >>
rect 140 635 2030 650
rect 140 155 155 635
rect 2015 155 2030 635
rect 140 140 2030 155
<< mimcapcontact >>
rect 155 155 2015 635
<< metal4 >>
rect 0 780 315 790
rect 0 695 10 780
rect 95 695 220 780
rect 305 695 315 780
rect 0 685 315 695
rect 560 780 1610 790
rect 560 715 570 780
rect 635 715 650 780
rect 715 715 1455 780
rect 1520 715 1535 780
rect 1600 715 1610 780
rect 0 650 105 685
rect 0 565 10 650
rect 95 565 105 650
rect 560 645 1610 715
rect 1855 780 2170 790
rect 1855 695 1865 780
rect 1950 695 2075 780
rect 2160 695 2170 780
rect 1855 685 2170 695
rect 2065 650 2170 685
rect 0 555 105 565
rect 145 635 2025 645
rect 145 515 155 635
rect 0 505 155 515
rect 0 405 10 505
rect 75 405 155 505
rect 0 385 155 405
rect 0 285 10 385
rect 75 285 155 385
rect 0 275 155 285
rect 0 225 105 235
rect 0 140 10 225
rect 95 140 105 225
rect 145 155 155 275
rect 2015 515 2025 635
rect 2065 565 2075 650
rect 2160 565 2170 650
rect 2065 555 2170 565
rect 2015 505 2170 515
rect 2015 405 2095 505
rect 2160 405 2170 505
rect 2015 385 2170 405
rect 2015 285 2095 385
rect 2160 285 2170 385
rect 2015 275 2170 285
rect 2015 155 2025 275
rect 145 145 2025 155
rect 2065 225 2170 235
rect 0 105 105 140
rect 0 95 315 105
rect 0 10 10 95
rect 95 10 220 95
rect 305 10 315 95
rect 0 0 315 10
rect 560 75 1610 145
rect 2065 140 2075 225
rect 2160 140 2170 225
rect 2065 105 2170 140
rect 560 10 570 75
rect 635 10 650 75
rect 715 10 1455 75
rect 1520 10 1535 75
rect 1600 10 1610 75
rect 560 0 1610 10
rect 1855 95 2170 105
rect 1855 10 1865 95
rect 1950 10 2075 95
rect 2160 10 2170 95
rect 1855 0 2170 10
<< labels >>
flabel metal1 s 0 0 320 120 5 FreeSans 160 0 0 0 nmoscap_bot
port 1 s
flabel metal1 s 0 670 320 790 1 FreeSans 160 0 0 0 nmoscap_bot
port 1 n
flabel metal1 s 1850 0 2170 120 5 FreeSans 160 0 0 0 nmoscap_bot
port 1 s
flabel metal1 s 1850 670 2170 790 1 FreeSans 160 0 0 0 nmoscap_bot
port 1 n
flabel metal1 s 0 505 120 790 7 FreeSans 80 90 0 0 nmoscap_bot
port 1 w
flabel metal1 s 0 0 120 285 7 FreeSans 80 90 0 0 nmoscap_bot
port 1 w
flabel metal1 s 2050 0 2170 285 3 FreeSans 80 90 0 0 nmoscap_bot
port 1 e
flabel metal1 s 2050 505 2170 790 3 FreeSans 80 90 0 0 nmoscap_bot
port 1 e
flabel metal1 s 560 0 1610 120 5 FreeSans 160 0 0 0 nmoscap_top
port 2 s
flabel metal1 s 560 670 1610 790 1 FreeSans 160 0 0 0 nmoscap_top
port 2 n
flabel metal1 s 0 305 120 490 7 FreeSans 160 90 0 0 nmoscap_top
port 2 w
flabel metal1 s 2050 300 2170 485 3 FreeSans 160 90 0 0 nmoscap_top
port 2 e
flabel locali s 325 0 555 40 5 FreeSans 160 0 0 0 pwell
port 3 s
flabel locali s 1615 0 1845 40 5 FreeSans 160 0 0 0 pwell
port 3 s
flabel locali s 325 750 555 790 1 FreeSans 160 0 0 0 pwell
port 3 n
flabel locali s 1615 750 1845 790 1 FreeSans 160 0 0 0 pwell
port 3 n
flabel metal3 s 0 0 320 120 5 FreeSans 160 0 0 0 mimcap_bot
port 4 s
flabel metal3 s 1850 0 2170 120 5 FreeSans 160 0 0 0 mimcap_bot
port 4 s
flabel metal3 s 0 670 320 790 1 FreeSans 160 0 0 0 mimcap_bot
port 4 n
flabel metal3 s 1850 670 2170 790 1 FreeSans 160 0 0 0 mimcap_bot
port 4 n
flabel metal3 s 0 550 125 790 7 FreeSans 160 90 0 0 mimcap_bot
port 4 w
flabel metal3 s 0 0 125 240 7 FreeSans 160 90 0 0 mimcap_bot
port 4 w
flabel metal3 s 2045 0 2170 240 3 FreeSans 160 90 0 0 mimcap_bot
port 4 e
flabel metal3 s 2045 550 2170 790 3 FreeSans 160 90 0 0 mimcap_bot
port 4 e
flabel metal3 s 560 0 1610 85 5 FreeSans 160 0 0 0 mimcap_top
port 5 s
flabel metal3 s 560 705 1610 790 1 FreeSans 160 0 0 0 mimcap_top
port 5 n
flabel metal3 s 2085 275 2170 515 3 FreeSans 160 90 0 0 mimcap_top
port 5 e
flabel metal3 s 0 275 85 515 7 FreeSans 160 90 0 0 mimcap_top
port 5 w
<< properties >>
string FIXED_BBOX 0 0 2170 790
<< end >>
