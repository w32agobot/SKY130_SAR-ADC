* SPICE3 file created from adc_array_wafflecap_16(8)x295aF_28um2.ext - technology: sky130A

.subckt adc_array_wafflecap_16(8)x295aF_28um2 cbot ctop
C0 cbot ctop 2.37fF
C1 cfloating cbot 2.31fF
C2 cbot VSUBS 2.16fF
.ends
