* NGSPICE file created from adc_core_digital.ext - technology: sky130A

.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
.ends

.subckt sky130_fd_sc_hd__decap_8 VPWR VGND VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
.ends

.subckt sky130_fd_sc_hd__decap_3 VPWR VGND VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
.ends

.subckt sky130_fd_sc_hd__nand2_2 Y A B VGND VPWR VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N X A2_N B2 B1 VGND VPWR VNB VPB
X0 a_294_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VPWR A2_N a_295_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 VPWR B1 a_665_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 VGND a_84_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 X a_84_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_581_47# a_295_369# a_84_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR a_84_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_665_369# B2 a_84_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8 VGND B2 a_581_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_295_369# A2_N a_294_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 X a_84_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_84_21# a_295_369# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X12 a_295_369# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X13 a_581_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__xnor2_4 Y B A VGND VPWR VNB VPB
X0 VGND A a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y a_38_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_38_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_820_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR a_38_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND B a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND B a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y B a_820_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_38_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_38_297# B a_38_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND A a_38_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_902_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_820_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_902_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VPWR A a_38_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 Y a_38_297# a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 Y a_38_297# a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_38_47# B a_38_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_38_47# B a_38_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_38_297# B a_38_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 a_38_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 VPWR B a_38_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 a_38_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 a_902_47# a_38_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_902_47# a_38_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 Y B a_820_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_38_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_820_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VPWR A a_38_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 VGND A a_38_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 VPWR A a_820_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 a_902_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X33 a_820_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 Y a_38_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 a_902_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X36 a_38_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X37 VPWR A a_820_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 VPWR a_38_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X39 VPWR B a_38_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__or2_2 B X A VPWR VGND VNB VPB
X0 a_121_297# B a_39_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 X a_39_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR a_39_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_39_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND a_39_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR A a_121_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND A a_39_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_39_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_1 VGND VPWR X A VNB VPB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor2_2 B Y A VGND VPWR VNB VPB
X0 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__decap_6 VPWR VGND VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
.ends

.subckt sky130_fd_sc_hd__o21ai_4 Y B1 A2 A1 VPWR VGND VNB VPB
X0 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_115_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_115_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A1 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A2 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y B1 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND A1 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_32_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 Y B1 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y A2 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_32_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_32_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_32_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_115_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_32_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_32_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VGND A2 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VPWR A1 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 Y A2 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VGND A1 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_115_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__o21ai_2 B1 Y A2 A1 VGND VPWR VNB VPB
X0 VGND A2 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y B1 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A1 a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_29_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y A2 a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND A1 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_112_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_112_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_29_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_29_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and2_2 VPWR VGND A X B VNB VPB
X0 X a_61_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR a_61_75# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR B a_61_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VGND B a_147_75# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 X a_61_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND a_61_75# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_61_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_147_75# A a_61_75# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o31a_2 X A1 A2 B1 A3 VGND VPWR VNB VPB
X0 a_108_21# B1 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_346_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X a_108_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_108_21# A3 a_430_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_430_297# A2 a_346_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR a_108_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_346_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND A2 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 X a_108_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR B1 a_108_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VGND a_108_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_346_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor3_2 C Y A B VGND VPWR VNB VPB
X0 Y C a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_281_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_281_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_27_297# B a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__xnor2_2 VGND VPWR Y A B VNB VPB
X0 a_27_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_560_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND B a_560_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y B a_474_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y a_27_297# a_560_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_474_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND A a_560_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_27_47# B a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_27_297# B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_474_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_560_47# a_27_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VPWR A a_474_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 Y a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VPWR a_27_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_560_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__o211ai_4 A1 B1 A2 C1 Y VGND VPWR VNB VPB
X0 VPWR A1 a_110_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A2 a_110_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_806_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_110_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_110_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_110_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR A1 a_110_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_27_47# B1 a_1314_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 Y A2 a_110_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 Y C1 a_978_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 Y C1 a_806_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 a_27_47# B1 a_806_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_110_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 a_806_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 a_978_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X28 a_1314_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_4 VPWR VGND X A VNB VPB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a31o_2 X B1 A3 A1 A2 VGND VPWR VNB VPB
X0 VPWR A2 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_277_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_79_21# B1 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_277_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_361_47# A2 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_277_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VGND B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_79_21# A1 a_361_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o21bai_4 Y B1_N A1 A2 VGND VPWR VNB VPB
X0 Y a_33_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_225_47# a_33_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR a_33_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_33_297# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y a_33_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y A2 a_561_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y a_33_297# a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y a_33_297# a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VGND A2 a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VGND A2 a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_561_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_225_47# a_33_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VPWR A1 a_561_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_225_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_225_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_225_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_225_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VPWR A1 a_561_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_561_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VPWR B1_N a_33_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_561_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 VGND A1 a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 Y A2 a_561_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VGND A1 a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 a_561_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 VPWR a_33_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__mux2_1 VGND VPWR S A1 A0 X VNB VPB
X0 VPWR a_505_21# a_535_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_505_21# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_218_374# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VGND a_505_21# a_439_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_76_199# A0 a_218_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_505_21# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_439_47# A0 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_535_374# A1 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_76_199# A1 a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_218_47# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__dfrtp_2 Q RESET_B D CLK VGND VPWR VNB VPB
X0 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X4 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X10 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X12 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X15 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X22 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X26 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o22a_2 A2 X B1 A1 B2 VGND VPWR VNB VPB
X0 a_301_47# B2 a_81_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VGND A2 a_301_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_383_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_301_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 X a_81_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 X a_81_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR A1 a_579_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_81_21# B1 a_301_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_579_297# A2 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_81_21# B2 a_383_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__inv_2 A Y VPWR VGND VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__a21oi_4 B1 A2 A1 Y VGND VPWR VNB VPB
X0 a_28_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_462_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y B1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_462_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_28_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_462_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y B1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y A1 a_462_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_28_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VPWR A2 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VGND A2 a_462_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_28_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VPWR A1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_28_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 VGND A2 a_462_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 VPWR A2 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_28_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 Y A1 a_462_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 a_462_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 VPWR A1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__o221a_2 B2 A2 X B1 C1 A1 VGND VPWR VNB VPB
X0 VPWR a_38_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR A1 a_497_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 X a_38_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_141_47# B2 a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_497_297# A2 a_38_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A1 a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR C1 a_38_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_237_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_38_47# B2 a_237_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_225_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 X a_38_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_141_47# C1 a_38_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND a_38_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_225_47# B1 a_141_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand2_8 A B Y VGND VPWR VNB VPB
X0 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_6 VPWR VGND X A VNB VPB
X0 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_161_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A a_161_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VPWR A a_161_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_161_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__a21bo_2 B1_N A2 X A1 VGND VPWR VNB VPB
X0 VPWR A1 a_485_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_485_297# a_297_93# a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_297_93# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_581_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_79_21# a_297_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND A2 a_581_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_297_93# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_485_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__inv_6 Y A VPWR VGND VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a221o_2 X B1 A1 B2 A2 VGND VPWR C1 VNB VPB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_465_47# A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_109_297# B1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_205_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR A2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_193_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_27_47# B1 a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_109_297# C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and2b_2 VPWR VGND X B A_N VNB VPB
X0 VPWR a_212_413# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_297_47# a_27_413# a_212_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 X a_212_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_212_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_212_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR B a_212_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VGND a_212_413# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_2 VPWR VGND X A VNB VPB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__xor2_4 X B A VGND VPWR VNB VPB
X0 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_806_47# B X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_806_47# B X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_112_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_297# B a_112_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_806_297# a_112_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND a_112_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 X B a_806_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 X a_112_47# a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_112_47# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_806_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND A a_806_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 X B a_806_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND A a_806_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_806_297# a_112_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND A a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_112_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VGND A a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_806_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VPWR B a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 VGND B a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 VGND B a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 VPWR B a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 a_806_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_806_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 a_27_297# B a_112_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_112_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X28 VGND a_112_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 a_806_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 a_112_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 a_112_47# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 VPWR A a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 X a_112_47# a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 a_806_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X37 X a_112_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X38 X a_112_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X39 VPWR A a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__and3_2 B X A C VPWR VGND VNB VPB
X0 VPWR a_29_311# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X a_29_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A a_29_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VGND a_29_311# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_184_53# B a_112_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR C a_29_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 X a_29_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_112_53# A a_29_311# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_29_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VGND C a_184_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o21a_2 A1 B1 A2 X VGND VPWR VNB VPB
X0 VPWR A1 a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_470_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_384_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_384_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a21oi_2 B1 A2 A1 Y VGND VPWR VNB VPB
X0 VGND A2 a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y A1 a_114_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_114_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_285_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a21o_2 X B1 A1 A2 VGND VPWR VNB VPB
X0 VPWR a_80_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X a_80_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND a_80_199# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_386_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_80_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_80_199# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_386_297# B1 a_80_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_458_47# A1 a_80_199# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR A1 a_386_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND A2 a_458_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a2bb2o_2 VGND VPWR B1 A1_N A2_N X B2 VNB VPB
X0 VPWR a_82_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_646_47# B2 a_82_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_574_369# a_313_47# a_82_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 a_574_369# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 VGND a_82_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR B2 a_574_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6 X a_82_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 X a_82_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_313_47# A2_N a_313_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X9 a_313_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_313_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X11 VGND A2_N a_313_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_82_21# a_313_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VGND B1 a_646_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o22a_4 B2 B1 X A1 A2 VGND VPWR VNB VPB
X0 VPWR B1 a_566_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_484_47# B1 a_96_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X a_96_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR a_96_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_96_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_566_297# B2 a_96_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR a_96_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X a_96_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VGND a_96_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_96_21# B2 a_566_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR A1 a_918_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_484_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_566_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_484_47# B2 a_96_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_96_21# A2 a_918_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_918_297# A2 a_96_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_484_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_918_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_96_21# B1 a_484_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 VGND A2 a_484_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_96_21# B2 a_484_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VGND A1 a_484_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 X a_96_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VGND a_96_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__dfstp_4 Q D VPWR SET_B CLK VGND VNB VPB
X0 a_1178_261# a_1028_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1 VGND a_652_21# a_586_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VPWR a_1028_413# a_1598_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 a_1178_261# a_1028_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=540000u l=150000u
X4 VGND a_1598_47# Q VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_956_413# a_476_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_1136_413# a_193_47# a_1028_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR a_1598_47# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR a_476_47# a_652_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_586_47# a_193_47# a_476_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X10 VGND a_1598_47# Q VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X12 Q a_1598_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_476_47# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X14 a_1056_47# a_476_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X16 a_652_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_1224_47# a_27_47# a_1028_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 a_562_413# a_27_47# a_476_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 a_1028_413# a_193_47# a_1056_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 a_476_47# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 Q a_1598_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_1296_47# a_1178_261# a_1224_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 VGND a_1028_413# a_1598_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 VPWR a_652_21# a_562_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 VPWR a_1598_47# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 VGND SET_B a_1296_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 Q a_1598_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 a_1028_413# a_27_47# a_956_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 VPWR a_1178_261# a_1136_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X31 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X32 Q a_1598_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 a_796_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X34 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X35 Q a_1598_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X36 Q a_1598_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X37 a_652_21# a_476_47# a_796_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X38 VPWR SET_B a_1028_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X39 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o211a_2 C1 B1 A2 A1 X VPWR VGND VNB VPB
X0 a_27_47# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A1 a_373_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_182_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_182_47# B1 a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_373_297# A2 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_110_47# C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND A1 a_182_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o221ai_2 B1 B2 Y A2 A1 C1 VGND VPWR VNB VPB
X0 Y A2 a_734_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_300_47# B2 a_28_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_300_47# B1 a_28_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_300_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_300_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_734_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_28_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y C1 a_28_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR B1 a_382_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_382_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_28_47# B1 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_28_47# B2 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VGND A1 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 Y B2 a_382_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VPWR A1 a_734_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VGND A2 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_382_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_734_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand2_4 Y A B VGND VPWR VNB VPB
X0 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a211o_2 X A2 A1 B1 C1 VGND VPWR VNB VPB
X0 a_79_21# A1 a_348_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_79_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_79_21# C1 a_585_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR A2 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_299_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_585_297# B1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_348_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a211o_4 VGND VPWR C1 B1 X A2 A1 VNB VPB
X0 X a_79_204# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR A1 a_473_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_473_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_79_204# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND C1 a_79_204# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_79_204# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR a_79_204# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_473_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_473_297# B1 a_727_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X a_79_204# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND B1 a_79_204# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_79_204# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND a_79_204# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_1123_47# A1 a_79_204# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_555_297# B1 a_473_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VPWR A2 a_473_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VGND A2 a_1123_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_951_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VPWR a_79_204# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND a_79_204# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_79_204# A1 a_951_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 a_79_204# C1 a_555_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_727_297# C1 a_79_204# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 X a_79_204# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__and2_4 X B A VGND VPWR VNB VPB
X0 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND B a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_110_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or4_2 C A X B D VPWR VGND VNB VPB
X0 a_27_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_27_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_277_297# B a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR A a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_205_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR a_27_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND a_27_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND C a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_109_297# D a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VGND A a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a211oi_4 A2 A1 C1 Y B1 VPWR VGND VNB VPB
X0 Y A1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND A2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_949_297# B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 Y C1 a_949_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_781_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_27_297# B1 a_781_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND A2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 Y A1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_781_297# B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_1301_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 Y C1 a_781_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_109_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_109_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_109_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_27_297# B1 a_1301_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 a_109_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or3_4 A X B C VPWR VGND VNB VPB
X0 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR A a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_193_297# B a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_109_297# C a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VGND C a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__dfrtp_4 Q RESET_B D CLK VGND VPWR VNB VPB
X0 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X3 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X12 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X16 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X24 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X29 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X31 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X32 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X33 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and4bb_2 VGND VPWR A_N C B_N X D VNB VPB
X0 a_174_21# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_174_21# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_476_47# a_27_47# a_174_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR a_174_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_174_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_548_47# a_505_280# a_476_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 X a_174_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR D a_174_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VGND D a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VPWR a_505_280# a_174_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_505_280# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 VGND a_174_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_505_280# B_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_639_47# C a_548_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a22oi_4 A2 B2 A1 B1 Y VGND VPWR VNB VPB
X0 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y A1 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 Y A1 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND A2 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_27_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_27_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_803_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_803_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_803_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_803_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 VGND B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 VGND A2 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 VGND B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a21boi_4 Y A1 B1_N A2 VGND VPWR VNB VPB
X0 a_223_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A1 a_658_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR B1_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_223_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Y a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND A2 a_658_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_223_297# a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR A2 a_223_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_658_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VPWR A1 a_223_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_223_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_658_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 Y a_27_47# a_223_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_223_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VPWR A2 a_223_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VPWR A1 a_223_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_658_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VGND B1_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_223_297# a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_658_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VGND A2 a_658_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 VGND a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 VGND a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 Y A1 a_658_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 Y a_27_47# a_223_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__xor2_2 VPWR VGND X B A VNB VPB
X0 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_470_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_470_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_112_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_470_47# B X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND A a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_112_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VGND B a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_470_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 X a_112_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VPWR B a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VGND a_112_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VGND A a_470_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_27_297# B a_112_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 X a_112_47# a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_470_297# a_112_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 X B a_470_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_112_47# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor2_4 Y A B VGND VPWR VNB VPB
X0 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__or2_4 X A B VGND VPWR VNB VPB
X0 a_121_297# B a_35_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR a_35_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 X a_35_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_35_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 X a_35_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR a_35_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 X a_35_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR A a_121_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND A a_35_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_35_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor4b_4 B A D_N C Y VGND VPWR VNB VPB
X0 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND D_N a_1191_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_803_297# a_1191_21# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_445_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y a_1191_21# a_803_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_803_297# a_1191_21# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 Y a_1191_21# a_803_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 Y a_1191_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VPWR D_N a_1191_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_27_297# B a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 VGND a_1191_21# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VGND a_1191_21# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 a_445_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 a_803_297# C a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 a_27_297# B a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_445_297# C a_803_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 a_803_297# C a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 Y a_1191_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 a_445_297# C a_803_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or2b_2 A B_N X VPWR VGND VNB VPB
X0 VPWR A a_300_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_218_297# a_27_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND B_N a_27_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_300_297# a_27_53# a_218_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 X a_218_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR a_218_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 X a_218_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND a_218_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_27_53# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VGND A a_218_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o32a_2 B1 B2 A3 A2 A1 X VGND VPWR VNB VPB
X0 a_429_297# A2 a_345_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A2 a_345_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_345_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_345_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_629_297# B2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR B1 a_629_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_79_21# B2 a_345_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_345_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_79_21# A3 a_429_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_345_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or4_4 B C A D X VPWR VGND VNB VPB
X0 VPWR A a_304_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_304_297# B a_220_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND C a_32_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_220_297# C a_114_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_32_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_32_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR a_32_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X a_32_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND A a_32_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR a_32_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 X a_32_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 X a_32_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 X a_32_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_114_297# D a_32_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VGND a_32_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VGND a_32_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 Y B2 VGND VPWR VNB VPB
X0 a_1224_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR A1 a_1224_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_27_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_806_297# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_806_297# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 Y A3 a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_27_47# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_27_47# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 Y A3 a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 a_27_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 a_806_297# A2 a_1224_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 Y B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 VPWR B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 a_1224_297# A2 a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 a_1224_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 a_806_297# A2 a_1224_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 VPWR A1 a_1224_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X36 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X37 a_1224_297# A2 a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 Y B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X39 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor4_4 A C Y D B VGND VPWR VNB VPB
X0 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_807_297# D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y D a_807_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 Y D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_27_297# B a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_449_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_807_297# C a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 VGND D Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 VGND D Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_807_297# C a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_449_297# C a_807_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_449_297# C a_807_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 a_27_297# B a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_807_297# D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_449_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 Y D a_807_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__conb_1 LO HI VPB VNB VGND VPWR
R0 HI VPWR sky130_fd_pr__res_generic_po w=480000u l=45000u
R1 VGND LO sky130_fd_pr__res_generic_po w=480000u l=45000u
.ends

.subckt sky130_fd_sc_hd__or4b_2 C A X B D_N VPWR VGND VNB VPB
X0 a_176_21# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VGND D_N a_27_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND a_176_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 X a_176_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR a_176_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_555_297# C a_483_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_176_21# a_27_53# a_555_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 X a_176_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_387_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_483_297# B a_387_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VGND B a_176_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VGND a_27_53# a_176_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 VPWR D_N a_27_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 a_176_21# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a311o_4 VGND VPWR C1 A1 A2 A3 X B1 VNB VPB
X0 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_277_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_861_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_297# B1 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_1059_47# A2 a_861_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_1059_47# A1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_277_297# B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_27_297# C1 a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND A3 a_861_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND C1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_109_47# A1 a_1059_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_109_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 VPWR A3 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 VPWR A2 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_109_47# C1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR A1 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 a_277_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 a_277_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 a_109_47# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 a_861_47# A2 a_1059_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o211a_4 A1 X C1 A2 B1 VGND VPWR VNB VPB
X0 VGND A1 a_474_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A1 a_1122_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR C1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_950_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_557_47# B1 a_474_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_474_47# B1 a_748_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND A2 a_474_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_79_21# C1 a_557_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_474_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_79_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_748_47# C1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_474_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 VPWR B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_79_21# A2 a_950_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_1122_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or3b_2 A B C_N X VPWR VGND VNB VPB
X0 a_388_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VPWR C_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND a_176_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 X a_176_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR a_176_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND B a_176_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 X a_176_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_176_21# a_27_47# a_472_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_472_297# B a_388_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_176_21# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_176_21# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VGND C_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or3b_4 A B C_N X VGND VPWR VNB VPB
X0 a_176_21# a_27_47# a_626_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_626_297# B a_542_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR C_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VGND a_176_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_542_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR a_176_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 X a_176_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X a_176_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 X a_176_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_176_21# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VPWR a_176_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 X a_176_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_176_21# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND a_176_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VGND B a_176_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VGND C_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or3_2 A B X C VGND VPWR VNB VPB
X0 VPWR a_30_53# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND a_30_53# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X a_30_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_112_297# C a_30_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 X a_30_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND A a_30_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_30_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND C a_30_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_184_297# B a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VPWR A a_184_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__inv_4 Y A VPWR VGND VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a2111o_2 D1 A1 B1 C1 X A2 VGND VPWR VNB VPB
X0 VPWR a_86_235# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND C1 a_86_235# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X a_86_235# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_86_235# D1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 X a_86_235# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_715_47# A1 a_86_235# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND A2 a_715_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_499_297# C1 a_427_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND a_86_235# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_86_235# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_607_297# B1 a_499_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_427_297# D1 a_86_235# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VPWR A1 a_607_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_607_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor2_8 Y A B VGND VPWR VNB VPB
X0 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__or4b_4 D_N B C A X VGND VPWR VNB VPB
X0 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND a_215_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR a_215_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_109_93# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_215_297# a_109_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND C a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND A a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_215_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_109_93# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VPWR A a_487_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND a_215_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_487_297# B a_403_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_403_297# C a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VPWR a_215_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_297_297# a_109_93# a_215_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__o31a_4 X B1 A3 A2 A1 VGND VPWR VNB VPB
X0 VPWR A1 a_926_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A1 a_496_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_926_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND A3 a_496_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND a_102_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND A2 a_496_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_926_297# A2 a_672_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_102_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_496_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 X a_102_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_102_21# B1 a_496_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR a_102_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 X a_102_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 X a_102_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VPWR a_102_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_672_297# A3 a_102_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_496_47# B1 a_102_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_102_21# A3 a_672_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 VGND a_102_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 X a_102_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_496_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VPWR B1 a_102_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_496_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_672_297# A2 a_926_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__a22o_2 A1 A2 X B2 B1 VPWR VGND VNB VPB
X0 VPWR a_27_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A2 a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_27_297# B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_27_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND a_27_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_381_47# A1 a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_109_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and4_2 X C A B D VGND VPWR VNB VPB
X0 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VGND D a_304_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_198_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_304_47# C a_198_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VPWR D a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand3b_2 Y C A_N B VGND VPWR VNB VPB
X0 a_408_47# B a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_408_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y a_27_47# a_408_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VGND C a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_218_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_218_47# B a_408_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__mux2_2 VGND VPWR A1 A0 S X VNB VPB
X0 VPWR S a_591_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 a_591_369# A0 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_79_21# A1 a_306_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND S a_578_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_306_369# a_257_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X7 a_79_21# A0 a_288_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_288_47# a_257_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_257_199# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_578_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_257_199# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X13 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a21o_4 A2 A1 X B1 VGND VPWR VNB VPB
X0 VGND B1 a_84_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_741_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_84_21# A1 a_741_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND A2 a_901_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR a_84_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR A2 a_483_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_483_297# B1 a_84_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X a_84_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_84_21# B1 a_483_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND a_84_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VPWR a_84_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_483_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VPWR A1 a_483_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VGND a_84_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 X a_84_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_84_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_483_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 X a_84_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_901_47# A1 a_84_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 X a_84_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__a32o_2 B2 X A2 A3 A1 B1 VGND VPWR VNB VPB
X0 VPWR A3 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_299_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_352_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_549_47# A1 a_21_199# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 X a_21_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND a_21_199# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_665_47# A2 a_549_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR A1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_299_297# B1 a_21_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_21_199# B2 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VGND A3 a_665_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR a_21_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 X a_21_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_21_199# B1 a_352_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o311a_2 X A2 A3 A1 B1 C1 VPWR VGND VNB VPB
X0 X a_91_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_91_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_360_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR B1 a_91_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_360_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A2 a_360_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_360_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR a_91_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND a_91_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 X a_91_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_677_47# B1 a_360_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_460_297# A2 a_360_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_91_21# C1 a_677_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_91_21# A3 a_460_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_8 A X VGND VPWR VNB VPB
X0 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a2111oi_4 D1 C1 B1 A2 A1 Y VGND VPWR VNB VPB
X0 Y D1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_455_297# B1 a_821_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_28_297# D1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_821_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_28_297# C1 a_455_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_455_297# C1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND D1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR A2 a_821_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 Y D1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND D1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 Y D1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_821_297# B1 a_455_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 Y D1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_1205_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_28_297# C1 a_455_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_1205_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 a_821_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 Y A1 a_1205_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 VPWR A1 a_821_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 Y A1 a_1205_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 a_1205_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X28 a_28_297# D1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VGND A2 a_1205_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 a_455_297# B1 a_821_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 a_821_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 a_1205_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X33 VGND A2 a_1205_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X34 VPWR A1 a_821_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 a_821_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 VPWR A2 a_821_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X37 a_455_297# C1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 a_821_297# B1 a_455_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X39 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o31ai_2 A1 Y B1 A3 A2 VGND VPWR VNB VPB
X0 a_281_297# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_281_297# A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 Y A3 a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_27_297# A2 a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__a41o_2 B1 A1 X A2 A4 A3 VGND VPWR VNB VPB
X0 a_381_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR A2 a_381_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_465_47# A4 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_549_47# A3 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_665_47# A2 a_549_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_381_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR A4 a_381_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_381_297# B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_79_21# A1 a_665_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and4b_2 VPWR VGND X A_N D C B VNB VPB
X0 VPWR a_193_413# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_297_47# a_27_413# a_193_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_369_47# B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X a_193_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR D a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND D a_469_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND a_193_413# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR B a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_193_413# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 X a_193_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_193_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_469_47# C a_369_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a31o_4 B1 A2 A3 A1 X VGND VPWR VNB VPB
X0 VPWR a_277_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X a_277_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 X a_277_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_277_47# B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND a_277_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND a_277_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_193_47# A2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_361_47# A1 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 X a_277_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VGND A3 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 X a_277_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_277_47# A1 a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_445_47# A2 a_361_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VGND B1 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_27_297# B1 a_277_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 VPWR a_277_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_109_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_277_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a2111oi_2 D1 C1 A2 A1 Y B1 VGND VPWR VNB VPB
X0 a_467_297# B1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_287_297# D1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A2 a_467_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_923_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_28_297# B1 a_467_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_28_297# C1 a_287_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Y A1 a_923_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VGND A2 a_684_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y D1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 Y D1 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_467_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VGND D1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VPWR A1 a_467_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_115_297# C1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_467_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_684_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o21bai_2 B1_N Y A2 A1 VGND VPWR VNB VPB
X0 a_397_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR B1_N a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 Y A2 a_397_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND A2 a_229_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND A1 a_229_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_28_297# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 Y a_28_297# a_229_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR a_28_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_397_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_229_47# a_28_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y a_28_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_229_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_229_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VPWR A1 a_397_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__a221oi_4 A2 Y C1 A1 B2 B1 VPWR VGND VNB VPB
X0 Y A1 a_1241_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_453_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y B1 a_453_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y A1 a_1241_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y C1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_471_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y B1 a_453_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND A2 a_1241_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_27_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR A2 a_471_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_453_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_471_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VGND B2 a_453_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_1241_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_27_297# B2 a_471_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_453_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_1241_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_1241_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 VPWR A2 a_471_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 a_471_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 a_471_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 a_471_297# B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 VPWR A1 a_471_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 Y C1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_27_297# B1 a_471_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VGND A2 a_1241_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 a_471_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 a_27_297# B1 a_471_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 a_1241_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X33 a_471_297# B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 VPWR A1 a_471_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 a_27_297# B2 a_471_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 a_471_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X37 a_27_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 a_453_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X39 VGND B2 a_453_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a311o_2 VGND VPWR X C1 B1 A1 A2 A3 VNB VPB
X0 a_79_21# C1 a_635_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR A2 a_319_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_417_47# A2 a_319_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_79_21# A1 a_417_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_319_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_319_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_319_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_79_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_635_297# B1 a_319_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 Y VPWR VGND VNB VPB
X0 a_109_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_467_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_467_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y A1 a_467_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_109_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND A2 a_467_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_27_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VPWR A1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_109_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and3b_2 VGND VPWR B X A_N C VNB VPB
X0 a_109_53# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 X a_215_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_109_53# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VGND C a_373_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VGND a_215_311# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR C a_215_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR a_215_311# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X a_215_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_301_53# a_109_53# a_215_311# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_215_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_373_53# B a_301_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VPWR a_109_53# a_215_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o2bb2a_4 A2_N A1_N X B2 B1 VGND VPWR VNB VPB
X0 a_27_47# a_415_21# a_193_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VPWR A2_N a_415_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_415_21# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_415_21# A2_N a_717_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_193_297# a_415_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR a_193_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X a_193_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_109_297# B2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X a_193_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_717_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_717_47# A2_N a_415_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 X a_193_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_27_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_27_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VGND a_193_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VGND A1_N a_717_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VGND a_193_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 VGND B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_193_297# a_415_21# a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VPWR a_193_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VPWR a_415_21# a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 X a_193_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 VPWR A1_N a_415_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 a_109_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 a_415_21# A2_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 VGND B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor3b_2 C_N Y A B VGND VPWR VNB VPB
X0 a_281_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND a_531_21# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR C_N a_531_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_281_297# a_531_21# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 Y a_531_21# a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND C_N a_531_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_27_297# B a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 Y a_531_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a31oi_2 A3 B1 Y A1 A2 VPWR VGND VNB VPB
X0 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_277_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_27_47# A2 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_277_47# A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 Y A1 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__mux2_8 S A1 VPWR VGND A0 X VNB VPB
X0 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_79_21# A0 a_792_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_1259_199# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_1302_47# A0 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_792_297# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_1259_199# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND a_1259_199# a_1302_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X14 a_79_21# A1 a_792_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X15 a_79_21# A0 a_1302_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X16 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VPWR S a_792_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_792_297# A0 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_1302_47# a_1259_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X23 VPWR a_1259_199# a_1302_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_1302_297# a_1259_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 a_792_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X27 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_1302_297# A1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VGND S a_792_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X30 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 a_79_21# A1 a_1302_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X33 a_792_47# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a31oi_4 Y B1 A1 A3 A2 VPWR VGND VNB VPB
X0 a_27_47# A2 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_27_47# A2 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_445_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_445_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 Y A1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 Y A1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_445_47# A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_445_47# A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X28 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 Y VGND VPWR VNB VPB
X0 a_27_47# C1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_803_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_27_47# C1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND A2 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_1163_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND A2 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Y A2 a_1163_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_1163_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_445_47# B1 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR D1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_445_47# B1 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 Y D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VPWR A1 a_1163_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_27_47# D1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_27_47# D1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VGND A1 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_1163_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_803_47# B1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 VPWR A1 a_1163_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 a_803_47# B1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 Y D1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_445_47# C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 a_803_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 a_1163_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 Y A2 a_1163_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 a_445_47# C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X34 a_803_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X35 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 a_803_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X37 VPWR D1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 Y D1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X39 VGND A1 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a22o_4 B1 B2 X A2 A1 VGND VPWR VNB VPB
X0 a_484_297# B2 a_96_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND B2 a_566_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X a_96_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR a_96_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_96_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_96_21# B1 a_484_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR a_96_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X a_96_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VGND a_96_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_484_297# B1 a_96_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_484_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND A2 a_918_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_96_21# B2 a_484_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_96_21# B1 a_566_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_484_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VPWR A1 a_484_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_96_21# A1 a_918_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VPWR A2 a_484_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_566_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_918_47# A1 a_96_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_566_47# B1 a_96_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 a_918_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 X a_96_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VGND a_96_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand3_4 Y A B C VGND VPWR VNB VPB
X0 a_27_47# B a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_27_47# B a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Y A a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y A a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_27_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_27_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_445_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_445_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND C a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_445_47# B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_445_47# B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VGND C a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 X VGND VPWR VNB VPB
X0 VGND A2 a_393_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_496_297# A4 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_393_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A1 a_697_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND A4 a_393_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_697_297# A2 a_597_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_393_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_393_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_597_297# A3 a_496_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 X VPWR VGND VNB VPB
X0 X a_80_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_475_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X a_80_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_762_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_475_47# B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND A2 a_475_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X a_80_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_80_21# A2 a_762_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_80_21# B1 a_475_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_80_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_475_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 X a_80_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VPWR A1 a_934_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_934_297# A2 a_80_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VPWR B1 a_80_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND A1 a_475_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o21ba_2 B1_N A1 X A2 VGND VPWR VNB VPB
X0 VGND B1_N a_27_93# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VGND A2 a_478_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_478_47# a_27_93# a_174_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_478_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 X a_174_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR a_174_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 X a_174_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR A1 a_574_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND a_174_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR B1_N a_27_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_574_297# A2 a_174_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_174_21# a_27_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_12 A X VGND VPWR VNB VPB
X0 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR A a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_109_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VPWR A a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND A a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VGND A a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_109_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_109_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 a_109_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a221o_4 A1 B1 C1 B2 X A2 VPWR VGND VNB VPB
X0 VGND A2 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VGND B2 a_1053_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_804_297# B1 a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_79_21# A1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_445_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_804_297# C1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_445_297# B1 a_804_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_1053_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_79_21# C1 a_804_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_1053_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_445_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND C1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_804_297# B2 a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_79_21# B1 a_1053_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_79_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_445_297# B2 a_804_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 a_445_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_445_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 VPWR A2 a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 VPWR A1 a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and3_4 A B C X VGND VPWR VNB VPB
X0 VPWR A a_94_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_294_47# B a_185_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_185_47# A a_94_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR a_94_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND C a_294_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_94_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 X a_94_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X a_94_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR C a_94_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X a_94_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND a_94_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR a_94_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND a_94_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 X a_94_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__and4bb_4 C A_N D X B_N VGND VPWR VNB VPB
X0 VPWR a_174_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_174_21# a_832_21# a_766_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X a_174_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_832_21# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_766_47# a_27_47# a_652_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR a_174_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 X a_174_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR B_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_652_47# C a_556_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_832_21# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 X a_174_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 X a_174_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_556_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_174_21# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VPWR C a_174_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND a_174_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VGND a_174_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VPWR a_832_21# a_174_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_174_21# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND B_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a41o_4 X A4 A3 A2 A1 B1 VGND VPWR VNB VPB
X0 a_639_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_639_47# A2 a_889_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A3 a_467_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_889_47# A2 a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_889_47# A3 a_1079_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_467_297# A4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_467_297# B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_467_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VPWR A4 a_467_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_1079_47# A3 a_889_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_79_21# B1 a_467_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_79_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_1079_47# A4 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 VPWR A2 a_467_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 a_467_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_79_21# A1 a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 VPWR A1 a_467_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 a_467_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 VGND A4 a_1079_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand4_4 A D C B Y VPWR VGND VNB VPB
X0 a_27_47# C a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_27_47# C a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_445_47# B a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_445_47# B a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_27_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_27_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 Y A a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 Y A a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_803_47# B a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_803_47# B a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VGND D a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_445_47# C a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_803_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 a_445_47# C a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_803_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 VGND D a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VPWR VPB VNB
D0 VNB DIODE sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06u area=4.347e+11p
.ends

.subckt sky130_fd_sc_hd__nor3_4 A C B Y VGND VPWR VNB VPB
X0 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_449_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_27_297# B a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y C a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_449_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y C a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_449_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_27_297# B a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 a_449_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__or2b_4 A B_N X VGND VPWR VNB VPB
X0 VPWR a_219_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND B_N a_27_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VPWR A a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_27_53# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 X a_219_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_301_297# a_27_53# a_219_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 X a_219_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND A a_219_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR a_219_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND a_219_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 X a_219_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND a_219_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_219_297# a_27_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 X a_219_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt adc_core_digital VGND VPWR clk_dig_in comparator_in config_1_in[0] config_1_in[10]
+ config_1_in[11] config_1_in[12] config_1_in[13] config_1_in[14] config_1_in[15]
+ config_1_in[1] config_1_in[2] config_1_in[3] config_1_in[4] config_1_in[5] config_1_in[6]
+ config_1_in[7] config_1_in[8] config_1_in[9] config_2_in[0] config_2_in[10] config_2_in[11]
+ config_2_in[12] config_2_in[13] config_2_in[14] config_2_in[15] config_2_in[1] config_2_in[2]
+ config_2_in[3] config_2_in[4] config_2_in[5] config_2_in[6] config_2_in[7] config_2_in[8]
+ config_2_in[9] conv_finished_out enable_loop_out nmatrix_bincap_out_n[0] nmatrix_bincap_out_n[1]
+ nmatrix_bincap_out_n[2] nmatrix_c0_out_n nmatrix_col_out_n[0] nmatrix_col_out_n[10]
+ nmatrix_col_out_n[11] nmatrix_col_out_n[12] nmatrix_col_out_n[13] nmatrix_col_out_n[14]
+ nmatrix_col_out_n[15] nmatrix_col_out_n[16] nmatrix_col_out_n[17] nmatrix_col_out_n[18]
+ nmatrix_col_out_n[19] nmatrix_col_out_n[1] nmatrix_col_out_n[20] nmatrix_col_out_n[21]
+ nmatrix_col_out_n[22] nmatrix_col_out_n[23] nmatrix_col_out_n[24] nmatrix_col_out_n[25]
+ nmatrix_col_out_n[26] nmatrix_col_out_n[27] nmatrix_col_out_n[28] nmatrix_col_out_n[29]
+ nmatrix_col_out_n[2] nmatrix_col_out_n[30] nmatrix_col_out_n[31] nmatrix_col_out_n[3]
+ nmatrix_col_out_n[4] nmatrix_col_out_n[5] nmatrix_col_out_n[6] nmatrix_col_out_n[7]
+ nmatrix_col_out_n[8] nmatrix_col_out_n[9] nmatrix_row_out_n[0] nmatrix_row_out_n[10]
+ nmatrix_row_out_n[11] nmatrix_row_out_n[12] nmatrix_row_out_n[13] nmatrix_row_out_n[14]
+ nmatrix_row_out_n[15] nmatrix_row_out_n[1] nmatrix_row_out_n[2] nmatrix_row_out_n[3]
+ nmatrix_row_out_n[4] nmatrix_row_out_n[5] nmatrix_row_out_n[6] nmatrix_row_out_n[7]
+ nmatrix_row_out_n[8] nmatrix_row_out_n[9] nmatrix_rowon_out_n[0] nmatrix_rowon_out_n[10]
+ nmatrix_rowon_out_n[11] nmatrix_rowon_out_n[12] nmatrix_rowon_out_n[13] nmatrix_rowon_out_n[14]
+ nmatrix_rowon_out_n[15] nmatrix_rowon_out_n[1] nmatrix_rowon_out_n[2] nmatrix_rowon_out_n[3]
+ nmatrix_rowon_out_n[4] nmatrix_rowon_out_n[5] nmatrix_rowon_out_n[6] nmatrix_rowon_out_n[7]
+ nmatrix_rowon_out_n[8] nmatrix_rowon_out_n[9] pmatrix_bincap_out_n[0] pmatrix_bincap_out_n[1]
+ pmatrix_bincap_out_n[2] pmatrix_c0_out_n pmatrix_col_out_n[0] pmatrix_col_out_n[10]
+ pmatrix_col_out_n[11] pmatrix_col_out_n[12] pmatrix_col_out_n[13] pmatrix_col_out_n[14]
+ pmatrix_col_out_n[15] pmatrix_col_out_n[16] pmatrix_col_out_n[17] pmatrix_col_out_n[18]
+ pmatrix_col_out_n[19] pmatrix_col_out_n[1] pmatrix_col_out_n[20] pmatrix_col_out_n[21]
+ pmatrix_col_out_n[22] pmatrix_col_out_n[23] pmatrix_col_out_n[24] pmatrix_col_out_n[25]
+ pmatrix_col_out_n[26] pmatrix_col_out_n[27] pmatrix_col_out_n[28] pmatrix_col_out_n[29]
+ pmatrix_col_out_n[2] pmatrix_col_out_n[30] pmatrix_col_out_n[31] pmatrix_col_out_n[3]
+ pmatrix_col_out_n[4] pmatrix_col_out_n[5] pmatrix_col_out_n[6] pmatrix_col_out_n[7]
+ pmatrix_col_out_n[8] pmatrix_col_out_n[9] pmatrix_row_out_n[0] pmatrix_row_out_n[10]
+ pmatrix_row_out_n[11] pmatrix_row_out_n[12] pmatrix_row_out_n[13] pmatrix_row_out_n[14]
+ pmatrix_row_out_n[15] pmatrix_row_out_n[1] pmatrix_row_out_n[2] pmatrix_row_out_n[3]
+ pmatrix_row_out_n[4] pmatrix_row_out_n[5] pmatrix_row_out_n[6] pmatrix_row_out_n[7]
+ pmatrix_row_out_n[8] pmatrix_row_out_n[9] pmatrix_rowon_out_n[0] pmatrix_rowon_out_n[10]
+ pmatrix_rowon_out_n[11] pmatrix_rowon_out_n[12] pmatrix_rowon_out_n[13] pmatrix_rowon_out_n[14]
+ pmatrix_rowon_out_n[15] pmatrix_rowon_out_n[1] pmatrix_rowon_out_n[2] pmatrix_rowon_out_n[3]
+ pmatrix_rowon_out_n[4] pmatrix_rowon_out_n[5] pmatrix_rowon_out_n[6] pmatrix_rowon_out_n[7]
+ pmatrix_rowon_out_n[8] pmatrix_rowon_out_n[9] result_out[0] result_out[10] result_out[11]
+ result_out[12] result_out[13] result_out[14] result_out[15] result_out[1] result_out[2]
+ result_out[3] result_out[4] result_out[5] result_out[6] result_out[7] result_out[8]
+ result_out[9] rst_n sample_matrix_out sample_matrix_out_n sample_switch_out sample_switch_out_n
XFILLER_45_258 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_144 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_73 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_67 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1270_ _1270_/Y _1276_/C _1270_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
XFILLER_36_214 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1606_ _1601_/X _1742_/D _1604_/Y _1605_/X _1604_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__o2bb2a_2
X_0985_ _1151_/B _1117_/S _1116_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__xnor2_4
X_1399_ _1770_/Q _1407_/A _1724_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
X_1537_ VGND VPWR _1706_/D _1537_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1468_ _1803_/A _1777_/A _1501_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_27_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_10 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_280 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0770_ _1420_/A _1602_/B _0768_/X _1689_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__o21ai_4
X_1322_ _1718_/Q _1328_/A _1764_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
X_1253_ _1132_/X _1253_/Y _1270_/B _1287_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__o21ai_2
X_1184_ VPWR VGND _1205_/A _1185_/A _1184_/B VGND VPWR sky130_fd_sc_hd__and2_2
X_0968_ _0968_/X _1062_/B _0916_/B _1671_/Q _0916_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__o31a_2
X_0899_ _0899_/C _0908_/B _0912_/A _0899_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nor3_2
XFILLER_0_79 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_66 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0822_ VGND VPWR _0823_/B _1750_/Q _1749_/Q VGND VPWR sky130_fd_sc_hd__xnor2_2
X_1305_ _1306_/B _1713_/Q _1410_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1236_ _1255_/A _1243_/A _1129_/X _1235_/Y _1236_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__o211ai_4
X_1167_ VPWR VGND _1221_/A _1276_/B VGND VPWR sky130_fd_sc_hd__buf_4
X_1098_ _1098_/X _1097_/X _1087_/X _1067_/X _1096_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_2
XFILLER_34_74 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_95 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1021_ _1033_/B _0908_/D _1076_/A _0925_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o21bai_4
X_1785_ VGND VPWR _1785_/X _1785_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_0805_ VGND VPWR _1754_/D input2/X _0805_/B VGND VPWR sky130_fd_sc_hd__xnor2_2
X_1219_ _1219_/B _1219_/Y _1219_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_37_183 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_293 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1570_ VGND VPWR _1626_/S _1718_/D _1716_/D _1570_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_1004_ VPWR VGND _1004_/A _1038_/B _1004_/B VGND VPWR sky130_fd_sc_hd__and2_2
X_1768_ _1768_/Q fanout176/X _1768_/D _1770_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1699_ _1699_/Q fanout178/X _1699_/D _1758_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_40_123 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xoutput31 VPWR VGND nmatrix_col_out_n[24] _1294_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput42 VPWR VGND nmatrix_col_out_n[5] _1262_/Y VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput75 VPWR VGND nmatrix_rowon_out_n[8] _1785_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput64 VPWR VGND nmatrix_rowon_out_n[11] _1788_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput20 VPWR VGND nmatrix_col_out_n[14] _1278_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput53 VPWR VGND nmatrix_row_out_n[1] _1777_/A VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput86 VPWR VGND pmatrix_col_out_n[15] _1204_/Y VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_48_289 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xoutput97 VPWR VGND pmatrix_col_out_n[25] _1236_/Y VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_16_186 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1622_ _1569_/B _1622_/X _1621_/X _1729_/D _1604_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__o22a_2
X_1553_ _1615_/C _1565_/A _1604_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1484_ _1797_/A _1786_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_22_156 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_178 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_57 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_226 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0984_ _0983_/X _0981_/X _0973_/X _1117_/S VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_4
X_1605_ _1569_/B _1720_/D _1605_/X _1726_/D _1563_/X _1620_/A VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__o221a_2
X_1536_ VGND VPWR _1542_/S _1706_/Q _1707_/Q _1537_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_1398_ _1401_/B _1724_/Q _1770_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1467_ _1467_/A _1487_/B _1803_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_8
XFILLER_37_52 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_240 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1321_ _1717_/D _1321_/B _1763_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__xnor2_4
X_1252_ _1265_/B _1252_/X _1252_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
X_1183_ VPWR VGND _1183_/X _1183_/A VGND VPWR sky130_fd_sc_hd__buf_4
X_0967_ VPWR VGND _1116_/A _0967_/A VGND VPWR sky130_fd_sc_hd__buf_6
X_0898_ VGND VPWR _1699_/Q _0897_/X _0896_/Y _0899_/C VGND VPWR sky130_fd_sc_hd__mux2_1
X_1519_ _1663_/B _1542_/S _1697_/D _1697_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__a21bo_2
XFILLER_23_10 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_188 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_295 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0821_ _1749_/D _1749_/Q _1542_/S VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
XFILLER_43_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1304_ _1410_/B _1420_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_6
X_1235_ _1235_/Y _1270_/B _1255_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1166_ _1166_/X _1255_/B _1255_/A _1164_/X _1256_/A VGND VPWR _1165_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_2
X_1097_ VPWR VGND _1097_/X _1487_/A _1680_/Q VGND VPWR sky130_fd_sc_hd__and2b_2
XFILLER_34_20 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_41 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_64 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1020_ _1677_/Q _1050_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
X_1784_ VPWR VGND _1784_/X _1784_/A VGND VPWR sky130_fd_sc_hd__buf_2
X_0804_ _0805_/B _1754_/Q _1542_/S VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1218_ _1219_/B _1471_/A _1265_/A _1221_/A _1152_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__o31a_2
X_1149_ _1149_/X _1140_/X _1217_/A _1255_/B _1255_/A VGND VPWR _1148_/Y VGND VPWR
+ sky130_fd_sc_hd__a221o_2
XFILLER_43_132 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_261 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1003_ _1016_/A _1035_/B _1676_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__xnor2_4
XFILLER_22_305 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1767_ _1767_/Q fanout176/X _1767_/D _1770_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1698_ _1698_/Q fanout179/X _1698_/D _1766_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_31_32 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xoutput54 VPWR VGND nmatrix_row_out_n[2] _1778_/A VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_0_220 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xoutput43 VPWR VGND nmatrix_col_out_n[6] _1264_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput10 VPWR VGND conv_finished_out _1463_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput21 VPWR VGND nmatrix_col_out_n[15] _1279_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput32 VPWR VGND nmatrix_col_out_n[25] _1295_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput65 VPWR VGND nmatrix_rowon_out_n[12] _1789_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput76 VPWR VGND nmatrix_rowon_out_n[9] _1786_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput87 VPWR VGND pmatrix_col_out_n[16] _1207_/Y VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput98 VPWR VGND pmatrix_col_out_n[26] _1238_/X VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_48_246 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1552_ _1584_/S _1558_/B _1604_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_8
X_1621_ VGND VPWR _1626_/S _1727_/D _1725_/D _1621_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_1483_ _1784_/A _1487_/B _1496_/A _1797_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_39_235 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_10 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_43 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_0983_ _0983_/X _0948_/X _1672_/Q _0980_/C _0975_/A VGND VPWR _0982_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_2
X_1604_ _1604_/B _1604_/Y _1604_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1535_ VGND VPWR _1705_/D _1535_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1397_ _1593_/A _1724_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
X_1466_ _1487_/B _1466_/B _1680_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__xor2_4
XFILLER_12_78 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_75 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_42 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1320_ _1321_/B _1410_/B _1319_/X _1318_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__o21ai_4
X_1251_ _1124_/X _1255_/B _1140_/X _1251_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_4
X_1182_ VPWR VGND _1205_/A _1183_/A _1287_/B VGND VPWR sky130_fd_sc_hd__and2_2
X_0966_ _0993_/B _0967_/A _0993_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
X_0897_ _1703_/Q _0897_/X _1701_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
XFILLER_32_285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1449_ _1449_/B _1449_/X _1691_/Q _1451_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
X_1518_ VPWR VGND _1663_/B _1665_/S VGND VPWR sky130_fd_sc_hd__buf_4
X_0820_ _0818_/Y _1542_/S _0819_/X _1758_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__o21a_2
X_1303_ _1233_/A _1203_/X _1255_/B _1303_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_2
X_1234_ _1234_/Y _1234_/A _1243_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1165_ _1265_/A _1165_/X _1276_/C _1258_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
X_1096_ _1096_/X _1093_/X _1090_/X _1092_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
X_0949_ _0974_/B _0949_/Y _0980_/C _0975_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor3_2
XFILLER_7_237 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1783_ VGND VPWR _1783_/X _1783_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_0803_ VPWR VGND _1542_/S _1546_/S VGND VPWR sky130_fd_sc_hd__buf_6
X_1217_ _1217_/B _1219_/A _1217_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1148_ _1178_/B _1237_/B _1144_/X _1148_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_2
X_1079_ VGND VPWR _1035_/B _1677_/Q _1048_/B _1079_/X _1035_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_2
XFILLER_20_56 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_10 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_185 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_155 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1002_ _1076_/A _0925_/X _1035_/B _0929_/C _0915_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__o22a_4
X_1766_ _1766_/Q fanout173/X _1766_/D _1766_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1697_ _1697_/Q fanout179/X _1697_/D _1766_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_31_44 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xoutput55 VPWR VGND nmatrix_row_out_n[3] _1779_/A VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput44 VPWR VGND nmatrix_col_out_n[7] _1266_/X VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_0_276 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xoutput99 VPWR VGND pmatrix_col_out_n[27] _1241_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput66 VPWR VGND nmatrix_rowon_out_n[13] _1790_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput11 VPWR VGND enable_loop_out _1809_/A VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput88 VPWR VGND pmatrix_col_out_n[17] _1212_/Y VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput77 VPWR VGND pmatrix_bincap_out_n[0] _0879_/A VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput33 VPWR VGND nmatrix_col_out_n[26] _1296_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput22 VPWR VGND nmatrix_col_out_n[16] _1280_/X VGND VPWR sky130_fd_sc_hd__buf_4
X_1482_ _1798_/A _1785_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
X_1620_ _1723_/D _1620_/X _1620_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
X_1551_ _1551_/Y _1733_/Q _1596_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
XFILLER_22_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_191 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1749_ _1749_/Q _1749_/D VPWR fanout178/X _1765_/CLK VGND VGND VPWR sky130_fd_sc_hd__dfstp_4
XFILLER_26_22 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_107 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_10 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0982_ _1672_/Q _0980_/D _0974_/B _0980_/C _0982_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o211a_2
X_1603_ _1604_/B _1602_/Y _1615_/A _1742_/Q _1596_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_2
X_1534_ VGND VPWR _1538_/S _1706_/Q _0989_/A _1535_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_1465_ _1497_/A _1501_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
X_1396_ _1593_/A _1396_/B _1770_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__xnor2_4
XFILLER_50_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_10 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1181_ _1175_/X _1140_/X _1181_/Y _1129_/X _1144_/X _1179_/Y VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__o221ai_2
X_1250_ _1237_/A _1233_/A _1129_/X _1250_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o21a_2
X_0965_ _0993_/B _0989_/A _1013_/B _1014_/B _1007_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__o31a_2
X_0896_ VGND VPWR _0896_/Y _1701_/Q _1703_/Q VGND VPWR sky130_fd_sc_hd__xnor2_2
X_1448_ _1449_/B _1451_/C _1691_/Q _1448_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_2
X_1517_ _1665_/S _1698_/Q _1524_/S VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_4
X_1379_ _1768_/Q _1385_/A _1722_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
XFILLER_46_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_264 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1302_ _1302_/X _1203_/X _1248_/X _1221_/B _1301_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__a211o_2
X_1233_ _1243_/A _1233_/A _1256_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_4
X_1164_ VPWR VGND _1164_/X _1164_/A VGND VPWR sky130_fd_sc_hd__buf_4
X_1095_ _1094_/Y _1083_/B _1095_/X _1088_/Y _1487_/A _1083_/A VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__o221a_2
XFILLER_20_278 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0948_ _0974_/B _0948_/X _0975_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
X_0879_ _0879_/A _0879_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_18_67 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_249 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0802_ VPWR VGND _1546_/S _0887_/B _1524_/S VGND VPWR sky130_fd_sc_hd__and2b_2
X_1782_ VGND VPWR _1782_/X _1782_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1216_ _1221_/A _1471_/A _1273_/A _1217_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_2
XFILLER_29_109 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1147_ VPWR VGND _1178_/B _1287_/B VGND VPWR sky130_fd_sc_hd__buf_6
X_1078_ _1078_/B _1078_/Y _1078_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_28_197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_10 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1001_ _1676_/Q _1035_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_34_167 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1765_ _1765_/Q fanout178/X _1765_/D _1765_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1696_ _1808_/A _1696_/D VPWR fanout172/X _1765_/CLK VGND VGND VPWR sky130_fd_sc_hd__dfstp_4
XFILLER_15_68 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_104 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xoutput23 VPWR VGND nmatrix_col_out_n[17] _1282_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput34 VPWR VGND nmatrix_col_out_n[27] _1297_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput12 VPWR VGND nmatrix_bincap_out_n[0] _0879_/Y VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput67 VPWR VGND nmatrix_rowon_out_n[14] _1791_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput45 VPWR VGND nmatrix_col_out_n[8] _1267_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput89 VPWR VGND pmatrix_col_out_n[18] _1215_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput78 VPWR VGND pmatrix_bincap_out_n[1] _0920_/A VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput56 VPWR VGND nmatrix_row_out_n[4] _1780_/A VGND VPWR sky130_fd_sc_hd__buf_4
X_1550_ VPWR VGND _1596_/C _1615_/A VGND VPWR sky130_fd_sc_hd__buf_4
X_1481_ _1784_/A _1487_/B _1497_/A _1798_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_47_281 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1748_ _1748_/Q fanout170/X _1748_/D _1748_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1679_ _1679_/Q fanout175/X _1679_/D _1769_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_26_67 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_22 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0981_ VGND VPWR _0980_/X _0979_/X _0981_/X _0975_/Y _0974_/X VGND VPWR sky130_fd_sc_hd__a211o_4
X_1602_ _1602_/B _1602_/Y _1602_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1464_ _1497_/A _1496_/A _1471_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__and2_4
X_1395_ _1393_/Y _1410_/B _1394_/X _1396_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__o21a_2
X_1533_ VGND VPWR _1704_/D _1533_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_35_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_265 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_295 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_276 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1180_ _1179_/Y _1180_/Y _1175_/X _1173_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__o21ai_2
X_0964_ _0964_/C _1013_/A _1007_/B _1013_/C _0964_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_2
X_1516_ _1696_/D _1682_/D _1507_/S _1542_/S VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
X_0895_ _1697_/Q _1698_/Q _0899_/B _1700_/Q _1808_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_2
X_1447_ _1692_/Q _1449_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
X_1378_ _1767_/Q _1381_/B _1721_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
XFILLER_23_79 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_232 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1232_ _1255_/B _1234_/A _1270_/B _1173_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__o21ai_2
X_1301_ _1301_/X _1276_/B _1246_/B _1255_/A _1246_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__o31a_2
X_1163_ _1246_/C _1164_/A _1246_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
X_1094_ _1093_/X _1092_/Y _1090_/X _1094_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_2
X_0947_ _0946_/X _0944_/X _0859_/B _0974_/B _1013_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__a211oi_4
X_0878_ _0919_/A _0879_/A _0878_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_7_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_305 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1781_ VGND VPWR _1781_/X _1781_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_0801_ _1699_/Q _0887_/B _1698_/Q _0946_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or3_4
X_1215_ _1215_/X _1214_/Y _1140_/X _1287_/A _1213_/Y VGND VPWR _1255_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_2
XFILLER_37_143 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1146_ _1258_/A _1158_/B _1158_/A _1237_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_4
X_1077_ _1078_/B _1076_/X _1035_/B _1035_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_4_209 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_154 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1000_ _1809_/A _0999_/X _1261_/C _1070_/A _1675_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__o211a_2
X_1764_ _1764_/Q fanout173/X _1764_/D _1765_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1695_ _1695_/Q fanout170/X _1695_/D _1748_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1129_ VPWR VGND _1129_/X _1129_/A VGND VPWR sky130_fd_sc_hd__buf_6
XFILLER_31_24 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xoutput24 VPWR VGND nmatrix_col_out_n[18] _1283_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput57 VPWR VGND nmatrix_row_out_n[5] _1781_/A VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput13 VPWR VGND nmatrix_bincap_out_n[1] _0920_/Y VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput46 VPWR VGND nmatrix_col_out_n[9] _1269_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput35 VPWR VGND nmatrix_col_out_n[28] _1298_/X VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_48_238 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xoutput68 VPWR VGND nmatrix_rowon_out_n[1] _1778_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput79 VPWR VGND pmatrix_bincap_out_n[2] _0939_/A VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_8_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1480_ _1800_/A _1783_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_47_293 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_260 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1747_ _1747_/Q fanout177/X _1747_/D _1462_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1678_ _1678_/Q fanout175/X _1678_/D _1769_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_45_219 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0980_ VGND VPWR _1672_/Q _0980_/C _0974_/B _0980_/X _0980_/D VGND VPWR sky130_fd_sc_hd__and4bb_2
XFILLER_8_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1601_ VGND VPWR _1626_/S _1593_/A _1376_/A _1601_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_1532_ VGND VPWR _1542_/S _1012_/B _0989_/A _1533_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_1463_ VGND VPWR _1463_/X _1463_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1394_ _1394_/B _1394_/X _1724_/Q _1394_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
XFILLER_50_222 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_277 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_123 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_0963_ VGND VPWR _0964_/D _1012_/B _1708_/Q VGND VPWR sky130_fd_sc_hd__xnor2_2
X_0894_ _1809_/A _1808_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_6
X_1515_ VGND VPWR _1686_/D _1515_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1446_ _1446_/B _1691_/D _1683_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1377_ _1381_/A _1721_/Q _1767_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
XFILLER_0_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_49 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1231_ VGND VPWR _1231_/X _1231_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1162_ _1157_/Y _1162_/X _1161_/Y _1256_/A _1132_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o22a_2
X_1300_ _1246_/X _1240_/X _1233_/A _1299_/Y _1300_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a22oi_4
X_1093_ _1093_/B _1093_/X _1093_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
XFILLER_9_281 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0946_ _0946_/A _0946_/X _1073_/B _0946_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__or3_4
X_0877_ _0919_/A _0873_/X _1670_/Q _0876_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__a21boi_4
X_1429_ VPWR VGND _1430_/B _1429_/B _1731_/Q VGND VPWR sky130_fd_sc_hd__xor2_2
XFILLER_28_303 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_35 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_303 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_314 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_177 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1780_ VGND VPWR _1780_/X _1780_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_0800_ _1701_/Q _0946_/A _1700_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
X_1214_ _1214_/Y _1276_/C _1237_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1145_ _1258_/A _1151_/A _1151_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_4
X_1076_ _1076_/X _1076_/A _1076_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__or2_4
X_0929_ _1073_/A _1706_/Q _1707_/Q _0929_/C _0975_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor4b_4
XFILLER_6_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_210 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_136 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1694_ _1694_/Q fanout174/X _1694_/D _1745_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1763_ _1763_/Q fanout179/X _1763_/D _1763_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1128_ _1130_/A _1129_/A _1151_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
X_1059_ _1064_/A _1059_/B _1679_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__xor2_4
XFILLER_33_191 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xoutput14 VPWR VGND nmatrix_bincap_out_n[2] _0939_/Y VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput25 VPWR VGND nmatrix_col_out_n[19] _1284_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput47 VPWR VGND nmatrix_row_out_n[10] _1786_/A VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput36 VPWR VGND nmatrix_col_out_n[29] _1300_/Y VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput69 VPWR VGND nmatrix_rowon_out_n[2] _1779_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput58 VPWR VGND nmatrix_row_out_n[6] _1782_/A VGND VPWR sky130_fd_sc_hd__buf_4
XPHY_0 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_272 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1746_ _1746_/Q fanout176/X _1746_/D _1746_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1677_ _1677_/Q fanout181/X _1677_/D _1769_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_53_220 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_305 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_80 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1462_ VPWR VGND _1462_/A _1463_/A _1683_/Q VGND VPWR sky130_fd_sc_hd__and2_2
X_1600_ _1741_/D _1640_/B _1763_/Q _1596_/X _1599_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__a211o_2
X_1531_ VGND VPWR _1703_/D _1531_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1393_ _1724_/Q _1394_/C _1394_/B _1393_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_2
XFILLER_50_234 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_220 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1729_ _1729_/Q fanout174/X _1729_/D _1745_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_53_23 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0962_ _1073_/A _0961_/X _0959_/X _0993_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_4
X_0893_ _1808_/A _0892_/X _0890_/X _1670_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_2
X_1445_ VGND VPWR _1446_/B _1691_/Q _1451_/C VGND VPWR sky130_fd_sc_hd__xnor2_2
X_1514_ VGND VPWR _1514_/S input8/X _1686_/Q _1515_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_1376_ _1376_/A _1722_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_2_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1161_ _1237_/A _1198_/B _1265_/A _1161_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_2
X_1230_ _1230_/A _1229_/X _1231_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or2b_2
XFILLER_49_142 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1092_ _1116_/B _1092_/Y _1061_/C _1116_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__o21ai_2
XFILLER_20_204 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_293 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0876_ _0875_/X _0849_/A _0874_/X _0859_/D _1073_/A _0876_/X VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__o32a_2
X_0945_ VGND VPWR _0946_/C _1703_/Q _1702_/Q VGND VPWR sky130_fd_sc_hd__xnor2_2
X_1428_ _1429_/B _1730_/Q _1428_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1359_ _1402_/C _1359_/X _1717_/Q _1402_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
XFILLER_11_237 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1213_ _1471_/A _1213_/Y _1276_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1144_ VPWR VGND _1144_/X _1276_/B VGND VPWR sky130_fd_sc_hd__buf_6
X_1075_ _1093_/A _1083_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
X_0859_ _0859_/B _0859_/C _1073_/A _0859_/D _0859_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_4
X_0928_ _1013_/C _0912_/A _0923_/X _0927_/X _0980_/D _1076_/A VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__o32ai_4
XFILLER_34_104 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_181 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1693_ _1693_/Q fanout171/X _1693_/D _1742_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1762_ _1762_/Q fanout179/X _1762_/D _1766_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1058_ _1058_/A _1058_/C _1059_/B _1058_/D _1058_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nor4_4
X_1127_ _1151_/A _1127_/B _1127_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__xnor2_4
Xoutput48 VPWR VGND nmatrix_row_out_n[11] _1787_/A VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput26 VPWR VGND nmatrix_col_out_n[1] _1251_/Y VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput15 VPWR VGND nmatrix_col_out_n[0] _1250_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput37 VPWR VGND nmatrix_col_out_n[2] _1254_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput59 VPWR VGND nmatrix_row_out_n[7] _1783_/A VGND VPWR sky130_fd_sc_hd__buf_4
XPHY_1 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1745_ _1745_/Q fanout174/X _1745_/D _1745_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1676_ _1676_/Q fanout181/X _1676_/D _1769_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_38_262 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xadc_core_digital_191 nmatrix_c0_out_n adc_core_digital_191/HI VPWR VGND VGND VPWR
+ sky130_fd_sc_hd__conb_1
XFILLER_53_276 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1461_ VGND VPWR _1682_/D _1461_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1392_ _1394_/C _1769_/Q _1392_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1530_ VGND VPWR _1538_/S _1012_/B _1703_/Q _1531_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_50_246 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1728_ _1728_/Q fanout174/X _1728_/D _1745_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_12_39 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1659_ VGND VPWR _1665_/S _1767_/Q _1678_/D _1660_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_232 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_0961_ _1007_/A _1026_/B _0961_/X _0964_/C _1012_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__or4b_2
X_0892_ _0892_/X _0876_/X _0873_/X _1070_/A _1670_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__a211o_2
X_1444_ VPWR VGND _1690_/Q _1451_/C _1444_/B VGND VPWR sky130_fd_sc_hd__and2_2
X_1513_ VGND VPWR _1685_/D _1513_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1375_ _1376_/A _1375_/B _1768_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__xnor2_4
X_1091_ VGND VPWR _1079_/X _1078_/A _1078_/B _1116_/B _1076_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_2
X_1160_ _1198_/B _1151_/A _1138_/A _1138_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
XFILLER_9_261 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0944_ _1013_/A _0944_/X _1013_/B _0944_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__or3_4
X_0875_ _0875_/C _1073_/C _0875_/X _1005_/B _0875_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_2
X_1427_ _1427_/B _1730_/D _1514_/S VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1358_ _1358_/X _1717_/Q _1402_/C _1402_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
X_1289_ VGND VPWR _1288_/X _1151_/A _1151_/B _1221_/B _1289_/X _1219_/A VGND VPWR
+ sky130_fd_sc_hd__a311o_4
XFILLER_11_249 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1212_ _1212_/Y _1211_/Y _1209_/X _1129_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o21ai_4
X_1143_ VPWR VGND _1255_/B _1143_/A VGND VPWR sky130_fd_sc_hd__buf_6
X_1074_ VGND VPWR _1712_/Q _1085_/C _1058_/B _1093_/A _1074_/D VGND VPWR sky130_fd_sc_hd__and4bb_2
X_0927_ _1084_/A _0927_/X _0926_/X _0924_/Y _0925_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o211a_4
X_0858_ _0858_/B _0859_/D _0989_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_0789_ _1667_/Q _1668_/Q _1669_/Q _0789_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__or3b_2
XFILLER_29_37 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1761_ _1761_/Q fanout181/X _1761_/D _1769_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1692_ _1692_/Q fanout171/X _1692_/D _1748_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1126_ VPWR VGND _1237_/A _1126_/A VGND VPWR sky130_fd_sc_hd__buf_6
X_1057_ _1809_/A _1056_/X _1287_/B _1070_/A _1678_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__o211a_2
Xoutput38 VPWR VGND nmatrix_col_out_n[30] _1302_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput49 VPWR VGND nmatrix_row_out_n[12] _1788_/A VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput16 VPWR VGND nmatrix_col_out_n[10] _1271_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput27 VPWR VGND nmatrix_col_out_n[20] _1286_/X VGND VPWR sky130_fd_sc_hd__buf_4
XPHY_100 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_182 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_2 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1744_ _1744_/Q fanout175/X _1744_/D _1746_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_30_141 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1675_ _1675_/Q fanout181/X _1675_/D _1769_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
Xadc_core_digital_192 nmatrix_row_out_n[0] adc_core_digital_192/HI VPWR VGND VGND
+ VPWR sky130_fd_sc_hd__conb_1
X_1109_ _1116_/A _1117_/S _1108_/X _1111_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__or3b_4
XFILLER_44_299 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1391_ _1723_/Q _1394_/B _1392_/B _1769_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__o21ai_2
X_1460_ VPWR VGND _1697_/Q _1461_/A _1548_/S VGND VPWR sky130_fd_sc_hd__and2_2
X_1727_ _1727_/Q fanout174/X _1727_/D _1745_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1658_ VGND VPWR _1766_/D _1658_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1589_ _1589_/X _1588_/X _1596_/C _1739_/Q _1596_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_2
X_0960_ _0989_/A _1014_/B _1007_/A _1013_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__or3_2
XFILLER_32_247 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1512_ VGND VPWR _1514_/S input7/X _1584_/S _1513_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_0891_ _1070_/A _1043_/S VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_4
X_1443_ _1443_/B _1690_/D _1683_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1374_ _1372_/Y _1410_/B _1373_/X _1375_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__o21a_2
XFILLER_23_247 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1090_ _1090_/X _0981_/X _0973_/X _0983_/X _1115_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__a211o_2
XFILLER_9_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0874_ _1707_/Q _0989_/A _1073_/C _1005_/B _0874_/X _0990_/A VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__a2111o_2
X_0943_ VGND VPWR _0944_/C _0989_/A _1012_/B VGND VPWR sky130_fd_sc_hd__xnor2_2
X_1426_ VGND VPWR _1427_/B _1730_/Q _1428_/B VGND VPWR sky130_fd_sc_hd__xnor2_2
X_1357_ _1764_/Q _1602_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
X_1288_ _1288_/X _1292_/B _1276_/B _1151_/B _1273_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_2
XFILLER_50_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1142_ _1276_/B _1143_/A _1276_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1211_ _1287_/A _1211_/Y _1210_/Y _1270_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__o21ai_2
X_1073_ _1073_/C _1085_/C _1073_/A _1073_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nor3_2
XFILLER_20_18 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0857_ VPWR VGND _0858_/B _1706_/Q _1012_/B VGND VPWR sky130_fd_sc_hd__xor2_2
X_0926_ _1050_/B _1058_/B _0926_/X _1708_/Q _1074_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__or4b_2
X_0788_ _1683_/D _1435_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_6
X_1409_ _1409_/C _1725_/Q _1410_/C _1409_/B _1409_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_2
XFILLER_51_150 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_191 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1691_ _1691_/Q fanout171/X _1691_/D _1742_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1760_ _1760_/Q fanout179/X _1760_/D _1766_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1125_ _1276_/B _1126_/A _1205_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
X_1056_ _1101_/B _1056_/X _1678_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
Xoutput17 VPWR VGND nmatrix_col_out_n[11] _1272_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput28 VPWR VGND nmatrix_col_out_n[21] _1289_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput39 VPWR VGND nmatrix_col_out_n[31] _1303_/Y VGND VPWR sky130_fd_sc_hd__buf_4
X_0909_ VGND VPWR _0909_/Y _1699_/Q _1701_/Q VGND VPWR sky130_fd_sc_hd__xnor2_2
XFILLER_0_249 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_101 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_61 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_80 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1743_ _1743_/Q fanout172/X _1743_/D _1743_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1674_ _1674_/Q fanout181/X _1674_/D _1769_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
Xadc_core_digital_193 pmatrix_row_out_n[0] adc_core_digital_193/HI VPWR VGND VGND
+ VPWR sky130_fd_sc_hd__conb_1
X_1039_ _1046_/B _1116_/A _1039_/X _1039_/B _1039_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_2
X_1108_ VGND VPWR _1116_/B _1107_/Y _1190_/A _1108_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_44_267 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1390_ _1723_/D _1390_/B _1769_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__xnor2_4
X_1726_ _1726_/Q fanout171/X _1726_/D _1742_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1588_ VPWR VGND _1761_/Q _1588_/X _1640_/B VGND VPWR sky130_fd_sc_hd__and2_2
X_1657_ VGND VPWR _1665_/S _1766_/Q _1677_/D _1658_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_17_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0890_ _1670_/Q _1101_/B _0890_/X _0869_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__a21bo_2
X_1442_ VGND VPWR _1443_/B _1690_/Q _1444_/B VGND VPWR sky130_fd_sc_hd__xnor2_2
X_1511_ VGND VPWR _1684_/D _1511_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1373_ _1373_/B _1373_/X _1722_/Q _1373_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
X_1709_ _1709_/Q fanout182/X _1709_/D _1770_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_48_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_248 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_101 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_0873_ _0871_/X _1058_/D _0912_/A _0836_/X _0946_/A _0873_/X VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__o32a_2
X_0942_ VPWR VGND _0980_/C _1673_/Q VGND VPWR sky130_fd_sc_hd__buf_6
X_1425_ _1729_/Q _1428_/B _1728_/Q _1432_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
X_1356_ VGND VPWR _1716_/D _1762_/Q _1356_/B VGND VPWR sky130_fd_sc_hd__xnor2_2
X_1287_ _1287_/B _1292_/B _1287_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_11_218 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_222 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_277 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_60 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1072_ _1072_/B _1680_/D _1507_/S VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1210_ _1210_/Y _1276_/A _1276_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1141_ VPWR VGND _1276_/A _1205_/A VGND VPWR sky130_fd_sc_hd__buf_6
XFILLER_37_126 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0787_ _1435_/B _1607_/B _1563_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_8
X_0856_ _0859_/C _1707_/Q _0989_/A _0990_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
X_0925_ _1710_/Q _1708_/Q _1709_/Q _1074_/D _0925_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__or4b_4
X_1408_ _1418_/C _1725_/Q _1409_/D _1409_/C _1409_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__o31a_4
X_1339_ _1339_/X _1765_/Q _1328_/B _1719_/Q _1328_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_2
XFILLER_28_126 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_137 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_61 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_151 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1690_ _1690_/Q fanout174/X _1690_/D _1745_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1124_ _1124_/X _1276_/C _1131_/A _1130_/A _1173_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__o31a_4
X_1055_ VPWR VGND _1287_/B _1170_/S VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput18 VPWR VGND nmatrix_col_out_n[12] _1274_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput29 VPWR VGND nmatrix_col_out_n[22] _1290_/X VGND VPWR sky130_fd_sc_hd__buf_4
X_0839_ _1084_/A _1074_/D _1058_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__or2_4
X_0908_ _1062_/B _1671_/Q _0918_/A _0908_/B _0908_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_2
XPHY_102 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_4 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_162 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1742_ _1742_/Q fanout172/X _1742_/D _1742_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1673_ _1673_/Q fanout179/X _1673_/D _1766_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
Xadc_core_digital_194 adc_core_digital_194/LO nmatrix_rowon_out_n[15] VPWR VGND VGND
+ VPWR sky130_fd_sc_hd__conb_1
XFILLER_26_29 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1107_ _1190_/A _1037_/B _1016_/A _1107_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_2
X_1038_ VPWR VGND _1039_/D _1038_/B _1037_/A VGND VPWR sky130_fd_sc_hd__and2b_2
X_1725_ _1725_/Q fanout175/X _1725_/D _1746_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1587_ _1559_/B _1569_/B _1587_/X _1584_/X _1586_/X _1723_/D VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__o221a_2
X_1656_ VGND VPWR _1765_/D _1656_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_17_257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_10 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1441_ _1688_/Q _1444_/B _1687_/Q _1689_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
XFILLER_4_183 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1510_ VGND VPWR _1514_/S input6/X _1626_/S _1511_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_1372_ _1722_/Q _1373_/C _1373_/B _1372_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_2
XFILLER_16_290 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1708_ _1708_/Q fanout181/X _1708_/D _1770_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1639_ _1726_/D _1639_/X _1732_/D _1620_/A _1569_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__o22a_2
XFILLER_1_164 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0941_ _1809_/A _0940_/X _0939_/A _1070_/A _1672_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__o211a_2
X_0872_ _1013_/A _1058_/D _1013_/C _1073_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__or3_4
X_1424_ _1514_/S _1423_/Y _1422_/X _1729_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_2
X_1355_ _1410_/B _1356_/B _1354_/X _1353_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__o21ai_2
X_1286_ _1169_/A _1209_/X _1286_/X _1273_/A _1285_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__a22o_2
XFILLER_6_234 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_289 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_8 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1140_ VPWR VGND _1140_/X _1140_/A VGND VPWR sky130_fd_sc_hd__buf_4
X_1071_ _1072_/B _1071_/B _1680_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__xnor2_4
X_0924_ VGND VPWR _0924_/Y _1708_/Q _1050_/B VGND VPWR sky130_fd_sc_hd__xnor2_2
X_0786_ _1563_/A _1615_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_4
X_0855_ _1706_/Q _0990_/A _1012_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
X_1407_ VPWR VGND _1407_/A _1409_/D _1407_/B VGND VPWR sky130_fd_sc_hd__and2_2
X_1338_ _1382_/B _1338_/C _1338_/A _1403_/A _1338_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__and4_2
XFILLER_45_39 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1269_ _1269_/X _1186_/X _1169_/A _1268_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
XFILLER_3_237 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1123_ VPWR VGND _1276_/C _1471_/A VGND VPWR sky130_fd_sc_hd__buf_6
X_1054_ VGND VPWR _1170_/S _1061_/B _1122_/B VGND VPWR sky130_fd_sc_hd__xnor2_2
X_0907_ _1073_/A _1012_/B _0933_/B _0914_/C _0908_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__nor4b_4
X_0769_ input7/X _1602_/B input6/X input8/X VPWR VGND VGND VPWR sky130_fd_sc_hd__or3_4
X_0838_ VPWR VGND _1058_/B _1710_/Q VGND VPWR sky130_fd_sc_hd__buf_6
Xoutput19 VPWR VGND nmatrix_col_out_n[13] _1275_/X VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_24_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_103 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_200 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_5 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_130 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_196 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1741_ _1741_/Q fanout173/X _1741_/D _1742_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_30_166 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1672_ _1672_/Q fanout181/X _1672_/D _1769_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1106_ _1106_/A _1104_/Y _1111_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__or2b_2
Xadc_core_digital_195 adc_core_digital_195/LO pmatrix_c0_out_n VPWR VGND VGND VPWR
+ sky130_fd_sc_hd__conb_1
X_1037_ _1037_/A _1037_/B _1037_/X _1078_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__or3_2
XFILLER_44_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_159 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_100 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_280 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_51 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1724_ _1724_/Q fanout175/X _1724_/D _1746_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1586_ _1586_/B _1586_/X _1719_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
X_1655_ VGND VPWR _1663_/B _1765_/Q _1676_/D _1656_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_40_261 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_22 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1440_ _1440_/B _1689_/D _1683_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1371_ _1373_/C _1767_/Q _1371_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1638_ _1637_/X _1638_/Y _1615_/B _1626_/S VGND VPWR VGND VPWR sky130_fd_sc_hd__o21ai_2
X_1707_ _1707_/Q fanout180/X _1707_/D _1707_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1569_ _1569_/B _1569_/X _1720_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
XFILLER_14_239 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_176 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_261 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0940_ _1101_/B _0940_/X _1672_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
X_0871_ _1026_/B _1027_/D _0871_/X _1005_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__or3_2
X_1423_ _1423_/Y _1728_/Q _1729_/Q _1432_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__nand3b_2
X_1354_ _1354_/B _1354_/X _1354_/A _1354_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
X_1285_ _1285_/X _1221_/B _1144_/X _1258_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
XFILLER_48_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_29 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_117 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_246 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1070_ _1466_/B _1071_/B _1070_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_0854_ VPWR VGND _1012_/B _1704_/Q VGND VPWR sky130_fd_sc_hd__buf_6
X_0923_ VGND VPWR _0897_/X _0896_/Y _1700_/Q _0923_/X VGND VPWR sky130_fd_sc_hd__mux2_2
X_0785_ _1420_/A _0785_/C _0785_/A _0785_/D _1615_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_4
X_1406_ _1401_/B _1405_/X _1407_/B _1404_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__a21bo_2
X_1337_ _1338_/D _1765_/Q _1719_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1268_ _1255_/A _1268_/Y _1270_/B _1173_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__o21ai_2
X_1199_ _1199_/X _1287_/B _1246_/B _1221_/A _1246_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__o31a_2
XFILLER_3_249 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_50 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_131 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1122_ _1471_/A _1122_/B _1122_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__xnor2_4
X_1053_ _1047_/Y _1040_/S _1122_/B _1052_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_4
X_0837_ VPWR VGND _1074_/D _1711_/Q VGND VPWR sky130_fd_sc_hd__buf_4
X_0906_ _1014_/C _0933_/B _1058_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_0768_ _0775_/B _1691_/Q _0768_/X _1695_/Q _0768_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_2
XPHY_104 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_6 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1740_ _1740_/Q fanout172/X _1740_/D _1742_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1671_ _1671_/Q fanout179/X _1671_/D _1766_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
Xadc_core_digital_196 adc_core_digital_196/LO pmatrix_rowon_out_n[15] VPWR VGND VGND
+ VPWR sky130_fd_sc_hd__conb_1
XFILLER_53_248 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1105_ _1111_/B _1040_/S _1113_/A _1104_/Y _0993_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__a211o_2
X_1036_ _1022_/X _1106_/A _1004_/B _1078_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_44_248 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1723_ _1723_/Q fanout175/X _1723_/D _1746_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1654_ VGND VPWR _1764_/D _1654_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1585_ _1586_/B _1633_/A _1585_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
XFILLER_41_218 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1019_ _1019_/B _1676_/D _1507_/S VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_1_303 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_207 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1370_ _1721_/Q _1373_/B _1371_/B _1767_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__o21ai_2
X_1637_ _1637_/X _1633_/A _1514_/S _1585_/B _1427_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__o31a_2
X_1706_ _1706_/Q fanout181/X _1706_/D _1770_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1568_ _1735_/Q _1735_/D _1563_/X _1567_/X _1620_/A _1435_/B VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__a32o_2
X_1499_ _1779_/A _1804_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_48_29 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_188 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0870_ _1084_/A _1073_/B _1702_/Q _1058_/C _0912_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_4
X_1422_ _1729_/Q _1432_/C _1422_/X _1728_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__a21bo_2
X_1353_ _1354_/A _1354_/C _1354_/B _1353_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_2
X_1284_ _1284_/X _1221_/B _1237_/B _1224_/Y _1248_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__a211o_2
XFILLER_48_192 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0999_ _1101_/B _0999_/X _1675_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
XFILLER_10_265 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_72 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0853_ VPWR VGND _0989_/A _1705_/Q VGND VPWR sky130_fd_sc_hd__buf_6
X_0922_ _1809_/A _0921_/X _0920_/A _1070_/A _1671_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__o211a_2
X_0784_ _1686_/Q _0783_/X _0780_/X _0785_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__o21a_2
X_1405_ _1405_/X _1723_/Q _1385_/B _1769_/Q _1385_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_2
X_1267_ _1267_/X _1129_/X _1144_/X _1183_/X _1178_/B VGND VPWR _1292_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_2
X_1198_ VPWR VGND _1265_/A _1198_/X _1198_/B VGND VPWR sky130_fd_sc_hd__and2_2
X_1336_ _1719_/Q _1338_/C _1765_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
Xinput1 VGND VPWR input1/X clk_dig_in VGND VPWR sky130_fd_sc_hd__buf_1
X_1121_ _1131_/A _1205_/A _1276_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1052_ _1052_/X _1051_/Y _1049_/Y _1024_/X _1025_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_2
X_0767_ _1693_/Q _1687_/Q _0768_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__or2b_2
X_0905_ _0989_/A _1074_/D _1014_/C _1058_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__or3_2
X_0836_ _1013_/C _0836_/X _0836_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
X_1319_ _1402_/C _1319_/X _1319_/A _1402_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
XPHY_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_10 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_7 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_45 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_67 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1670_ _1670_/Q fanout179/X _1670_/D _1766_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_23_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1035_ _1035_/B _1037_/A _1035_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1104_ VGND VPWR _1104_/Y _1190_/A _1115_/A VGND VPWR sky130_fd_sc_hd__xnor2_2
XFILLER_21_113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1799_ VGND VPWR _1799_/X _1799_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_0819_ _0819_/B _0819_/X _1757_/Q _0819_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
XFILLER_12_179 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1584_ VGND VPWR _1584_/S _1721_/D _1717_/D _1584_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_1722_ _1722_/Q fanout176/X _1722_/D _1746_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1653_ VGND VPWR _1663_/B _1764_/Q _1675_/D _1654_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_26_249 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_271 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1018_ VGND VPWR _1043_/S _1205_/A _1035_/A _1019_/B VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_40_274 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_197 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1705_ _1705_/Q fanout180/X _1705_/D _1707_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1636_ _1747_/D _1569_/B _1632_/X _1731_/D _1634_/X _1635_/X VPWR VGND VGND VPWR
+ sky130_fd_sc_hd__o311a_2
X_1567_ VGND VPWR _1585_/B _1566_/X _1719_/D _1567_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_1498_ _1788_/A _1795_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_38_52 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_296 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1421_ _1615_/B _1728_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
X_1283_ _1283_/X _1221_/B _1140_/X _1219_/B _1248_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__a211o_2
X_1352_ _1716_/Q _1354_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
X_0998_ _1261_/C _1190_/B _1190_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__xor2_4
X_1619_ _1744_/D _1619_/A _1619_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
XFILLER_10_277 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0921_ _1101_/B _0921_/X _1671_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
X_0783_ _0783_/X _0782_/X _0781_/Y _1558_/B _1693_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__a211o_2
X_0852_ _0852_/A _1073_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__buf_8
XFILLER_5_281 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1404_ _1404_/X _1769_/Q _1385_/A _1385_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
X_1335_ _1720_/Q _1403_/A _1766_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
X_1266_ _1266_/X _1255_/Y _1248_/X _1265_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
Xinput2 VPWR VGND input2/X comparator_in VGND VPWR sky130_fd_sc_hd__buf_4
X_1197_ _1196_/X _1197_/Y _1195_/X _1276_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__o21ai_2
XFILLER_19_10 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_262 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1051_ _1076_/B _1051_/Y _1076_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1120_ _1158_/A _1158_/B _1130_/A _1138_/B _1138_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__a22o_2
X_0904_ VGND VPWR _0914_/C _1707_/Q _1706_/Q VGND VPWR sky130_fd_sc_hd__xnor2_2
X_0766_ _1692_/Q _1688_/Q _0775_/B _1690_/Q _1694_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_2
X_0835_ VPWR VGND _1013_/C _0865_/C VGND VPWR sky130_fd_sc_hd__buf_6
X_1318_ _1319_/A _1402_/D _1402_/C _1318_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_2
XPHY_106 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1249_ _1132_/X _1203_/X _1248_/X _1249_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_47_236 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_52 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_8 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1103_ _1784_/A _1799_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
X_1034_ _1031_/Y _1030_/Y _1039_/B _1034_/Y _1037_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__a211oi_4
X_0818_ _0819_/B _0819_/C _1757_/Q _0818_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_2
X_1798_ VGND VPWR _1798_/X _1798_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_29_203 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1721_ _1721_/Q fanout176/X _1721_/D _1721_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1583_ _1738_/D _1579_/X _1760_/Q _1581_/X _1640_/B VGND VPWR _1582_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_2
X_1652_ VGND VPWR _1763_/D _1652_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1017_ VPWR VGND _1205_/A _1208_/A VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_43_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1704_ _1704_/Q fanout180/X _1704_/D _1707_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1497_ _1788_/A _1794_/A _1497_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1635_ _1683_/D _1747_/Q _1632_/X _1725_/D _1620_/A _1635_/X VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__o32a_2
X_1566_ VGND VPWR _1626_/S _1717_/D _1715_/D _1566_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_13_89 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1420_ _1420_/B _1615_/B _1420_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
X_1351_ VPWR VGND _1714_/D _1351_/B _1760_/Q VGND VPWR sky130_fd_sc_hd__xor2_2
X_1282_ _1237_/A _1281_/X _1209_/X _1270_/B _1282_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o211a_2
X_1618_ _1596_/C _1633_/A _1604_/A _1617_/Y _1619_/B _1593_/A VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__a2111o_2
X_0997_ _0993_/A _1040_/S _1113_/A _1190_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_4
X_1549_ VGND VPWR _1712_/D _1549_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_10_201 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_289 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_44 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_10 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_109 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_0920_ _0920_/A _0920_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
X_0782_ _1584_/S _1580_/S _0782_/X _1687_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__or3_2
X_0851_ _1013_/C _0852_/A _1013_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
XFILLER_5_293 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1265_ _1265_/Y _1265_/A _1265_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1403_ _1403_/B _1409_/C _1403_/A _1403_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
X_1334_ _1338_/A _1766_/Q _1720_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
Xinput3 VGND VPWR input3/X config_1_in[0] VGND VPWR sky130_fd_sc_hd__buf_1
X_1196_ _1196_/X _1221_/A _1158_/B _1178_/B _1158_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_2
XFILLER_27_120 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_274 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1050_ _1050_/C _1074_/D _1076_/B _1050_/B _1050_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_2
X_0903_ _0866_/A _1026_/B _0902_/X _0901_/Y _1058_/A _1062_/B VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__a2111oi_4
X_0834_ _1697_/Q _1699_/Q _0865_/C _1698_/Q _1808_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_2
X_0765_ VGND VPWR _1689_/Q _0764_/X _0762_/X _0785_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_1317_ _1717_/Q _1319_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
X_1248_ VPWR VGND _1248_/X _1292_/A VGND VPWR sky130_fd_sc_hd__buf_6
X_1179_ _1179_/Y _1287_/A _1179_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
XFILLER_24_167 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_107 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_9 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_248 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1102_ _1808_/A _1681_/D _1101_/X _1467_/A _1070_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__o31ai_2
XFILLER_38_248 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1033_ _1033_/B _1039_/B _1676_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1797_ VPWR VGND _1797_/X _1797_/A VGND VPWR sky130_fd_sc_hd__buf_2
X_0817_ _1758_/Q _0819_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_16_56 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_67 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1720_ _1720_/Q fanout173/X _1720_/D _1743_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1651_ VGND VPWR _1663_/B _1763_/Q _1674_/D _1652_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_1582_ _1596_/B _1582_/X _1738_/Q _1615_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
X_1016_ VPWR VGND _1208_/A _1016_/B _1016_/A VGND VPWR sky130_fd_sc_hd__xor2_2
XFILLER_4_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_155 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1634_ _1632_/X _1626_/S _1604_/A _1633_/X _1634_/X _1729_/D VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__a2111o_2
X_1703_ _1703_/Q fanout180/X _1703_/D _1758_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_31_298 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1565_ VPWR VGND _1620_/A _1565_/A VGND VPWR sky130_fd_sc_hd__buf_4
X_1496_ _1793_/A _1496_/A _1788_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_13_35 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_221 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_287 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1350_ _1350_/B _1351_/B _1420_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1281_ _1144_/X _1151_/A _1281_/X _1276_/C _1246_/C _1246_/B VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__a41o_2
XFILLER_48_162 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_0996_ _0981_/X _0938_/B _1040_/S _0995_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_4
X_1617_ _1726_/D _1617_/Y _1633_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1479_ _1800_/A _1784_/A _1495_/A _1487_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__o21ai_4
X_1548_ VGND VPWR _1548_/S _1507_/S _1712_/Q _1549_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_10_213 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_22 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0850_ _1701_/Q _1703_/Q _1700_/Q _1702_/Q _1013_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_4
X_0781_ _1687_/Q _0781_/Y _1580_/S _1584_/S VGND VPWR VGND VPWR sky130_fd_sc_hd__o21ai_2
XFILLER_5_261 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1402_ VPWR VGND _1409_/B _1382_/Y _1402_/D _1402_/C _1403_/C VGND VPWR sky130_fd_sc_hd__and4b_2
X_1264_ _1248_/X _1164_/X _1264_/X _1233_/A _1263_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__a22o_2
Xinput4 VGND VPWR input4/X config_1_in[1] VGND VPWR sky130_fd_sc_hd__buf_1
X_1333_ _1719_/D _1333_/B _1765_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__xnor2_4
X_1195_ _1195_/X _1191_/A _1287_/B _1221_/A _1194_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__o31a_2
XFILLER_36_176 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0979_ _0975_/A _0976_/Y _0979_/X _0980_/D _0978_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__a22o_2
XFILLER_35_66 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_286 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0902_ _1058_/B _1074_/D _1050_/B _0902_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o21a_2
X_0833_ _1703_/Q _0836_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
X_0764_ _1565_/A _0764_/X _1691_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
X_1316_ _1716_/Q _1354_/B _1354_/C _1762_/Q _1402_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_4
X_1178_ _1179_/B _1276_/A _1178_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1247_ _1247_/X _1246_/X _1255_/B _1178_/B _1203_/X VGND VPWR _1213_/Y VGND VPWR
+ sky130_fd_sc_hd__a221o_2
Xoutput160 VPWR VGND sample_switch_out _1808_/X VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_46_10 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_43 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1101_ _1808_/A _1101_/B _1681_/Q _1101_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__or3b_2
X_1032_ _1037_/B _1048_/B _1050_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__xnor2_4
XFILLER_38_205 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1796_ VGND VPWR _1796_/X _1796_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_0816_ _0816_/B _1757_/D _1538_/S VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_35_208 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1581_ _1581_/B _1581_/X _1604_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
X_1650_ VGND VPWR _1762_/D _1650_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1015_ _1010_/Y _1016_/B _1011_/X _1014_/X _1013_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o2bb2a_2
X_1779_ VPWR VGND _1779_/X _1779_/A VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_17_219 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_101 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_288 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1564_ _1734_/Q _1435_/B _1734_/D _1563_/X _1562_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__a22o_2
X_1633_ VPWR VGND _1633_/A _1633_/X _1727_/D VGND VPWR sky130_fd_sc_hd__and2_2
X_1702_ _1702_/Q fanout180/X _1702_/D _1758_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1495_ _1792_/A _1495_/A _1788_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_22_211 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_303 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_237 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1280_ _1129_/X _1169_/A _1209_/X _1280_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o21a_2
X_0995_ _0995_/X _0977_/X _0980_/C _0933_/X _0974_/B VGND VPWR _0994_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_2
X_1616_ _1619_/A _1596_/C _1376_/A _1620_/A _1614_/Y _1615_/X VPWR VGND VGND VPWR
+ sky130_fd_sc_hd__o311a_2
X_1547_ VGND VPWR _1711_/D _1547_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1478_ _1801_/A _1782_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_10_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_79 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_10 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0780_ _0779_/X _1687_/Q _0768_/D _1580_/S _1584_/S _0780_/X VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__o32a_2
XFILLER_5_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1401_ _1403_/C _1407_/A _1401_/A _1401_/B _1401_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__and4_2
X_1263_ _1263_/X _1237_/A _1265_/A _1265_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
X_1332_ _1420_/A _1332_/B _1367_/B _1333_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__or3b_4
Xinput5 VGND VPWR input5/X config_1_in[2] VGND VPWR sky130_fd_sc_hd__buf_1
X_1194_ _1173_/A _1138_/B _1138_/A _1194_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_2
X_0978_ _1013_/C _0859_/B _0946_/X _0944_/X _0978_/Y _0977_/X VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__a2111oi_2
XFILLER_2_221 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0763_ _1565_/A _1560_/A _0763_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_0832_ _0830_/Y _1542_/S _0831_/X _1753_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__o21a_2
X_0901_ VGND VPWR _0901_/Y _1058_/B _1050_/B VGND VPWR sky130_fd_sc_hd__xnor2_2
X_1315_ _1354_/C _1354_/B _1402_/C _1762_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_2_71 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1246_ _1246_/A _1246_/B _1246_/X _1246_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__or3_2
X_1177_ VPWR VGND _1287_/A _1246_/A VGND VPWR sky130_fd_sc_hd__buf_6
Xoutput150 VPWR VGND result_out[2] _1735_/Q VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput161 VPWR VGND sample_switch_out_n _1809_/X VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_46_22 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_106 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1100_ VPWR VGND _1100_/X _1467_/A VGND VPWR sky130_fd_sc_hd__buf_6
X_1031_ _1038_/B _1031_/Y _1025_/B _1113_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__o21bai_2
X_1795_ VGND VPWR _1795_/X _1795_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_0815_ VGND VPWR _0816_/B _1757_/Q _0819_/C VGND VPWR sky130_fd_sc_hd__xnor2_2
XFILLER_16_47 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_231 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1229_ _1229_/X _1209_/X _1252_/A _1265_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
XFILLER_43_231 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1580_ VGND VPWR _1580_/S _1720_/D _1718_/D _1581_/B VGND VPWR sky130_fd_sc_hd__mux2_1
X_1014_ _1014_/C _1050_/B _1014_/X _1014_/B _1026_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__or4b_2
X_1778_ VPWR VGND _1778_/X _1778_/A VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_27_13 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1701_ _1701_/Q fanout180/X _1701_/D _1758_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1494_ VPWR VGND _1791_/A _1494_/A VGND VPWR sky130_fd_sc_hd__buf_2
X_1632_ _1769_/Q _1615_/A _1602_/B _1632_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o21a_2
X_1563_ VPWR VGND _1563_/X _1563_/A VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_9_249 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0994_ _1672_/Q _0980_/D _0974_/B _0980_/C _0994_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o211a_2
X_1615_ _1615_/A _1615_/B _1615_/X _1615_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__or3_2
X_1477_ _1801_/A _1784_/A _1487_/B _1496_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__o21ai_4
X_1546_ VGND VPWR _1546_/S _1074_/D _1712_/Q _1547_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_27_315 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_237 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_22 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1331_ _1367_/B _1719_/Q _1331_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1400_ VPWR VGND _1401_/D _1769_/Q _1723_/Q VGND VPWR sky130_fd_sc_hd__xor2_2
X_1193_ _1179_/Y _1193_/Y _1192_/X _1273_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__o21ai_2
X_1262_ _1256_/A _1262_/Y _1261_/X _1276_/C _1164_/X _1143_/A VPWR VGND VGND VPWR
+ sky130_fd_sc_hd__a221oi_4
Xinput6 VPWR VGND input6/X config_1_in[3] VGND VPWR sky130_fd_sc_hd__buf_2
X_0977_ _1673_/Q _0977_/X _1672_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
X_1529_ VGND VPWR _1702_/D _1529_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_42_104 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_233 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_90 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_0900_ _1074_/D _1058_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_33_148 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_0762_ _0759_/X _0762_/X _0763_/B _1560_/A _1691_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__o22a_2
X_0831_ _1752_/Q _0831_/X _0831_/A _0831_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
X_1314_ _1354_/C _1715_/Q _1761_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_44_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1245_ _1245_/X _1244_/X _1255_/B _1178_/B _1157_/Y VGND VPWR _1213_/Y VGND VPWR
+ sky130_fd_sc_hd__a221o_2
XFILLER_49_281 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1176_ _1029_/Y _1040_/X _1034_/Y _1246_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__o21a_2
Xoutput151 VPWR VGND result_out[3] _1736_/Q VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput140 VPWR VGND pmatrix_rowon_out_n[8] _1800_/X VGND VPWR sky130_fd_sc_hd__buf_4
X_1030_ _1030_/Y _1676_/Q _1033_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_0814_ VPWR VGND _1756_/Q _0819_/C _0814_/B VGND VPWR sky130_fd_sc_hd__and2_2
X_1794_ VGND VPWR _1794_/X _1794_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1228_ VGND VPWR _1228_/X _1227_/X _1230_/A _1173_/A _1287_/A _1157_/Y VGND VPWR
+ sky130_fd_sc_hd__a311o_2
XFILLER_52_287 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_243 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1159_ VPWR VGND _1265_/A _1252_/A VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_20_173 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_100 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1013_ _1013_/C _1013_/A _1013_/X _1013_/B _1013_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_2
X_1777_ VGND VPWR _1777_/X _1777_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_27_25 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_254 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1631_ _1746_/D _1630_/X _1628_/X _1563_/X _1627_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_2
X_1700_ _1700_/Q fanout178/X _1700_/D _1758_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_33_90 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1493_ _1788_/A _1494_/A _1495_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
X_1562_ _1593_/B _1562_/X _0763_/B _1716_/D _1584_/S _1718_/D VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__a32o_2
XFILLER_9_206 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0993_ _1113_/A _0993_/A _0993_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_4
X_1614_ _1766_/Q _1640_/B _1435_/B _1744_/Q _1614_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__a22oi_2
X_1476_ _1802_/A _1781_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
X_1545_ VGND VPWR _1710_/D _1545_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_24_15 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_165 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_209 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_249 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_34 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_157 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1330_ _1331_/B _1332_/B _1719_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1261_ VGND VPWR _1471_/A _1261_/X _1194_/Y _1261_/C VGND VPWR sky130_fd_sc_hd__and3b_2
X_1192_ _1221_/A _1175_/X _1152_/C _1192_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o21a_2
Xinput7 VPWR VGND input7/X config_1_in[4] VGND VPWR sky130_fd_sc_hd__buf_2
X_0976_ _0980_/C _0976_/Y _1672_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1459_ _1459_/B _1695_/D _1683_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1528_ VGND VPWR _1542_/S _1702_/Q _1703_/Q _1529_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_51_57 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0830_ _0831_/A _0831_/C _1752_/Q _0830_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_2
XPHY_91 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_80 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_0761_ _1686_/Q _0763_/B _1633_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1313_ _1715_/Q _1761_/Q _1354_/B _1310_/C _1310_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__a22o_2
X_1244_ _1287_/A _1246_/B _1198_/B _1244_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__or3b_2
XFILLER_49_293 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1175_ VPWR VGND _1175_/X _1175_/A VGND VPWR sky130_fd_sc_hd__buf_4
X_0959_ _1073_/B _0964_/C _0959_/X _0959_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__or3_2
Xoutput141 VPWR VGND pmatrix_rowon_out_n[9] _1801_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput152 VPWR VGND result_out[4] _1737_/Q VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput130 VPWR VGND pmatrix_rowon_out_n[12] _1804_/X VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_47_219 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0813_ _0813_/B _1756_/D _1538_/S VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1793_ VGND VPWR _1793_/X _1793_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1227_ _1246_/B _1213_/Y _1246_/C _1227_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o21a_2
X_1158_ VPWR VGND _1158_/A _1252_/A _1158_/B VGND VPWR sky130_fd_sc_hd__and2_2
X_1089_ _1079_/X _1076_/X _1115_/A _1078_/A _1078_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__o2bb2a_4
XFILLER_32_15 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_263 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_123 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1012_ _1012_/B _1013_/D _1712_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
XFILLER_27_37 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_277 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1630_ _1630_/X _1629_/X _1596_/C _1746_/Q _1596_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_2
X_1561_ _1585_/B _1593_/B _1561_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1492_ VPWR VGND _1790_/A _1492_/A VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_39_314 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1759_ _1759_/Q fanout179/X _1759_/D _1766_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_13_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_218 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_177 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0992_ _1190_/A _1004_/B _1004_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__xnor2_4
X_1613_ VGND VPWR _1743_/D _1613_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1544_ VGND VPWR _1546_/S _1058_/B _1074_/D _1545_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_1475_ _1802_/A _1784_/A _1487_/B _1497_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_49_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xinput8 VPWR VGND input8/X config_1_in[5] VGND VPWR sky130_fd_sc_hd__buf_2
X_1260_ _1260_/X _1255_/Y _1273_/A _1259_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
X_1191_ VPWR VGND _1273_/A _1191_/A VGND VPWR sky130_fd_sc_hd__buf_4
X_0975_ _1672_/Q _0975_/Y _0975_/A _0980_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__nor3b_2
X_1527_ VGND VPWR _1701_/D _1527_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1458_ VPWR VGND _1459_/B _1458_/B _1695_/Q VGND VPWR sky130_fd_sc_hd__xor2_2
X_1389_ _1420_/A _1389_/B _1388_/Y _1390_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__or3b_4
XFILLER_35_15 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_37 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0760_ _1684_/Q _1633_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XPHY_92 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_70 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1312_ VGND VPWR _1715_/D _1761_/Q _1312_/B VGND VPWR sky130_fd_sc_hd__xnor2_2
X_1174_ _1287_/B _1175_/A _1205_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
X_1243_ _1243_/Y _1243_/A _1243_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
XFILLER_24_106 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_0958_ _0959_/C _1026_/B _1674_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_0889_ VPWR VGND _1101_/B _1043_/S VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput142 VPWR VGND result_out[0] _1733_/Q VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput120 VPWR VGND pmatrix_row_out_n[3] _1794_/A VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput131 VPWR VGND pmatrix_rowon_out_n[13] _1805_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput153 VPWR VGND result_out[5] _1738_/Q VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_7_305 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1792_ VGND VPWR _1792_/X _1792_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_0812_ VGND VPWR _0813_/B _1756_/Q _0814_/B VGND VPWR sky130_fd_sc_hd__xnor2_2
X_1226_ _1225_/X _1226_/Y _1223_/X _1151_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__o21ai_2
X_1157_ _1246_/C _1157_/Y _1246_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1088_ _1679_/Q _1088_/Y _1062_/B _1678_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__o21ai_2
XFILLER_43_289 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_220 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1011_ _1011_/X _1008_/Y _0938_/B _1675_/Q _0981_/X VGND VPWR _0995_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_2
XFILLER_43_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1209_ VPWR VGND _1209_/X _1209_/A VGND VPWR sky130_fd_sc_hd__buf_4
X_1560_ _1585_/B _1560_/A _1686_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_4
X_1491_ _1788_/A _1492_/A _1496_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
X_1689_ _1689_/Q fanout174/X _1689_/D _1745_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1758_ _1758_/Q fanout178/X _1758_/D _1758_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_38_15 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_237 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_185 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0991_ _1073_/A _0990_/X _1004_/B _1076_/A _0927_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o22a_4
X_1474_ _1803_/A _1780_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
X_1612_ VPWR VGND _1612_/A _1613_/A _1612_/B VGND VPWR sky130_fd_sc_hd__and2_2
X_1543_ VGND VPWR _1709_/D _1543_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_39_123 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xinput9 VGND VPWR input9/X rst_n VGND VPWR sky130_fd_sc_hd__buf_1
X_1190_ VGND VPWR _1191_/A _1190_/A _1190_/B VGND VPWR sky130_fd_sc_hd__xnor2_2
XFILLER_36_115 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0974_ VPWR VGND _0974_/X _0974_/B _0980_/C VGND VPWR sky130_fd_sc_hd__xor2_2
X_1457_ _1458_/B _1694_/Q _1457_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1526_ VGND VPWR _1538_/S _1702_/Q _1701_/Q _1527_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_1388_ _1388_/Y _1723_/Q _1392_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
XFILLER_51_26 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_60 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_93 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1311_ _1420_/A _1311_/B _1312_/B _1311_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__or3_2
XFILLER_2_20 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1173_ _1270_/B _1173_/Y _1173_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1242_ _1243_/B _1273_/A _1255_/A _1153_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
XFILLER_24_118 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_184 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xoutput121 VPWR VGND pmatrix_row_out_n[4] _1795_/A VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput110 VPWR VGND pmatrix_col_out_n[8] _1180_/Y VGND VPWR sky130_fd_sc_hd__buf_4
X_0957_ _1710_/Q _1712_/Q _0964_/C _1711_/Q _1709_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_2
Xoutput132 VPWR VGND pmatrix_rowon_out_n[14] _1806_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput143 VPWR VGND result_out[10] _1743_/Q VGND VPWR sky130_fd_sc_hd__buf_4
X_0888_ _0887_/Y _0887_/B _0885_/X _1524_/S _1043_/S VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_4
Xoutput154 VPWR VGND result_out[6] _1739_/Q VGND VPWR sky130_fd_sc_hd__buf_4
X_1509_ VPWR VGND _1626_/S _1580_/S VGND VPWR sky130_fd_sc_hd__buf_6
XFILLER_15_107 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_265 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_92 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1791_ VGND VPWR _1791_/X _1791_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_0811_ input2/X _0814_/B _1754_/Q _1755_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
XFILLER_16_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1225_ _1255_/A _1225_/X _1224_/Y _1144_/X _1276_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__o22a_2
X_1087_ VPWR VGND _1087_/X _1680_/Q _1487_/A VGND VPWR sky130_fd_sc_hd__and2b_2
XFILLER_37_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_210 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1156_ _1132_/X _1256_/A _1156_/X _1261_/C _1155_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__a22o_2
X_1010_ _1010_/B _1010_/Y _1038_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1208_ _1471_/A _1209_/A _1208_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
X_1139_ VPWR VGND _1246_/B _1140_/A _1246_/C VGND VPWR sky130_fd_sc_hd__and2_2
XFILLER_25_235 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_27 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1490_ VGND VPWR _1789_/A _1490_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_15_290 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1688_ _1688_/Q fanout170/X _1688_/D _1745_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1757_ _1757_/Q fanout182/X _1757_/D _1758_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_13_249 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_260 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1611_ _1612_/B _1609_/X _1585_/B _1610_/X _1596_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__a211o_2
X_0990_ _1005_/B _0990_/A _0990_/X _1073_/C _1005_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_2
X_1473_ VPWR VGND _1779_/A _1473_/A VGND VPWR sky130_fd_sc_hd__buf_2
X_1542_ VGND VPWR _1542_/S _1050_/B _1058_/B _1543_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_39_179 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1809_ VGND VPWR _1809_/X _1809_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_40_39 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_0973_ VGND VPWR _0972_/Y _1670_/Q _0869_/B _0917_/B _0973_/X _0968_/X VGND VPWR
+ sky130_fd_sc_hd__a311o_4
X_1456_ _1456_/B _1694_/D _1683_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1387_ _1392_/B _1389_/B _1723_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1525_ VGND VPWR _1700_/D _1525_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_51_38 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_50 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_61 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_94 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1310_ _1310_/B _1311_/C _1715_/Q _1310_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
X_1241_ VGND VPWR _1240_/X _1255_/A _1239_/X _1241_/X _1217_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_2
X_1172_ _1169_/Y _1172_/X _1171_/Y _1217_/A _1132_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o22a_2
X_0956_ _1674_/Q _1014_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
Xoutput100 VPWR VGND pmatrix_col_out_n[28] _1243_/Y VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput111 VPWR VGND pmatrix_col_out_n[9] _1181_/Y VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput155 VPWR VGND result_out[7] _1740_/Q VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput122 VPWR VGND pmatrix_row_out_n[5] _1796_/A VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput144 VPWR VGND result_out[11] _1744_/Q VGND VPWR sky130_fd_sc_hd__buf_4
X_0887_ _0887_/B _0887_/Y _0887_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
Xoutput133 VPWR VGND pmatrix_rowon_out_n[1] _1793_/X VGND VPWR sky130_fd_sc_hd__buf_4
X_1439_ VPWR VGND _1440_/B _1439_/B _1689_/Q VGND VPWR sky130_fd_sc_hd__xor2_2
X_1508_ VGND VPWR _1669_/D _1508_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_46_277 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1790_ VGND VPWR _1790_/X _1790_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_0810_ _0810_/B _1755_/D _1538_/S VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1224_ _1287_/A _1178_/B _1261_/C _1224_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_2
XFILLER_35_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1086_ VGND VPWR _1487_/A _1681_/Q _1086_/B VGND VPWR sky130_fd_sc_hd__xnor2_2
X_1155_ _1237_/A _1155_/Y _1152_/C _1178_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__o21ai_2
XFILLER_20_100 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0939_ _0939_/A _0939_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_28_222 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_203 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_148 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xfanout190 VPWR VGND _1770_/CLK input1/X VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_19_277 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_53 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_192 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1207_ _1169_/A _1221_/B _1173_/Y _1207_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_4
X_1069_ _1064_/B _1068_/X _1059_/B _1067_/X _1466_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__a22oi_4
XFILLER_43_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1138_ _1138_/A _1138_/B _1246_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_8
XFILLER_16_236 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_247 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1756_ _1756_/Q fanout182/X _1756_/D _1758_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1687_ _1687_/Q _1687_/D VPWR fanout170/X _1748_/CLK VGND VGND VPWR sky130_fd_sc_hd__dfstp_4
XFILLER_8_265 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1610_ _1561_/A _1721_/D _1610_/X _1593_/B _1727_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__a22o_2
XFILLER_5_87 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1472_ _1487_/B _1473_/A _1784_/A _1495_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
X_1541_ VGND VPWR _1708_/D _1541_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1739_ _1739_/Q fanout176/X _1739_/D _1746_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1808_ VGND VPWR _1808_/X _1808_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_14_85 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_95 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0972_ _0970_/X _0971_/Y _0972_/Y _0859_/X _0849_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__a31oi_2
X_1524_ VGND VPWR _1524_/S _1701_/Q _1700_/Q _1525_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_1455_ VGND VPWR _1456_/B _1694_/Q _1457_/B VGND VPWR sky130_fd_sc_hd__xnor2_2
X_1386_ VGND VPWR _1385_/X _1383_/X _1392_/B _1401_/A _1342_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_50_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_40 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_84 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1171_ _1169_/A _1265_/B _1265_/A _1171_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_2
X_1240_ _1240_/X _1287_/B _1158_/B _1287_/A _1158_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_2
X_0955_ VPWR VGND _1507_/S _1808_/A VGND VPWR sky130_fd_sc_hd__buf_6
X_0886_ input2/X _0887_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_32_164 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xoutput145 VPWR VGND result_out[12] _1745_/Q VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput134 VPWR VGND pmatrix_rowon_out_n[2] _1794_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput101 VPWR VGND pmatrix_col_out_n[29] _1245_/X VGND VPWR sky130_fd_sc_hd__buf_4
X_1507_ VGND VPWR _1507_/S input5/X _1669_/Q _1508_/A VGND VPWR sky130_fd_sc_hd__mux2_1
Xoutput123 VPWR VGND pmatrix_row_out_n[6] _1797_/A VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput156 VPWR VGND result_out[8] _1741_/Q VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput112 VPWR VGND pmatrix_row_out_n[10] _1801_/A VGND VPWR sky130_fd_sc_hd__buf_4
X_1438_ _1439_/B _1687_/Q _1688_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1369_ _1720_/D _1369_/B _1766_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__xnor2_4
XFILLER_23_164 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_289 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_234 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1223_ _1221_/A _1223_/X _1209_/X _1273_/A _1151_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__o22a_2
XFILLER_28_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1154_ _1132_/X _1256_/A _1154_/X _1261_/C _1153_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__a22o_2
X_1085_ _1085_/B _1086_/B _1712_/Q _1085_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
X_0938_ _0939_/A _0938_/B _0938_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__xor2_4
X_0869_ _0869_/B _0878_/A _1670_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_51_281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xfanout180 VPWR VGND fanout180/X fanout182/X VGND VPWR sky130_fd_sc_hd__buf_6
X_1206_ VPWR VGND _1221_/B _1206_/A VGND VPWR sky130_fd_sc_hd__buf_6
X_1137_ _1246_/B _1158_/A _1158_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_4
X_1068_ _1093_/B _1040_/S _1052_/X _1059_/B _1068_/X _1047_/Y VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__a2111o_2
XFILLER_31_207 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_163 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1686_ _1686_/Q fanout170/X _1686_/D _1748_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1755_ _1755_/Q fanout180/X _1755_/D _1758_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_38_29 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_277 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1540_ VGND VPWR _1548_/S _1050_/B _1026_/B _1541_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_1471_ _1495_/A _1471_/A _1496_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__or2_4
X_1807_ VGND VPWR _1807_/X _1809_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1738_ _1738_/Q fanout175/X _1738_/D _1746_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1669_ _1669_/Q fanout178/X _1669_/D _1765_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_14_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_151 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_151 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0971_ _0971_/Y _1670_/Q _1671_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1454_ VPWR VGND _1693_/Q _1457_/B _1454_/B VGND VPWR sky130_fd_sc_hd__and2_2
X_1523_ VGND VPWR _1699_/D _1523_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1385_ VPWR VGND _1385_/A _1385_/X _1385_/B VGND VPWR sky130_fd_sc_hd__and2_2
XFILLER_23_313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_30 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_232 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1170_ _1170_/S _1152_/C VPWR VGND _1258_/A _1265_/B VGND VPWR sky130_fd_sc_hd__mux2_8
X_0885_ VGND VPWR _0885_/S _0884_/X _1755_/Q _0885_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_0954_ _1809_/A _0953_/X _1173_/A _1070_/A _1673_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__o211a_2
Xoutput135 VPWR VGND pmatrix_rowon_out_n[3] _1795_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput102 VPWR VGND pmatrix_col_out_n[2] _1149_/X VGND VPWR sky130_fd_sc_hd__buf_4
X_1437_ _1437_/B _1688_/D _1683_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1506_ VGND VPWR _1668_/D _1506_/A VGND VPWR sky130_fd_sc_hd__buf_1
Xoutput157 VPWR VGND result_out[9] _1742_/Q VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput146 VPWR VGND result_out[13] _1746_/Q VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput113 VPWR VGND pmatrix_row_out_n[11] _1802_/A VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput124 VPWR VGND pmatrix_row_out_n[7] _1798_/A VGND VPWR sky130_fd_sc_hd__buf_4
X_1368_ _1369_/B _1410_/B _1367_/X _1366_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__o21ai_4
X_1299_ _1299_/Y _1276_/A _1151_/A _1246_/C _1276_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__a31oi_4
XFILLER_11_305 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_10 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_246 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1222_ _1222_/X _1230_/A _1261_/C _1220_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
X_1153_ _1153_/Y _1233_/A _1153_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1084_ _1084_/A _1085_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_37_246 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0868_ _0836_/X _0843_/X _0849_/X _0859_/X _0867_/X _0869_/B VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__o2111ai_4
X_0937_ _0918_/A _0919_/A _0938_/B _0936_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_4
X_0799_ _0793_/X _0798_/X _1524_/S _0789_/X _1753_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__a22o_4
Xfanout170 VPWR VGND fanout170/X fanout183/X VGND VPWR sky130_fd_sc_hd__buf_6
Xfanout181 VPWR VGND fanout181/X fanout182/X VGND VPWR sky130_fd_sc_hd__buf_6
XFILLER_18_290 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1205_ VPWR VGND _1205_/A _1206_/A _1471_/A VGND VPWR sky130_fd_sc_hd__and2_2
X_1136_ VPWR VGND _1255_/A _1471_/A VGND VPWR sky130_fd_sc_hd__buf_6
X_1067_ _1678_/Q _1679_/Q _1062_/B _1067_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o21a_2
XFILLER_0_304 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_53 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_63 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1685_ _1685_/Q fanout170/X _1685_/D _1748_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1754_ _1754_/Q fanout180/X _1754_/D _1758_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1119_ _1138_/B _1122_/A _1119_/B _1119_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__nand3_4
XFILLER_12_230 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_67 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_289 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1470_ VPWR VGND _1778_/A _1470_/A VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_35_300 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1806_ VGND VPWR _1806_/X _1806_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1737_ _1737_/Q fanout172/X _1737_/D _1742_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1599_ _1563_/X _1598_/X _1597_/X _1604_/A _1599_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o211a_2
X_1668_ _1668_/Q fanout172/X _1668_/D _1765_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_5_237 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0970_ _0969_/X _1073_/A _0912_/A _0836_/X _0946_/A _0970_/X VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__o32a_2
X_1453_ _1453_/B _1693_/D _1683_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_4_270 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1522_ VGND VPWR _1524_/S _1700_/Q _1699_/Q _1523_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_1384_ _1721_/Q _1767_/Q _1385_/B _1768_/Q _1722_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__a22o_2
XPHY_20 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_163 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_53 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_74 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_75 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_244 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xoutput114 VPWR VGND pmatrix_row_out_n[12] _1803_/A VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput125 VPWR VGND pmatrix_row_out_n[8] _1799_/A VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput103 VPWR VGND pmatrix_col_out_n[30] _1247_/X VGND VPWR sky130_fd_sc_hd__buf_4
X_0884_ VGND VPWR _1668_/Q _0883_/X _0881_/X _0884_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_0953_ _1101_/B _0953_/X _0980_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
Xoutput158 VPWR VGND sample_matrix_out _1808_/A VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput136 VPWR VGND pmatrix_rowon_out_n[4] _1796_/X VGND VPWR sky130_fd_sc_hd__buf_4
X_1436_ VGND VPWR _1437_/B _1687_/Q _1688_/Q VGND VPWR sky130_fd_sc_hd__xnor2_2
Xoutput147 VPWR VGND result_out[14] _1747_/Q VGND VPWR sky130_fd_sc_hd__buf_4
X_1505_ VGND VPWR _1507_/S input4/X _1668_/Q _1506_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_1367_ _1367_/B _1367_/X _1720_/Q _1367_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
X_1298_ _1256_/Y _1132_/X _1292_/B _1221_/B _1273_/A _1298_/X VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__o32a_2
X_1221_ _1221_/B _1230_/A _1221_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1152_ _1205_/A _1276_/B _1153_/B _1152_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__or3_2
X_1083_ _1083_/B _1083_/Y _1083_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_20_136 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_291 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0936_ _0936_/X _0908_/B _1062_/B _1671_/Q _0908_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__o31a_2
X_0867_ _1076_/A _1026_/B _0867_/X _1027_/D _1084_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_2
X_0798_ _0797_/X _0796_/X _0789_/X _1753_/Q _0798_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o211a_2
X_1419_ VGND VPWR _1420_/B _1728_/Q _1432_/C VGND VPWR sky130_fd_sc_hd__xnor2_2
XFILLER_51_261 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xfanout171 VPWR VGND fanout171/X fanout183/X VGND VPWR sky130_fd_sc_hd__buf_2
Xfanout182 VPWR VGND fanout182/X fanout183/X VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_47_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1770_ _1770_/Q fanout176/X _1770_/D _1770_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_42_272 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1204_ _1169_/A _1183_/X _1203_/X _1204_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_2
XFILLER_33_3 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1066_ _1809_/A _1065_/Y _1101_/B _1679_/Q _1679_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__o211a_2
X_1135_ _1205_/A _1217_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
X_0919_ _0920_/A _0919_/B _0919_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__xor2_4
XFILLER_17_10 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_154 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_198 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1753_ _1753_/Q fanout178/X _1753_/D _1763_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1684_ _1684_/Q fanout170/X _1684_/D _1748_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1049_ _1049_/A _1049_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
X_1118_ _1119_/C _1119_/B _1138_/A _1122_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_0_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_224 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_242 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1805_ VGND VPWR _1805_/X _1805_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1736_ _1736_/Q fanout171/X _1736_/D _1742_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1598_ _1719_/D _1598_/X _1725_/D _1620_/A _1615_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__o22a_2
X_1667_ _1667_/Q fanout172/X _1667_/D _1765_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_5_205 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_249 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_10 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_41 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1452_ VGND VPWR _1453_/B _1693_/Q _1454_/B VGND VPWR sky130_fd_sc_hd__xnor2_2
XFILLER_4_282 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1383_ VPWR VGND _1383_/X _1382_/Y _1401_/A _1402_/C _1402_/D VGND VPWR sky130_fd_sc_hd__and4b_2
X_1521_ VGND VPWR _1698_/D _1521_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_50_156 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1719_ _1719_/Q fanout173/X _1719_/D _1743_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XPHY_10 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_43 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_54 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_145 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_76 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_53 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_164 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_256 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0952_ _1173_/A _1127_/B _1127_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__xor2_4
Xoutput159 VPWR VGND sample_matrix_out_n _1807_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput115 VPWR VGND pmatrix_row_out_n[13] _1804_/A VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput126 VPWR VGND pmatrix_row_out_n[9] _1800_/A VGND VPWR sky130_fd_sc_hd__buf_4
X_1504_ VGND VPWR _1667_/D _1504_/A VGND VPWR sky130_fd_sc_hd__buf_1
Xoutput104 VPWR VGND pmatrix_col_out_n[31] _1249_/Y VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput148 VPWR VGND result_out[15] _1748_/Q VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput137 VPWR VGND pmatrix_rowon_out_n[5] _1797_/X VGND VPWR sky130_fd_sc_hd__buf_4
X_0883_ VGND VPWR _1669_/Q input2/X _0882_/X _0883_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_1435_ _1687_/D _1687_/Q _1435_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1366_ _1720_/Q _1367_/C _1367_/B _1366_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_2
XFILLER_23_134 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1297_ VGND VPWR _1248_/X _1233_/A _1237_/Y _1297_/X _1265_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_2
X_1220_ _1209_/X _1220_/Y _1152_/C _1144_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o21ai_2
X_1151_ _1152_/C _1151_/B _1151_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_45_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_270 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1082_ _1116_/A _1117_/S _1061_/B _1061_/C _1081_/X _1083_/B VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__o41a_2
X_0866_ VPWR VGND _1076_/A _0866_/A VGND VPWR sky130_fd_sc_hd__buf_6
X_0935_ _0938_/A _0935_/A _0935_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_4
X_0797_ _0831_/C _1669_/Q _0797_/X _1752_/Q _1668_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__or4b_2
X_1418_ _1727_/Q _1432_/C _1726_/Q _1418_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
X_1349_ VPWR VGND _1350_/B _1349_/B _1714_/Q VGND VPWR sky130_fd_sc_hd__xor2_2
XFILLER_51_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_108 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xfanout172 VPWR VGND fanout172/X fanout173/X VGND VPWR sky130_fd_sc_hd__buf_6
Xfanout183 VPWR VGND fanout183/X input9/X VGND VPWR sky130_fd_sc_hd__buf_4
X_1134_ _1133_/Y _1134_/Y _1129_/X _1237_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__o21ai_2
X_1203_ VPWR VGND _1203_/X _1203_/A VGND VPWR sky130_fd_sc_hd__buf_4
X_1065_ _1065_/Y _1101_/B _1496_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_0849_ _0859_/B _0875_/C _0849_/A _0875_/D _0849_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_4
X_0918_ VPWR VGND _0918_/A _0919_/B _0918_/B VGND VPWR sky130_fd_sc_hd__and2_2
X_1683_ _1683_/Q fanout174/X _1683_/D _1462_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1752_ _1752_/Q fanout178/X _1752_/D _1763_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_30_232 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1117_ VGND VPWR _1116_/Y _1115_/X _1117_/S _1119_/C VGND VPWR sky130_fd_sc_hd__mux2_2
X_1048_ _1048_/B _1049_/A _1677_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_48_107 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_64 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_236 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_265 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1735_ _1735_/Q fanout170/X _1735_/D _1748_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1666_ VGND VPWR _1770_/D _1666_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1804_ VGND VPWR _1804_/X _1804_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1597_ VGND VPWR _1626_/S _1723_/D _1721_/D _1597_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_67 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_53 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1520_ VGND VPWR _1524_/S _1699_/Q _1698_/Q _1521_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_1451_ _1692_/Q _1454_/B _1691_/Q _1451_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
XFILLER_4_294 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1382_ _1382_/Y _1382_/A _1382_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
XFILLER_2_209 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1718_ _1718_/Q fanout172/X _1718_/D _1743_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1649_ VGND VPWR _1663_/B _1762_/Q _1673_/D _1650_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XPHY_11 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_99 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_55 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_124 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_98 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_275 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_176 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_268 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0882_ VGND VPWR _1667_/Q _1757_/Q _1756_/Q _0882_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_0951_ _0935_/B _0938_/B _0931_/A _1127_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__o21a_4
Xoutput116 VPWR VGND pmatrix_row_out_n[14] _1805_/A VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput149 VPWR VGND result_out[1] _1734_/Q VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput127 VPWR VGND pmatrix_rowon_out_n[0] _1792_/X VGND VPWR sky130_fd_sc_hd__buf_4
X_1503_ VGND VPWR _1507_/S input3/X _1667_/Q _1504_/A VGND VPWR sky130_fd_sc_hd__mux2_1
Xoutput138 VPWR VGND pmatrix_rowon_out_n[6] _1798_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput105 VPWR VGND pmatrix_col_out_n[3] _1154_/X VGND VPWR sky130_fd_sc_hd__buf_4
X_1434_ _1434_/B _1732_/D _1514_/S VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1365_ _1765_/Q _1367_/C _1331_/B _1719_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__o21ai_2
X_1296_ _1209_/X _1235_/Y _1239_/X _1255_/A _1296_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o211a_2
XFILLER_23_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_10 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1150_ VPWR VGND _1233_/A _1287_/B VGND VPWR sky130_fd_sc_hd__buf_6
XFILLER_52_219 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1081_ _1093_/B _1078_/Y _1081_/X _1080_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o21ba_2
XFILLER_9_194 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0865_ _1013_/B _0865_/C _1013_/A _0865_/D _0866_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_4
X_0934_ _0933_/X _1672_/Q _0980_/D _0935_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__o21a_2
X_1417_ _1417_/B _1727_/D _1420_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_0796_ _1752_/Q _0831_/C _0796_/X _0789_/X _0795_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__a22o_2
X_1348_ _1349_/B _1713_/Q _1759_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1279_ _1175_/X _1169_/A _1265_/Y _1279_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o21a_2
Xfanout173 VPWR VGND fanout173/X fanout183/X VGND VPWR sky130_fd_sc_hd__buf_4
Xfanout162 _1100_/X _1784_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__buf_12
Xfanout184 VPWR VGND _1765_/CLK _1763_/CLK VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_6_120 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_197 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1064_ _1496_/A _1064_/B _1064_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__xnor2_4
X_1133_ _1132_/X _1133_/Y _1256_/A _1270_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__o21ai_2
X_1202_ VPWR VGND _1252_/A _1203_/A _1265_/B VGND VPWR sky130_fd_sc_hd__and2_2
XFILLER_33_274 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0779_ _0779_/X _1584_/S _1633_/A _0778_/X _1693_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__o31a_2
X_0848_ VGND VPWR _0875_/D _1698_/Q _1702_/Q VGND VPWR sky130_fd_sc_hd__xnor2_2
X_0917_ _0918_/B _1671_/Q _0917_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
XFILLER_15_252 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1682_ _1682_/Q fanout172/X _1682_/D _1765_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1751_ _1751_/Q fanout178/X _1751_/D _1765_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1047_ _1061_/C _1047_/Y _1116_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1116_ _1116_/Y _1116_/A _1116_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
XFILLER_28_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_248 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_277 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1803_ VGND VPWR _1803_/X _1803_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_7_281 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1734_ _1734_/Q fanout170/X _1734_/D _1748_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1596_ _1596_/B _1596_/X _1741_/Q _1596_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
X_1665_ VGND VPWR _1665_/S _1770_/Q _1681_/D _1666_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_38_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_188 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_10 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1450_ _1448_/Y _1435_/B _1449_/X _1692_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__o21a_2
X_1381_ _1401_/A _1385_/A _1381_/A _1381_/B _1381_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__and4_2
X_1579_ _1569_/B _1716_/D _1579_/X _1722_/D _1563_/A _1620_/A VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__o221a_2
X_1717_ _1717_/Q fanout172/X _1717_/D _1743_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1648_ VGND VPWR _1761_/D _1648_/A VGND VPWR sky130_fd_sc_hd__buf_1
XPHY_12 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_89 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_221 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_214 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_0881_ VGND VPWR _0881_/S _1758_/Q input2/X _0881_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_0950_ _0949_/Y _0948_/X _0980_/C _1127_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_4
Xoutput128 VPWR VGND pmatrix_rowon_out_n[10] _1802_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput117 VPWR VGND pmatrix_row_out_n[15] _1806_/A VGND VPWR sky130_fd_sc_hd__buf_4
X_1433_ VGND VPWR _1434_/B _1732_/Q _1433_/B VGND VPWR sky130_fd_sc_hd__xnor2_2
Xoutput106 VPWR VGND pmatrix_col_out_n[4] _1156_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput139 VPWR VGND pmatrix_rowon_out_n[7] _1799_/X VGND VPWR sky130_fd_sc_hd__buf_4
X_1502_ VPWR VGND _1806_/A _1502_/A VGND VPWR sky130_fd_sc_hd__buf_2
X_1364_ VPWR VGND _1718_/D _1364_/A VGND VPWR sky130_fd_sc_hd__buf_2
X_1295_ _1270_/B _1248_/X _1295_/X _1132_/X _1234_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__a22o_2
XFILLER_39_291 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1080_ _1080_/X _1061_/B _1076_/X _1079_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
XFILLER_52_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0864_ _1712_/Q _1705_/Q _0865_/D _1704_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__or3_2
X_0933_ _0933_/B _0933_/X _1707_/Q _0933_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
X_0795_ _0795_/Y _1667_/Q _1669_/Q _1668_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__nand3b_2
X_1416_ VPWR VGND _1417_/B _1416_/B _1727_/Q VGND VPWR sky130_fd_sc_hd__xor2_2
X_1347_ _1721_/D _1347_/B _1767_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__xnor2_4
X_1278_ _1277_/X _1276_/X _1164_/X _1175_/X _1278_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o211a_2
XFILLER_22_68 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xfanout174 VPWR VGND fanout174/X fanout177/X VGND VPWR sky130_fd_sc_hd__buf_6
Xfanout163 VPWR VGND _1748_/CLK _1742_/CLK VGND VPWR sky130_fd_sc_hd__buf_4
Xfanout185 VPWR VGND _1766_/CLK _1763_/CLK VGND VPWR sky130_fd_sc_hd__buf_2
X_1201_ _1164_/X _1165_/X _1201_/X _1179_/B _1256_/A _1287_/A VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__o221a_2
X_1132_ VPWR VGND _1132_/X _1276_/C VGND VPWR sky130_fd_sc_hd__buf_6
X_1063_ _1122_/A _1061_/Y _1093_/B _1040_/S _1064_/B _1052_/X VPWR VGND VGND VPWR
+ sky130_fd_sc_hd__a221o_4
X_0916_ _1062_/B _0916_/B _0917_/B _0916_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__or3_2
X_0778_ _0778_/X _1560_/A _0776_/X _0777_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
X_0847_ _1697_/Q _1699_/Q _0875_/C _1703_/Q _1808_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_2
XFILLER_17_79 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_34 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_231 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1750_ _1750_/Q fanout178/X _1750_/D _1765_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1681_ _1681_/Q fanout181/X _1681_/D _1770_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_31_3 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_304 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1046_ _1190_/A _1046_/B _1016_/A _1061_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__or3b_4
X_1115_ _1115_/A _1116_/A _1061_/C _1115_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__or3b_2
XFILLER_12_289 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_315 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1802_ VGND VPWR _1802_/X _1802_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1733_ _1733_/Q fanout170/X _1733_/D _1748_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_7_293 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1595_ _1740_/D _1592_/X _1762_/Q _1593_/Y _1640_/B VGND VPWR _1594_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_2
X_1664_ _1507_/S _1769_/D _1663_/Y _1663_/B _1072_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__o31ai_2
X_1029_ _1046_/B _1025_/X _1024_/X _1029_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_2
XFILLER_29_153 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_175 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1380_ _1381_/D _1722_/Q _1768_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1716_ _1716_/Q fanout173/X _1716_/D _1742_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1578_ _1737_/D _1573_/X _1759_/Q _1575_/X _1640_/B VGND VPWR _1577_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_2
X_1647_ VGND VPWR _1663_/B _1761_/Q _1672_/D _1648_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XPHY_13 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_255 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xoutput107 VPWR VGND pmatrix_col_out_n[5] _1162_/X VGND VPWR sky130_fd_sc_hd__buf_4
X_0880_ VPWR VGND _0881_/S _1669_/Q _1667_/Q VGND VPWR sky130_fd_sc_hd__and2b_2
X_1432_ _1433_/B _1432_/C _1728_/Q _1729_/Q _1432_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__and4_2
X_1363_ _1364_/A _1362_/Y _1361_/Y _1602_/A _1410_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_2
Xoutput118 VPWR VGND pmatrix_row_out_n[1] _1792_/A VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput129 VPWR VGND pmatrix_rowon_out_n[11] _1803_/X VGND VPWR sky130_fd_sc_hd__buf_4
X_1501_ _1803_/A _1502_/A _1501_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
X_1294_ _1132_/X _1237_/A _1294_/X _1248_/X _1129_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__a22o_2
X_0932_ _0990_/A _0933_/C _1073_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_9_163 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0863_ _1706_/Q _1013_/B _1707_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
X_0794_ _1751_/Q _1750_/Q _1749_/Q _0831_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__and3_4
X_1415_ _1416_/B _1726_/Q _1418_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1346_ _1420_/A _1347_/B _1346_/B _1346_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__or3_4
X_1277_ _1277_/X _1144_/X _1210_/Y _1265_/A _1265_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_2
Xfanout164 VPWR VGND _1742_/CLK _1721_/CLK VGND VPWR sky130_fd_sc_hd__buf_4
Xfanout175 VPWR VGND fanout175/X fanout177/X VGND VPWR sky130_fd_sc_hd__buf_6
Xfanout186 VPWR VGND _1763_/CLK _1707_/CLK VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_6_155 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1200_ _1183_/X _1198_/X _1292_/A _1200_/Y _1199_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__a211oi_4
X_1131_ _1131_/A _1256_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__buf_8
X_1062_ VPWR VGND _1678_/Q _1093_/B _1062_/B VGND VPWR sky130_fd_sc_hd__and2_2
X_0915_ _0915_/B _0916_/C _0929_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_0777_ _0777_/Y _1580_/S _1693_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_0846_ _0859_/B _1073_/C _1005_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__or2_4
X_1329_ _1331_/B _1328_/X _1382_/A _1402_/C _1402_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_2
X_1680_ _1680_/Q fanout181/X _1680_/D _1769_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1114_ VGND VPWR _1113_/Y _1112_/Y _1117_/S _1119_/B VGND VPWR sky130_fd_sc_hd__mux2_2
X_1045_ _1061_/B _1062_/B _1678_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__xnor2_4
X_0829_ _1753_/Q _0831_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_28_68 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_121 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1801_ VGND VPWR _1801_/X _1801_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_7_261 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1732_ _1732_/Q fanout174/X _1732_/D _1745_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1663_ _1663_/Y _1769_/Q _1663_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1594_ _1596_/B _1594_/X _1740_/Q _1615_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
XFILLER_53_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1028_ VGND VPWR _1046_/B _1677_/Q _1048_/B VGND VPWR sky130_fd_sc_hd__xnor2_2
XFILLER_30_36 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_58 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_165 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_93 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1715_ _1715_/Q fanout175/X _1715_/D _1746_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1646_ VGND VPWR _1760_/D _1646_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1577_ _1596_/B _1577_/X _1737_/Q _1596_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
XPHY_14 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_57 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_160 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1500_ _1778_/A _1805_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
Xoutput119 VPWR VGND pmatrix_row_out_n[2] _1793_/A VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput108 VPWR VGND pmatrix_col_out_n[6] _1166_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput90 VPWR VGND pmatrix_col_out_n[19] _1219_/Y VGND VPWR sky130_fd_sc_hd__buf_4
X_1431_ VPWR VGND _1730_/Q _1432_/D _1731_/Q VGND VPWR sky130_fd_sc_hd__and2_2
X_1362_ _1602_/A _1361_/Y _1410_/B _1362_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_2
X_1293_ VGND VPWR _1293_/X _1293_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_11_49 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1629_ VPWR VGND _1768_/Q _1629_/X _1640_/B VGND VPWR sky130_fd_sc_hd__and2_2
XFILLER_52_56 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0862_ _1050_/B _1027_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
X_0931_ _0931_/A _0935_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
X_0793_ _0793_/X _0792_/X _0791_/X _1752_/Q _1751_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__a211o_2
X_1414_ _1414_/B _1726_/D _1514_/S VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1345_ VPWR VGND _1721_/Q _1346_/C _1371_/B VGND VPWR sky130_fd_sc_hd__and2_2
X_1276_ _1276_/A _1276_/B _1276_/X _1276_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__or3_2
Xfanout165 VGND VPWR _1743_/CLK _1721_/CLK VGND VPWR sky130_fd_sc_hd__buf_1
Xfanout176 VPWR VGND fanout176/X fanout177/X VGND VPWR sky130_fd_sc_hd__buf_4
Xfanout187 VPWR VGND _1758_/CLK _1707_/CLK VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_10_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1130_ VPWR VGND _1270_/B _1130_/A VGND VPWR sky130_fd_sc_hd__buf_6
X_1061_ _1061_/C _1061_/Y _1116_/A _1061_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nor3_2
X_0845_ _1712_/Q _1005_/B _1711_/Q _1710_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__or3_4
X_0914_ _1013_/A _1013_/C _0915_/B _0914_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__or3_2
X_0776_ _1684_/Q _1693_/Q _1691_/Q _0776_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__or3b_2
X_1259_ _1259_/X _1292_/A _1178_/B _1258_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
X_1328_ VPWR VGND _1328_/A _1328_/X _1328_/B VGND VPWR sky130_fd_sc_hd__and2_2
XFILLER_15_244 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_181 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1113_ _1113_/Y _1113_/A _1115_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1044_ _1044_/B _1677_/D _1507_/S VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_0759_ _1580_/S _1691_/Q _1686_/Q _0759_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o21a_2
X_0828_ _0828_/B _1752_/D _1538_/S VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_18_80 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1800_ VGND VPWR _1800_/X _1800_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1731_ _1731_/Q fanout177/X _1731_/D _1462_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_7_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1662_ VGND VPWR _1768_/D _1662_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1593_ _1593_/Y _1593_/A _1593_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
XFILLER_53_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1027_ _1058_/A _1076_/A _1027_/D _1048_/B _1050_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__and4bb_4
XFILLER_44_103 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_221 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_61 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1714_ _1714_/Q fanout174/X _1714_/D _1745_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1576_ VPWR VGND _1596_/B _1602_/B VGND VPWR sky130_fd_sc_hd__buf_4
X_1645_ VGND VPWR _1663_/B _1760_/Q _1671_/D _1646_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XPHY_15 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1430_ _1430_/B _1731_/D _1514_/S VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
Xoutput109 VPWR VGND pmatrix_col_out_n[7] _1172_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput80 VPWR VGND pmatrix_col_out_n[0] _1124_/X VGND VPWR sky130_fd_sc_hd__buf_4
X_1361_ VGND VPWR _1361_/Y _1718_/Q _1361_/B VGND VPWR sky130_fd_sc_hd__xnor2_2
X_1292_ _1292_/A _1292_/B _1293_/A _1292_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__or3_2
Xoutput91 VPWR VGND pmatrix_col_out_n[1] _1134_/Y VGND VPWR sky130_fd_sc_hd__buf_4
X_1559_ _1559_/B _1561_/A _1584_/S VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1628_ _1561_/A _1628_/X _1593_/A _1569_/B _1730_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__o2bb2a_2
XFILLER_10_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_128 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0861_ VPWR VGND _1050_/B _1709_/Q VGND VPWR sky130_fd_sc_hd__buf_6
X_0930_ _1672_/Q _0980_/D _0931_/A _0975_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__or3_2
X_0792_ _0885_/S _0792_/X _1750_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
X_1413_ VGND VPWR _1414_/B _1726_/Q _1418_/C VGND VPWR sky130_fd_sc_hd__xnor2_2
XFILLER_3_84 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1344_ _1371_/B _1346_/B _1721_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1275_ _1275_/X _1183_/X _1157_/Y _1195_/X _1248_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__a211o_2
XFILLER_11_109 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xfanout166 VPWR VGND _1745_/CLK _1721_/CLK VGND VPWR sky130_fd_sc_hd__buf_4
Xfanout177 VPWR VGND fanout177/X fanout183/X VGND VPWR sky130_fd_sc_hd__buf_4
Xfanout188 VPWR VGND _1707_/CLK input1/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_47_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_29 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1060_ _1122_/A _1062_/B _1678_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__xor2_4
X_0775_ _0775_/A _0775_/B _0774_/X _0785_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__or3b_2
X_0913_ _1012_/B _1073_/C _1705_/Q _1005_/B _0929_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_4
X_0844_ _1073_/C _1708_/Q _1709_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__or2_4
X_1327_ _1763_/Q _1717_/Q _1328_/B _1718_/Q _1764_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__a22o_2
X_1189_ VGND VPWR _1189_/X _1189_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1258_ _1258_/A _1258_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_3_127 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1112_ _1112_/Y _1116_/A _1115_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1043_ VGND VPWR _1043_/S _1276_/B _1050_/C _1044_/B VGND VPWR sky130_fd_sc_hd__mux2_1
X_0758_ VPWR VGND _1580_/S _1684_/Q VGND VPWR sky130_fd_sc_hd__buf_4
X_0827_ VGND VPWR _0828_/B _1752_/Q _0831_/C VGND VPWR sky130_fd_sc_hd__xnor2_2
XFILLER_28_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_304 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_315 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1730_ _1730_/Q fanout177/X _1730_/D _1462_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_11_281 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1592_ _1592_/X _1560_/A _1559_/B _1591_/X _1722_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__o31a_2
X_1661_ VGND VPWR _1665_/S _1768_/Q _1679_/D _1662_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_1026_ VGND VPWR _1050_/D _1058_/B _1026_/B VGND VPWR sky130_fd_sc_hd__xnor2_2
XFILLER_38_156 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_192 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_233 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1713_ _1713_/Q fanout175/X _1713_/D _1746_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1575_ _1575_/B _1575_/X _1604_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
X_1644_ VGND VPWR _1759_/D _1644_/A VGND VPWR sky130_fd_sc_hd__buf_1
XPHY_16 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1009_ _1675_/Q _1010_/B _1008_/Y _0993_/A _0993_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__o2bb2a_2
XFILLER_1_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_184 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xoutput70 VPWR VGND nmatrix_rowon_out_n[3] _1780_/X VGND VPWR sky130_fd_sc_hd__buf_4
X_1360_ _1359_/X _1358_/X _1763_/Q _1361_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_2
Xoutput92 VPWR VGND pmatrix_col_out_n[20] _1222_/X VGND VPWR sky130_fd_sc_hd__buf_4
X_1291_ _1292_/C _1151_/A _1246_/B _1221_/B _1246_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__o31a_2
Xoutput81 VPWR VGND pmatrix_col_out_n[10] _1189_/X VGND VPWR sky130_fd_sc_hd__buf_4
X_1558_ _1559_/B _1580_/S _1558_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1627_ _1585_/B _1627_/Y _1626_/X _1514_/S VGND VPWR VGND VPWR sky130_fd_sc_hd__o21ai_2
X_1489_ _1788_/A _1490_/A _1497_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
XFILLER_52_36 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_81 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_122 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_195 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0860_ VPWR VGND _1026_/B _1708_/Q VGND VPWR sky130_fd_sc_hd__buf_4
X_0791_ _0791_/X _1749_/Q _1750_/Q _0885_/S VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
X_1412_ VPWR VGND _1514_/S _1420_/A VGND VPWR sky130_fd_sc_hd__buf_6
X_1343_ _1371_/B _1382_/B _1382_/A _1402_/D _1402_/C _1342_/X VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__a41o_4
X_1274_ _1198_/X _1183_/X _1274_/X _1169_/A _1273_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__a22o_2
X_0989_ VGND VPWR _1005_/C _0989_/A _1707_/Q VGND VPWR sky130_fd_sc_hd__xnor2_2
Xfanout167 VGND VPWR _1462_/A _1721_/CLK VGND VPWR sky130_fd_sc_hd__buf_1
Xfanout189 VPWR VGND _1769_/CLK _1770_/CLK VGND VPWR sky130_fd_sc_hd__buf_2
Xfanout178 VPWR VGND fanout178/X fanout180/X VGND VPWR sky130_fd_sc_hd__buf_6
XFILLER_27_243 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_276 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_298 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_136 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0912_ _0912_/B _0916_/B _0912_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_0774_ _1558_/B _1685_/Q _0774_/X _1684_/Q _1695_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_2
X_0843_ _0849_/A _1702_/Q _0843_/X _1084_/A _1058_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_2
X_1326_ _1382_/A _1326_/C _1328_/A _1326_/B _1326_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__and4_2
X_1257_ _1255_/Y _1257_/X _1256_/Y _1273_/A _1233_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__o22a_2
X_1188_ VPWR VGND _1189_/A _1188_/B _1186_/X VGND VPWR sky130_fd_sc_hd__and2b_2
XFILLER_47_305 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_249 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1042_ VPWR VGND _1276_/B _1184_/B VGND VPWR sky130_fd_sc_hd__buf_6
X_1111_ _1122_/A _1111_/D _1111_/C _1111_/B _1158_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__nand4_4
X_0757_ _1685_/Q _1560_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
X_0826_ _0826_/B _1751_/D _1538_/S VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1309_ _1715_/Q _1310_/C _1310_/B _1311_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_2
XFILLER_44_15 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_293 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1591_ _1586_/B _1718_/D _1591_/X _1720_/D _1563_/A _1565_/A VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__o221a_2
X_1660_ VGND VPWR _1767_/D _1660_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_38_135 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1025_ _1025_/B _1025_/X _1033_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
X_0809_ VPWR VGND _0810_/B _0809_/B _1755_/Q VGND VPWR sky130_fd_sc_hd__xor2_2
X_1789_ VGND VPWR _1789_/X _1789_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_29_113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_116 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1 _1243_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_1712_ _1712_/Q fanout179/X _1712_/D _1766_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1643_ VGND VPWR _1663_/B _1759_/Q _1670_/D _1644_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_1574_ VGND VPWR _1580_/S _1719_/D _1717_/D _1575_/B VGND VPWR sky130_fd_sc_hd__mux2_1
XPHY_17 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1008_ _1008_/Y _1008_/A _1106_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
XFILLER_41_38 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xoutput71 VPWR VGND nmatrix_rowon_out_n[4] _1781_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput93 VPWR VGND pmatrix_col_out_n[21] _1226_/Y VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput82 VPWR VGND pmatrix_col_out_n[11] _1193_/Y VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput60 VPWR VGND nmatrix_row_out_n[8] _1100_/X VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_0_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1290_ _1164_/X _1221_/B _1290_/X _1169_/A _1229_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__a22o_2
XFILLER_48_230 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1626_ VGND VPWR _1626_/S _1420_/B _1414_/B _1626_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_1557_ _1640_/B _1555_/X _1551_/Y _1733_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_2
X_1488_ VPWR VGND _1788_/A _1488_/A VGND VPWR sky130_fd_sc_hd__buf_6
XFILLER_52_48 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_244 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_0790_ _1668_/Q _1669_/Q _1667_/Q _0885_/S VPWR VGND VGND VPWR sky130_fd_sc_hd__or3b_2
X_1411_ VPWR VGND _1725_/D _1411_/A VGND VPWR sky130_fd_sc_hd__buf_2
X_1273_ _1273_/A _1276_/A _1273_/X _1287_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__or3_2
X_1342_ VPWR VGND _1403_/A _1342_/X _1403_/B VGND VPWR sky130_fd_sc_hd__and2_2
XFILLER_51_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0988_ _1675_/Q _1004_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
X_1609_ VGND VPWR _1626_/S _1725_/D _1723_/D _1609_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xfanout168 VPWR VGND _1746_/CLK _1721_/CLK VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_27_200 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xfanout179 VPWR VGND fanout179/X fanout180/X VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_10_188 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_0842_ _1712_/Q _1058_/C _1708_/Q _1709_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__or3_4
X_0911_ _0910_/X _1013_/C _0909_/Y _0899_/B _1703_/Q _0912_/B VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__o32a_2
XFILLER_33_247 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_0773_ _0775_/A _1584_/S _1580_/S _1695_/Q _1558_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__o31a_2
X_1325_ _1717_/Q _1326_/D _1763_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
X_1256_ _1258_/A _1256_/Y _1256_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1187_ _1144_/X _1188_/B _1237_/B _1178_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__o21ai_2
XFILLER_3_107 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1110_ _1122_/A _1111_/C _1111_/D _1111_/B _1158_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_4
X_1041_ _1040_/X _1184_/B _1034_/Y _1029_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__o21ai_2
X_0825_ VPWR VGND _0826_/B _0825_/B _1751_/Q VGND VPWR sky130_fd_sc_hd__xor2_2
X_0756_ input7/X input8/X input6/X _1607_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nor3_4
X_1308_ _1310_/C _1714_/Q _1759_/Q _1760_/Q _1713_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_2
X_1239_ _1265_/A _1221_/A _1265_/B _1239_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o21a_2
XFILLER_47_158 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_261 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1590_ _1739_/D _1589_/X _1563_/X _1587_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
XFILLER_50_70 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1024_ _1024_/X _1676_/Q _1033_/B _1025_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
X_1788_ VGND VPWR _1788_/X _1788_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_0808_ _0809_/B _1754_/Q input2/X VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
XFILLER_6_75 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1642_ _1748_/D _1641_/X _1639_/X _1563_/X _1638_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_2
XANTENNA_2 _1172_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_1711_ _1711_/Q fanout182/X _1711_/D _1770_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1573_ _1569_/B _1715_/D _1573_/X _1721_/D _1563_/A _1620_/A VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__o221a_2
XPHY_18 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1007_ _1106_/A _1007_/A _1007_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_1_205 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_305 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_40 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_84 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xoutput61 VPWR VGND nmatrix_row_out_n[9] _1785_/A VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput72 VPWR VGND nmatrix_rowon_out_n[5] _1782_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput83 VPWR VGND pmatrix_col_out_n[12] _1197_/Y VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput94 VPWR VGND pmatrix_col_out_n[22] _1228_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput50 VPWR VGND nmatrix_row_out_n[13] _1789_/A VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_48_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1625_ _1745_/D _1624_/X _1622_/X _1563_/X _1620_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_2
X_1556_ VPWR VGND _1640_/B _1607_/B VGND VPWR sky130_fd_sc_hd__buf_4
X_1487_ _1487_/B _1488_/A _1487_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
XFILLER_22_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_146 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_131 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1410_ VGND VPWR _1410_/B _1411_/A _1418_/C _1410_/C VGND VPWR sky130_fd_sc_hd__and3b_2
XFILLER_3_10 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1341_ _1338_/A _1340_/X _1403_/B _1339_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__a21bo_2
X_1272_ _1188_/B _1196_/X _1272_/X _1276_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__a21bo_2
XFILLER_51_215 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_237 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0987_ _0987_/B _1674_/D _1507_/S VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1608_ _1596_/B _1612_/A _1563_/X _1765_/Q _1607_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o22a_2
X_1539_ VGND VPWR _1707_/D _1539_/A VGND VPWR sky130_fd_sc_hd__buf_1
Xfanout169 VPWR VGND _1721_/CLK _1682_/Q VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_27_212 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_85 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_93 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_0772_ _1558_/B _1686_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_4
X_0841_ _1073_/B _0849_/A _0946_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
X_0910_ _1700_/Q _1701_/Q _1703_/Q _0910_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__or3b_2
X_1255_ _1255_/B _1255_/Y _1255_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1324_ _1326_/C _1763_/Q _1717_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1186_ _1186_/X _1292_/A _1130_/A _1183_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
XFILLER_31_9 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1040_ VGND VPWR _1040_/S _1039_/X _1037_/X _1040_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_0824_ _0825_/B _1750_/Q _1749_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1307_ _1310_/B _1760_/Q _1713_/Q _1759_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
X_1169_ _1233_/A _1169_/Y _1169_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1238_ _1256_/A _1238_/X _1237_/Y _1140_/X _1233_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__o22a_2
XFILLER_12_218 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_60 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_192 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1023_ _1022_/X _1106_/A _1008_/A _1025_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_2
X_1787_ VGND VPWR _1787_/X _1787_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_0807_ VPWR VGND _1538_/S _1548_/S VGND VPWR sky130_fd_sc_hd__buf_6
XFILLER_4_258 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_3 _1802_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_1572_ _1736_/Q _1435_/B _1736_/D _1571_/X _1569_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__a22o_2
X_1641_ _1641_/X _1640_/X _1596_/C _1748_/Q _1596_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_2
X_1710_ _1710_/Q fanout182/X _1710_/D _1770_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XPHY_19 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_107 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1006_ _0927_/X _1076_/A _1005_/X _0990_/A _1073_/A _1008_/A VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__o32a_2
XFILLER_15_52 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xoutput73 VPWR VGND nmatrix_rowon_out_n[6] _1783_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput95 VPWR VGND pmatrix_col_out_n[23] _1231_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput84 VPWR VGND pmatrix_col_out_n[13] _1200_/Y VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput40 VPWR VGND nmatrix_col_out_n[3] _1257_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput51 VPWR VGND nmatrix_row_out_n[14] _1790_/A VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput62 VPWR VGND nmatrix_rowon_out_n[0] _1777_/X VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_48_265 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1555_ _1615_/A _1569_/B _1717_/D _1555_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__or3b_2
X_1624_ _1624_/X _1623_/X _1596_/C _1745_/Q _1596_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_2
X_1486_ _1796_/A _1787_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_9_169 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_22 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1340_ _1340_/X _1719_/Q _1328_/A _1328_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
X_1271_ _1144_/X _1252_/X _1292_/A _1183_/X _1271_/X _1270_/Y VPWR VGND VGND VPWR
+ sky130_fd_sc_hd__a221o_4
XFILLER_51_249 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0986_ VGND VPWR _1101_/B _1151_/B _1014_/B _0987_/B VGND VPWR sky130_fd_sc_hd__mux2_1
X_1469_ _1784_/A _1470_/A _1496_/A _1487_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
X_1607_ _1607_/B _1607_/X _1743_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
X_1538_ VGND VPWR _1538_/S _1026_/B _1707_/Q _1539_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_10_135 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0771_ VPWR VGND _1584_/S _1685_/Q VGND VPWR sky130_fd_sc_hd__buf_6
X_0840_ _1704_/Q _1707_/Q _1705_/Q _1706_/Q _1073_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_5_194 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1323_ _1326_/B _1764_/Q _1718_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
XFILLER_38_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1185_ VPWR VGND _1292_/A _1185_/A VGND VPWR sky130_fd_sc_hd__buf_4
X_1254_ _1175_/X _1253_/Y _1252_/X _1237_/A _1254_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o211a_2
X_0969_ _1073_/B _1026_/B _0969_/X _1027_/D _1005_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_2
XFILLER_2_197 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_71 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_10 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_219 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0823_ _0823_/B _1750_/D _1538_/S VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1306_ VGND VPWR _1713_/D _1759_/Q _1306_/B VGND VPWR sky130_fd_sc_hd__xnor2_2
X_1168_ VPWR VGND _1169_/A _1221_/A VGND VPWR sky130_fd_sc_hd__buf_6
X_1237_ _1237_/B _1237_/Y _1237_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1099_ VGND VPWR _1098_/X _1095_/X _1467_/A _1087_/X _1083_/Y VGND VPWR sky130_fd_sc_hd__a211o_4
X_1022_ _1050_/B _1076_/A _1084_/A _0959_/C _1004_/A _1022_/X VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__o41a_2
X_1786_ VGND VPWR _1786_/X _1786_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_0806_ _1524_/S _0887_/B _1548_/S VGND VPWR VGND VPWR sky130_fd_sc_hd__or2b_4
XFILLER_52_163 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_4 _0920_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_3_281 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1571_ _1570_/X _1714_/D _1571_/X _1604_/A _1563_/X _1620_/A VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__o221a_2
X_1640_ VPWR VGND _1770_/Q _1640_/X _1640_/B VGND VPWR sky130_fd_sc_hd__and2_2
X_1005_ _1073_/C _1005_/B _1005_/X _1005_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__or3_2
X_1769_ _1769_/Q fanout175/X _1769_/D _1769_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_25_196 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xoutput41 VPWR VGND nmatrix_col_out_n[4] _1260_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput52 VPWR VGND nmatrix_row_out_n[15] _1791_/A VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput30 VPWR VGND nmatrix_col_out_n[23] _1293_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput63 VPWR VGND nmatrix_rowon_out_n[10] _1787_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput74 VPWR VGND nmatrix_rowon_out_n[7] _1784_/X VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_48_277 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xoutput96 VPWR VGND pmatrix_col_out_n[24] _1234_/Y VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput85 VPWR VGND pmatrix_col_out_n[14] _1201_/X VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_31_100 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1554_ VPWR VGND _1569_/B _1615_/C VGND VPWR sky130_fd_sc_hd__buf_4
X_1623_ VPWR VGND _1767_/Q _1623_/X _1640_/B VGND VPWR sky130_fd_sc_hd__and2_2
X_1485_ _1784_/A _1495_/A _1487_/B _1796_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_4
.ends

