magic
tech sky130A
timestamp 1664100429
<< nwell >>
rect 117 474 521 661
<< nmos >>
rect 254 390 304 440
rect 333 390 383 440
<< pmos >>
rect 189 493 289 593
rect 348 493 448 593
<< ndiff >>
rect 225 434 254 440
rect 225 396 231 434
rect 248 396 254 434
rect 225 390 254 396
rect 304 434 333 440
rect 304 396 310 434
rect 327 396 333 434
rect 304 390 333 396
rect 383 434 412 440
rect 383 396 389 434
rect 406 396 412 434
rect 383 390 412 396
<< pdiff >>
rect 160 587 189 593
rect 160 499 166 587
rect 183 499 189 587
rect 160 493 189 499
rect 289 587 348 593
rect 289 499 296 587
rect 342 499 348 587
rect 289 493 348 499
rect 448 587 477 593
rect 448 499 454 587
rect 471 499 477 587
rect 448 493 477 499
<< ndiffc >>
rect 231 396 248 434
rect 310 396 327 434
rect 389 396 406 434
<< pdiffc >>
rect 166 499 183 587
rect 296 499 342 587
rect 454 499 471 587
<< psubdiff >>
rect 161 295 173 312
rect 190 295 203 312
rect 403 295 415 312
rect 432 295 451 312
rect 468 295 480 312
<< nsubdiff >>
rect 162 640 255 643
rect 162 623 174 640
rect 191 623 226 640
rect 243 623 255 640
rect 162 620 255 623
rect 389 640 480 643
rect 389 623 401 640
rect 418 623 448 640
rect 465 623 480 640
rect 389 620 480 623
<< psubdiffcont >>
rect 173 295 190 312
rect 415 295 432 312
rect 451 295 468 312
<< nsubdiffcont >>
rect 174 623 191 640
rect 226 623 243 640
rect 401 623 418 640
rect 448 623 465 640
<< poly >>
rect 189 593 289 606
rect 348 593 448 606
rect 189 480 289 493
rect 348 480 448 493
rect 189 422 207 480
rect 254 440 304 453
rect 333 440 383 453
rect 172 414 207 422
rect 172 395 180 414
rect 199 395 207 414
rect 172 378 207 395
rect 430 422 448 480
rect 430 414 465 422
rect 430 395 438 414
rect 457 395 465 414
rect 172 359 180 378
rect 199 359 207 378
rect 254 377 304 390
rect 333 377 383 390
rect 254 362 383 377
rect 430 378 465 395
rect 172 351 207 359
rect 189 340 207 351
rect 189 325 270 340
rect 235 315 270 325
rect 235 296 243 315
rect 262 296 270 315
rect 235 288 270 296
rect 345 315 380 362
rect 430 359 438 378
rect 457 359 465 378
rect 430 351 465 359
rect 345 296 353 315
rect 372 296 380 315
rect 345 288 380 296
<< polycont >>
rect 180 395 199 414
rect 438 395 457 414
rect 180 359 199 378
rect 243 296 262 315
rect 438 359 457 378
rect 353 296 372 315
<< locali >>
rect 127 354 144 664
rect 162 640 255 643
rect 162 623 174 640
rect 191 623 226 640
rect 243 623 255 640
rect 162 620 255 623
rect 389 640 480 643
rect 389 623 401 640
rect 418 623 448 640
rect 465 623 480 640
rect 389 620 480 623
rect 166 587 183 595
rect 166 473 183 499
rect 296 587 342 596
rect 296 491 342 499
rect 454 587 471 595
rect 166 456 248 473
rect 231 434 248 456
rect 180 414 199 422
rect 180 382 199 395
rect 180 351 199 359
rect 231 358 248 396
rect 310 434 327 491
rect 454 473 471 499
rect 310 388 327 396
rect 389 456 471 473
rect 389 434 406 456
rect 389 358 406 396
rect 231 340 406 358
rect 438 414 457 422
rect 438 384 457 395
rect 438 351 457 359
rect 127 285 144 337
rect 243 315 262 323
rect 161 295 173 312
rect 190 295 203 312
rect 243 288 262 296
rect 244 285 261 288
rect 280 285 297 340
rect 353 315 372 323
rect 353 288 372 296
rect 403 295 415 312
rect 432 295 451 312
rect 468 295 480 312
rect 354 285 371 288
rect 497 285 514 664
<< viali >>
rect 174 623 191 640
rect 226 623 243 640
rect 401 623 418 640
rect 448 623 465 640
rect 307 531 335 565
rect 127 337 144 354
rect 180 378 199 382
rect 180 364 199 378
rect 438 378 457 384
rect 438 364 457 378
rect 173 295 190 312
rect 415 295 432 312
rect 451 295 468 312
<< metal1 >>
rect 117 640 521 648
rect 117 623 174 640
rect 191 623 226 640
rect 243 623 401 640
rect 418 623 448 640
rect 465 623 521 640
rect 117 620 521 623
rect 117 591 521 606
rect 304 565 338 571
rect 304 531 307 565
rect 335 531 338 565
rect 304 512 338 531
rect 117 477 521 491
rect 117 436 521 450
rect 117 408 521 422
rect 174 382 206 387
rect 174 364 180 382
rect 199 378 206 382
rect 432 384 463 387
rect 432 378 438 384
rect 199 364 438 378
rect 457 364 463 384
rect 124 354 147 360
rect 174 359 463 364
rect 124 345 127 354
rect 117 337 127 345
rect 144 345 147 354
rect 144 337 521 345
rect 117 331 521 337
rect 117 312 521 317
rect 117 295 173 312
rect 190 295 415 312
rect 432 295 451 312
rect 468 295 521 312
rect 117 289 521 295
<< via1 >>
rect 308 531 334 565
<< metal2 >>
rect 307 565 335 571
rect 307 526 335 531
<< via2 >>
rect 307 531 308 565
rect 308 531 334 565
rect 334 531 335 565
<< metal3 >>
rect 304 565 338 587
rect 304 531 305 565
rect 337 531 338 565
rect 304 512 338 531
<< via3 >>
rect 305 531 307 565
rect 307 531 335 565
rect 335 531 337 565
<< metal4 >>
rect 305 570 337 587
rect 304 565 338 570
rect 304 531 305 565
rect 337 531 338 565
rect 304 527 338 531
rect 305 512 337 527
<< labels >>
rlabel metal1 117 436 117 450 7 col_n
port 6 w
rlabel metal1 117 477 117 491 7 colon_n
port 7 w
rlabel metal1 117 331 117 345 7 vcom
port 3 w
rlabel metal1 117 591 117 606 7 sample_n
port 5 w
rlabel metal1 117 408 117 422 7 sample
port 4 w
rlabel metal1 117 289 117 317 7 VSS
port 2 w
rlabel metal1 117 620 117 648 7 VDD
port 1 w
rlabel locali 497 285 514 285 5 row_n
port 8 s
rlabel locali 244 285 261 285 5 sw_n
port 9 s
rlabel locali 354 285 371 285 5 sw
port 11 s
rlabel metal4 305 587 337 587 1 out
port 12 n
rlabel locali 280 285 297 285 5 in
port 10 s
<< end >>
