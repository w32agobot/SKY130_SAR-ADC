magic
tech sky130A
magscale 1 2
timestamp 1662452629
<< nwell >>
rect -38 244 1690 582
<< pwell >>
rect -38 -18 1690 244
<< nmos >>
rect 56 80 856 164
rect 1050 80 1080 164
rect 1146 80 1176 164
rect 1350 80 1380 164
rect 1446 80 1476 164
<< pmos >>
rect 1028 308 1058 468
rect 1124 308 1154 468
rect 1444 308 1474 468
rect 1540 308 1570 468
<< pmoslvt >>
rect 56 304 856 472
<< ndiff >>
rect -2 152 56 164
rect -2 92 10 152
rect 44 92 56 152
rect -2 80 56 92
rect 856 152 914 164
rect 856 92 868 152
rect 902 92 914 152
rect 856 80 914 92
rect 990 152 1050 164
rect 990 92 1000 152
rect 1034 92 1050 152
rect 990 80 1050 92
rect 1080 152 1146 164
rect 1080 92 1096 152
rect 1130 92 1146 152
rect 1080 80 1146 92
rect 1176 152 1234 164
rect 1176 92 1192 152
rect 1226 92 1234 152
rect 1176 80 1234 92
rect 1288 152 1350 164
rect 1288 92 1300 152
rect 1334 92 1350 152
rect 1288 80 1350 92
rect 1380 152 1446 164
rect 1380 92 1396 152
rect 1430 92 1446 152
rect 1380 80 1446 92
rect 1476 152 1538 164
rect 1476 92 1492 152
rect 1526 92 1538 152
rect 1476 80 1538 92
<< pdiff >>
rect -2 460 56 472
rect -2 316 10 460
rect 44 316 56 460
rect -2 304 56 316
rect 856 460 914 472
rect 856 316 868 460
rect 902 316 914 460
rect 856 304 914 316
rect 968 456 1028 468
rect 968 320 978 456
rect 1012 320 1028 456
rect 968 308 1028 320
rect 1058 456 1124 468
rect 1058 320 1074 456
rect 1108 320 1124 456
rect 1058 308 1124 320
rect 1154 456 1214 468
rect 1154 320 1170 456
rect 1204 320 1214 456
rect 1154 308 1214 320
rect 1382 456 1444 468
rect 1382 320 1394 456
rect 1428 320 1444 456
rect 1382 308 1444 320
rect 1474 456 1540 468
rect 1474 320 1490 456
rect 1524 320 1540 456
rect 1474 308 1540 320
rect 1570 456 1632 468
rect 1570 320 1586 456
rect 1620 320 1632 456
rect 1570 308 1632 320
<< ndiffc >>
rect 10 92 44 152
rect 868 92 902 152
rect 1000 92 1034 152
rect 1096 92 1130 152
rect 1192 92 1226 152
rect 1300 92 1334 152
rect 1396 92 1430 152
rect 1492 92 1526 152
<< pdiffc >>
rect 10 316 44 460
rect 868 316 902 460
rect 978 320 1012 456
rect 1074 320 1108 456
rect 1170 320 1204 456
rect 1394 320 1428 456
rect 1490 320 1524 456
rect 1586 320 1620 456
<< psubdiff >>
rect 94 -18 1594 26
<< poly >>
rect 56 472 856 498
rect 1028 468 1058 494
rect 1124 468 1154 494
rect 1444 468 1474 494
rect 1540 468 1570 494
rect 56 278 856 304
rect 1028 282 1058 308
rect 1124 282 1154 308
rect 56 266 182 278
rect -32 256 182 266
rect -32 210 -16 256
rect 32 210 182 256
rect -32 200 182 210
rect 898 248 986 258
rect 1028 252 1176 282
rect 1028 248 1080 252
rect 898 246 1080 248
rect 898 212 936 246
rect 970 212 1080 246
rect 898 206 1080 212
rect 898 202 986 206
rect 56 190 182 200
rect 56 164 856 190
rect 1050 164 1080 206
rect 1146 164 1176 252
rect 1236 252 1302 262
rect 1236 218 1252 252
rect 1286 220 1302 252
rect 1444 220 1474 308
rect 1540 220 1570 308
rect 1286 218 1570 220
rect 1236 190 1570 218
rect 1350 164 1380 190
rect 1446 164 1476 190
rect 56 54 856 80
rect 1050 54 1080 80
rect 1146 54 1176 80
rect 1350 54 1380 80
rect 1446 54 1476 80
<< polycont >>
rect -16 210 32 256
rect 936 212 970 246
rect 1252 218 1286 252
<< locali >>
rect 0 561 1652 562
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 1652 561
rect 0 526 1652 527
rect 10 460 44 476
rect 10 300 44 316
rect 868 460 902 476
rect -32 256 48 260
rect -32 210 -16 256
rect 32 210 48 256
rect -32 206 48 210
rect 868 258 902 316
rect 978 456 1012 526
rect 978 304 1012 320
rect 1074 456 1108 472
rect 1074 304 1108 320
rect 1170 456 1204 472
rect 1170 304 1204 320
rect 1320 270 1354 526
rect 1388 456 1428 472
rect 1388 320 1394 456
rect 1388 304 1428 320
rect 1490 456 1524 472
rect 868 246 986 258
rect 868 212 914 246
rect 970 212 986 246
rect 868 202 986 212
rect 1252 252 1286 268
rect 1320 236 1430 270
rect 1252 202 1286 218
rect 10 152 44 168
rect 10 76 44 92
rect 868 152 902 202
rect 868 76 902 92
rect 1000 152 1034 168
rect 1000 18 1034 92
rect 1096 152 1130 168
rect 1096 76 1130 92
rect 1192 76 1226 92
rect 1300 152 1334 168
rect 1300 76 1334 92
rect 1396 152 1430 236
rect 1490 236 1524 320
rect 1586 456 1626 472
rect 1620 320 1626 456
rect 1586 304 1626 320
rect 1490 202 1594 236
rect 1396 76 1430 92
rect 1492 152 1526 168
rect 1492 76 1526 92
rect 1560 18 1594 202
rect 0 -18 28 18
rect 64 17 1652 18
rect 64 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 1365 17
rect 1399 -17 1457 17
rect 1491 -17 1549 17
rect 1583 -17 1652 17
rect 64 -18 1652 -17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 10 316 44 460
rect 868 316 902 446
rect 1074 320 1108 456
rect 1170 320 1204 376
rect 1394 340 1428 456
rect 914 212 936 246
rect 936 212 970 246
rect 1252 218 1286 252
rect 10 92 44 152
rect 1096 92 1130 152
rect 1192 152 1226 178
rect 1192 144 1226 152
rect 1300 92 1334 132
rect 1586 340 1620 456
rect 1492 92 1526 132
rect 28 -18 64 18
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 1365 -17 1399 17
rect 1457 -17 1491 17
rect 1549 -17 1583 17
<< metal1 >>
rect 0 561 1652 594
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 1652 561
rect 0 496 1652 527
rect 4 460 50 496
rect 4 316 10 460
rect 44 316 50 460
rect 4 304 50 316
rect 862 446 908 468
rect 862 316 868 446
rect 902 316 908 446
rect 862 258 908 316
rect 1068 456 1626 468
rect 1068 320 1074 456
rect 1108 434 1394 456
rect 1108 320 1114 434
rect 1068 308 1114 320
rect 1164 376 1210 406
rect 1164 320 1170 376
rect 1204 320 1210 376
rect 1388 340 1394 434
rect 1428 434 1586 456
rect 1428 340 1434 434
rect 1388 328 1434 340
rect 1580 340 1586 434
rect 1620 340 1626 456
rect 1580 328 1626 340
rect 862 256 986 258
rect 862 204 914 256
rect 970 204 986 256
rect 1164 248 1210 320
rect 1246 252 1292 264
rect 1246 248 1252 252
rect 1164 220 1252 248
rect 862 202 986 204
rect 1186 218 1252 220
rect 1286 248 1292 252
rect 1286 220 1652 248
rect 1286 218 1292 220
rect 1186 206 1292 218
rect 1186 178 1232 206
rect 4 152 50 164
rect 4 92 10 152
rect 44 92 50 152
rect 1090 152 1136 164
rect 4 48 50 92
rect 864 110 968 118
rect 864 58 884 110
rect 948 58 968 110
rect 1090 92 1096 152
rect 1130 104 1136 152
rect 1186 144 1192 178
rect 1226 144 1232 178
rect 1186 132 1232 144
rect 1294 132 1340 144
rect 1294 104 1300 132
rect 1130 92 1300 104
rect 1334 104 1340 132
rect 1486 132 1532 144
rect 1486 104 1492 132
rect 1334 92 1492 104
rect 1526 92 1532 132
rect 1090 76 1532 92
rect 864 48 968 58
rect 0 18 1652 48
rect 0 -18 28 18
rect 64 17 1652 18
rect 64 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 1365 17
rect 1399 -17 1457 17
rect 1491 -17 1549 17
rect 1583 -17 1652 17
rect 64 -18 1652 -17
rect 0 -48 1652 -18
<< via1 >>
rect 914 246 970 256
rect 914 212 970 246
rect 914 204 970 212
rect 884 58 948 110
<< metal2 >>
rect 910 260 984 290
rect 910 258 920 260
rect 898 256 920 258
rect 898 204 914 256
rect 898 202 920 204
rect 976 202 984 260
rect 910 168 984 202
rect 864 116 968 118
rect 864 58 884 116
rect 948 58 968 116
rect 864 48 968 58
<< via2 >>
rect 920 256 976 260
rect 920 204 970 256
rect 970 204 976 256
rect 920 202 976 204
rect 884 110 948 116
rect 884 60 948 110
<< metal3 >>
rect 54 122 850 496
rect 910 264 986 318
rect 910 200 916 264
rect 980 200 986 264
rect 910 182 986 200
rect 1046 122 1652 496
rect 54 116 1652 122
rect 54 60 884 116
rect 948 60 1652 116
rect 54 54 1652 60
<< via3 >>
rect 916 260 980 264
rect 916 202 920 260
rect 920 202 976 260
rect 976 202 980 260
rect 916 200 980 202
<< mimcap >>
rect 86 264 822 468
rect 86 200 736 264
rect 800 200 822 264
rect 86 82 822 200
rect 1074 264 1600 468
rect 1074 200 1124 264
rect 1188 200 1600 264
rect 1074 82 1600 200
<< mimcapcontact >>
rect 736 200 800 264
rect 1124 200 1188 264
<< metal4 >>
rect 910 268 992 290
rect 732 264 1198 268
rect 732 200 736 264
rect 800 200 916 264
rect 980 200 1124 264
rect 1188 200 1198 264
rect 732 194 1198 200
rect 910 168 992 194
<< labels >>
rlabel locali -16 210 32 256 7 in
port 2 w
rlabel metal1 1622 220 1652 248 3 out
port 3 e
rlabel metal1 0 496 1652 594 7 VPWR
port 1 w
rlabel nwell 28 526 64 562 7 VPB
port 6 w
rlabel metal1 0 -48 1652 48 7 VGND
port 7 w
rlabel psubdiff 120 -18 156 18 7 VNB
port 8 w
rlabel locali 868 172 902 172 1 cap_top
<< end >>
