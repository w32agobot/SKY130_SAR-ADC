VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO adc_comp_latch
  CLASS BLOCK ;
  FOREIGN adc_comp_latch ;
  ORIGIN 0.000 0.000 ;
  SIZE 42.000 BY 129.000 ;
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 27.590 68.020 35.500 68.040 ;
        RECT 15.800 66.000 35.500 68.020 ;
        RECT 15.800 65.910 27.260 66.000 ;
        RECT 18.430 65.900 19.640 65.910 ;
        RECT 21.470 64.160 27.260 65.910 ;
        RECT 30.450 65.760 35.500 66.000 ;
        RECT 13.440 62.070 15.650 64.060 ;
        RECT 31.250 62.300 33.820 62.560 ;
        RECT 27.770 60.280 33.820 62.300 ;
      LAYER li1 ;
        RECT 27.600 67.650 30.340 68.140 ;
        RECT 30.890 67.690 35.120 67.860 ;
        RECT 14.910 67.190 20.270 67.430 ;
        RECT 22.490 67.240 26.110 67.480 ;
        RECT 14.910 64.060 15.340 67.190 ;
        RECT 16.050 67.100 20.060 67.190 ;
        RECT 16.050 66.390 16.220 67.100 ;
        RECT 17.010 66.390 17.180 67.100 ;
        RECT 17.970 66.390 18.140 67.100 ;
        RECT 18.930 66.390 19.100 67.100 ;
        RECT 19.890 66.390 20.060 67.100 ;
        RECT 24.170 67.070 24.620 67.240 ;
        RECT 23.320 66.900 25.410 67.070 ;
        RECT 23.320 64.640 23.490 66.900 ;
        RECT 24.280 64.640 24.450 66.900 ;
        RECT 25.240 64.640 25.410 66.900 ;
        RECT 28.490 66.290 28.660 67.650 ;
        RECT 29.450 66.290 29.620 67.650 ;
        RECT 13.310 63.860 15.340 64.060 ;
        RECT 13.310 62.940 13.490 63.860 ;
        RECT 13.750 63.700 14.170 63.860 ;
        RECT 14.440 62.940 14.660 63.860 ;
        RECT 14.920 63.700 15.340 63.860 ;
        RECT 13.310 62.750 14.190 62.940 ;
        RECT 14.440 62.750 15.360 62.940 ;
        RECT 28.490 60.650 28.660 62.010 ;
        RECT 29.450 60.650 29.620 62.010 ;
        RECT 30.060 60.650 30.340 67.650 ;
        RECT 31.650 66.250 31.820 67.690 ;
        RECT 34.130 66.250 34.300 67.690 ;
        RECT 27.610 60.630 30.340 60.650 ;
        RECT 32.450 60.630 32.620 62.070 ;
        RECT 27.610 60.460 33.440 60.630 ;
      LAYER mcon ;
        RECT 28.070 67.860 28.250 68.040 ;
        RECT 28.450 67.860 28.630 68.040 ;
        RECT 28.830 67.860 29.010 68.040 ;
        RECT 29.210 67.860 29.390 68.040 ;
        RECT 29.590 67.860 29.770 68.040 ;
        RECT 29.970 67.860 30.150 68.040 ;
        RECT 14.970 67.220 15.140 67.400 ;
        RECT 15.360 67.220 15.530 67.400 ;
        RECT 15.720 67.220 15.890 67.400 ;
        RECT 16.140 67.220 16.310 67.390 ;
        RECT 16.560 67.220 16.730 67.390 ;
        RECT 16.980 67.220 17.150 67.390 ;
        RECT 17.400 67.220 17.570 67.390 ;
        RECT 17.820 67.220 17.990 67.390 ;
        RECT 18.240 67.220 18.410 67.390 ;
        RECT 18.660 67.220 18.830 67.390 ;
        RECT 19.080 67.220 19.250 67.390 ;
        RECT 19.500 67.220 19.670 67.390 ;
        RECT 19.950 67.220 20.120 67.390 ;
        RECT 22.680 67.270 22.850 67.440 ;
        RECT 23.100 67.270 23.270 67.440 ;
        RECT 23.520 67.270 23.690 67.440 ;
        RECT 23.940 67.270 24.110 67.440 ;
        RECT 24.360 67.270 24.530 67.440 ;
        RECT 24.780 67.270 24.950 67.440 ;
        RECT 25.200 67.270 25.370 67.440 ;
        RECT 25.620 67.270 25.790 67.440 ;
        RECT 13.870 63.890 14.050 64.060 ;
        RECT 15.040 63.890 15.220 64.060 ;
      LAYER met1 ;
        RECT 8.010 67.700 40.330 68.850 ;
        RECT 14.910 67.190 20.270 67.700 ;
        RECT 22.490 67.240 26.110 67.700 ;
        RECT 13.710 63.860 14.200 64.090 ;
        RECT 14.880 63.860 15.370 64.090 ;
      LAYER via ;
        RECT 8.330 67.790 9.730 68.740 ;
        RECT 38.830 67.790 40.230 68.740 ;
      LAYER met2 ;
        RECT 8.240 67.700 9.840 68.850 ;
        RECT 38.730 67.700 40.330 68.850 ;
      LAYER via2 ;
        RECT 8.330 67.790 9.730 68.740 ;
        RECT 38.830 67.790 40.230 68.740 ;
      LAYER met3 ;
        RECT 8.240 67.700 9.840 68.850 ;
        RECT 38.730 67.700 40.330 68.850 ;
      LAYER via3 ;
        RECT 8.330 67.790 9.730 68.740 ;
        RECT 38.830 67.790 40.230 68.740 ;
      LAYER met4 ;
        RECT 8.240 50.000 9.840 77.980 ;
        RECT 38.730 50.000 40.330 77.980 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 16.530 75.990 18.930 76.890 ;
        RECT 29.430 75.990 31.830 76.890 ;
        RECT 14.230 75.590 20.480 75.990 ;
        RECT 23.730 75.590 24.630 75.990 ;
        RECT 27.880 75.590 34.130 75.990 ;
        RECT 14.230 70.290 34.130 75.590 ;
        RECT 14.230 69.890 20.480 70.290 ;
        RECT 23.730 69.890 24.630 70.290 ;
        RECT 27.880 69.890 34.130 70.290 ;
        RECT 16.530 68.990 18.930 69.890 ;
        RECT 29.430 68.990 31.830 69.890 ;
        RECT 16.530 58.040 18.930 58.940 ;
        RECT 29.430 58.040 31.830 58.940 ;
        RECT 14.230 57.640 20.480 58.040 ;
        RECT 23.730 57.640 24.630 58.040 ;
        RECT 27.880 57.640 34.130 58.040 ;
        RECT 14.230 52.340 34.130 57.640 ;
        RECT 14.230 51.940 20.480 52.340 ;
        RECT 23.730 51.940 24.630 52.340 ;
        RECT 27.880 51.940 34.130 52.340 ;
        RECT 16.530 51.040 18.930 51.940 ;
        RECT 29.430 51.040 31.830 51.940 ;
      LAYER li1 ;
        RECT 12.150 76.990 36.540 77.980 ;
        RECT 12.150 74.540 13.330 76.990 ;
        RECT 16.580 76.490 18.880 76.990 ;
        RECT 29.480 76.490 31.780 76.990 ;
        RECT 13.730 76.090 34.630 76.490 ;
        RECT 12.150 50.990 13.140 74.540 ;
        RECT 13.730 69.790 14.130 76.090 ;
        RECT 16.580 76.040 18.880 76.090 ;
        RECT 29.480 76.040 31.780 76.090 ;
        RECT 14.930 74.890 33.430 75.490 ;
        RECT 17.530 74.290 17.880 74.890 ;
        RECT 15.280 74.090 17.880 74.290 ;
        RECT 17.530 73.490 17.880 74.090 ;
        RECT 15.280 73.290 17.880 73.490 ;
        RECT 18.480 73.390 18.680 74.890 ;
        RECT 19.280 73.390 19.480 74.890 ;
        RECT 20.080 73.390 20.280 74.890 ;
        RECT 20.880 73.390 21.080 74.890 ;
        RECT 21.680 73.390 21.880 74.890 ;
        RECT 22.480 73.390 22.680 74.890 ;
        RECT 23.280 73.390 23.480 74.890 ;
        RECT 24.080 73.390 24.280 74.890 ;
        RECT 24.880 73.390 25.080 74.890 ;
        RECT 25.680 73.390 25.880 74.890 ;
        RECT 26.480 73.390 26.680 74.890 ;
        RECT 27.280 73.390 27.480 74.890 ;
        RECT 28.080 73.390 28.280 74.890 ;
        RECT 28.880 73.390 29.080 74.890 ;
        RECT 29.680 73.390 29.880 74.890 ;
        RECT 30.480 74.290 30.830 74.890 ;
        RECT 30.480 74.090 33.080 74.290 ;
        RECT 30.480 73.490 30.830 74.090 ;
        RECT 30.480 73.290 33.030 73.490 ;
        RECT 15.280 72.390 17.880 72.590 ;
        RECT 17.530 71.790 17.880 72.390 ;
        RECT 15.280 71.590 17.880 71.790 ;
        RECT 17.530 70.990 17.880 71.590 ;
        RECT 18.480 70.990 18.680 72.490 ;
        RECT 19.280 70.990 19.480 72.490 ;
        RECT 20.080 70.990 20.280 72.490 ;
        RECT 20.880 70.990 21.080 72.490 ;
        RECT 21.680 70.990 21.880 72.490 ;
        RECT 22.480 70.990 22.680 72.490 ;
        RECT 23.280 70.990 23.480 72.490 ;
        RECT 24.080 70.990 24.280 72.490 ;
        RECT 24.880 70.990 25.080 72.490 ;
        RECT 25.680 70.990 25.880 72.490 ;
        RECT 26.480 70.990 26.680 72.490 ;
        RECT 27.280 70.990 27.480 72.490 ;
        RECT 28.080 70.990 28.280 72.490 ;
        RECT 28.880 70.990 29.080 72.490 ;
        RECT 29.680 70.990 29.880 72.490 ;
        RECT 30.480 72.390 33.030 72.590 ;
        RECT 30.480 71.790 30.830 72.390 ;
        RECT 30.480 71.590 33.080 71.790 ;
        RECT 30.480 70.990 30.830 71.590 ;
        RECT 14.930 70.390 33.430 70.990 ;
        RECT 16.580 69.790 18.880 69.840 ;
        RECT 29.480 69.790 31.780 69.840 ;
        RECT 34.230 69.790 34.630 76.090 ;
        RECT 13.730 69.390 34.630 69.790 ;
        RECT 16.580 68.990 18.880 69.390 ;
        RECT 29.480 68.990 31.780 69.390 ;
        RECT 28.490 64.410 28.660 65.200 ;
        RECT 29.450 64.410 29.620 65.200 ;
        RECT 31.170 64.740 31.340 65.440 ;
        RECT 33.650 64.740 33.820 65.440 ;
        RECT 35.550 64.740 36.540 76.990 ;
        RECT 31.040 64.480 36.540 64.740 ;
        RECT 27.950 64.320 29.730 64.410 ;
        RECT 27.270 63.980 29.730 64.320 ;
        RECT 13.730 61.060 14.190 61.230 ;
        RECT 14.900 61.060 15.360 61.230 ;
        RECT 13.750 60.530 14.170 61.060 ;
        RECT 14.920 60.530 15.340 61.060 ;
        RECT 16.530 60.310 16.700 61.570 ;
        RECT 17.490 60.310 17.660 61.560 ;
        RECT 18.450 60.310 18.620 61.560 ;
        RECT 19.410 60.310 19.580 61.560 ;
        RECT 23.320 60.450 23.490 63.030 ;
        RECT 24.280 60.450 24.450 63.030 ;
        RECT 25.240 60.450 25.410 63.030 ;
        RECT 27.270 62.350 27.610 63.980 ;
        RECT 27.950 63.890 29.730 63.980 ;
        RECT 28.490 63.100 28.660 63.890 ;
        RECT 29.450 63.100 29.620 63.890 ;
        RECT 31.850 63.590 32.280 64.480 ;
        RECT 31.970 62.880 32.140 63.590 ;
        RECT 26.920 62.010 27.610 62.350 ;
        RECT 16.530 60.240 19.580 60.310 ;
        RECT 23.290 60.260 25.550 60.450 ;
        RECT 26.920 60.260 27.320 62.010 ;
        RECT 15.960 60.030 20.050 60.240 ;
        RECT 16.580 58.540 18.880 60.030 ;
        RECT 26.920 59.910 31.780 60.260 ;
        RECT 29.480 58.540 31.780 59.910 ;
        RECT 13.730 58.140 34.630 58.540 ;
        RECT 13.730 51.840 14.130 58.140 ;
        RECT 16.580 58.090 18.880 58.140 ;
        RECT 29.480 58.090 31.780 58.140 ;
        RECT 14.930 56.940 33.430 57.540 ;
        RECT 17.530 56.340 17.880 56.940 ;
        RECT 15.280 56.140 17.880 56.340 ;
        RECT 17.530 55.540 17.880 56.140 ;
        RECT 15.280 55.340 17.880 55.540 ;
        RECT 18.480 55.440 18.680 56.940 ;
        RECT 19.280 55.440 19.480 56.940 ;
        RECT 20.080 55.440 20.280 56.940 ;
        RECT 20.880 55.440 21.080 56.940 ;
        RECT 21.680 55.440 21.880 56.940 ;
        RECT 22.480 55.440 22.680 56.940 ;
        RECT 23.280 55.440 23.480 56.940 ;
        RECT 24.080 55.440 24.280 56.940 ;
        RECT 24.880 55.440 25.080 56.940 ;
        RECT 25.680 55.440 25.880 56.940 ;
        RECT 26.480 55.440 26.680 56.940 ;
        RECT 27.280 55.440 27.480 56.940 ;
        RECT 28.080 55.440 28.280 56.940 ;
        RECT 28.880 55.440 29.080 56.940 ;
        RECT 29.680 55.440 29.880 56.940 ;
        RECT 30.480 56.340 30.830 56.940 ;
        RECT 30.480 56.140 33.080 56.340 ;
        RECT 30.480 55.540 30.830 56.140 ;
        RECT 30.480 55.340 33.030 55.540 ;
        RECT 15.280 54.440 17.880 54.640 ;
        RECT 17.530 53.840 17.880 54.440 ;
        RECT 15.280 53.640 17.880 53.840 ;
        RECT 17.530 53.040 17.880 53.640 ;
        RECT 18.480 53.040 18.680 54.540 ;
        RECT 19.280 53.040 19.480 54.540 ;
        RECT 20.080 53.040 20.280 54.540 ;
        RECT 20.880 53.040 21.080 54.540 ;
        RECT 21.680 53.040 21.880 54.540 ;
        RECT 22.480 53.040 22.680 54.540 ;
        RECT 23.280 53.040 23.480 54.540 ;
        RECT 24.080 53.040 24.280 54.540 ;
        RECT 24.880 53.040 25.080 54.540 ;
        RECT 25.680 53.040 25.880 54.540 ;
        RECT 26.480 53.040 26.680 54.540 ;
        RECT 27.280 53.040 27.480 54.540 ;
        RECT 28.080 53.040 28.280 54.540 ;
        RECT 28.880 53.040 29.080 54.540 ;
        RECT 29.680 53.040 29.880 54.540 ;
        RECT 30.480 54.440 33.030 54.640 ;
        RECT 30.480 53.840 30.830 54.440 ;
        RECT 30.480 53.640 33.080 53.840 ;
        RECT 30.480 53.040 30.830 53.640 ;
        RECT 14.930 52.440 33.430 53.040 ;
        RECT 16.580 51.840 18.880 51.890 ;
        RECT 29.480 51.840 31.780 51.890 ;
        RECT 34.230 51.840 34.630 58.140 ;
        RECT 13.730 51.440 34.630 51.840 ;
        RECT 16.580 50.990 18.880 51.440 ;
        RECT 29.480 50.990 31.780 51.440 ;
        RECT 35.550 50.990 36.540 64.480 ;
        RECT 12.150 50.000 36.540 50.990 ;
      LAYER mcon ;
        RECT 12.330 74.740 12.980 76.740 ;
        RECT 12.250 71.840 12.930 74.040 ;
        RECT 12.250 69.090 13.030 71.240 ;
        RECT 15.030 74.990 15.630 75.490 ;
        RECT 15.830 74.990 16.430 75.490 ;
        RECT 16.630 74.990 17.230 75.490 ;
        RECT 17.430 74.990 18.030 75.490 ;
        RECT 30.330 74.990 30.930 75.490 ;
        RECT 31.130 74.990 31.730 75.490 ;
        RECT 31.930 74.990 32.530 75.490 ;
        RECT 32.730 74.990 33.330 75.490 ;
        RECT 15.030 70.390 15.630 70.890 ;
        RECT 15.830 70.390 16.430 70.890 ;
        RECT 16.630 70.390 17.230 70.890 ;
        RECT 17.430 70.390 18.030 70.890 ;
        RECT 30.330 70.390 30.930 70.890 ;
        RECT 31.130 70.390 31.730 70.890 ;
        RECT 31.930 70.390 32.530 70.890 ;
        RECT 32.730 70.390 33.330 70.890 ;
        RECT 12.230 60.610 12.400 60.780 ;
        RECT 12.590 60.610 12.760 60.780 ;
        RECT 12.950 60.610 13.120 60.780 ;
        RECT 13.870 60.560 14.050 60.730 ;
        RECT 15.040 60.560 15.220 60.730 ;
        RECT 12.230 60.250 12.400 60.420 ;
        RECT 12.590 60.250 12.760 60.420 ;
        RECT 12.950 60.250 13.120 60.420 ;
        RECT 23.410 60.270 23.590 60.450 ;
        RECT 23.870 60.270 24.050 60.450 ;
        RECT 24.330 60.270 24.510 60.450 ;
        RECT 24.790 60.270 24.970 60.450 ;
        RECT 25.250 60.270 25.430 60.450 ;
        RECT 35.620 60.610 35.790 60.780 ;
        RECT 35.980 60.610 36.150 60.780 ;
        RECT 36.340 60.610 36.510 60.780 ;
        RECT 12.230 59.890 12.400 60.060 ;
        RECT 12.590 59.890 12.760 60.060 ;
        RECT 12.950 59.890 13.120 60.060 ;
        RECT 16.080 60.050 16.260 60.230 ;
        RECT 16.670 60.050 16.850 60.230 ;
        RECT 17.260 60.050 17.440 60.230 ;
        RECT 17.850 60.050 18.030 60.230 ;
        RECT 18.440 60.050 18.620 60.230 ;
        RECT 19.030 60.050 19.210 60.230 ;
        RECT 19.620 60.050 19.800 60.230 ;
        RECT 12.230 59.530 12.400 59.700 ;
        RECT 12.590 59.530 12.760 59.700 ;
        RECT 12.950 59.530 13.120 59.700 ;
        RECT 12.220 59.170 12.390 59.340 ;
        RECT 12.580 59.170 12.750 59.340 ;
        RECT 12.940 59.170 13.110 59.340 ;
        RECT 12.240 56.690 13.030 58.840 ;
        RECT 26.960 59.980 27.140 60.160 ;
        RECT 27.330 59.990 27.510 60.170 ;
        RECT 27.730 59.990 27.910 60.170 ;
        RECT 28.130 59.990 28.310 60.170 ;
        RECT 28.530 59.990 28.710 60.170 ;
        RECT 35.620 60.250 35.790 60.420 ;
        RECT 35.980 60.250 36.150 60.420 ;
        RECT 36.340 60.250 36.510 60.420 ;
        RECT 35.620 59.890 35.790 60.060 ;
        RECT 35.980 59.890 36.150 60.060 ;
        RECT 36.340 59.890 36.510 60.060 ;
        RECT 35.620 59.530 35.790 59.700 ;
        RECT 35.980 59.530 36.150 59.700 ;
        RECT 36.340 59.530 36.510 59.700 ;
        RECT 35.620 59.170 35.790 59.340 ;
        RECT 35.980 59.170 36.150 59.340 ;
        RECT 36.340 59.170 36.510 59.340 ;
        RECT 12.280 53.890 12.930 56.090 ;
        RECT 12.280 51.190 13.080 53.240 ;
        RECT 15.030 57.040 15.630 57.540 ;
        RECT 15.830 57.040 16.430 57.540 ;
        RECT 16.630 57.040 17.230 57.540 ;
        RECT 17.430 57.040 18.030 57.540 ;
        RECT 30.330 57.040 30.930 57.540 ;
        RECT 31.130 57.040 31.730 57.540 ;
        RECT 31.930 57.040 32.530 57.540 ;
        RECT 32.730 57.040 33.330 57.540 ;
        RECT 15.030 52.440 15.630 52.940 ;
        RECT 15.830 52.440 16.430 52.940 ;
        RECT 16.630 52.440 17.230 52.940 ;
        RECT 17.430 52.440 18.030 52.940 ;
        RECT 30.330 52.440 30.930 52.940 ;
        RECT 31.130 52.440 31.730 52.940 ;
        RECT 31.930 52.440 32.530 52.940 ;
        RECT 32.730 52.440 33.330 52.940 ;
      LAYER met1 ;
        RECT 12.150 75.690 16.530 76.890 ;
        RECT 31.830 75.690 35.030 76.890 ;
        RECT 12.150 75.540 15.630 75.690 ;
        RECT 32.730 75.540 35.030 75.690 ;
        RECT 12.150 75.390 23.730 75.540 ;
        RECT 24.630 75.390 35.030 75.540 ;
        RECT 12.150 74.940 18.130 75.390 ;
        RECT 30.230 74.940 35.030 75.390 ;
        RECT 12.150 74.540 14.530 74.940 ;
        RECT 14.980 74.890 23.730 74.940 ;
        RECT 12.150 71.740 13.030 74.140 ;
        RECT 13.330 74.040 14.530 74.540 ;
        RECT 15.130 73.540 15.280 74.890 ;
        RECT 15.730 73.540 15.880 74.890 ;
        RECT 16.330 73.540 16.480 74.890 ;
        RECT 16.930 73.540 17.080 74.890 ;
        RECT 17.530 74.790 23.730 74.890 ;
        RECT 24.630 74.890 33.380 74.940 ;
        RECT 24.630 74.790 30.830 74.890 ;
        RECT 17.530 74.340 18.130 74.790 ;
        RECT 30.230 74.340 30.830 74.790 ;
        RECT 17.530 74.190 23.730 74.340 ;
        RECT 24.630 74.190 30.830 74.340 ;
        RECT 17.530 73.740 18.130 74.190 ;
        RECT 30.230 73.740 30.830 74.190 ;
        RECT 17.530 73.590 23.730 73.740 ;
        RECT 24.630 73.590 30.830 73.740 ;
        RECT 17.530 73.390 18.130 73.590 ;
        RECT 30.230 73.390 30.830 73.590 ;
        RECT 31.280 73.540 31.430 74.890 ;
        RECT 31.880 73.540 32.030 74.890 ;
        RECT 32.480 73.540 32.630 74.890 ;
        RECT 33.080 73.540 33.230 74.890 ;
        RECT 33.830 74.040 35.030 74.940 ;
        RECT 13.330 71.340 14.530 71.840 ;
        RECT 12.150 70.940 14.530 71.340 ;
        RECT 15.130 70.990 15.280 72.290 ;
        RECT 15.730 70.990 15.880 72.290 ;
        RECT 16.330 70.990 16.480 72.290 ;
        RECT 16.930 70.990 17.080 72.290 ;
        RECT 17.530 72.140 23.730 72.290 ;
        RECT 24.630 72.140 30.830 72.290 ;
        RECT 17.530 71.690 18.130 72.140 ;
        RECT 30.230 71.690 30.830 72.140 ;
        RECT 17.530 71.540 23.730 71.690 ;
        RECT 24.630 71.540 30.830 71.690 ;
        RECT 17.530 71.090 18.130 71.540 ;
        RECT 30.230 71.090 30.830 71.540 ;
        RECT 17.530 70.990 23.730 71.090 ;
        RECT 14.980 70.940 23.730 70.990 ;
        RECT 24.630 70.990 30.830 71.090 ;
        RECT 31.280 70.990 31.430 72.290 ;
        RECT 31.880 70.990 32.030 72.290 ;
        RECT 32.480 70.990 32.630 72.290 ;
        RECT 33.080 70.990 33.230 72.290 ;
        RECT 24.630 70.940 33.380 70.990 ;
        RECT 33.830 70.940 35.030 71.840 ;
        RECT 12.150 70.490 18.130 70.940 ;
        RECT 30.230 70.490 35.030 70.940 ;
        RECT 12.150 70.340 23.730 70.490 ;
        RECT 24.630 70.340 35.030 70.490 ;
        RECT 12.150 70.190 15.630 70.340 ;
        RECT 32.730 70.190 35.030 70.340 ;
        RECT 12.150 68.990 16.530 70.190 ;
        RECT 31.830 68.990 35.030 70.190 ;
        RECT 12.150 60.780 13.150 60.880 ;
        RECT 12.150 60.260 15.420 60.780 ;
        RECT 23.290 60.260 25.550 60.480 ;
        RECT 35.550 60.260 36.540 60.880 ;
        RECT 8.010 59.100 38.380 60.260 ;
        RECT 12.140 57.740 16.530 58.940 ;
        RECT 31.830 57.740 35.030 58.940 ;
        RECT 12.140 57.590 15.630 57.740 ;
        RECT 32.730 57.590 35.030 57.740 ;
        RECT 12.140 57.440 23.730 57.590 ;
        RECT 24.630 57.440 35.030 57.590 ;
        RECT 12.140 56.990 18.130 57.440 ;
        RECT 30.230 56.990 35.030 57.440 ;
        RECT 12.140 56.590 14.530 56.990 ;
        RECT 14.980 56.940 23.730 56.990 ;
        RECT 12.150 53.790 13.030 56.190 ;
        RECT 13.330 56.090 14.530 56.590 ;
        RECT 15.130 55.590 15.280 56.940 ;
        RECT 15.730 55.590 15.880 56.940 ;
        RECT 16.330 55.590 16.480 56.940 ;
        RECT 16.930 55.590 17.080 56.940 ;
        RECT 17.530 56.840 23.730 56.940 ;
        RECT 24.630 56.940 33.380 56.990 ;
        RECT 24.630 56.840 30.830 56.940 ;
        RECT 17.530 56.390 18.130 56.840 ;
        RECT 30.230 56.390 30.830 56.840 ;
        RECT 17.530 56.240 23.730 56.390 ;
        RECT 24.630 56.240 30.830 56.390 ;
        RECT 17.530 55.790 18.130 56.240 ;
        RECT 30.230 55.790 30.830 56.240 ;
        RECT 17.530 55.640 23.730 55.790 ;
        RECT 24.630 55.640 30.830 55.790 ;
        RECT 17.530 55.440 18.130 55.640 ;
        RECT 30.230 55.440 30.830 55.640 ;
        RECT 31.280 55.590 31.430 56.940 ;
        RECT 31.880 55.590 32.030 56.940 ;
        RECT 32.480 55.590 32.630 56.940 ;
        RECT 33.080 55.590 33.230 56.940 ;
        RECT 33.830 56.090 35.030 56.990 ;
        RECT 13.330 53.390 14.530 53.890 ;
        RECT 12.150 52.990 14.530 53.390 ;
        RECT 15.130 53.040 15.280 54.340 ;
        RECT 15.730 53.040 15.880 54.340 ;
        RECT 16.330 53.040 16.480 54.340 ;
        RECT 16.930 53.040 17.080 54.340 ;
        RECT 17.530 54.190 23.730 54.340 ;
        RECT 24.630 54.190 30.830 54.340 ;
        RECT 17.530 53.740 18.130 54.190 ;
        RECT 30.230 53.740 30.830 54.190 ;
        RECT 17.530 53.590 23.730 53.740 ;
        RECT 24.630 53.590 30.830 53.740 ;
        RECT 17.530 53.140 18.130 53.590 ;
        RECT 30.230 53.140 30.830 53.590 ;
        RECT 17.530 53.040 23.730 53.140 ;
        RECT 14.980 52.990 23.730 53.040 ;
        RECT 24.630 53.040 30.830 53.140 ;
        RECT 31.280 53.040 31.430 54.340 ;
        RECT 31.880 53.040 32.030 54.340 ;
        RECT 32.480 53.040 32.630 54.340 ;
        RECT 33.080 53.040 33.230 54.340 ;
        RECT 24.630 52.990 33.380 53.040 ;
        RECT 33.830 52.990 35.030 53.890 ;
        RECT 12.150 52.540 18.130 52.990 ;
        RECT 30.230 52.540 35.030 52.990 ;
        RECT 12.150 52.390 23.730 52.540 ;
        RECT 24.630 52.390 35.030 52.540 ;
        RECT 12.150 52.240 15.630 52.390 ;
        RECT 32.730 52.240 35.030 52.390 ;
        RECT 12.150 51.040 16.530 52.240 ;
        RECT 31.830 51.040 35.030 52.240 ;
      LAYER via ;
        RECT 12.330 74.740 12.980 76.740 ;
        RECT 13.430 75.790 14.430 76.790 ;
        RECT 15.430 75.790 16.430 76.790 ;
        RECT 31.930 75.790 32.930 76.790 ;
        RECT 33.930 75.790 34.930 76.790 ;
        RECT 13.430 74.190 14.430 75.190 ;
        RECT 12.250 71.840 12.930 74.040 ;
        RECT 33.930 74.190 34.930 75.190 ;
        RECT 13.430 70.690 14.430 71.690 ;
        RECT 33.930 70.690 34.930 71.690 ;
        RECT 13.430 69.090 14.430 70.090 ;
        RECT 15.430 69.090 16.430 70.090 ;
        RECT 31.930 69.090 32.930 70.090 ;
        RECT 33.930 69.090 34.930 70.090 ;
        RECT 10.330 59.190 11.730 60.140 ;
        RECT 13.430 59.290 16.210 60.120 ;
        RECT 36.880 59.190 38.280 60.140 ;
        RECT 13.430 57.840 14.430 58.840 ;
        RECT 15.430 57.840 16.430 58.840 ;
        RECT 31.930 57.840 32.930 58.840 ;
        RECT 33.930 57.840 34.930 58.840 ;
        RECT 13.430 56.240 14.430 57.240 ;
        RECT 12.280 53.890 12.930 56.090 ;
        RECT 33.930 56.240 34.930 57.240 ;
        RECT 12.280 51.190 12.940 53.240 ;
        RECT 13.430 52.740 14.430 53.740 ;
        RECT 33.930 52.740 34.930 53.740 ;
        RECT 13.430 51.140 14.430 52.140 ;
        RECT 15.430 51.140 16.430 52.140 ;
        RECT 31.930 51.140 32.930 52.140 ;
        RECT 33.930 51.140 34.930 52.140 ;
      LAYER met2 ;
        RECT 12.150 75.690 16.530 76.890 ;
        RECT 31.830 75.690 35.030 76.890 ;
        RECT 12.150 74.740 15.280 75.690 ;
        RECT 33.080 74.740 35.030 75.690 ;
        RECT 12.150 74.590 17.280 74.740 ;
        RECT 12.150 74.540 15.280 74.590 ;
        RECT 13.330 74.140 15.280 74.540 ;
        RECT 12.150 71.740 13.030 74.140 ;
        RECT 13.330 74.040 17.280 74.140 ;
        RECT 14.730 73.990 17.280 74.040 ;
        RECT 14.730 73.390 15.280 73.990 ;
        RECT 14.730 73.090 17.280 73.390 ;
        RECT 17.880 73.090 18.030 74.740 ;
        RECT 18.480 73.090 18.630 74.740 ;
        RECT 19.080 73.090 19.230 74.740 ;
        RECT 19.680 73.090 19.830 74.740 ;
        RECT 20.280 73.090 20.430 74.740 ;
        RECT 20.880 73.090 21.030 74.740 ;
        RECT 21.480 73.090 21.630 74.740 ;
        RECT 22.080 73.090 22.230 74.740 ;
        RECT 22.680 73.090 22.830 74.740 ;
        RECT 23.280 73.090 23.430 74.740 ;
        RECT 23.880 73.090 24.480 74.740 ;
        RECT 24.930 73.090 25.080 74.740 ;
        RECT 25.530 73.090 25.680 74.740 ;
        RECT 26.130 73.090 26.280 74.740 ;
        RECT 26.730 73.090 26.880 74.740 ;
        RECT 27.330 73.090 27.480 74.740 ;
        RECT 27.930 73.090 28.080 74.740 ;
        RECT 28.530 73.090 28.680 74.740 ;
        RECT 29.130 73.090 29.280 74.740 ;
        RECT 29.730 73.090 29.880 74.740 ;
        RECT 30.330 73.090 30.480 74.740 ;
        RECT 31.080 74.590 35.030 74.740 ;
        RECT 33.080 74.140 35.030 74.590 ;
        RECT 31.080 74.040 35.030 74.140 ;
        RECT 31.080 73.990 33.630 74.040 ;
        RECT 33.080 73.390 33.630 73.990 ;
        RECT 31.080 73.090 33.630 73.390 ;
        RECT 14.730 72.790 33.630 73.090 ;
        RECT 14.730 72.340 17.280 72.790 ;
        RECT 14.730 71.890 15.280 72.340 ;
        RECT 14.730 71.840 17.280 71.890 ;
        RECT 13.330 71.740 17.280 71.840 ;
        RECT 13.330 71.290 15.280 71.740 ;
        RECT 13.330 71.140 17.280 71.290 ;
        RECT 17.880 71.140 18.030 72.790 ;
        RECT 18.480 71.140 18.630 72.790 ;
        RECT 19.080 71.140 19.230 72.790 ;
        RECT 19.680 71.140 19.830 72.790 ;
        RECT 20.280 71.140 20.430 72.790 ;
        RECT 20.880 71.140 21.030 72.790 ;
        RECT 21.480 71.140 21.630 72.790 ;
        RECT 22.080 71.140 22.230 72.790 ;
        RECT 22.680 71.140 22.830 72.790 ;
        RECT 23.280 71.140 23.430 72.790 ;
        RECT 23.880 71.140 24.480 72.790 ;
        RECT 24.930 71.140 25.080 72.790 ;
        RECT 25.530 71.140 25.680 72.790 ;
        RECT 26.130 71.140 26.280 72.790 ;
        RECT 26.730 71.140 26.880 72.790 ;
        RECT 27.330 71.140 27.480 72.790 ;
        RECT 27.930 71.140 28.080 72.790 ;
        RECT 28.530 71.140 28.680 72.790 ;
        RECT 29.130 71.140 29.280 72.790 ;
        RECT 29.730 71.140 29.880 72.790 ;
        RECT 30.330 71.140 30.480 72.790 ;
        RECT 31.080 72.340 33.630 72.790 ;
        RECT 33.080 71.890 33.630 72.340 ;
        RECT 31.080 71.840 33.630 71.890 ;
        RECT 31.080 71.740 35.030 71.840 ;
        RECT 33.080 71.290 35.030 71.740 ;
        RECT 31.080 71.140 35.030 71.290 ;
        RECT 13.330 70.190 15.280 71.140 ;
        RECT 33.080 70.190 35.030 71.140 ;
        RECT 13.330 68.990 16.530 70.190 ;
        RECT 31.830 68.990 35.030 70.190 ;
        RECT 10.220 59.100 11.820 60.260 ;
        RECT 13.290 59.260 16.440 60.260 ;
        RECT 13.330 58.940 16.480 59.260 ;
        RECT 36.780 59.100 38.380 60.260 ;
        RECT 13.330 57.740 16.530 58.940 ;
        RECT 31.830 57.740 35.030 58.940 ;
        RECT 13.330 56.790 15.280 57.740 ;
        RECT 33.080 56.790 35.030 57.740 ;
        RECT 13.330 56.640 17.280 56.790 ;
        RECT 13.330 56.190 15.280 56.640 ;
        RECT 12.150 53.790 13.030 56.190 ;
        RECT 13.330 56.090 17.280 56.190 ;
        RECT 14.730 56.040 17.280 56.090 ;
        RECT 14.730 55.440 15.280 56.040 ;
        RECT 14.730 55.140 17.280 55.440 ;
        RECT 17.880 55.140 18.030 56.790 ;
        RECT 18.480 55.140 18.630 56.790 ;
        RECT 19.080 55.140 19.230 56.790 ;
        RECT 19.680 55.140 19.830 56.790 ;
        RECT 20.280 55.140 20.430 56.790 ;
        RECT 20.880 55.140 21.030 56.790 ;
        RECT 21.480 55.140 21.630 56.790 ;
        RECT 22.080 55.140 22.230 56.790 ;
        RECT 22.680 55.140 22.830 56.790 ;
        RECT 23.280 55.140 23.430 56.790 ;
        RECT 23.880 55.140 24.480 56.790 ;
        RECT 24.930 55.140 25.080 56.790 ;
        RECT 25.530 55.140 25.680 56.790 ;
        RECT 26.130 55.140 26.280 56.790 ;
        RECT 26.730 55.140 26.880 56.790 ;
        RECT 27.330 55.140 27.480 56.790 ;
        RECT 27.930 55.140 28.080 56.790 ;
        RECT 28.530 55.140 28.680 56.790 ;
        RECT 29.130 55.140 29.280 56.790 ;
        RECT 29.730 55.140 29.880 56.790 ;
        RECT 30.330 55.140 30.480 56.790 ;
        RECT 31.080 56.640 35.030 56.790 ;
        RECT 33.080 56.190 35.030 56.640 ;
        RECT 31.080 56.090 35.030 56.190 ;
        RECT 31.080 56.040 33.630 56.090 ;
        RECT 33.080 55.440 33.630 56.040 ;
        RECT 31.080 55.140 33.630 55.440 ;
        RECT 14.730 54.840 33.630 55.140 ;
        RECT 14.730 54.390 17.280 54.840 ;
        RECT 14.730 53.940 15.280 54.390 ;
        RECT 14.730 53.890 17.280 53.940 ;
        RECT 13.330 53.790 17.280 53.890 ;
        RECT 13.330 53.390 15.280 53.790 ;
        RECT 12.150 53.340 15.280 53.390 ;
        RECT 12.150 53.190 17.280 53.340 ;
        RECT 17.880 53.190 18.030 54.840 ;
        RECT 18.480 53.190 18.630 54.840 ;
        RECT 19.080 53.190 19.230 54.840 ;
        RECT 19.680 53.190 19.830 54.840 ;
        RECT 20.280 53.190 20.430 54.840 ;
        RECT 20.880 53.190 21.030 54.840 ;
        RECT 21.480 53.190 21.630 54.840 ;
        RECT 22.080 53.190 22.230 54.840 ;
        RECT 22.680 53.190 22.830 54.840 ;
        RECT 23.280 53.190 23.430 54.840 ;
        RECT 23.880 53.190 24.480 54.840 ;
        RECT 24.930 53.190 25.080 54.840 ;
        RECT 25.530 53.190 25.680 54.840 ;
        RECT 26.130 53.190 26.280 54.840 ;
        RECT 26.730 53.190 26.880 54.840 ;
        RECT 27.330 53.190 27.480 54.840 ;
        RECT 27.930 53.190 28.080 54.840 ;
        RECT 28.530 53.190 28.680 54.840 ;
        RECT 29.130 53.190 29.280 54.840 ;
        RECT 29.730 53.190 29.880 54.840 ;
        RECT 30.330 53.190 30.480 54.840 ;
        RECT 31.080 54.390 33.630 54.840 ;
        RECT 33.080 53.940 33.630 54.390 ;
        RECT 31.080 53.890 33.630 53.940 ;
        RECT 31.080 53.790 35.030 53.890 ;
        RECT 33.080 53.340 35.030 53.790 ;
        RECT 31.080 53.190 35.030 53.340 ;
        RECT 12.150 52.240 15.280 53.190 ;
        RECT 33.080 52.240 35.030 53.190 ;
        RECT 12.150 51.040 16.530 52.240 ;
        RECT 31.830 51.040 35.030 52.240 ;
      LAYER via2 ;
        RECT 12.330 74.740 12.980 76.740 ;
        RECT 12.250 71.840 12.930 74.040 ;
        RECT 10.330 59.190 11.730 60.140 ;
        RECT 13.430 59.290 16.210 60.120 ;
        RECT 36.880 59.190 38.280 60.140 ;
        RECT 12.280 53.890 12.930 56.090 ;
        RECT 12.280 51.190 12.940 53.240 ;
      LAYER met3 ;
        RECT 12.150 74.540 13.020 76.890 ;
        RECT 13.330 75.640 16.530 76.890 ;
        RECT 18.930 76.040 29.430 76.890 ;
        RECT 31.830 75.640 35.030 76.890 ;
        RECT 13.330 74.490 35.030 75.640 ;
        RECT 12.150 71.740 13.030 74.140 ;
        RECT 13.330 71.740 14.180 74.140 ;
        RECT 14.580 71.390 33.780 74.490 ;
        RECT 34.180 71.740 35.030 74.140 ;
        RECT 13.330 70.240 35.030 71.390 ;
        RECT 13.330 68.990 16.530 70.240 ;
        RECT 18.930 68.990 29.430 69.840 ;
        RECT 31.830 68.990 35.030 70.240 ;
        RECT 10.220 59.100 11.820 60.260 ;
        RECT 13.290 59.260 16.440 60.260 ;
        RECT 36.780 59.100 38.380 60.260 ;
        RECT 13.330 57.690 16.530 58.940 ;
        RECT 18.930 58.090 29.430 58.940 ;
        RECT 31.830 57.690 35.030 58.940 ;
        RECT 13.330 56.540 35.030 57.690 ;
        RECT 12.150 53.790 13.030 56.190 ;
        RECT 13.330 53.790 14.180 56.190 ;
        RECT 14.580 53.440 33.780 56.540 ;
        RECT 34.180 53.790 35.030 56.190 ;
        RECT 12.150 51.040 13.010 53.390 ;
        RECT 13.330 52.290 35.030 53.440 ;
        RECT 13.330 51.040 16.530 52.290 ;
        RECT 18.930 51.040 29.430 51.890 ;
        RECT 31.830 51.040 35.030 52.290 ;
      LAYER via3 ;
        RECT 12.330 74.740 12.980 76.740 ;
        RECT 13.430 75.940 14.280 76.790 ;
        RECT 15.530 75.940 16.380 76.790 ;
        RECT 19.030 76.140 19.680 76.790 ;
        RECT 19.830 76.140 20.480 76.790 ;
        RECT 27.880 76.140 28.530 76.790 ;
        RECT 28.680 76.140 29.330 76.790 ;
        RECT 31.980 75.940 32.830 76.790 ;
        RECT 34.080 75.940 34.930 76.790 ;
        RECT 13.430 74.640 14.280 75.490 ;
        RECT 34.080 74.640 34.930 75.490 ;
        RECT 12.250 71.840 12.930 74.040 ;
        RECT 13.430 73.040 14.080 74.040 ;
        RECT 13.430 71.840 14.080 72.840 ;
        RECT 34.280 73.040 34.930 74.040 ;
        RECT 34.280 71.840 34.930 72.840 ;
        RECT 13.430 70.390 14.280 71.240 ;
        RECT 34.080 70.390 34.930 71.240 ;
        RECT 13.430 69.090 14.280 69.940 ;
        RECT 15.530 69.090 16.380 69.940 ;
        RECT 19.030 69.090 19.680 69.740 ;
        RECT 19.830 69.090 20.480 69.740 ;
        RECT 27.880 69.090 28.530 69.740 ;
        RECT 28.680 69.090 29.330 69.740 ;
        RECT 31.980 69.090 32.830 69.940 ;
        RECT 34.080 69.090 34.930 69.940 ;
        RECT 10.330 59.190 11.730 60.140 ;
        RECT 36.880 59.190 38.280 60.140 ;
        RECT 13.430 57.990 14.280 58.840 ;
        RECT 15.530 57.990 16.380 58.840 ;
        RECT 19.030 58.190 19.680 58.840 ;
        RECT 19.830 58.190 20.480 58.840 ;
        RECT 27.880 58.190 28.530 58.840 ;
        RECT 28.680 58.190 29.330 58.840 ;
        RECT 31.980 57.990 32.830 58.840 ;
        RECT 34.080 57.990 34.930 58.840 ;
        RECT 13.430 56.690 14.280 57.540 ;
        RECT 34.080 56.690 34.930 57.540 ;
        RECT 12.280 53.890 12.930 56.090 ;
        RECT 13.430 55.090 14.080 56.090 ;
        RECT 13.430 53.890 14.080 54.890 ;
        RECT 34.280 55.090 34.930 56.090 ;
        RECT 34.280 53.890 34.930 54.890 ;
        RECT 12.280 51.190 12.940 53.240 ;
        RECT 13.430 52.440 14.280 53.290 ;
        RECT 34.080 52.440 34.930 53.290 ;
        RECT 13.430 51.140 14.280 51.990 ;
        RECT 15.530 51.140 16.380 51.990 ;
        RECT 19.030 51.140 19.680 51.790 ;
        RECT 19.830 51.140 20.480 51.790 ;
        RECT 27.880 51.140 28.530 51.790 ;
        RECT 28.680 51.140 29.330 51.790 ;
        RECT 31.980 51.140 32.830 51.990 ;
        RECT 34.080 51.140 34.930 51.990 ;
      LAYER met4 ;
        RECT 10.220 50.000 11.820 77.980 ;
        RECT 12.150 75.840 16.480 76.890 ;
        RECT 12.150 74.540 14.380 75.840 ;
        RECT 18.930 75.440 29.430 76.890 ;
        RECT 31.880 75.840 35.030 76.890 ;
        RECT 14.780 74.140 33.580 75.440 ;
        RECT 33.980 74.540 35.030 75.840 ;
        RECT 12.150 71.740 35.030 74.140 ;
        RECT 13.330 70.040 14.380 71.340 ;
        RECT 14.780 70.440 33.580 71.740 ;
        RECT 13.330 68.990 16.480 70.040 ;
        RECT 18.930 68.990 29.430 70.440 ;
        RECT 33.980 70.040 35.030 71.340 ;
        RECT 31.880 68.990 35.030 70.040 ;
        RECT 13.330 57.890 16.480 58.940 ;
        RECT 13.330 56.590 14.380 57.890 ;
        RECT 18.930 57.490 29.430 58.940 ;
        RECT 31.880 57.890 35.030 58.940 ;
        RECT 14.780 56.190 33.580 57.490 ;
        RECT 33.980 56.590 35.030 57.890 ;
        RECT 12.150 53.790 35.030 56.190 ;
        RECT 12.150 52.090 14.380 53.390 ;
        RECT 14.780 52.490 33.580 53.790 ;
        RECT 12.150 51.040 16.480 52.090 ;
        RECT 18.930 51.040 29.430 52.490 ;
        RECT 33.980 52.090 35.030 53.390 ;
        RECT 31.880 51.040 35.030 52.090 ;
        RECT 36.780 50.000 38.380 77.980 ;
    END
  END VGND
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.189000 ;
    PORT
      LAYER li1 ;
        RECT 13.310 61.790 13.580 62.120 ;
      LAYER mcon ;
        RECT 13.390 61.870 13.560 62.040 ;
      LAYER met1 ;
        RECT 13.280 62.030 13.590 62.120 ;
        RECT 8.010 61.890 13.590 62.030 ;
        RECT 13.280 61.790 13.590 61.890 ;
    END
  END clk
  PIN inp
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.200000 ;
    PORT
      LAYER li1 ;
        RECT 18.840 65.220 19.200 65.520 ;
      LAYER mcon ;
        RECT 18.920 65.270 19.120 65.470 ;
      LAYER met1 ;
        RECT 8.010 65.410 19.200 65.550 ;
        RECT 18.840 65.220 19.200 65.410 ;
    END
  END inp
  PIN inn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.200000 ;
    PORT
      LAYER li1 ;
        RECT 16.880 64.970 17.240 65.270 ;
      LAYER mcon ;
        RECT 16.960 65.020 17.160 65.220 ;
      LAYER met1 ;
        RECT 8.010 65.130 17.240 65.270 ;
        RECT 16.880 64.970 17.240 65.130 ;
    END
  END inn
  PIN comp_trig
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.756400 ;
    PORT
      LAYER li1 ;
        RECT 31.490 61.230 31.660 63.340 ;
        RECT 32.450 62.880 32.720 63.340 ;
        RECT 32.550 62.780 32.720 62.880 ;
        RECT 32.550 62.590 34.580 62.780 ;
        RECT 33.410 61.230 33.580 62.590 ;
        RECT 33.900 62.540 34.580 62.590 ;
      LAYER mcon ;
        RECT 31.490 62.960 31.660 63.260 ;
        RECT 32.450 62.960 32.620 63.260 ;
        RECT 33.960 62.570 34.140 62.750 ;
        RECT 34.340 62.570 34.520 62.750 ;
      LAYER met1 ;
        RECT 31.460 63.180 31.690 63.320 ;
        RECT 32.420 63.180 32.650 63.320 ;
        RECT 31.460 63.040 32.650 63.180 ;
        RECT 31.460 62.900 31.690 63.040 ;
        RECT 32.420 62.900 32.650 63.040 ;
        RECT 33.900 62.730 34.580 62.780 ;
        RECT 33.900 62.590 40.330 62.730 ;
        RECT 33.900 62.540 34.580 62.590 ;
    END
  END comp_trig
  PIN latch_qn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.303000 ;
    ANTENNADIFFAREA 0.756400 ;
    PORT
      LAYER li1 ;
        RECT 31.270 65.810 31.600 66.070 ;
        RECT 33.170 64.980 33.340 67.090 ;
        RECT 35.090 65.730 35.260 67.090 ;
        RECT 34.230 65.540 35.380 65.730 ;
        RECT 34.230 65.440 34.400 65.540 ;
        RECT 34.710 65.490 35.380 65.540 ;
        RECT 34.130 64.980 34.400 65.440 ;
      LAYER mcon ;
        RECT 31.350 65.860 31.520 66.030 ;
        RECT 34.770 65.520 34.950 65.700 ;
        RECT 35.140 65.520 35.320 65.700 ;
        RECT 33.170 65.060 33.340 65.360 ;
        RECT 34.130 65.060 34.300 65.360 ;
      LAYER met1 ;
        RECT 31.270 66.050 31.600 66.070 ;
        RECT 30.610 65.870 32.400 66.050 ;
        RECT 31.270 65.810 31.600 65.870 ;
        RECT 32.220 65.310 32.400 65.870 ;
        RECT 34.710 65.680 35.380 65.730 ;
        RECT 34.710 65.540 40.330 65.680 ;
        RECT 34.710 65.490 35.380 65.540 ;
        RECT 33.140 65.310 33.370 65.420 ;
        RECT 32.220 65.280 33.370 65.310 ;
        RECT 34.100 65.280 34.330 65.420 ;
        RECT 32.220 65.140 34.330 65.280 ;
        RECT 32.220 65.130 33.370 65.140 ;
        RECT 33.140 65.000 33.370 65.130 ;
        RECT 34.100 65.000 34.330 65.140 ;
    END
  END latch_qn
  PIN latch_q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.303000 ;
    ANTENNADIFFAREA 0.756400 ;
    PORT
      LAYER li1 ;
        RECT 30.690 64.980 30.860 67.090 ;
        RECT 32.610 65.780 32.780 67.090 ;
        RECT 33.750 65.810 34.080 66.070 ;
        RECT 32.610 65.730 32.850 65.780 ;
        RECT 31.750 65.540 32.850 65.730 ;
        RECT 31.750 65.440 31.920 65.540 ;
        RECT 31.650 64.980 31.920 65.440 ;
      LAYER mcon ;
        RECT 33.830 65.860 34.000 66.030 ;
        RECT 32.650 65.580 32.820 65.750 ;
        RECT 30.690 65.060 30.860 65.360 ;
        RECT 31.650 65.060 31.820 65.360 ;
      LAYER met1 ;
        RECT 33.750 66.060 34.080 66.070 ;
        RECT 33.690 66.050 35.280 66.060 ;
        RECT 32.670 66.020 35.280 66.050 ;
        RECT 32.670 65.880 40.330 66.020 ;
        RECT 32.670 65.870 34.080 65.880 ;
        RECT 32.670 65.810 32.850 65.870 ;
        RECT 33.750 65.810 34.080 65.870 ;
        RECT 32.610 65.520 32.850 65.810 ;
        RECT 30.660 65.280 30.890 65.420 ;
        RECT 31.620 65.280 31.850 65.420 ;
        RECT 30.660 65.140 31.850 65.280 ;
        RECT 30.660 65.000 30.890 65.140 ;
        RECT 31.620 65.000 31.850 65.140 ;
    END
  END latch_q
  OBS
      LAYER li1 ;
        RECT 14.530 74.490 17.330 74.690 ;
        RECT 14.530 73.890 15.080 74.490 ;
        RECT 14.530 73.690 17.330 73.890 ;
        RECT 14.530 73.090 15.080 73.690 ;
        RECT 18.080 73.140 18.280 74.690 ;
        RECT 18.880 73.140 19.080 74.690 ;
        RECT 19.680 73.140 19.880 74.690 ;
        RECT 20.480 73.140 20.680 74.690 ;
        RECT 21.280 73.140 21.480 74.690 ;
        RECT 22.080 73.140 22.280 74.690 ;
        RECT 22.880 73.140 23.080 74.690 ;
        RECT 23.680 73.140 23.880 74.690 ;
        RECT 24.480 73.140 24.680 74.690 ;
        RECT 25.280 73.140 25.480 74.690 ;
        RECT 26.080 73.140 26.280 74.690 ;
        RECT 26.880 73.140 27.080 74.690 ;
        RECT 27.680 73.140 27.880 74.690 ;
        RECT 28.480 73.140 28.680 74.690 ;
        RECT 29.280 73.140 29.480 74.690 ;
        RECT 30.080 73.140 30.280 74.690 ;
        RECT 31.030 74.490 33.830 74.690 ;
        RECT 33.280 73.890 33.830 74.490 ;
        RECT 31.030 73.690 33.830 73.890 ;
        RECT 18.080 73.090 30.280 73.140 ;
        RECT 33.280 73.090 33.830 73.690 ;
        RECT 14.530 72.790 33.830 73.090 ;
        RECT 14.530 72.190 15.080 72.790 ;
        RECT 18.080 72.740 30.280 72.790 ;
        RECT 14.530 71.990 17.330 72.190 ;
        RECT 14.530 71.390 15.080 71.990 ;
        RECT 14.530 71.190 17.330 71.390 ;
        RECT 18.080 71.190 18.280 72.740 ;
        RECT 18.880 71.190 19.080 72.740 ;
        RECT 19.680 71.190 19.880 72.740 ;
        RECT 20.480 71.190 20.680 72.740 ;
        RECT 21.280 71.190 21.480 72.740 ;
        RECT 22.080 71.190 22.280 72.740 ;
        RECT 22.880 71.190 23.080 72.740 ;
        RECT 23.680 71.240 23.880 72.740 ;
        RECT 24.480 71.240 24.680 72.740 ;
        RECT 25.280 71.190 25.480 72.740 ;
        RECT 26.080 71.190 26.280 72.740 ;
        RECT 26.880 71.190 27.080 72.740 ;
        RECT 27.680 71.190 27.880 72.740 ;
        RECT 28.480 71.190 28.680 72.740 ;
        RECT 29.280 71.190 29.480 72.740 ;
        RECT 30.080 71.190 30.280 72.740 ;
        RECT 33.280 72.190 33.830 72.790 ;
        RECT 31.030 71.990 33.830 72.190 ;
        RECT 33.280 71.390 33.830 71.990 ;
        RECT 31.030 71.190 33.830 71.390 ;
        RECT 16.530 66.090 16.700 66.930 ;
        RECT 17.490 66.090 17.660 66.930 ;
        RECT 16.530 65.920 17.660 66.090 ;
        RECT 18.450 66.090 18.620 66.930 ;
        RECT 19.410 66.090 19.580 66.930 ;
        RECT 20.530 66.290 21.480 67.240 ;
        RECT 21.710 66.850 22.840 67.020 ;
        RECT 18.450 65.920 19.580 66.090 ;
        RECT 15.510 65.620 15.840 65.910 ;
        RECT 13.750 63.400 14.170 63.430 ;
        RECT 14.920 63.400 15.340 63.430 ;
        RECT 13.730 63.210 14.190 63.400 ;
        RECT 14.900 63.210 15.360 63.400 ;
        RECT 13.730 62.310 14.190 62.480 ;
        RECT 14.900 62.310 15.360 62.480 ;
        RECT 13.750 62.070 14.170 62.310 ;
        RECT 14.480 62.070 14.750 62.120 ;
        RECT 13.750 61.840 14.750 62.070 ;
        RECT 13.750 61.670 14.170 61.840 ;
        RECT 14.480 61.790 14.750 61.840 ;
        RECT 14.920 62.070 15.340 62.310 ;
        RECT 15.610 62.070 15.840 65.620 ;
        RECT 16.530 64.800 16.700 65.920 ;
        RECT 17.420 64.800 17.660 65.100 ;
        RECT 16.530 64.630 17.660 64.800 ;
        RECT 14.920 61.920 15.840 62.070 ;
        RECT 16.050 62.150 16.220 64.360 ;
        RECT 16.530 62.320 16.700 64.630 ;
        RECT 17.010 62.150 17.180 64.360 ;
        RECT 17.490 62.320 17.660 64.630 ;
        RECT 18.450 64.810 18.620 65.920 ;
        RECT 18.450 64.640 20.830 64.810 ;
        RECT 17.970 62.150 18.140 64.360 ;
        RECT 18.450 62.320 18.620 64.640 ;
        RECT 18.930 62.150 19.100 64.360 ;
        RECT 19.410 62.320 19.580 64.640 ;
        RECT 19.890 62.150 20.060 64.360 ;
        RECT 20.450 64.190 20.830 64.640 ;
        RECT 21.060 64.360 21.440 66.290 ;
        RECT 20.450 63.130 21.440 64.190 ;
        RECT 21.710 64.050 21.880 66.850 ;
        RECT 22.190 64.390 22.360 66.680 ;
        RECT 22.670 64.640 22.840 66.850 ;
        RECT 25.890 66.850 27.020 67.020 ;
        RECT 23.800 64.390 23.970 66.680 ;
        RECT 22.190 64.220 23.970 64.390 ;
        RECT 24.760 64.390 24.930 66.680 ;
        RECT 25.890 64.640 26.060 66.850 ;
        RECT 26.370 64.390 26.540 66.680 ;
        RECT 24.760 64.220 26.540 64.390 ;
        RECT 26.850 65.950 27.020 66.850 ;
        RECT 26.850 65.260 27.840 65.950 ;
        RECT 28.010 65.900 28.180 67.330 ;
        RECT 28.010 65.560 28.800 65.900 ;
        RECT 28.970 65.720 29.140 67.330 ;
        RECT 30.690 67.260 31.020 67.520 ;
        RECT 33.170 67.260 33.500 67.520 ;
        RECT 31.170 66.250 31.340 67.090 ;
        RECT 32.130 66.250 32.300 67.090 ;
        RECT 33.650 66.250 33.820 67.090 ;
        RECT 34.610 66.250 34.780 67.090 ;
        RECT 29.510 65.720 29.810 65.770 ;
        RECT 26.850 64.050 27.020 65.260 ;
        RECT 28.010 64.660 28.180 65.560 ;
        RECT 28.970 65.530 29.880 65.720 ;
        RECT 28.970 64.660 29.140 65.530 ;
        RECT 29.510 65.470 29.810 65.530 ;
        RECT 21.630 63.880 23.690 64.050 ;
        RECT 23.870 63.880 27.080 64.050 ;
        RECT 23.520 63.710 23.690 63.880 ;
        RECT 23.520 63.540 24.870 63.710 ;
        RECT 16.050 61.970 20.060 62.150 ;
        RECT 14.920 61.840 15.880 61.920 ;
        RECT 14.920 61.670 15.340 61.840 ;
        RECT 13.730 61.500 14.190 61.670 ;
        RECT 14.900 61.500 15.360 61.670 ;
        RECT 15.550 61.650 15.880 61.840 ;
        RECT 13.750 61.470 14.170 61.500 ;
        RECT 14.920 61.470 15.340 61.500 ;
        RECT 16.050 61.020 16.220 61.970 ;
        RECT 17.010 61.020 17.180 61.970 ;
        RECT 17.970 61.020 18.140 61.970 ;
        RECT 18.930 61.020 19.100 61.970 ;
        RECT 19.890 61.020 20.060 61.970 ;
        RECT 21.060 61.840 21.440 63.130 ;
        RECT 21.030 60.890 21.980 61.840 ;
        RECT 23.800 60.990 23.970 63.540 ;
        RECT 25.090 63.370 25.260 63.880 ;
        RECT 24.760 63.200 25.260 63.370 ;
        RECT 26.140 63.210 26.750 63.550 ;
        RECT 24.760 60.990 24.930 63.200 ;
        RECT 28.010 62.740 28.180 63.640 ;
        RECT 28.970 62.770 29.140 63.640 ;
        RECT 29.530 62.770 29.830 62.820 ;
        RECT 28.010 62.400 28.800 62.740 ;
        RECT 28.970 62.580 29.890 62.770 ;
        RECT 28.010 60.970 28.180 62.400 ;
        RECT 28.970 60.970 29.140 62.580 ;
        RECT 29.530 62.520 29.830 62.580 ;
        RECT 30.510 61.060 30.750 64.730 ;
        RECT 30.920 62.280 31.160 64.260 ;
        RECT 32.070 62.250 32.400 62.510 ;
        RECT 31.970 61.230 32.140 62.070 ;
        RECT 32.930 61.230 33.100 62.070 ;
        RECT 30.510 60.800 31.820 61.060 ;
        RECT 22.390 60.400 23.110 60.670 ;
        RECT 14.530 56.540 17.330 56.740 ;
        RECT 14.530 55.940 15.080 56.540 ;
        RECT 14.530 55.740 17.330 55.940 ;
        RECT 14.530 55.140 15.080 55.740 ;
        RECT 18.080 55.190 18.280 56.740 ;
        RECT 18.880 55.190 19.080 56.740 ;
        RECT 19.680 55.190 19.880 56.740 ;
        RECT 20.480 55.190 20.680 56.740 ;
        RECT 21.280 55.190 21.480 56.740 ;
        RECT 22.080 55.190 22.280 56.740 ;
        RECT 22.880 55.190 23.080 56.740 ;
        RECT 23.680 55.190 23.880 56.740 ;
        RECT 24.480 55.190 24.680 56.740 ;
        RECT 25.280 55.190 25.480 56.740 ;
        RECT 26.080 55.190 26.280 56.740 ;
        RECT 26.880 55.190 27.080 56.740 ;
        RECT 27.680 55.190 27.880 56.740 ;
        RECT 28.480 55.190 28.680 56.740 ;
        RECT 29.280 55.190 29.480 56.740 ;
        RECT 30.080 55.190 30.280 56.740 ;
        RECT 31.030 56.540 33.830 56.740 ;
        RECT 33.280 55.940 33.830 56.540 ;
        RECT 31.030 55.740 33.830 55.940 ;
        RECT 18.080 55.140 30.280 55.190 ;
        RECT 33.280 55.140 33.830 55.740 ;
        RECT 14.530 54.840 33.830 55.140 ;
        RECT 14.530 54.240 15.080 54.840 ;
        RECT 18.080 54.790 30.280 54.840 ;
        RECT 14.530 54.040 17.330 54.240 ;
        RECT 14.530 53.440 15.080 54.040 ;
        RECT 14.530 53.240 17.330 53.440 ;
        RECT 18.080 53.240 18.280 54.790 ;
        RECT 18.880 53.240 19.080 54.790 ;
        RECT 19.680 53.240 19.880 54.790 ;
        RECT 20.480 53.240 20.680 54.790 ;
        RECT 21.280 53.240 21.480 54.790 ;
        RECT 22.080 53.240 22.280 54.790 ;
        RECT 22.880 53.240 23.080 54.790 ;
        RECT 23.680 53.290 23.880 54.790 ;
        RECT 24.480 53.290 24.680 54.790 ;
        RECT 25.280 53.240 25.480 54.790 ;
        RECT 26.080 53.240 26.280 54.790 ;
        RECT 26.880 53.240 27.080 54.790 ;
        RECT 27.680 53.240 27.880 54.790 ;
        RECT 28.480 53.240 28.680 54.790 ;
        RECT 29.280 53.240 29.480 54.790 ;
        RECT 30.080 53.240 30.280 54.790 ;
        RECT 33.280 54.240 33.830 54.840 ;
        RECT 31.030 54.040 33.830 54.240 ;
        RECT 33.280 53.440 33.830 54.040 ;
        RECT 31.030 53.240 33.830 53.440 ;
      LAYER mcon ;
        RECT 14.630 73.540 14.880 73.790 ;
        RECT 14.630 73.090 14.880 73.340 ;
        RECT 33.480 73.490 33.730 73.740 ;
        RECT 33.480 73.040 33.730 73.290 ;
        RECT 14.630 72.590 14.880 72.840 ;
        RECT 14.630 72.140 14.880 72.390 ;
        RECT 33.480 72.540 33.730 72.790 ;
        RECT 33.480 72.090 33.730 72.340 ;
        RECT 20.630 66.390 21.380 67.140 ;
        RECT 13.810 63.220 14.110 63.390 ;
        RECT 14.980 63.220 15.280 63.390 ;
        RECT 13.810 62.310 14.110 62.480 ;
        RECT 14.980 62.310 15.280 62.480 ;
        RECT 14.560 61.870 14.730 62.040 ;
        RECT 17.450 64.890 17.630 65.070 ;
        RECT 21.160 65.240 21.340 65.420 ;
        RECT 21.160 64.870 21.340 65.050 ;
        RECT 21.160 64.500 21.340 64.680 ;
        RECT 21.160 63.950 21.340 64.130 ;
        RECT 27.630 65.700 27.810 65.870 ;
        RECT 27.630 65.340 27.810 65.510 ;
        RECT 33.250 67.320 33.420 67.490 ;
        RECT 29.540 65.530 29.720 65.710 ;
        RECT 21.160 63.570 21.340 63.750 ;
        RECT 21.160 63.200 21.340 63.380 ;
        RECT 21.130 60.990 21.880 61.740 ;
        RECT 26.170 63.290 26.350 63.470 ;
        RECT 26.540 63.290 26.720 63.470 ;
        RECT 29.570 62.580 29.740 62.760 ;
        RECT 30.540 62.640 30.720 62.820 ;
        RECT 30.950 64.020 31.130 64.200 ;
        RECT 30.950 62.340 31.130 62.520 ;
        RECT 32.150 62.290 32.320 62.460 ;
        RECT 22.470 60.450 22.640 60.620 ;
        RECT 22.860 60.450 23.030 60.620 ;
        RECT 14.630 55.590 14.880 55.840 ;
        RECT 14.630 55.140 14.880 55.390 ;
        RECT 33.480 55.540 33.730 55.790 ;
        RECT 33.480 55.090 33.730 55.340 ;
        RECT 14.630 54.640 14.880 54.890 ;
        RECT 14.630 54.190 14.880 54.440 ;
        RECT 33.480 54.590 33.730 54.840 ;
        RECT 33.480 54.140 33.730 54.390 ;
      LAYER met1 ;
        RECT 18.930 75.690 29.430 76.890 ;
        RECT 23.880 75.240 24.480 75.690 ;
        RECT 18.280 75.090 30.080 75.240 ;
        RECT 13.330 73.240 14.980 73.890 ;
        RECT 15.430 73.240 15.580 74.740 ;
        RECT 16.030 73.240 16.180 74.740 ;
        RECT 16.630 73.240 16.780 74.740 ;
        RECT 17.230 73.240 17.380 74.740 ;
        RECT 23.880 74.640 24.480 75.090 ;
        RECT 18.280 74.490 30.080 74.640 ;
        RECT 23.880 74.040 24.480 74.490 ;
        RECT 18.280 73.890 30.080 74.040 ;
        RECT 23.880 73.440 24.480 73.890 ;
        RECT 18.280 73.290 30.080 73.440 ;
        RECT 13.330 73.140 17.380 73.240 ;
        RECT 23.880 73.140 24.480 73.290 ;
        RECT 30.980 73.240 31.130 74.740 ;
        RECT 31.580 73.240 31.730 74.740 ;
        RECT 32.180 73.240 32.330 74.740 ;
        RECT 32.780 73.240 32.930 74.740 ;
        RECT 33.380 73.240 35.030 73.840 ;
        RECT 30.980 73.140 35.030 73.240 ;
        RECT 13.330 72.440 35.030 73.140 ;
        RECT 13.330 72.040 14.980 72.440 ;
        RECT 15.430 71.140 15.580 72.440 ;
        RECT 16.030 71.140 16.180 72.440 ;
        RECT 16.630 71.140 16.780 72.440 ;
        RECT 17.230 71.140 17.380 72.440 ;
        RECT 23.880 71.990 24.480 72.440 ;
        RECT 18.280 71.840 30.080 71.990 ;
        RECT 23.880 71.390 24.480 71.840 ;
        RECT 18.280 71.240 30.080 71.390 ;
        RECT 23.880 70.790 24.480 71.240 ;
        RECT 30.980 71.140 31.130 72.440 ;
        RECT 31.580 71.140 31.730 72.440 ;
        RECT 32.180 71.140 32.330 72.440 ;
        RECT 32.780 71.140 32.930 72.440 ;
        RECT 33.380 71.990 35.030 72.440 ;
        RECT 18.280 70.640 30.080 70.790 ;
        RECT 23.880 70.190 24.480 70.640 ;
        RECT 18.930 68.990 29.430 70.190 ;
        RECT 29.810 67.520 31.030 67.550 ;
        RECT 29.810 67.380 33.480 67.520 ;
        RECT 20.530 66.290 21.480 67.240 ;
        RECT 17.390 65.080 17.660 65.100 ;
        RECT 21.100 65.080 21.400 65.470 ;
        RECT 27.560 65.250 27.840 65.950 ;
        RECT 29.810 65.770 29.990 67.380 ;
        RECT 33.170 67.290 33.480 67.380 ;
        RECT 29.510 65.470 29.990 65.770 ;
        RECT 17.390 65.010 21.400 65.080 ;
        RECT 17.380 64.820 21.400 65.010 ;
        RECT 21.100 64.470 21.400 64.820 ;
        RECT 29.810 64.260 29.990 65.470 ;
        RECT 13.770 62.250 14.160 63.460 ;
        RECT 14.940 62.250 15.330 63.460 ;
        RECT 21.100 63.390 21.400 64.160 ;
        RECT 29.810 64.070 31.160 64.260 ;
        RECT 30.920 63.960 31.160 64.070 ;
        RECT 26.120 63.390 26.770 63.550 ;
        RECT 21.100 63.210 26.770 63.390 ;
        RECT 21.100 63.170 21.400 63.210 ;
        RECT 29.530 62.770 29.830 62.820 ;
        RECT 30.510 62.770 30.750 62.880 ;
        RECT 29.530 62.580 30.750 62.770 ;
        RECT 29.530 62.520 29.830 62.580 ;
        RECT 30.920 62.450 31.160 62.580 ;
        RECT 32.070 62.450 32.400 62.510 ;
        RECT 30.920 62.270 32.400 62.450 ;
        RECT 30.920 62.260 31.410 62.270 ;
        RECT 32.070 62.250 32.400 62.270 ;
        RECT 14.480 61.950 14.760 62.120 ;
        RECT 14.480 61.790 15.780 61.950 ;
        RECT 15.570 60.670 15.780 61.790 ;
        RECT 21.030 60.890 21.980 61.840 ;
        RECT 15.570 60.400 23.110 60.670 ;
        RECT 18.930 57.740 29.430 58.940 ;
        RECT 23.880 57.290 24.480 57.740 ;
        RECT 18.280 57.140 30.080 57.290 ;
        RECT 13.330 55.290 14.980 55.940 ;
        RECT 15.430 55.290 15.580 56.790 ;
        RECT 16.030 55.290 16.180 56.790 ;
        RECT 16.630 55.290 16.780 56.790 ;
        RECT 17.230 55.290 17.380 56.790 ;
        RECT 23.880 56.690 24.480 57.140 ;
        RECT 18.280 56.540 30.080 56.690 ;
        RECT 23.880 56.090 24.480 56.540 ;
        RECT 18.280 55.940 30.080 56.090 ;
        RECT 23.880 55.490 24.480 55.940 ;
        RECT 18.280 55.340 30.080 55.490 ;
        RECT 13.330 55.190 17.380 55.290 ;
        RECT 23.880 55.190 24.480 55.340 ;
        RECT 30.980 55.290 31.130 56.790 ;
        RECT 31.580 55.290 31.730 56.790 ;
        RECT 32.180 55.290 32.330 56.790 ;
        RECT 32.780 55.290 32.930 56.790 ;
        RECT 33.380 55.290 35.030 55.890 ;
        RECT 30.980 55.190 35.030 55.290 ;
        RECT 13.330 54.490 35.030 55.190 ;
        RECT 13.330 54.090 14.980 54.490 ;
        RECT 15.430 53.190 15.580 54.490 ;
        RECT 16.030 53.190 16.180 54.490 ;
        RECT 16.630 53.190 16.780 54.490 ;
        RECT 17.230 53.190 17.380 54.490 ;
        RECT 23.880 54.040 24.480 54.490 ;
        RECT 18.280 53.890 30.080 54.040 ;
        RECT 23.880 53.440 24.480 53.890 ;
        RECT 18.280 53.290 30.080 53.440 ;
        RECT 23.880 52.840 24.480 53.290 ;
        RECT 30.980 53.190 31.130 54.490 ;
        RECT 31.580 53.190 31.730 54.490 ;
        RECT 32.180 53.190 32.330 54.490 ;
        RECT 32.780 53.190 32.930 54.490 ;
        RECT 33.380 54.040 35.030 54.490 ;
        RECT 18.280 52.690 30.080 52.840 ;
        RECT 23.880 52.240 24.480 52.690 ;
        RECT 18.930 51.040 29.430 52.240 ;
      LAYER via ;
        RECT 19.030 75.790 20.030 76.790 ;
        RECT 20.130 75.790 21.130 76.790 ;
        RECT 23.730 75.790 24.630 76.790 ;
        RECT 27.230 75.790 28.230 76.790 ;
        RECT 28.330 75.790 29.330 76.790 ;
        RECT 13.430 73.190 14.430 73.740 ;
        RECT 33.930 73.190 34.930 73.740 ;
        RECT 13.430 72.140 14.430 72.690 ;
        RECT 33.930 72.140 34.930 72.690 ;
        RECT 19.030 69.090 20.030 70.090 ;
        RECT 20.130 69.090 21.130 70.090 ;
        RECT 23.730 69.090 24.630 70.090 ;
        RECT 27.230 69.090 28.230 70.090 ;
        RECT 28.330 69.090 29.330 70.090 ;
        RECT 20.630 66.390 21.380 67.140 ;
        RECT 21.130 60.990 21.880 61.740 ;
        RECT 19.030 57.840 20.030 58.840 ;
        RECT 20.130 57.840 21.130 58.840 ;
        RECT 23.730 57.840 24.630 58.840 ;
        RECT 27.230 57.840 28.230 58.840 ;
        RECT 28.330 57.840 29.330 58.840 ;
        RECT 13.430 55.240 14.430 55.790 ;
        RECT 33.930 55.240 34.930 55.790 ;
        RECT 13.430 54.190 14.430 54.740 ;
        RECT 33.930 54.190 34.930 54.740 ;
        RECT 19.030 51.140 20.030 52.140 ;
        RECT 20.130 51.140 21.130 52.140 ;
        RECT 23.730 51.140 24.630 52.140 ;
        RECT 27.230 51.140 28.230 52.140 ;
        RECT 28.330 51.140 29.330 52.140 ;
      LAYER met2 ;
        RECT 18.930 75.490 29.430 76.890 ;
        RECT 15.430 74.890 32.930 75.490 ;
        RECT 17.430 74.440 17.730 74.890 ;
        RECT 15.430 74.290 17.730 74.440 ;
        RECT 17.430 73.840 17.730 74.290 ;
        RECT 13.330 72.040 14.530 73.840 ;
        RECT 15.430 73.690 17.730 73.840 ;
        RECT 17.430 73.240 17.730 73.690 ;
        RECT 18.180 73.240 18.330 74.890 ;
        RECT 18.780 73.240 18.930 74.890 ;
        RECT 19.380 73.240 19.530 74.890 ;
        RECT 19.980 73.240 20.130 74.890 ;
        RECT 20.580 73.240 20.730 74.890 ;
        RECT 21.180 73.240 21.330 74.890 ;
        RECT 21.780 73.240 21.930 74.890 ;
        RECT 22.380 73.240 22.530 74.890 ;
        RECT 22.980 73.240 23.130 74.890 ;
        RECT 23.580 73.240 23.730 74.890 ;
        RECT 24.630 73.240 24.780 74.890 ;
        RECT 25.230 73.240 25.380 74.890 ;
        RECT 25.830 73.240 25.980 74.890 ;
        RECT 26.430 73.240 26.580 74.890 ;
        RECT 27.030 73.240 27.180 74.890 ;
        RECT 27.630 73.240 27.780 74.890 ;
        RECT 28.230 73.240 28.380 74.890 ;
        RECT 28.830 73.240 28.980 74.890 ;
        RECT 29.430 73.240 29.580 74.890 ;
        RECT 30.030 73.240 30.180 74.890 ;
        RECT 30.630 74.440 30.930 74.890 ;
        RECT 30.630 74.290 32.930 74.440 ;
        RECT 30.630 73.840 30.930 74.290 ;
        RECT 30.630 73.690 32.930 73.840 ;
        RECT 30.630 73.240 30.930 73.690 ;
        RECT 17.430 72.190 17.730 72.640 ;
        RECT 15.430 72.040 17.730 72.190 ;
        RECT 17.430 71.590 17.730 72.040 ;
        RECT 15.430 71.440 17.730 71.590 ;
        RECT 17.430 70.990 17.730 71.440 ;
        RECT 18.180 70.990 18.330 72.640 ;
        RECT 18.780 70.990 18.930 72.640 ;
        RECT 19.380 70.990 19.530 72.640 ;
        RECT 19.980 70.990 20.130 72.640 ;
        RECT 20.580 70.990 20.730 72.640 ;
        RECT 21.180 70.990 21.330 72.640 ;
        RECT 21.780 70.990 21.930 72.640 ;
        RECT 22.380 70.990 22.530 72.640 ;
        RECT 22.980 70.990 23.130 72.640 ;
        RECT 23.580 70.990 23.730 72.640 ;
        RECT 24.630 70.990 24.780 72.640 ;
        RECT 25.230 70.990 25.380 72.640 ;
        RECT 25.830 70.990 25.980 72.640 ;
        RECT 26.430 70.990 26.580 72.640 ;
        RECT 27.030 70.990 27.180 72.640 ;
        RECT 27.630 70.990 27.780 72.640 ;
        RECT 28.230 70.990 28.380 72.640 ;
        RECT 28.830 70.990 28.980 72.640 ;
        RECT 29.430 70.990 29.580 72.640 ;
        RECT 30.030 70.990 30.180 72.640 ;
        RECT 30.630 72.190 30.930 72.640 ;
        RECT 30.630 72.040 32.930 72.190 ;
        RECT 33.830 72.040 35.030 73.840 ;
        RECT 30.630 71.590 30.930 72.040 ;
        RECT 30.630 71.440 32.930 71.590 ;
        RECT 30.630 70.990 30.930 71.440 ;
        RECT 15.430 70.390 32.930 70.990 ;
        RECT 18.930 68.990 29.430 70.390 ;
        RECT 20.530 66.290 21.480 68.990 ;
        RECT 21.030 58.940 21.980 61.840 ;
        RECT 18.930 57.540 29.430 58.940 ;
        RECT 15.430 56.940 32.930 57.540 ;
        RECT 17.430 56.490 17.730 56.940 ;
        RECT 15.430 56.340 17.730 56.490 ;
        RECT 17.430 55.890 17.730 56.340 ;
        RECT 13.330 54.090 14.530 55.890 ;
        RECT 15.430 55.740 17.730 55.890 ;
        RECT 17.430 55.290 17.730 55.740 ;
        RECT 18.180 55.290 18.330 56.940 ;
        RECT 18.780 55.290 18.930 56.940 ;
        RECT 19.380 55.290 19.530 56.940 ;
        RECT 19.980 55.290 20.130 56.940 ;
        RECT 20.580 55.290 20.730 56.940 ;
        RECT 21.180 55.290 21.330 56.940 ;
        RECT 21.780 55.290 21.930 56.940 ;
        RECT 22.380 55.290 22.530 56.940 ;
        RECT 22.980 55.290 23.130 56.940 ;
        RECT 23.580 55.290 23.730 56.940 ;
        RECT 24.630 55.290 24.780 56.940 ;
        RECT 25.230 55.290 25.380 56.940 ;
        RECT 25.830 55.290 25.980 56.940 ;
        RECT 26.430 55.290 26.580 56.940 ;
        RECT 27.030 55.290 27.180 56.940 ;
        RECT 27.630 55.290 27.780 56.940 ;
        RECT 28.230 55.290 28.380 56.940 ;
        RECT 28.830 55.290 28.980 56.940 ;
        RECT 29.430 55.290 29.580 56.940 ;
        RECT 30.030 55.290 30.180 56.940 ;
        RECT 30.630 56.490 30.930 56.940 ;
        RECT 30.630 56.340 32.930 56.490 ;
        RECT 30.630 55.890 30.930 56.340 ;
        RECT 30.630 55.740 32.930 55.890 ;
        RECT 30.630 55.290 30.930 55.740 ;
        RECT 17.430 54.240 17.730 54.690 ;
        RECT 15.430 54.090 17.730 54.240 ;
        RECT 17.430 53.640 17.730 54.090 ;
        RECT 15.430 53.490 17.730 53.640 ;
        RECT 17.430 53.040 17.730 53.490 ;
        RECT 18.180 53.040 18.330 54.690 ;
        RECT 18.780 53.040 18.930 54.690 ;
        RECT 19.380 53.040 19.530 54.690 ;
        RECT 19.980 53.040 20.130 54.690 ;
        RECT 20.580 53.040 20.730 54.690 ;
        RECT 21.180 53.040 21.330 54.690 ;
        RECT 21.780 53.040 21.930 54.690 ;
        RECT 22.380 53.040 22.530 54.690 ;
        RECT 22.980 53.040 23.130 54.690 ;
        RECT 23.580 53.040 23.730 54.690 ;
        RECT 24.630 53.040 24.780 54.690 ;
        RECT 25.230 53.040 25.380 54.690 ;
        RECT 25.830 53.040 25.980 54.690 ;
        RECT 26.430 53.040 26.580 54.690 ;
        RECT 27.030 53.040 27.180 54.690 ;
        RECT 27.630 53.040 27.780 54.690 ;
        RECT 28.230 53.040 28.380 54.690 ;
        RECT 28.830 53.040 28.980 54.690 ;
        RECT 29.430 53.040 29.580 54.690 ;
        RECT 30.030 53.040 30.180 54.690 ;
        RECT 30.630 54.240 30.930 54.690 ;
        RECT 30.630 54.090 32.930 54.240 ;
        RECT 33.830 54.090 35.030 55.890 ;
        RECT 30.630 53.640 30.930 54.090 ;
        RECT 30.630 53.490 32.930 53.640 ;
        RECT 30.630 53.040 30.930 53.490 ;
        RECT 15.430 52.440 32.930 53.040 ;
        RECT 18.930 51.040 29.430 52.440 ;
  END
END adc_comp_latch
END LIBRARY

