magic
tech sky130A
magscale 1 2
timestamp 1673796976
<< nwell >>
rect 6253 13313 6283 13555
rect 3046 12966 3205 13221
rect 3619 12966 3722 13221
rect 4120 12966 4309 13189
rect 2867 12812 2898 12903
rect 2494 12785 2898 12812
rect 2494 12772 2884 12785
rect 2460 12722 2884 12772
rect 2448 12681 2884 12722
rect 2448 12652 2504 12681
rect 2456 12617 2504 12652
rect 2456 12440 2484 12617
rect 2622 12588 2884 12681
rect 2610 12550 2884 12588
rect 2622 12440 2884 12550
rect 2456 12414 2884 12440
rect 5814 12056 6961 12472
<< locali >>
rect 6517 12976 6891 13030
rect 2488 12755 2578 12826
rect 2752 12756 2842 12826
rect 2488 12721 2634 12755
rect 2752 12721 2910 12756
rect 2598 12588 2634 12721
rect 2874 12588 2910 12721
rect 2564 12550 2634 12588
rect 2840 12550 2910 12588
<< viali >>
rect 2488 12366 2550 12408
rect 2764 12366 2824 12405
<< metal1 >>
rect 6155 13457 6213 13466
rect 6155 13395 6156 13457
rect 6155 13386 6213 13395
rect 2756 13201 2946 13277
rect 7390 13225 7396 13249
rect 2756 12826 2842 13201
rect 7285 13197 7396 13225
rect 7452 13197 7458 13249
rect 6294 13010 6358 13011
rect 6185 12982 6300 13010
rect 6294 12957 6300 12982
rect 6352 12957 6358 13010
rect 2488 12772 2842 12826
rect 6275 12781 6477 12809
rect 6275 12722 6303 12781
rect 6185 12694 6303 12722
rect 2756 12668 2834 12681
rect 6329 12677 6477 12678
rect 6329 12624 6335 12677
rect 6387 12650 6477 12677
rect 6387 12624 6393 12650
rect 6245 12567 6297 12573
rect 6233 12515 6245 12538
rect 6233 12510 6297 12515
rect 6245 12509 6297 12510
rect 2382 12419 2445 12426
rect 2434 12367 2445 12419
rect 2382 12359 2445 12367
rect 2476 12408 2560 12420
rect 2476 12366 2488 12408
rect 2550 12404 2560 12408
rect 2666 12404 2718 12426
rect 2550 12366 2718 12404
rect 2476 12358 2718 12366
rect 2752 12405 2836 12418
rect 2752 12366 2764 12405
rect 2824 12404 2836 12405
rect 2824 12366 2932 12404
rect 2752 12358 2932 12366
rect 2666 12352 2718 12358
rect 2430 12052 2857 12156
rect 2885 12134 2932 12358
rect 2885 12080 4100 12134
rect 2628 12050 2857 12052
<< via1 >>
rect 6156 13395 6213 13457
rect 7396 13197 7452 13249
rect 6300 12957 6352 13010
rect 6335 12624 6387 12677
rect 6245 12515 6297 12567
rect 2382 12367 2434 12419
<< metal2 >>
rect 6155 13457 6213 13466
rect 6155 13395 6156 13457
rect 6155 13386 6213 13395
rect 6238 13309 6295 13318
rect 6238 13238 6295 13247
rect 6238 12573 6266 13238
rect 7387 13197 7396 13253
rect 7452 13197 7461 13253
rect 7285 13128 7349 13137
rect 7285 13111 7292 13128
rect 7283 13097 7292 13111
rect 7292 13057 7349 13066
rect 6294 13010 6358 13011
rect 6294 12957 6300 13010
rect 6352 12957 6358 13010
rect 6329 12678 6358 12957
rect 6915 12909 6972 12913
rect 6908 12904 6972 12909
rect 6908 12881 6915 12904
rect 6915 12833 6972 12842
rect 6329 12677 6393 12678
rect 6329 12624 6335 12677
rect 6387 12624 6393 12677
rect 6238 12567 6297 12573
rect 6238 12515 6245 12567
rect 6238 12509 6297 12515
rect 2382 12421 2445 12426
rect 2358 12365 2367 12421
rect 2434 12365 2445 12421
rect 2382 12359 2445 12365
<< via2 >>
rect 6156 13395 6213 13457
rect 6238 13247 6295 13309
rect 7396 13249 7452 13253
rect 7396 13197 7452 13249
rect 7292 13066 7349 13128
rect 6915 12842 6972 12904
rect 2367 12419 2434 12421
rect 2367 12367 2382 12419
rect 2382 12367 2434 12419
rect 2367 12365 2434 12367
<< metal3 >>
rect 2237 13554 3752 13614
rect 2237 13434 3367 13494
rect 3307 13039 3367 13434
rect 3288 12979 3367 13039
rect 3691 13022 3752 13554
rect 6151 13457 6219 13462
rect 6151 13395 6156 13457
rect 6213 13449 6219 13457
rect 6213 13395 6313 13449
rect 6151 13389 6313 13395
rect 6233 13309 6313 13314
rect 6233 13247 6238 13309
rect 6295 13254 6313 13309
rect 6295 13247 6301 13254
rect 6233 13241 6301 13247
rect 7387 13253 7461 13258
rect 7387 13197 7396 13253
rect 7452 13252 7461 13253
rect 7452 13197 8066 13252
rect 7387 13192 8066 13197
rect 7285 13128 7362 13137
rect 7285 13066 7292 13128
rect 7349 13125 7362 13128
rect 7349 13066 8066 13125
rect 7285 13065 8066 13066
rect 7285 13057 7362 13065
rect 3691 12979 3768 13022
rect 3288 12845 3349 12979
rect 3708 12847 3768 12979
rect 6908 12904 6985 12913
rect 6908 12842 6915 12904
rect 6972 12893 6985 12904
rect 6972 12842 8066 12893
rect 6908 12833 8066 12842
rect 2358 12423 2439 12426
rect 2357 12422 2439 12423
rect 2237 12421 2439 12422
rect 2237 12365 2367 12421
rect 2434 12365 2439 12421
rect 2237 12362 2439 12365
rect 2358 12359 2439 12362
<< metal4 >>
rect 7356 10000 7676 15596
rect 7746 10000 8066 15596
use adc_comp_circuit  adc_comp_circuit_0
timestamp 1673796976
transform 1 0 3088 0 1 13378
box -686 -3378 4978 2218
use adc_inverter  adc_inverter_1
timestamp 1673727735
transform 1 0 2690 0 1 12236
box -29 -130 220 582
use adc_inverter  adc_inverter_2
timestamp 1673727735
transform 1 0 2414 0 1 12236
box -29 -130 220 582
use adc_nor  adc_nor_0
timestamp 1673698727
transform 1 0 6455 0 -1 12762
box -8 -214 506 390
use adc_nor_latch  adc_nor_latch_0
timestamp 1673708941
transform 1 0 6123 0 1 12820
box 160 210 1202 814
<< labels >>
flabel metal4 7746 10000 8066 15596 0 FreeSans 1600 90 0 0 VDD
port 1 nsew power bidirectional
flabel metal4 7356 10000 7676 15596 0 FreeSans 1600 90 0 0 VSS
port 2 nsew ground bidirectional
flabel metal3 7942 12833 8066 12893 0 FreeSans 160 0 0 0 comp_trig
port 6 nsew signal output
flabel metal3 7903 13192 8066 13252 0 FreeSans 160 0 0 0 latch_qn
port 7 nsew signal output
flabel metal3 7903 13065 8066 13125 0 FreeSans 160 0 0 0 latch_q
port 8 nsew signal output
flabel metal3 s 2237 12362 2271 12422 7 FreeSans 160 0 0 0 clk
port 3 w signal input
flabel metal3 s 2237 13554 2271 13614 7 FreeSans 160 0 0 0 inp
port 4 w signal input
flabel metal3 s 2237 13434 2271 13494 7 FreeSans 160 0 0 0 inn
port 5 w signal input
<< properties >>
string FIXED_BBOX 0 0 8400 25800
string LEFclass BLOCK
string LEForigin 0 0
string LEFsource USER
<< end >>
