VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO adc_comp_latch
  CLASS BLOCK ;
  FOREIGN adc_comp_latch ;
  ORIGIN 2.790 -13.980 ;
  SIZE 30.050 BY 27.980 ;
  PIN latch_q
    ANTENNAGATEAREA 0.303000 ;
    ANTENNADIFFAREA 0.756400 ;
    PORT
      LAYER li1 ;
        RECT 18.690 28.960 18.860 31.070 ;
        RECT 20.610 29.760 20.780 31.070 ;
        RECT 21.750 29.790 22.080 30.050 ;
        RECT 20.610 29.710 20.850 29.760 ;
        RECT 19.750 29.520 20.850 29.710 ;
        RECT 19.750 29.420 19.920 29.520 ;
        RECT 19.650 28.960 19.920 29.420 ;
      LAYER mcon ;
        RECT 21.830 29.840 22.000 30.010 ;
        RECT 20.650 29.560 20.820 29.730 ;
        RECT 18.690 29.040 18.860 29.340 ;
        RECT 19.650 29.040 19.820 29.340 ;
      LAYER met1 ;
        RECT 21.750 30.040 22.080 30.050 ;
        RECT 21.690 30.030 23.280 30.040 ;
        RECT 20.670 30.000 23.280 30.030 ;
        RECT 20.670 29.860 27.260 30.000 ;
        RECT 20.670 29.850 22.080 29.860 ;
        RECT 20.670 29.790 20.850 29.850 ;
        RECT 21.750 29.790 22.080 29.850 ;
        RECT 20.610 29.500 20.850 29.790 ;
        RECT 18.660 29.260 18.890 29.400 ;
        RECT 19.620 29.260 19.850 29.400 ;
        RECT 18.660 29.120 19.850 29.260 ;
        RECT 18.660 28.980 18.890 29.120 ;
        RECT 19.620 28.980 19.850 29.120 ;
    END
  END latch_q
  PIN latch_qn
    ANTENNAGATEAREA 0.303000 ;
    ANTENNADIFFAREA 0.756400 ;
    PORT
      LAYER li1 ;
        RECT 19.270 29.790 19.600 30.050 ;
        RECT 21.170 28.960 21.340 31.070 ;
        RECT 23.090 29.710 23.260 31.070 ;
        RECT 22.230 29.520 23.380 29.710 ;
        RECT 22.230 29.420 22.400 29.520 ;
        RECT 22.710 29.470 23.380 29.520 ;
        RECT 22.130 28.960 22.400 29.420 ;
      LAYER mcon ;
        RECT 19.350 29.840 19.520 30.010 ;
        RECT 22.770 29.500 22.950 29.680 ;
        RECT 23.140 29.500 23.320 29.680 ;
        RECT 21.170 29.040 21.340 29.340 ;
        RECT 22.130 29.040 22.300 29.340 ;
      LAYER met1 ;
        RECT 19.270 30.030 19.600 30.050 ;
        RECT 18.610 29.850 20.400 30.030 ;
        RECT 19.270 29.790 19.600 29.850 ;
        RECT 20.220 29.290 20.400 29.850 ;
        RECT 22.710 29.660 23.380 29.710 ;
        RECT 22.710 29.520 27.260 29.660 ;
        RECT 22.710 29.470 23.380 29.520 ;
        RECT 21.140 29.290 21.370 29.400 ;
        RECT 20.220 29.260 21.370 29.290 ;
        RECT 22.100 29.260 22.330 29.400 ;
        RECT 20.220 29.120 22.330 29.260 ;
        RECT 20.220 29.110 21.370 29.120 ;
        RECT 21.140 28.980 21.370 29.110 ;
        RECT 22.100 28.980 22.330 29.120 ;
    END
  END latch_qn
  PIN comp_trig
    ANTENNADIFFAREA 0.756400 ;
    PORT
      LAYER li1 ;
        RECT 19.490 25.210 19.660 27.320 ;
        RECT 20.450 26.860 20.720 27.320 ;
        RECT 20.550 26.760 20.720 26.860 ;
        RECT 20.550 26.570 22.580 26.760 ;
        RECT 21.410 25.210 21.580 26.570 ;
        RECT 21.900 26.520 22.580 26.570 ;
      LAYER mcon ;
        RECT 19.490 26.940 19.660 27.240 ;
        RECT 20.450 26.940 20.620 27.240 ;
        RECT 21.960 26.550 22.140 26.730 ;
        RECT 22.340 26.550 22.520 26.730 ;
      LAYER met1 ;
        RECT 19.460 27.160 19.690 27.300 ;
        RECT 20.420 27.160 20.650 27.300 ;
        RECT 19.460 27.020 20.650 27.160 ;
        RECT 19.460 26.880 19.690 27.020 ;
        RECT 20.420 26.880 20.650 27.020 ;
        RECT 21.900 26.710 22.580 26.760 ;
        RECT 21.900 26.570 27.260 26.710 ;
        RECT 21.900 26.520 22.580 26.570 ;
    END
  END comp_trig
  PIN VSS
    ANTENNADIFFAREA 79.479301 ;
    PORT
      LAYER pwell ;
        RECT 4.530 39.970 6.930 40.870 ;
        RECT 17.430 39.970 19.830 40.870 ;
        RECT 2.230 39.570 8.480 39.970 ;
        RECT 11.730 39.570 12.630 39.970 ;
        RECT 15.880 39.570 22.130 39.970 ;
        RECT 2.230 34.270 22.130 39.570 ;
        RECT 2.230 33.870 8.480 34.270 ;
        RECT 11.730 33.870 12.630 34.270 ;
        RECT 15.880 33.870 22.130 34.270 ;
        RECT 4.530 32.970 6.930 33.870 ;
        RECT 17.430 32.970 19.830 33.870 ;
        RECT 4.530 22.020 6.930 22.920 ;
        RECT 17.430 22.020 19.830 22.920 ;
        RECT 2.230 21.620 8.480 22.020 ;
        RECT 11.730 21.620 12.630 22.020 ;
        RECT 15.880 21.620 22.130 22.020 ;
        RECT 2.230 16.320 22.130 21.620 ;
        RECT 2.230 15.920 8.480 16.320 ;
        RECT 11.730 15.920 12.630 16.320 ;
        RECT 15.880 15.920 22.130 16.320 ;
        RECT 4.530 15.020 6.930 15.920 ;
        RECT 17.430 15.020 19.830 15.920 ;
      LAYER li1 ;
        RECT 0.150 40.970 24.540 41.960 ;
        RECT 0.150 38.520 1.330 40.970 ;
        RECT 4.580 40.470 6.880 40.970 ;
        RECT 17.480 40.470 19.780 40.970 ;
        RECT 1.730 40.070 22.630 40.470 ;
        RECT 0.150 14.970 1.140 38.520 ;
        RECT 1.730 33.770 2.130 40.070 ;
        RECT 4.580 40.020 6.880 40.070 ;
        RECT 17.480 40.020 19.780 40.070 ;
        RECT 2.930 38.870 21.430 39.470 ;
        RECT 5.530 38.270 5.880 38.870 ;
        RECT 3.280 38.070 5.880 38.270 ;
        RECT 5.530 37.470 5.880 38.070 ;
        RECT 3.280 37.270 5.880 37.470 ;
        RECT 6.480 37.370 6.680 38.870 ;
        RECT 7.280 37.370 7.480 38.870 ;
        RECT 8.080 37.370 8.280 38.870 ;
        RECT 8.880 37.370 9.080 38.870 ;
        RECT 9.680 37.370 9.880 38.870 ;
        RECT 10.480 37.370 10.680 38.870 ;
        RECT 11.280 37.370 11.480 38.870 ;
        RECT 12.080 37.370 12.280 38.870 ;
        RECT 12.880 37.370 13.080 38.870 ;
        RECT 13.680 37.370 13.880 38.870 ;
        RECT 14.480 37.370 14.680 38.870 ;
        RECT 15.280 37.370 15.480 38.870 ;
        RECT 16.080 37.370 16.280 38.870 ;
        RECT 16.880 37.370 17.080 38.870 ;
        RECT 17.680 37.370 17.880 38.870 ;
        RECT 18.480 38.270 18.830 38.870 ;
        RECT 18.480 38.070 21.080 38.270 ;
        RECT 18.480 37.470 18.830 38.070 ;
        RECT 18.480 37.270 21.030 37.470 ;
        RECT 3.280 36.370 5.880 36.570 ;
        RECT 5.530 35.770 5.880 36.370 ;
        RECT 3.280 35.570 5.880 35.770 ;
        RECT 5.530 34.970 5.880 35.570 ;
        RECT 6.480 34.970 6.680 36.470 ;
        RECT 7.280 34.970 7.480 36.470 ;
        RECT 8.080 34.970 8.280 36.470 ;
        RECT 8.880 34.970 9.080 36.470 ;
        RECT 9.680 34.970 9.880 36.470 ;
        RECT 10.480 34.970 10.680 36.470 ;
        RECT 11.280 34.970 11.480 36.470 ;
        RECT 12.080 34.970 12.280 36.470 ;
        RECT 12.880 34.970 13.080 36.470 ;
        RECT 13.680 34.970 13.880 36.470 ;
        RECT 14.480 34.970 14.680 36.470 ;
        RECT 15.280 34.970 15.480 36.470 ;
        RECT 16.080 34.970 16.280 36.470 ;
        RECT 16.880 34.970 17.080 36.470 ;
        RECT 17.680 34.970 17.880 36.470 ;
        RECT 18.480 36.370 21.030 36.570 ;
        RECT 18.480 35.770 18.830 36.370 ;
        RECT 18.480 35.570 21.080 35.770 ;
        RECT 18.480 34.970 18.830 35.570 ;
        RECT 2.930 34.370 21.430 34.970 ;
        RECT 4.580 33.770 6.880 33.820 ;
        RECT 17.480 33.770 19.780 33.820 ;
        RECT 22.230 33.770 22.630 40.070 ;
        RECT 1.730 33.370 22.630 33.770 ;
        RECT 4.580 32.970 6.880 33.370 ;
        RECT 17.480 32.970 19.780 33.370 ;
        RECT 16.490 28.390 16.660 29.180 ;
        RECT 17.450 28.390 17.620 29.180 ;
        RECT 19.170 28.720 19.340 29.420 ;
        RECT 21.650 28.720 21.820 29.420 ;
        RECT 23.550 28.720 24.540 40.970 ;
        RECT 19.040 28.460 24.540 28.720 ;
        RECT 15.950 28.300 17.730 28.390 ;
        RECT 15.270 27.960 17.730 28.300 ;
        RECT 1.730 25.040 2.190 25.210 ;
        RECT 2.900 25.040 3.360 25.210 ;
        RECT 1.750 24.510 2.170 25.040 ;
        RECT 2.920 24.510 3.340 25.040 ;
        RECT 4.530 24.290 4.700 25.550 ;
        RECT 5.490 24.290 5.660 25.540 ;
        RECT 6.450 24.290 6.620 25.540 ;
        RECT 7.410 24.290 7.580 25.540 ;
        RECT 11.320 24.430 11.490 27.010 ;
        RECT 12.280 24.430 12.450 27.010 ;
        RECT 13.240 24.430 13.410 27.010 ;
        RECT 15.270 26.330 15.610 27.960 ;
        RECT 15.950 27.870 17.730 27.960 ;
        RECT 16.490 27.080 16.660 27.870 ;
        RECT 17.450 27.080 17.620 27.870 ;
        RECT 19.850 27.570 20.280 28.460 ;
        RECT 19.970 26.860 20.140 27.570 ;
        RECT 14.920 25.990 15.610 26.330 ;
        RECT 4.530 24.220 7.580 24.290 ;
        RECT 11.290 24.240 13.550 24.430 ;
        RECT 14.920 24.240 15.320 25.990 ;
        RECT 3.960 24.010 8.050 24.220 ;
        RECT 4.580 22.520 6.880 24.010 ;
        RECT 14.920 23.890 19.780 24.240 ;
        RECT 17.480 22.520 19.780 23.890 ;
        RECT 1.730 22.120 22.630 22.520 ;
        RECT 1.730 15.820 2.130 22.120 ;
        RECT 4.580 22.070 6.880 22.120 ;
        RECT 17.480 22.070 19.780 22.120 ;
        RECT 2.930 20.920 21.430 21.520 ;
        RECT 5.530 20.320 5.880 20.920 ;
        RECT 3.280 20.120 5.880 20.320 ;
        RECT 5.530 19.520 5.880 20.120 ;
        RECT 3.280 19.320 5.880 19.520 ;
        RECT 6.480 19.420 6.680 20.920 ;
        RECT 7.280 19.420 7.480 20.920 ;
        RECT 8.080 19.420 8.280 20.920 ;
        RECT 8.880 19.420 9.080 20.920 ;
        RECT 9.680 19.420 9.880 20.920 ;
        RECT 10.480 19.420 10.680 20.920 ;
        RECT 11.280 19.420 11.480 20.920 ;
        RECT 12.080 19.420 12.280 20.920 ;
        RECT 12.880 19.420 13.080 20.920 ;
        RECT 13.680 19.420 13.880 20.920 ;
        RECT 14.480 19.420 14.680 20.920 ;
        RECT 15.280 19.420 15.480 20.920 ;
        RECT 16.080 19.420 16.280 20.920 ;
        RECT 16.880 19.420 17.080 20.920 ;
        RECT 17.680 19.420 17.880 20.920 ;
        RECT 18.480 20.320 18.830 20.920 ;
        RECT 18.480 20.120 21.080 20.320 ;
        RECT 18.480 19.520 18.830 20.120 ;
        RECT 18.480 19.320 21.030 19.520 ;
        RECT 3.280 18.420 5.880 18.620 ;
        RECT 5.530 17.820 5.880 18.420 ;
        RECT 3.280 17.620 5.880 17.820 ;
        RECT 5.530 17.020 5.880 17.620 ;
        RECT 6.480 17.020 6.680 18.520 ;
        RECT 7.280 17.020 7.480 18.520 ;
        RECT 8.080 17.020 8.280 18.520 ;
        RECT 8.880 17.020 9.080 18.520 ;
        RECT 9.680 17.020 9.880 18.520 ;
        RECT 10.480 17.020 10.680 18.520 ;
        RECT 11.280 17.020 11.480 18.520 ;
        RECT 12.080 17.020 12.280 18.520 ;
        RECT 12.880 17.020 13.080 18.520 ;
        RECT 13.680 17.020 13.880 18.520 ;
        RECT 14.480 17.020 14.680 18.520 ;
        RECT 15.280 17.020 15.480 18.520 ;
        RECT 16.080 17.020 16.280 18.520 ;
        RECT 16.880 17.020 17.080 18.520 ;
        RECT 17.680 17.020 17.880 18.520 ;
        RECT 18.480 18.420 21.030 18.620 ;
        RECT 18.480 17.820 18.830 18.420 ;
        RECT 18.480 17.620 21.080 17.820 ;
        RECT 18.480 17.020 18.830 17.620 ;
        RECT 2.930 16.420 21.430 17.020 ;
        RECT 4.580 15.820 6.880 15.870 ;
        RECT 17.480 15.820 19.780 15.870 ;
        RECT 22.230 15.820 22.630 22.120 ;
        RECT 1.730 15.420 22.630 15.820 ;
        RECT 4.580 14.970 6.880 15.420 ;
        RECT 17.480 14.970 19.780 15.420 ;
        RECT 23.550 14.970 24.540 28.460 ;
        RECT 0.150 13.980 24.540 14.970 ;
      LAYER mcon ;
        RECT 0.330 38.720 0.980 40.720 ;
        RECT 0.250 35.820 0.930 38.020 ;
        RECT 0.250 33.070 1.030 35.220 ;
        RECT 3.030 38.970 3.630 39.470 ;
        RECT 3.830 38.970 4.430 39.470 ;
        RECT 4.630 38.970 5.230 39.470 ;
        RECT 5.430 38.970 6.030 39.470 ;
        RECT 18.330 38.970 18.930 39.470 ;
        RECT 19.130 38.970 19.730 39.470 ;
        RECT 19.930 38.970 20.530 39.470 ;
        RECT 20.730 38.970 21.330 39.470 ;
        RECT 3.030 34.370 3.630 34.870 ;
        RECT 3.830 34.370 4.430 34.870 ;
        RECT 4.630 34.370 5.230 34.870 ;
        RECT 5.430 34.370 6.030 34.870 ;
        RECT 18.330 34.370 18.930 34.870 ;
        RECT 19.130 34.370 19.730 34.870 ;
        RECT 19.930 34.370 20.530 34.870 ;
        RECT 20.730 34.370 21.330 34.870 ;
        RECT 0.230 24.590 0.400 24.760 ;
        RECT 0.590 24.590 0.760 24.760 ;
        RECT 0.950 24.590 1.120 24.760 ;
        RECT 1.870 24.540 2.050 24.710 ;
        RECT 3.040 24.540 3.220 24.710 ;
        RECT 0.230 24.230 0.400 24.400 ;
        RECT 0.590 24.230 0.760 24.400 ;
        RECT 0.950 24.230 1.120 24.400 ;
        RECT 11.410 24.250 11.590 24.430 ;
        RECT 11.870 24.250 12.050 24.430 ;
        RECT 12.330 24.250 12.510 24.430 ;
        RECT 12.790 24.250 12.970 24.430 ;
        RECT 13.250 24.250 13.430 24.430 ;
        RECT 23.620 24.590 23.790 24.760 ;
        RECT 23.980 24.590 24.150 24.760 ;
        RECT 24.340 24.590 24.510 24.760 ;
        RECT 0.230 23.870 0.400 24.040 ;
        RECT 0.590 23.870 0.760 24.040 ;
        RECT 0.950 23.870 1.120 24.040 ;
        RECT 4.080 24.030 4.260 24.210 ;
        RECT 4.670 24.030 4.850 24.210 ;
        RECT 5.260 24.030 5.440 24.210 ;
        RECT 5.850 24.030 6.030 24.210 ;
        RECT 6.440 24.030 6.620 24.210 ;
        RECT 7.030 24.030 7.210 24.210 ;
        RECT 7.620 24.030 7.800 24.210 ;
        RECT 0.230 23.510 0.400 23.680 ;
        RECT 0.590 23.510 0.760 23.680 ;
        RECT 0.950 23.510 1.120 23.680 ;
        RECT 0.220 23.150 0.390 23.320 ;
        RECT 0.580 23.150 0.750 23.320 ;
        RECT 0.940 23.150 1.110 23.320 ;
        RECT 0.240 20.670 1.030 22.820 ;
        RECT 14.960 23.960 15.140 24.140 ;
        RECT 15.330 23.970 15.510 24.150 ;
        RECT 15.730 23.970 15.910 24.150 ;
        RECT 16.130 23.970 16.310 24.150 ;
        RECT 16.530 23.970 16.710 24.150 ;
        RECT 23.620 24.230 23.790 24.400 ;
        RECT 23.980 24.230 24.150 24.400 ;
        RECT 24.340 24.230 24.510 24.400 ;
        RECT 23.620 23.870 23.790 24.040 ;
        RECT 23.980 23.870 24.150 24.040 ;
        RECT 24.340 23.870 24.510 24.040 ;
        RECT 23.620 23.510 23.790 23.680 ;
        RECT 23.980 23.510 24.150 23.680 ;
        RECT 24.340 23.510 24.510 23.680 ;
        RECT 23.620 23.150 23.790 23.320 ;
        RECT 23.980 23.150 24.150 23.320 ;
        RECT 24.340 23.150 24.510 23.320 ;
        RECT 0.280 17.870 0.930 20.070 ;
        RECT 0.280 15.170 1.080 17.220 ;
        RECT 3.030 21.020 3.630 21.520 ;
        RECT 3.830 21.020 4.430 21.520 ;
        RECT 4.630 21.020 5.230 21.520 ;
        RECT 5.430 21.020 6.030 21.520 ;
        RECT 18.330 21.020 18.930 21.520 ;
        RECT 19.130 21.020 19.730 21.520 ;
        RECT 19.930 21.020 20.530 21.520 ;
        RECT 20.730 21.020 21.330 21.520 ;
        RECT 3.030 16.420 3.630 16.920 ;
        RECT 3.830 16.420 4.430 16.920 ;
        RECT 4.630 16.420 5.230 16.920 ;
        RECT 5.430 16.420 6.030 16.920 ;
        RECT 18.330 16.420 18.930 16.920 ;
        RECT 19.130 16.420 19.730 16.920 ;
        RECT 19.930 16.420 20.530 16.920 ;
        RECT 20.730 16.420 21.330 16.920 ;
      LAYER met1 ;
        RECT 0.150 39.670 4.530 40.870 ;
        RECT 19.830 39.670 23.030 40.870 ;
        RECT 0.150 39.520 3.630 39.670 ;
        RECT 20.730 39.520 23.030 39.670 ;
        RECT 0.150 39.370 11.730 39.520 ;
        RECT 12.630 39.370 23.030 39.520 ;
        RECT 0.150 38.920 6.130 39.370 ;
        RECT 18.230 38.920 23.030 39.370 ;
        RECT 0.150 38.520 2.530 38.920 ;
        RECT 2.980 38.870 11.730 38.920 ;
        RECT 0.150 35.720 1.030 38.120 ;
        RECT 1.330 38.020 2.530 38.520 ;
        RECT 3.130 37.520 3.280 38.870 ;
        RECT 3.730 37.520 3.880 38.870 ;
        RECT 4.330 37.520 4.480 38.870 ;
        RECT 4.930 37.520 5.080 38.870 ;
        RECT 5.530 38.770 11.730 38.870 ;
        RECT 12.630 38.870 21.380 38.920 ;
        RECT 12.630 38.770 18.830 38.870 ;
        RECT 5.530 38.320 6.130 38.770 ;
        RECT 18.230 38.320 18.830 38.770 ;
        RECT 5.530 38.170 11.730 38.320 ;
        RECT 12.630 38.170 18.830 38.320 ;
        RECT 5.530 37.720 6.130 38.170 ;
        RECT 18.230 37.720 18.830 38.170 ;
        RECT 5.530 37.570 11.730 37.720 ;
        RECT 12.630 37.570 18.830 37.720 ;
        RECT 5.530 37.370 6.130 37.570 ;
        RECT 18.230 37.370 18.830 37.570 ;
        RECT 19.280 37.520 19.430 38.870 ;
        RECT 19.880 37.520 20.030 38.870 ;
        RECT 20.480 37.520 20.630 38.870 ;
        RECT 21.080 37.520 21.230 38.870 ;
        RECT 21.830 38.020 23.030 38.920 ;
        RECT 1.330 35.320 2.530 35.820 ;
        RECT 0.150 34.920 2.530 35.320 ;
        RECT 3.130 34.970 3.280 36.270 ;
        RECT 3.730 34.970 3.880 36.270 ;
        RECT 4.330 34.970 4.480 36.270 ;
        RECT 4.930 34.970 5.080 36.270 ;
        RECT 5.530 36.120 11.730 36.270 ;
        RECT 12.630 36.120 18.830 36.270 ;
        RECT 5.530 35.670 6.130 36.120 ;
        RECT 18.230 35.670 18.830 36.120 ;
        RECT 5.530 35.520 11.730 35.670 ;
        RECT 12.630 35.520 18.830 35.670 ;
        RECT 5.530 35.070 6.130 35.520 ;
        RECT 18.230 35.070 18.830 35.520 ;
        RECT 5.530 34.970 11.730 35.070 ;
        RECT 2.980 34.920 11.730 34.970 ;
        RECT 12.630 34.970 18.830 35.070 ;
        RECT 19.280 34.970 19.430 36.270 ;
        RECT 19.880 34.970 20.030 36.270 ;
        RECT 20.480 34.970 20.630 36.270 ;
        RECT 21.080 34.970 21.230 36.270 ;
        RECT 12.630 34.920 21.380 34.970 ;
        RECT 21.830 34.920 23.030 35.820 ;
        RECT 0.150 34.470 6.130 34.920 ;
        RECT 18.230 34.470 23.030 34.920 ;
        RECT 0.150 34.320 11.730 34.470 ;
        RECT 12.630 34.320 23.030 34.470 ;
        RECT 0.150 34.170 3.630 34.320 ;
        RECT 20.730 34.170 23.030 34.320 ;
        RECT 0.150 32.970 4.530 34.170 ;
        RECT 19.830 32.970 23.030 34.170 ;
        RECT 0.150 24.760 1.150 24.860 ;
        RECT 0.150 24.240 3.420 24.760 ;
        RECT 11.290 24.240 13.550 24.460 ;
        RECT 23.550 24.240 24.540 24.860 ;
        RECT -2.790 23.080 25.780 24.240 ;
        RECT 0.140 21.720 4.530 22.920 ;
        RECT 19.830 21.720 23.030 22.920 ;
        RECT 0.140 21.570 3.630 21.720 ;
        RECT 20.730 21.570 23.030 21.720 ;
        RECT 0.140 21.420 11.730 21.570 ;
        RECT 12.630 21.420 23.030 21.570 ;
        RECT 0.140 20.970 6.130 21.420 ;
        RECT 18.230 20.970 23.030 21.420 ;
        RECT 0.140 20.570 2.530 20.970 ;
        RECT 2.980 20.920 11.730 20.970 ;
        RECT 0.150 17.770 1.030 20.170 ;
        RECT 1.330 20.070 2.530 20.570 ;
        RECT 3.130 19.570 3.280 20.920 ;
        RECT 3.730 19.570 3.880 20.920 ;
        RECT 4.330 19.570 4.480 20.920 ;
        RECT 4.930 19.570 5.080 20.920 ;
        RECT 5.530 20.820 11.730 20.920 ;
        RECT 12.630 20.920 21.380 20.970 ;
        RECT 12.630 20.820 18.830 20.920 ;
        RECT 5.530 20.370 6.130 20.820 ;
        RECT 18.230 20.370 18.830 20.820 ;
        RECT 5.530 20.220 11.730 20.370 ;
        RECT 12.630 20.220 18.830 20.370 ;
        RECT 5.530 19.770 6.130 20.220 ;
        RECT 18.230 19.770 18.830 20.220 ;
        RECT 5.530 19.620 11.730 19.770 ;
        RECT 12.630 19.620 18.830 19.770 ;
        RECT 5.530 19.420 6.130 19.620 ;
        RECT 18.230 19.420 18.830 19.620 ;
        RECT 19.280 19.570 19.430 20.920 ;
        RECT 19.880 19.570 20.030 20.920 ;
        RECT 20.480 19.570 20.630 20.920 ;
        RECT 21.080 19.570 21.230 20.920 ;
        RECT 21.830 20.070 23.030 20.970 ;
        RECT 1.330 17.370 2.530 17.870 ;
        RECT 0.150 16.970 2.530 17.370 ;
        RECT 3.130 17.020 3.280 18.320 ;
        RECT 3.730 17.020 3.880 18.320 ;
        RECT 4.330 17.020 4.480 18.320 ;
        RECT 4.930 17.020 5.080 18.320 ;
        RECT 5.530 18.170 11.730 18.320 ;
        RECT 12.630 18.170 18.830 18.320 ;
        RECT 5.530 17.720 6.130 18.170 ;
        RECT 18.230 17.720 18.830 18.170 ;
        RECT 5.530 17.570 11.730 17.720 ;
        RECT 12.630 17.570 18.830 17.720 ;
        RECT 5.530 17.120 6.130 17.570 ;
        RECT 18.230 17.120 18.830 17.570 ;
        RECT 5.530 17.020 11.730 17.120 ;
        RECT 2.980 16.970 11.730 17.020 ;
        RECT 12.630 17.020 18.830 17.120 ;
        RECT 19.280 17.020 19.430 18.320 ;
        RECT 19.880 17.020 20.030 18.320 ;
        RECT 20.480 17.020 20.630 18.320 ;
        RECT 21.080 17.020 21.230 18.320 ;
        RECT 12.630 16.970 21.380 17.020 ;
        RECT 21.830 16.970 23.030 17.870 ;
        RECT 0.150 16.520 6.130 16.970 ;
        RECT 18.230 16.520 23.030 16.970 ;
        RECT 0.150 16.370 11.730 16.520 ;
        RECT 12.630 16.370 23.030 16.520 ;
        RECT 0.150 16.220 3.630 16.370 ;
        RECT 20.730 16.220 23.030 16.370 ;
        RECT 0.150 15.020 4.530 16.220 ;
        RECT 19.830 15.020 23.030 16.220 ;
      LAYER via ;
        RECT 0.330 38.720 0.980 40.720 ;
        RECT 1.430 39.770 2.430 40.770 ;
        RECT 3.430 39.770 4.430 40.770 ;
        RECT 19.930 39.770 20.930 40.770 ;
        RECT 21.930 39.770 22.930 40.770 ;
        RECT 1.430 38.170 2.430 39.170 ;
        RECT 0.250 35.820 0.930 38.020 ;
        RECT 21.930 38.170 22.930 39.170 ;
        RECT 1.430 34.670 2.430 35.670 ;
        RECT 21.930 34.670 22.930 35.670 ;
        RECT 1.430 33.070 2.430 34.070 ;
        RECT 3.430 33.070 4.430 34.070 ;
        RECT 19.930 33.070 20.930 34.070 ;
        RECT 21.930 33.070 22.930 34.070 ;
        RECT -1.070 23.170 -0.270 24.120 ;
        RECT 1.430 23.270 4.210 24.100 ;
        RECT 24.880 23.170 25.680 24.120 ;
        RECT 1.430 21.820 2.430 22.820 ;
        RECT 3.430 21.820 4.430 22.820 ;
        RECT 19.930 21.820 20.930 22.820 ;
        RECT 21.930 21.820 22.930 22.820 ;
        RECT 1.430 20.220 2.430 21.220 ;
        RECT 0.280 17.870 0.930 20.070 ;
        RECT 21.930 20.220 22.930 21.220 ;
        RECT 0.280 15.170 1.080 17.220 ;
        RECT 1.430 16.720 2.430 17.720 ;
        RECT 21.930 16.720 22.930 17.720 ;
        RECT 1.430 15.120 2.430 16.120 ;
        RECT 3.430 15.120 4.430 16.120 ;
        RECT 19.930 15.120 20.930 16.120 ;
        RECT 21.930 15.120 22.930 16.120 ;
      LAYER met2 ;
        RECT 0.150 39.670 4.530 40.870 ;
        RECT 19.830 39.670 23.030 40.870 ;
        RECT 0.150 38.720 3.280 39.670 ;
        RECT 21.080 38.720 23.030 39.670 ;
        RECT 0.150 38.570 5.280 38.720 ;
        RECT 0.150 38.520 3.280 38.570 ;
        RECT 1.330 38.120 3.280 38.520 ;
        RECT 0.150 35.720 1.030 38.120 ;
        RECT 1.330 38.020 5.280 38.120 ;
        RECT 2.730 37.970 5.280 38.020 ;
        RECT 2.730 37.370 3.280 37.970 ;
        RECT 2.730 37.070 5.280 37.370 ;
        RECT 5.880 37.070 6.030 38.720 ;
        RECT 6.480 37.070 6.630 38.720 ;
        RECT 7.080 37.070 7.230 38.720 ;
        RECT 7.680 37.070 7.830 38.720 ;
        RECT 8.280 37.070 8.430 38.720 ;
        RECT 8.880 37.070 9.030 38.720 ;
        RECT 9.480 37.070 9.630 38.720 ;
        RECT 10.080 37.070 10.230 38.720 ;
        RECT 10.680 37.070 10.830 38.720 ;
        RECT 11.280 37.070 11.430 38.720 ;
        RECT 11.880 37.070 12.480 38.720 ;
        RECT 12.930 37.070 13.080 38.720 ;
        RECT 13.530 37.070 13.680 38.720 ;
        RECT 14.130 37.070 14.280 38.720 ;
        RECT 14.730 37.070 14.880 38.720 ;
        RECT 15.330 37.070 15.480 38.720 ;
        RECT 15.930 37.070 16.080 38.720 ;
        RECT 16.530 37.070 16.680 38.720 ;
        RECT 17.130 37.070 17.280 38.720 ;
        RECT 17.730 37.070 17.880 38.720 ;
        RECT 18.330 37.070 18.480 38.720 ;
        RECT 19.080 38.570 23.030 38.720 ;
        RECT 21.080 38.120 23.030 38.570 ;
        RECT 19.080 38.020 23.030 38.120 ;
        RECT 19.080 37.970 21.630 38.020 ;
        RECT 21.080 37.370 21.630 37.970 ;
        RECT 19.080 37.070 21.630 37.370 ;
        RECT 2.730 36.770 21.630 37.070 ;
        RECT 2.730 36.320 5.280 36.770 ;
        RECT 2.730 35.870 3.280 36.320 ;
        RECT 2.730 35.820 5.280 35.870 ;
        RECT 1.330 35.720 5.280 35.820 ;
        RECT 1.330 35.270 3.280 35.720 ;
        RECT 1.330 35.120 5.280 35.270 ;
        RECT 5.880 35.120 6.030 36.770 ;
        RECT 6.480 35.120 6.630 36.770 ;
        RECT 7.080 35.120 7.230 36.770 ;
        RECT 7.680 35.120 7.830 36.770 ;
        RECT 8.280 35.120 8.430 36.770 ;
        RECT 8.880 35.120 9.030 36.770 ;
        RECT 9.480 35.120 9.630 36.770 ;
        RECT 10.080 35.120 10.230 36.770 ;
        RECT 10.680 35.120 10.830 36.770 ;
        RECT 11.280 35.120 11.430 36.770 ;
        RECT 11.880 35.120 12.480 36.770 ;
        RECT 12.930 35.120 13.080 36.770 ;
        RECT 13.530 35.120 13.680 36.770 ;
        RECT 14.130 35.120 14.280 36.770 ;
        RECT 14.730 35.120 14.880 36.770 ;
        RECT 15.330 35.120 15.480 36.770 ;
        RECT 15.930 35.120 16.080 36.770 ;
        RECT 16.530 35.120 16.680 36.770 ;
        RECT 17.130 35.120 17.280 36.770 ;
        RECT 17.730 35.120 17.880 36.770 ;
        RECT 18.330 35.120 18.480 36.770 ;
        RECT 19.080 36.320 21.630 36.770 ;
        RECT 21.080 35.870 21.630 36.320 ;
        RECT 19.080 35.820 21.630 35.870 ;
        RECT 19.080 35.720 23.030 35.820 ;
        RECT 21.080 35.270 23.030 35.720 ;
        RECT 19.080 35.120 23.030 35.270 ;
        RECT 1.330 34.170 3.280 35.120 ;
        RECT 21.080 34.170 23.030 35.120 ;
        RECT 1.330 32.970 4.530 34.170 ;
        RECT 19.830 32.970 23.030 34.170 ;
        RECT -1.180 23.080 -0.180 24.240 ;
        RECT 1.290 23.240 4.440 24.240 ;
        RECT 1.330 22.920 4.480 23.240 ;
        RECT 24.780 23.080 25.780 24.240 ;
        RECT 1.330 21.720 4.530 22.920 ;
        RECT 19.830 21.720 23.030 22.920 ;
        RECT 1.330 20.770 3.280 21.720 ;
        RECT 21.080 20.770 23.030 21.720 ;
        RECT 1.330 20.620 5.280 20.770 ;
        RECT 1.330 20.170 3.280 20.620 ;
        RECT 0.150 17.770 1.030 20.170 ;
        RECT 1.330 20.070 5.280 20.170 ;
        RECT 2.730 20.020 5.280 20.070 ;
        RECT 2.730 19.420 3.280 20.020 ;
        RECT 2.730 19.120 5.280 19.420 ;
        RECT 5.880 19.120 6.030 20.770 ;
        RECT 6.480 19.120 6.630 20.770 ;
        RECT 7.080 19.120 7.230 20.770 ;
        RECT 7.680 19.120 7.830 20.770 ;
        RECT 8.280 19.120 8.430 20.770 ;
        RECT 8.880 19.120 9.030 20.770 ;
        RECT 9.480 19.120 9.630 20.770 ;
        RECT 10.080 19.120 10.230 20.770 ;
        RECT 10.680 19.120 10.830 20.770 ;
        RECT 11.280 19.120 11.430 20.770 ;
        RECT 11.880 19.120 12.480 20.770 ;
        RECT 12.930 19.120 13.080 20.770 ;
        RECT 13.530 19.120 13.680 20.770 ;
        RECT 14.130 19.120 14.280 20.770 ;
        RECT 14.730 19.120 14.880 20.770 ;
        RECT 15.330 19.120 15.480 20.770 ;
        RECT 15.930 19.120 16.080 20.770 ;
        RECT 16.530 19.120 16.680 20.770 ;
        RECT 17.130 19.120 17.280 20.770 ;
        RECT 17.730 19.120 17.880 20.770 ;
        RECT 18.330 19.120 18.480 20.770 ;
        RECT 19.080 20.620 23.030 20.770 ;
        RECT 21.080 20.170 23.030 20.620 ;
        RECT 19.080 20.070 23.030 20.170 ;
        RECT 19.080 20.020 21.630 20.070 ;
        RECT 21.080 19.420 21.630 20.020 ;
        RECT 19.080 19.120 21.630 19.420 ;
        RECT 2.730 18.820 21.630 19.120 ;
        RECT 2.730 18.370 5.280 18.820 ;
        RECT 2.730 17.920 3.280 18.370 ;
        RECT 2.730 17.870 5.280 17.920 ;
        RECT 1.330 17.770 5.280 17.870 ;
        RECT 1.330 17.370 3.280 17.770 ;
        RECT 0.150 17.320 3.280 17.370 ;
        RECT 0.150 17.170 5.280 17.320 ;
        RECT 5.880 17.170 6.030 18.820 ;
        RECT 6.480 17.170 6.630 18.820 ;
        RECT 7.080 17.170 7.230 18.820 ;
        RECT 7.680 17.170 7.830 18.820 ;
        RECT 8.280 17.170 8.430 18.820 ;
        RECT 8.880 17.170 9.030 18.820 ;
        RECT 9.480 17.170 9.630 18.820 ;
        RECT 10.080 17.170 10.230 18.820 ;
        RECT 10.680 17.170 10.830 18.820 ;
        RECT 11.280 17.170 11.430 18.820 ;
        RECT 11.880 17.170 12.480 18.820 ;
        RECT 12.930 17.170 13.080 18.820 ;
        RECT 13.530 17.170 13.680 18.820 ;
        RECT 14.130 17.170 14.280 18.820 ;
        RECT 14.730 17.170 14.880 18.820 ;
        RECT 15.330 17.170 15.480 18.820 ;
        RECT 15.930 17.170 16.080 18.820 ;
        RECT 16.530 17.170 16.680 18.820 ;
        RECT 17.130 17.170 17.280 18.820 ;
        RECT 17.730 17.170 17.880 18.820 ;
        RECT 18.330 17.170 18.480 18.820 ;
        RECT 19.080 18.370 21.630 18.820 ;
        RECT 21.080 17.920 21.630 18.370 ;
        RECT 19.080 17.870 21.630 17.920 ;
        RECT 19.080 17.770 23.030 17.870 ;
        RECT 21.080 17.320 23.030 17.770 ;
        RECT 19.080 17.170 23.030 17.320 ;
        RECT 0.150 16.220 3.280 17.170 ;
        RECT 21.080 16.220 23.030 17.170 ;
        RECT 0.150 15.020 4.530 16.220 ;
        RECT 19.830 15.020 23.030 16.220 ;
      LAYER via2 ;
        RECT 0.330 38.720 0.980 40.720 ;
        RECT 0.250 35.820 0.930 38.020 ;
        RECT -1.070 23.170 -0.270 24.120 ;
        RECT 1.430 23.270 4.210 24.100 ;
        RECT 24.880 23.170 25.680 24.120 ;
        RECT 0.280 17.870 0.930 20.070 ;
        RECT 0.280 15.170 1.080 17.220 ;
      LAYER met3 ;
        RECT 0.150 39.620 4.530 40.870 ;
        RECT 6.930 40.020 17.430 40.870 ;
        RECT 19.830 39.620 23.030 40.870 ;
        RECT 0.150 38.520 23.030 39.620 ;
        RECT 1.330 38.470 23.030 38.520 ;
        RECT 0.150 35.720 1.030 38.120 ;
        RECT 1.330 35.720 2.180 38.120 ;
        RECT 2.580 35.370 21.780 38.470 ;
        RECT 22.180 35.720 23.030 38.120 ;
        RECT 1.330 34.220 23.030 35.370 ;
        RECT 1.330 32.970 4.530 34.220 ;
        RECT 6.930 32.970 17.430 33.820 ;
        RECT 19.830 32.970 23.030 34.220 ;
        RECT -1.180 23.080 -0.180 24.240 ;
        RECT 1.290 23.240 4.440 24.240 ;
        RECT 24.780 23.080 25.780 24.240 ;
        RECT 1.330 21.670 4.530 22.920 ;
        RECT 6.930 22.070 17.430 22.920 ;
        RECT 19.830 21.670 23.030 22.920 ;
        RECT 1.330 20.520 23.030 21.670 ;
        RECT 0.150 17.770 1.030 20.170 ;
        RECT 1.330 17.770 2.180 20.170 ;
        RECT 2.580 17.420 21.780 20.520 ;
        RECT 22.180 17.770 23.030 20.170 ;
        RECT 1.330 17.370 23.030 17.420 ;
        RECT 0.150 16.270 23.030 17.370 ;
        RECT 0.150 15.020 4.530 16.270 ;
        RECT 6.930 15.020 17.430 15.870 ;
        RECT 19.830 15.020 23.030 16.270 ;
      LAYER via3 ;
        RECT 0.330 38.720 0.980 40.720 ;
        RECT 1.430 39.920 2.280 40.770 ;
        RECT 3.530 39.920 4.380 40.770 ;
        RECT 7.030 40.120 7.680 40.770 ;
        RECT 7.830 40.120 8.480 40.770 ;
        RECT 15.880 40.120 16.530 40.770 ;
        RECT 16.680 40.120 17.330 40.770 ;
        RECT 19.980 39.920 20.830 40.770 ;
        RECT 22.080 39.920 22.930 40.770 ;
        RECT 1.430 38.620 2.280 39.470 ;
        RECT 22.080 38.620 22.930 39.470 ;
        RECT 0.250 35.820 0.930 38.020 ;
        RECT 1.430 37.020 2.080 38.020 ;
        RECT 1.430 35.820 2.080 36.820 ;
        RECT 22.280 37.020 22.930 38.020 ;
        RECT 22.280 35.820 22.930 36.820 ;
        RECT 1.430 34.370 2.280 35.220 ;
        RECT 22.080 34.370 22.930 35.220 ;
        RECT 1.430 33.070 2.280 33.920 ;
        RECT 3.530 33.070 4.380 33.920 ;
        RECT 7.030 33.070 7.680 33.720 ;
        RECT 7.830 33.070 8.480 33.720 ;
        RECT 15.880 33.070 16.530 33.720 ;
        RECT 16.680 33.070 17.330 33.720 ;
        RECT 19.980 33.070 20.830 33.920 ;
        RECT 22.080 33.070 22.930 33.920 ;
        RECT -1.070 23.170 -0.270 24.120 ;
        RECT 24.880 23.170 25.680 24.120 ;
        RECT 1.430 21.970 2.280 22.820 ;
        RECT 3.530 21.970 4.380 22.820 ;
        RECT 7.030 22.170 7.680 22.820 ;
        RECT 7.830 22.170 8.480 22.820 ;
        RECT 15.880 22.170 16.530 22.820 ;
        RECT 16.680 22.170 17.330 22.820 ;
        RECT 19.980 21.970 20.830 22.820 ;
        RECT 22.080 21.970 22.930 22.820 ;
        RECT 1.430 20.670 2.280 21.520 ;
        RECT 22.080 20.670 22.930 21.520 ;
        RECT 0.280 17.870 0.930 20.070 ;
        RECT 1.430 19.070 2.080 20.070 ;
        RECT 1.430 17.870 2.080 18.870 ;
        RECT 22.280 19.070 22.930 20.070 ;
        RECT 22.280 17.870 22.930 18.870 ;
        RECT 0.280 15.170 1.080 17.220 ;
        RECT 1.430 16.420 2.280 17.270 ;
        RECT 22.080 16.420 22.930 17.270 ;
        RECT 1.430 15.120 2.280 15.970 ;
        RECT 3.530 15.120 4.380 15.970 ;
        RECT 7.030 15.120 7.680 15.770 ;
        RECT 7.830 15.120 8.480 15.770 ;
        RECT 15.880 15.120 16.530 15.770 ;
        RECT 16.680 15.120 17.330 15.770 ;
        RECT 19.980 15.120 20.830 15.970 ;
        RECT 22.080 15.120 22.930 15.970 ;
      LAYER met4 ;
        RECT -1.180 13.980 -0.180 41.960 ;
        RECT 0.150 39.820 4.480 40.870 ;
        RECT 0.150 38.520 2.380 39.820 ;
        RECT 6.930 39.420 17.430 40.870 ;
        RECT 19.880 39.820 23.030 40.870 ;
        RECT 2.780 38.120 21.580 39.420 ;
        RECT 21.980 38.520 23.030 39.820 ;
        RECT 0.150 35.720 23.030 38.120 ;
        RECT 1.330 34.020 2.380 35.320 ;
        RECT 2.780 34.420 21.580 35.720 ;
        RECT 1.330 32.970 4.480 34.020 ;
        RECT 6.930 32.970 17.430 34.420 ;
        RECT 21.980 34.020 23.030 35.320 ;
        RECT 19.880 32.970 23.030 34.020 ;
        RECT 1.330 21.870 4.480 22.920 ;
        RECT 1.330 20.570 2.380 21.870 ;
        RECT 6.930 21.470 17.430 22.920 ;
        RECT 19.880 21.870 23.030 22.920 ;
        RECT 2.780 20.170 21.580 21.470 ;
        RECT 21.980 20.570 23.030 21.870 ;
        RECT 0.150 17.770 23.030 20.170 ;
        RECT 0.150 16.070 2.380 17.370 ;
        RECT 2.780 16.470 21.580 17.770 ;
        RECT 0.150 15.020 4.480 16.070 ;
        RECT 6.930 15.020 17.430 16.470 ;
        RECT 21.980 16.070 23.030 17.370 ;
        RECT 19.880 15.020 23.030 16.070 ;
        RECT 24.780 13.980 25.780 41.960 ;
    END
  END VSS
  PIN VDD
    ANTENNADIFFAREA 8.718300 ;
    PORT
      LAYER nwell ;
        RECT 15.590 32.000 23.500 32.020 ;
        RECT 3.800 29.980 23.500 32.000 ;
        RECT 3.800 29.890 15.260 29.980 ;
        RECT 6.430 29.880 7.640 29.890 ;
        RECT 9.470 28.140 15.260 29.890 ;
        RECT 18.450 29.740 23.500 29.980 ;
        RECT 1.440 26.050 3.650 28.040 ;
        RECT 19.250 26.280 21.820 26.540 ;
        RECT 15.770 24.260 21.820 26.280 ;
      LAYER li1 ;
        RECT 15.600 31.630 18.340 32.120 ;
        RECT 18.890 31.670 23.120 31.840 ;
        RECT 2.910 31.170 8.270 31.410 ;
        RECT 10.490 31.220 14.110 31.460 ;
        RECT 2.910 28.040 3.340 31.170 ;
        RECT 4.050 31.080 8.060 31.170 ;
        RECT 4.050 30.370 4.220 31.080 ;
        RECT 5.010 30.370 5.180 31.080 ;
        RECT 5.970 30.370 6.140 31.080 ;
        RECT 6.930 30.370 7.100 31.080 ;
        RECT 7.890 30.370 8.060 31.080 ;
        RECT 12.170 31.050 12.620 31.220 ;
        RECT 11.320 30.880 13.410 31.050 ;
        RECT 11.320 28.620 11.490 30.880 ;
        RECT 12.280 28.620 12.450 30.880 ;
        RECT 13.240 28.620 13.410 30.880 ;
        RECT 16.490 30.270 16.660 31.630 ;
        RECT 17.450 30.270 17.620 31.630 ;
        RECT 1.310 27.840 3.340 28.040 ;
        RECT 1.310 26.920 1.490 27.840 ;
        RECT 1.750 27.680 2.170 27.840 ;
        RECT 2.440 26.920 2.660 27.840 ;
        RECT 2.920 27.680 3.340 27.840 ;
        RECT 1.310 26.730 2.210 26.920 ;
        RECT 2.440 26.730 3.380 26.920 ;
        RECT 16.490 24.630 16.660 25.990 ;
        RECT 17.450 24.630 17.620 25.990 ;
        RECT 18.060 24.630 18.340 31.630 ;
        RECT 19.650 30.230 19.820 31.670 ;
        RECT 22.130 30.230 22.300 31.670 ;
        RECT 15.610 24.610 18.340 24.630 ;
        RECT 20.450 24.610 20.620 26.050 ;
        RECT 15.610 24.440 21.440 24.610 ;
      LAYER mcon ;
        RECT 16.070 31.840 16.250 32.020 ;
        RECT 16.450 31.840 16.630 32.020 ;
        RECT 16.830 31.840 17.010 32.020 ;
        RECT 17.210 31.840 17.390 32.020 ;
        RECT 17.590 31.840 17.770 32.020 ;
        RECT 17.970 31.840 18.150 32.020 ;
        RECT 2.970 31.200 3.140 31.380 ;
        RECT 3.360 31.200 3.530 31.380 ;
        RECT 3.720 31.200 3.890 31.380 ;
        RECT 4.140 31.200 4.310 31.370 ;
        RECT 4.560 31.200 4.730 31.370 ;
        RECT 4.980 31.200 5.150 31.370 ;
        RECT 5.400 31.200 5.570 31.370 ;
        RECT 5.820 31.200 5.990 31.370 ;
        RECT 6.240 31.200 6.410 31.370 ;
        RECT 6.660 31.200 6.830 31.370 ;
        RECT 7.080 31.200 7.250 31.370 ;
        RECT 7.500 31.200 7.670 31.370 ;
        RECT 7.950 31.200 8.120 31.370 ;
        RECT 10.680 31.250 10.850 31.420 ;
        RECT 11.100 31.250 11.270 31.420 ;
        RECT 11.520 31.250 11.690 31.420 ;
        RECT 11.940 31.250 12.110 31.420 ;
        RECT 12.360 31.250 12.530 31.420 ;
        RECT 12.780 31.250 12.950 31.420 ;
        RECT 13.200 31.250 13.370 31.420 ;
        RECT 13.620 31.250 13.790 31.420 ;
        RECT 1.870 27.870 2.050 28.040 ;
        RECT 3.040 27.870 3.220 28.040 ;
      LAYER met1 ;
        RECT -2.790 31.680 27.130 32.830 ;
        RECT 2.910 31.170 8.270 31.680 ;
        RECT 10.490 31.220 14.110 31.680 ;
        RECT 1.710 27.840 2.200 28.070 ;
        RECT 2.880 27.840 3.370 28.070 ;
      LAYER via ;
        RECT -2.470 31.770 -1.670 32.720 ;
        RECT 26.230 31.770 27.030 32.720 ;
      LAYER met2 ;
        RECT -2.560 31.680 -1.560 32.830 ;
        RECT 26.130 31.680 27.130 32.830 ;
      LAYER via2 ;
        RECT -2.470 31.770 -1.670 32.720 ;
        RECT 26.230 31.770 27.030 32.720 ;
      LAYER met3 ;
        RECT -2.560 31.680 -1.560 32.830 ;
        RECT 26.130 31.680 27.130 32.830 ;
      LAYER via3 ;
        RECT -2.470 31.770 -1.670 32.720 ;
        RECT 26.230 31.770 27.030 32.720 ;
      LAYER met4 ;
        RECT -2.560 13.980 -1.560 41.960 ;
        RECT 26.130 13.980 27.130 41.960 ;
    END
  END VDD
  PIN inn
    ANTENNAGATEAREA 1.200000 ;
    PORT
      LAYER li1 ;
        RECT 4.880 28.950 5.240 29.250 ;
      LAYER mcon ;
        RECT 4.960 29.000 5.160 29.200 ;
      LAYER met1 ;
        RECT -2.790 29.110 5.240 29.250 ;
        RECT 4.880 28.950 5.240 29.110 ;
    END
  END inn
  PIN inp
    ANTENNAGATEAREA 1.200000 ;
    PORT
      LAYER li1 ;
        RECT 6.840 29.200 7.200 29.500 ;
      LAYER mcon ;
        RECT 6.920 29.250 7.120 29.450 ;
      LAYER met1 ;
        RECT -2.790 29.390 7.200 29.530 ;
        RECT 6.840 29.200 7.200 29.390 ;
    END
  END inp
  PIN clk
    ANTENNAGATEAREA 0.195000 ;
    PORT
      LAYER li1 ;
        RECT 1.310 25.770 1.580 26.100 ;
      LAYER mcon ;
        RECT 1.390 25.850 1.560 26.020 ;
      LAYER met1 ;
        RECT 1.280 26.010 1.590 26.100 ;
        RECT -2.790 25.870 1.590 26.010 ;
        RECT 1.280 25.770 1.590 25.870 ;
    END
  END clk
  OBS
      LAYER li1 ;
        RECT 2.530 38.470 5.330 38.670 ;
        RECT 2.530 37.870 3.080 38.470 ;
        RECT 2.530 37.670 5.330 37.870 ;
        RECT 2.530 37.070 3.080 37.670 ;
        RECT 6.080 37.120 6.280 38.670 ;
        RECT 6.880 37.120 7.080 38.670 ;
        RECT 7.680 37.120 7.880 38.670 ;
        RECT 8.480 37.120 8.680 38.670 ;
        RECT 9.280 37.120 9.480 38.670 ;
        RECT 10.080 37.120 10.280 38.670 ;
        RECT 10.880 37.120 11.080 38.670 ;
        RECT 11.680 37.120 11.880 38.670 ;
        RECT 12.480 37.120 12.680 38.670 ;
        RECT 13.280 37.120 13.480 38.670 ;
        RECT 14.080 37.120 14.280 38.670 ;
        RECT 14.880 37.120 15.080 38.670 ;
        RECT 15.680 37.120 15.880 38.670 ;
        RECT 16.480 37.120 16.680 38.670 ;
        RECT 17.280 37.120 17.480 38.670 ;
        RECT 18.080 37.120 18.280 38.670 ;
        RECT 19.030 38.470 21.830 38.670 ;
        RECT 21.280 37.870 21.830 38.470 ;
        RECT 19.030 37.670 21.830 37.870 ;
        RECT 6.080 37.070 18.280 37.120 ;
        RECT 21.280 37.070 21.830 37.670 ;
        RECT 2.530 36.770 21.830 37.070 ;
        RECT 2.530 36.170 3.080 36.770 ;
        RECT 6.080 36.720 18.280 36.770 ;
        RECT 2.530 35.970 5.330 36.170 ;
        RECT 2.530 35.370 3.080 35.970 ;
        RECT 2.530 35.170 5.330 35.370 ;
        RECT 6.080 35.170 6.280 36.720 ;
        RECT 6.880 35.170 7.080 36.720 ;
        RECT 7.680 35.170 7.880 36.720 ;
        RECT 8.480 35.170 8.680 36.720 ;
        RECT 9.280 35.170 9.480 36.720 ;
        RECT 10.080 35.170 10.280 36.720 ;
        RECT 10.880 35.170 11.080 36.720 ;
        RECT 11.680 35.220 11.880 36.720 ;
        RECT 12.480 35.220 12.680 36.720 ;
        RECT 13.280 35.170 13.480 36.720 ;
        RECT 14.080 35.170 14.280 36.720 ;
        RECT 14.880 35.170 15.080 36.720 ;
        RECT 15.680 35.170 15.880 36.720 ;
        RECT 16.480 35.170 16.680 36.720 ;
        RECT 17.280 35.170 17.480 36.720 ;
        RECT 18.080 35.170 18.280 36.720 ;
        RECT 21.280 36.170 21.830 36.770 ;
        RECT 19.030 35.970 21.830 36.170 ;
        RECT 21.280 35.370 21.830 35.970 ;
        RECT 19.030 35.170 21.830 35.370 ;
        RECT 4.530 30.070 4.700 30.910 ;
        RECT 5.490 30.070 5.660 30.910 ;
        RECT 4.530 29.900 5.660 30.070 ;
        RECT 6.450 30.070 6.620 30.910 ;
        RECT 7.410 30.070 7.580 30.910 ;
        RECT 8.530 30.270 9.480 31.220 ;
        RECT 9.710 30.830 10.840 31.000 ;
        RECT 6.450 29.900 7.580 30.070 ;
        RECT 3.510 29.600 3.840 29.890 ;
        RECT 1.750 27.380 2.190 27.410 ;
        RECT 2.920 27.380 3.360 27.410 ;
        RECT 1.730 27.190 2.210 27.380 ;
        RECT 2.900 27.190 3.380 27.380 ;
        RECT 1.730 26.290 2.210 26.460 ;
        RECT 2.900 26.290 3.380 26.460 ;
        RECT 1.750 26.230 2.190 26.290 ;
        RECT 2.920 26.230 3.360 26.290 ;
        RECT 1.750 26.050 2.170 26.230 ;
        RECT 2.480 26.050 2.750 26.100 ;
        RECT 1.750 25.820 2.750 26.050 ;
        RECT 1.750 25.650 2.170 25.820 ;
        RECT 2.480 25.770 2.750 25.820 ;
        RECT 2.920 26.050 3.340 26.230 ;
        RECT 3.610 26.050 3.840 29.600 ;
        RECT 4.530 28.780 4.700 29.900 ;
        RECT 5.420 28.780 5.660 29.080 ;
        RECT 4.530 28.610 5.660 28.780 ;
        RECT 2.920 25.900 3.840 26.050 ;
        RECT 4.050 26.130 4.220 28.340 ;
        RECT 4.530 26.300 4.700 28.610 ;
        RECT 5.010 26.130 5.180 28.340 ;
        RECT 5.490 26.300 5.660 28.610 ;
        RECT 6.450 28.790 6.620 29.900 ;
        RECT 6.450 28.620 8.830 28.790 ;
        RECT 5.970 26.130 6.140 28.340 ;
        RECT 6.450 26.300 6.620 28.620 ;
        RECT 6.930 26.130 7.100 28.340 ;
        RECT 7.410 26.300 7.580 28.620 ;
        RECT 7.890 26.130 8.060 28.340 ;
        RECT 8.450 28.170 8.830 28.620 ;
        RECT 9.060 28.340 9.440 30.270 ;
        RECT 8.450 27.110 9.440 28.170 ;
        RECT 9.710 28.030 9.880 30.830 ;
        RECT 10.190 28.370 10.360 30.660 ;
        RECT 10.670 28.620 10.840 30.830 ;
        RECT 13.890 30.830 15.020 31.000 ;
        RECT 11.800 28.370 11.970 30.660 ;
        RECT 10.190 28.200 11.970 28.370 ;
        RECT 12.760 28.370 12.930 30.660 ;
        RECT 13.890 28.620 14.060 30.830 ;
        RECT 14.370 28.370 14.540 30.660 ;
        RECT 12.760 28.200 14.540 28.370 ;
        RECT 14.850 29.930 15.020 30.830 ;
        RECT 14.850 29.240 15.840 29.930 ;
        RECT 16.010 29.880 16.180 31.310 ;
        RECT 16.010 29.540 16.800 29.880 ;
        RECT 16.970 29.700 17.140 31.310 ;
        RECT 18.690 31.240 19.020 31.500 ;
        RECT 21.170 31.240 21.500 31.500 ;
        RECT 19.170 30.230 19.340 31.070 ;
        RECT 20.130 30.230 20.300 31.070 ;
        RECT 21.650 30.230 21.820 31.070 ;
        RECT 22.610 30.230 22.780 31.070 ;
        RECT 17.510 29.700 17.810 29.750 ;
        RECT 14.850 28.030 15.020 29.240 ;
        RECT 16.010 28.640 16.180 29.540 ;
        RECT 16.970 29.510 17.880 29.700 ;
        RECT 16.970 28.640 17.140 29.510 ;
        RECT 17.510 29.450 17.810 29.510 ;
        RECT 9.630 27.860 11.690 28.030 ;
        RECT 11.870 27.860 15.080 28.030 ;
        RECT 11.520 27.690 11.690 27.860 ;
        RECT 11.520 27.520 12.870 27.690 ;
        RECT 4.050 25.950 8.060 26.130 ;
        RECT 2.920 25.820 3.880 25.900 ;
        RECT 2.920 25.650 3.340 25.820 ;
        RECT 1.730 25.480 2.190 25.650 ;
        RECT 2.900 25.480 3.360 25.650 ;
        RECT 3.550 25.630 3.880 25.820 ;
        RECT 1.750 25.450 2.170 25.480 ;
        RECT 2.920 25.450 3.340 25.480 ;
        RECT 4.050 25.000 4.220 25.950 ;
        RECT 5.010 25.000 5.180 25.950 ;
        RECT 5.970 25.000 6.140 25.950 ;
        RECT 6.930 25.000 7.100 25.950 ;
        RECT 7.890 25.000 8.060 25.950 ;
        RECT 9.060 25.820 9.440 27.110 ;
        RECT 9.030 24.870 9.980 25.820 ;
        RECT 11.800 24.970 11.970 27.520 ;
        RECT 13.090 27.350 13.260 27.860 ;
        RECT 12.760 27.180 13.260 27.350 ;
        RECT 14.140 27.190 14.750 27.530 ;
        RECT 12.760 24.970 12.930 27.180 ;
        RECT 16.010 26.720 16.180 27.620 ;
        RECT 16.970 26.750 17.140 27.620 ;
        RECT 17.530 26.750 17.830 26.800 ;
        RECT 16.010 26.380 16.800 26.720 ;
        RECT 16.970 26.560 17.890 26.750 ;
        RECT 16.010 24.950 16.180 26.380 ;
        RECT 16.970 24.950 17.140 26.560 ;
        RECT 17.530 26.500 17.830 26.560 ;
        RECT 18.510 25.040 18.750 28.710 ;
        RECT 18.920 26.260 19.160 28.240 ;
        RECT 20.070 26.230 20.400 26.490 ;
        RECT 19.970 25.210 20.140 26.050 ;
        RECT 20.930 25.210 21.100 26.050 ;
        RECT 18.510 24.780 19.820 25.040 ;
        RECT 10.390 24.380 11.110 24.650 ;
        RECT 2.530 20.520 5.330 20.720 ;
        RECT 2.530 19.920 3.080 20.520 ;
        RECT 2.530 19.720 5.330 19.920 ;
        RECT 2.530 19.120 3.080 19.720 ;
        RECT 6.080 19.170 6.280 20.720 ;
        RECT 6.880 19.170 7.080 20.720 ;
        RECT 7.680 19.170 7.880 20.720 ;
        RECT 8.480 19.170 8.680 20.720 ;
        RECT 9.280 19.170 9.480 20.720 ;
        RECT 10.080 19.170 10.280 20.720 ;
        RECT 10.880 19.170 11.080 20.720 ;
        RECT 11.680 19.170 11.880 20.720 ;
        RECT 12.480 19.170 12.680 20.720 ;
        RECT 13.280 19.170 13.480 20.720 ;
        RECT 14.080 19.170 14.280 20.720 ;
        RECT 14.880 19.170 15.080 20.720 ;
        RECT 15.680 19.170 15.880 20.720 ;
        RECT 16.480 19.170 16.680 20.720 ;
        RECT 17.280 19.170 17.480 20.720 ;
        RECT 18.080 19.170 18.280 20.720 ;
        RECT 19.030 20.520 21.830 20.720 ;
        RECT 21.280 19.920 21.830 20.520 ;
        RECT 19.030 19.720 21.830 19.920 ;
        RECT 6.080 19.120 18.280 19.170 ;
        RECT 21.280 19.120 21.830 19.720 ;
        RECT 2.530 18.820 21.830 19.120 ;
        RECT 2.530 18.220 3.080 18.820 ;
        RECT 6.080 18.770 18.280 18.820 ;
        RECT 2.530 18.020 5.330 18.220 ;
        RECT 2.530 17.420 3.080 18.020 ;
        RECT 2.530 17.220 5.330 17.420 ;
        RECT 6.080 17.220 6.280 18.770 ;
        RECT 6.880 17.220 7.080 18.770 ;
        RECT 7.680 17.220 7.880 18.770 ;
        RECT 8.480 17.220 8.680 18.770 ;
        RECT 9.280 17.220 9.480 18.770 ;
        RECT 10.080 17.220 10.280 18.770 ;
        RECT 10.880 17.220 11.080 18.770 ;
        RECT 11.680 17.270 11.880 18.770 ;
        RECT 12.480 17.270 12.680 18.770 ;
        RECT 13.280 17.220 13.480 18.770 ;
        RECT 14.080 17.220 14.280 18.770 ;
        RECT 14.880 17.220 15.080 18.770 ;
        RECT 15.680 17.220 15.880 18.770 ;
        RECT 16.480 17.220 16.680 18.770 ;
        RECT 17.280 17.220 17.480 18.770 ;
        RECT 18.080 17.220 18.280 18.770 ;
        RECT 21.280 18.220 21.830 18.820 ;
        RECT 19.030 18.020 21.830 18.220 ;
        RECT 21.280 17.420 21.830 18.020 ;
        RECT 19.030 17.220 21.830 17.420 ;
      LAYER mcon ;
        RECT 2.630 37.520 2.880 37.770 ;
        RECT 2.630 37.070 2.880 37.320 ;
        RECT 21.480 37.470 21.730 37.720 ;
        RECT 21.480 37.020 21.730 37.270 ;
        RECT 2.630 36.570 2.880 36.820 ;
        RECT 2.630 36.120 2.880 36.370 ;
        RECT 21.480 36.520 21.730 36.770 ;
        RECT 21.480 36.070 21.730 36.320 ;
        RECT 8.630 30.370 9.380 31.120 ;
        RECT 1.810 27.200 2.110 27.370 ;
        RECT 2.980 27.200 3.280 27.370 ;
        RECT 1.810 26.290 2.110 26.460 ;
        RECT 2.980 26.290 3.280 26.460 ;
        RECT 2.560 25.850 2.730 26.020 ;
        RECT 5.450 28.870 5.630 29.050 ;
        RECT 9.160 29.220 9.340 29.400 ;
        RECT 9.160 28.850 9.340 29.030 ;
        RECT 9.160 28.480 9.340 28.660 ;
        RECT 9.160 27.930 9.340 28.110 ;
        RECT 15.630 29.680 15.810 29.850 ;
        RECT 15.630 29.320 15.810 29.490 ;
        RECT 21.250 31.300 21.420 31.470 ;
        RECT 17.540 29.510 17.720 29.690 ;
        RECT 9.160 27.550 9.340 27.730 ;
        RECT 9.160 27.180 9.340 27.360 ;
        RECT 9.130 24.970 9.880 25.720 ;
        RECT 14.170 27.270 14.350 27.450 ;
        RECT 14.540 27.270 14.720 27.450 ;
        RECT 17.560 26.560 17.740 26.740 ;
        RECT 18.540 26.620 18.720 26.800 ;
        RECT 18.950 28.000 19.130 28.180 ;
        RECT 18.950 26.320 19.130 26.500 ;
        RECT 20.150 26.270 20.320 26.440 ;
        RECT 10.470 24.430 10.640 24.600 ;
        RECT 10.860 24.430 11.030 24.600 ;
        RECT 2.630 19.570 2.880 19.820 ;
        RECT 2.630 19.120 2.880 19.370 ;
        RECT 21.480 19.520 21.730 19.770 ;
        RECT 21.480 19.070 21.730 19.320 ;
        RECT 2.630 18.620 2.880 18.870 ;
        RECT 2.630 18.170 2.880 18.420 ;
        RECT 21.480 18.570 21.730 18.820 ;
        RECT 21.480 18.120 21.730 18.370 ;
      LAYER met1 ;
        RECT 6.930 39.670 17.430 40.870 ;
        RECT 11.880 39.220 12.480 39.670 ;
        RECT 6.280 39.070 18.080 39.220 ;
        RECT 1.330 37.220 2.980 37.870 ;
        RECT 3.430 37.220 3.580 38.720 ;
        RECT 4.030 37.220 4.180 38.720 ;
        RECT 4.630 37.220 4.780 38.720 ;
        RECT 5.230 37.220 5.380 38.720 ;
        RECT 11.880 38.620 12.480 39.070 ;
        RECT 6.280 38.470 18.080 38.620 ;
        RECT 11.880 38.020 12.480 38.470 ;
        RECT 6.280 37.870 18.080 38.020 ;
        RECT 11.880 37.420 12.480 37.870 ;
        RECT 6.280 37.270 18.080 37.420 ;
        RECT 1.330 37.120 5.380 37.220 ;
        RECT 11.880 37.120 12.480 37.270 ;
        RECT 18.980 37.220 19.130 38.720 ;
        RECT 19.580 37.220 19.730 38.720 ;
        RECT 20.180 37.220 20.330 38.720 ;
        RECT 20.780 37.220 20.930 38.720 ;
        RECT 21.380 37.220 23.030 37.820 ;
        RECT 18.980 37.120 23.030 37.220 ;
        RECT 1.330 36.420 23.030 37.120 ;
        RECT 1.330 36.020 2.980 36.420 ;
        RECT 3.430 35.120 3.580 36.420 ;
        RECT 4.030 35.120 4.180 36.420 ;
        RECT 4.630 35.120 4.780 36.420 ;
        RECT 5.230 35.120 5.380 36.420 ;
        RECT 11.880 35.970 12.480 36.420 ;
        RECT 6.280 35.820 18.080 35.970 ;
        RECT 11.880 35.370 12.480 35.820 ;
        RECT 6.280 35.220 18.080 35.370 ;
        RECT 11.880 34.770 12.480 35.220 ;
        RECT 18.980 35.120 19.130 36.420 ;
        RECT 19.580 35.120 19.730 36.420 ;
        RECT 20.180 35.120 20.330 36.420 ;
        RECT 20.780 35.120 20.930 36.420 ;
        RECT 21.380 35.970 23.030 36.420 ;
        RECT 6.280 34.620 18.080 34.770 ;
        RECT 11.880 34.170 12.480 34.620 ;
        RECT 6.930 32.970 17.430 34.170 ;
        RECT 17.810 31.500 19.030 31.530 ;
        RECT 17.810 31.360 21.480 31.500 ;
        RECT 8.530 30.270 9.480 31.220 ;
        RECT 5.390 29.060 5.660 29.080 ;
        RECT 9.100 29.060 9.400 29.450 ;
        RECT 15.560 29.230 15.840 29.930 ;
        RECT 17.810 29.750 17.990 31.360 ;
        RECT 21.170 31.270 21.480 31.360 ;
        RECT 17.510 29.450 17.990 29.750 ;
        RECT 5.390 28.990 9.400 29.060 ;
        RECT 5.380 28.800 9.400 28.990 ;
        RECT 9.100 28.450 9.400 28.800 ;
        RECT 17.810 28.240 17.990 29.450 ;
        RECT 1.770 26.230 2.160 27.440 ;
        RECT 2.940 26.230 3.330 27.440 ;
        RECT 9.100 27.370 9.400 28.140 ;
        RECT 17.810 28.050 19.160 28.240 ;
        RECT 18.920 27.940 19.160 28.050 ;
        RECT 14.120 27.370 14.770 27.530 ;
        RECT 9.100 27.190 14.770 27.370 ;
        RECT 9.100 27.150 9.400 27.190 ;
        RECT 17.530 26.750 17.830 26.800 ;
        RECT 18.510 26.750 18.750 26.860 ;
        RECT 17.530 26.560 18.750 26.750 ;
        RECT 17.530 26.500 17.830 26.560 ;
        RECT 18.920 26.430 19.160 26.560 ;
        RECT 20.070 26.430 20.400 26.490 ;
        RECT 18.920 26.250 20.400 26.430 ;
        RECT 18.920 26.240 19.410 26.250 ;
        RECT 20.070 26.230 20.400 26.250 ;
        RECT 2.480 25.930 2.760 26.100 ;
        RECT 2.480 25.770 3.780 25.930 ;
        RECT 3.570 24.650 3.780 25.770 ;
        RECT 9.030 24.870 9.980 25.820 ;
        RECT 3.570 24.380 11.110 24.650 ;
        RECT 6.930 21.720 17.430 22.920 ;
        RECT 11.880 21.270 12.480 21.720 ;
        RECT 6.280 21.120 18.080 21.270 ;
        RECT 1.330 19.270 2.980 19.920 ;
        RECT 3.430 19.270 3.580 20.770 ;
        RECT 4.030 19.270 4.180 20.770 ;
        RECT 4.630 19.270 4.780 20.770 ;
        RECT 5.230 19.270 5.380 20.770 ;
        RECT 11.880 20.670 12.480 21.120 ;
        RECT 6.280 20.520 18.080 20.670 ;
        RECT 11.880 20.070 12.480 20.520 ;
        RECT 6.280 19.920 18.080 20.070 ;
        RECT 11.880 19.470 12.480 19.920 ;
        RECT 6.280 19.320 18.080 19.470 ;
        RECT 1.330 19.170 5.380 19.270 ;
        RECT 11.880 19.170 12.480 19.320 ;
        RECT 18.980 19.270 19.130 20.770 ;
        RECT 19.580 19.270 19.730 20.770 ;
        RECT 20.180 19.270 20.330 20.770 ;
        RECT 20.780 19.270 20.930 20.770 ;
        RECT 21.380 19.270 23.030 19.870 ;
        RECT 18.980 19.170 23.030 19.270 ;
        RECT 1.330 18.470 23.030 19.170 ;
        RECT 1.330 18.070 2.980 18.470 ;
        RECT 3.430 17.170 3.580 18.470 ;
        RECT 4.030 17.170 4.180 18.470 ;
        RECT 4.630 17.170 4.780 18.470 ;
        RECT 5.230 17.170 5.380 18.470 ;
        RECT 11.880 18.020 12.480 18.470 ;
        RECT 6.280 17.870 18.080 18.020 ;
        RECT 11.880 17.420 12.480 17.870 ;
        RECT 6.280 17.270 18.080 17.420 ;
        RECT 11.880 16.820 12.480 17.270 ;
        RECT 18.980 17.170 19.130 18.470 ;
        RECT 19.580 17.170 19.730 18.470 ;
        RECT 20.180 17.170 20.330 18.470 ;
        RECT 20.780 17.170 20.930 18.470 ;
        RECT 21.380 18.020 23.030 18.470 ;
        RECT 6.280 16.670 18.080 16.820 ;
        RECT 11.880 16.220 12.480 16.670 ;
        RECT 6.930 15.020 17.430 16.220 ;
      LAYER via ;
        RECT 7.030 39.770 8.030 40.770 ;
        RECT 8.130 39.770 9.130 40.770 ;
        RECT 11.730 39.770 12.630 40.770 ;
        RECT 15.230 39.770 16.230 40.770 ;
        RECT 16.330 39.770 17.330 40.770 ;
        RECT 1.430 37.170 2.430 37.720 ;
        RECT 21.930 37.170 22.930 37.720 ;
        RECT 1.430 36.120 2.430 36.670 ;
        RECT 21.930 36.120 22.930 36.670 ;
        RECT 7.030 33.070 8.030 34.070 ;
        RECT 8.130 33.070 9.130 34.070 ;
        RECT 11.730 33.070 12.630 34.070 ;
        RECT 15.230 33.070 16.230 34.070 ;
        RECT 16.330 33.070 17.330 34.070 ;
        RECT 8.630 30.370 9.380 31.120 ;
        RECT 9.130 24.970 9.880 25.720 ;
        RECT 7.030 21.820 8.030 22.820 ;
        RECT 8.130 21.820 9.130 22.820 ;
        RECT 11.730 21.820 12.630 22.820 ;
        RECT 15.230 21.820 16.230 22.820 ;
        RECT 16.330 21.820 17.330 22.820 ;
        RECT 1.430 19.220 2.430 19.770 ;
        RECT 21.930 19.220 22.930 19.770 ;
        RECT 1.430 18.170 2.430 18.720 ;
        RECT 21.930 18.170 22.930 18.720 ;
        RECT 7.030 15.120 8.030 16.120 ;
        RECT 8.130 15.120 9.130 16.120 ;
        RECT 11.730 15.120 12.630 16.120 ;
        RECT 15.230 15.120 16.230 16.120 ;
        RECT 16.330 15.120 17.330 16.120 ;
      LAYER met2 ;
        RECT 6.930 39.470 17.430 40.870 ;
        RECT 3.430 38.870 20.930 39.470 ;
        RECT 5.430 38.420 5.730 38.870 ;
        RECT 3.430 38.270 5.730 38.420 ;
        RECT 5.430 37.820 5.730 38.270 ;
        RECT 1.330 36.020 2.530 37.820 ;
        RECT 3.430 37.670 5.730 37.820 ;
        RECT 5.430 37.220 5.730 37.670 ;
        RECT 6.180 37.220 6.330 38.870 ;
        RECT 6.780 37.220 6.930 38.870 ;
        RECT 7.380 37.220 7.530 38.870 ;
        RECT 7.980 37.220 8.130 38.870 ;
        RECT 8.580 37.220 8.730 38.870 ;
        RECT 9.180 37.220 9.330 38.870 ;
        RECT 9.780 37.220 9.930 38.870 ;
        RECT 10.380 37.220 10.530 38.870 ;
        RECT 10.980 37.220 11.130 38.870 ;
        RECT 11.580 37.220 11.730 38.870 ;
        RECT 12.630 37.220 12.780 38.870 ;
        RECT 13.230 37.220 13.380 38.870 ;
        RECT 13.830 37.220 13.980 38.870 ;
        RECT 14.430 37.220 14.580 38.870 ;
        RECT 15.030 37.220 15.180 38.870 ;
        RECT 15.630 37.220 15.780 38.870 ;
        RECT 16.230 37.220 16.380 38.870 ;
        RECT 16.830 37.220 16.980 38.870 ;
        RECT 17.430 37.220 17.580 38.870 ;
        RECT 18.030 37.220 18.180 38.870 ;
        RECT 18.630 38.420 18.930 38.870 ;
        RECT 18.630 38.270 20.930 38.420 ;
        RECT 18.630 37.820 18.930 38.270 ;
        RECT 18.630 37.670 20.930 37.820 ;
        RECT 18.630 37.220 18.930 37.670 ;
        RECT 5.430 36.170 5.730 36.620 ;
        RECT 3.430 36.020 5.730 36.170 ;
        RECT 5.430 35.570 5.730 36.020 ;
        RECT 3.430 35.420 5.730 35.570 ;
        RECT 5.430 34.970 5.730 35.420 ;
        RECT 6.180 34.970 6.330 36.620 ;
        RECT 6.780 34.970 6.930 36.620 ;
        RECT 7.380 34.970 7.530 36.620 ;
        RECT 7.980 34.970 8.130 36.620 ;
        RECT 8.580 34.970 8.730 36.620 ;
        RECT 9.180 34.970 9.330 36.620 ;
        RECT 9.780 34.970 9.930 36.620 ;
        RECT 10.380 34.970 10.530 36.620 ;
        RECT 10.980 34.970 11.130 36.620 ;
        RECT 11.580 34.970 11.730 36.620 ;
        RECT 12.630 34.970 12.780 36.620 ;
        RECT 13.230 34.970 13.380 36.620 ;
        RECT 13.830 34.970 13.980 36.620 ;
        RECT 14.430 34.970 14.580 36.620 ;
        RECT 15.030 34.970 15.180 36.620 ;
        RECT 15.630 34.970 15.780 36.620 ;
        RECT 16.230 34.970 16.380 36.620 ;
        RECT 16.830 34.970 16.980 36.620 ;
        RECT 17.430 34.970 17.580 36.620 ;
        RECT 18.030 34.970 18.180 36.620 ;
        RECT 18.630 36.170 18.930 36.620 ;
        RECT 18.630 36.020 20.930 36.170 ;
        RECT 21.830 36.020 23.030 37.820 ;
        RECT 18.630 35.570 18.930 36.020 ;
        RECT 18.630 35.420 20.930 35.570 ;
        RECT 18.630 34.970 18.930 35.420 ;
        RECT 3.430 34.370 20.930 34.970 ;
        RECT 6.930 32.970 17.430 34.370 ;
        RECT 8.530 30.270 9.480 32.970 ;
        RECT 9.030 22.920 9.980 25.820 ;
        RECT 6.930 21.520 17.430 22.920 ;
        RECT 3.430 20.920 20.930 21.520 ;
        RECT 5.430 20.470 5.730 20.920 ;
        RECT 3.430 20.320 5.730 20.470 ;
        RECT 5.430 19.870 5.730 20.320 ;
        RECT 1.330 18.070 2.530 19.870 ;
        RECT 3.430 19.720 5.730 19.870 ;
        RECT 5.430 19.270 5.730 19.720 ;
        RECT 6.180 19.270 6.330 20.920 ;
        RECT 6.780 19.270 6.930 20.920 ;
        RECT 7.380 19.270 7.530 20.920 ;
        RECT 7.980 19.270 8.130 20.920 ;
        RECT 8.580 19.270 8.730 20.920 ;
        RECT 9.180 19.270 9.330 20.920 ;
        RECT 9.780 19.270 9.930 20.920 ;
        RECT 10.380 19.270 10.530 20.920 ;
        RECT 10.980 19.270 11.130 20.920 ;
        RECT 11.580 19.270 11.730 20.920 ;
        RECT 12.630 19.270 12.780 20.920 ;
        RECT 13.230 19.270 13.380 20.920 ;
        RECT 13.830 19.270 13.980 20.920 ;
        RECT 14.430 19.270 14.580 20.920 ;
        RECT 15.030 19.270 15.180 20.920 ;
        RECT 15.630 19.270 15.780 20.920 ;
        RECT 16.230 19.270 16.380 20.920 ;
        RECT 16.830 19.270 16.980 20.920 ;
        RECT 17.430 19.270 17.580 20.920 ;
        RECT 18.030 19.270 18.180 20.920 ;
        RECT 18.630 20.470 18.930 20.920 ;
        RECT 18.630 20.320 20.930 20.470 ;
        RECT 18.630 19.870 18.930 20.320 ;
        RECT 18.630 19.720 20.930 19.870 ;
        RECT 18.630 19.270 18.930 19.720 ;
        RECT 5.430 18.220 5.730 18.670 ;
        RECT 3.430 18.070 5.730 18.220 ;
        RECT 5.430 17.620 5.730 18.070 ;
        RECT 3.430 17.470 5.730 17.620 ;
        RECT 5.430 17.020 5.730 17.470 ;
        RECT 6.180 17.020 6.330 18.670 ;
        RECT 6.780 17.020 6.930 18.670 ;
        RECT 7.380 17.020 7.530 18.670 ;
        RECT 7.980 17.020 8.130 18.670 ;
        RECT 8.580 17.020 8.730 18.670 ;
        RECT 9.180 17.020 9.330 18.670 ;
        RECT 9.780 17.020 9.930 18.670 ;
        RECT 10.380 17.020 10.530 18.670 ;
        RECT 10.980 17.020 11.130 18.670 ;
        RECT 11.580 17.020 11.730 18.670 ;
        RECT 12.630 17.020 12.780 18.670 ;
        RECT 13.230 17.020 13.380 18.670 ;
        RECT 13.830 17.020 13.980 18.670 ;
        RECT 14.430 17.020 14.580 18.670 ;
        RECT 15.030 17.020 15.180 18.670 ;
        RECT 15.630 17.020 15.780 18.670 ;
        RECT 16.230 17.020 16.380 18.670 ;
        RECT 16.830 17.020 16.980 18.670 ;
        RECT 17.430 17.020 17.580 18.670 ;
        RECT 18.030 17.020 18.180 18.670 ;
        RECT 18.630 18.220 18.930 18.670 ;
        RECT 18.630 18.070 20.930 18.220 ;
        RECT 21.830 18.070 23.030 19.870 ;
        RECT 18.630 17.620 18.930 18.070 ;
        RECT 18.630 17.470 20.930 17.620 ;
        RECT 18.630 17.020 18.930 17.470 ;
        RECT 3.430 16.420 20.930 17.020 ;
        RECT 6.930 15.020 17.430 16.420 ;
  END
END adc_comp_latch
END LIBRARY

