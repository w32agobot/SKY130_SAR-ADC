magic
tech sky130A
timestamp 1658400657
<< nwell >>
rect 0 400 680 660
<< nmos >>
rect 130 160 148 202
rect 178 160 196 202
rect 330 160 348 202
rect 378 160 396 202
rect 426 160 444 202
<< pmos >>
rect 120 440 138 530
rect 188 440 206 530
rect 332 440 350 530
rect 400 440 418 530
rect 468 440 486 530
<< ndiff >>
rect 100 189 130 202
rect 100 172 106 189
rect 124 172 130 189
rect 100 160 130 172
rect 148 189 178 202
rect 148 172 154 189
rect 172 172 178 189
rect 148 160 178 172
rect 196 189 226 202
rect 196 172 202 189
rect 220 172 226 189
rect 196 160 226 172
rect 300 189 330 202
rect 300 172 306 189
rect 324 172 330 189
rect 300 160 330 172
rect 348 189 378 202
rect 348 172 354 189
rect 372 172 378 189
rect 348 160 378 172
rect 396 189 426 202
rect 396 172 402 189
rect 420 172 426 189
rect 396 160 426 172
rect 444 189 473 202
rect 444 172 450 189
rect 468 172 473 189
rect 444 160 473 172
<< pdiff >>
rect 70 509 120 530
rect 70 492 86 509
rect 104 492 120 509
rect 70 468 120 492
rect 70 451 86 468
rect 104 451 120 468
rect 70 440 120 451
rect 138 509 188 530
rect 138 492 154 509
rect 172 492 188 509
rect 138 468 188 492
rect 138 451 154 468
rect 172 451 188 468
rect 138 440 188 451
rect 206 509 251 530
rect 206 492 222 509
rect 240 492 251 509
rect 206 468 251 492
rect 206 451 222 468
rect 240 451 251 468
rect 206 440 251 451
rect 282 509 332 530
rect 282 492 298 509
rect 316 492 332 509
rect 282 468 332 492
rect 282 451 298 468
rect 316 451 332 468
rect 282 440 332 451
rect 350 509 400 530
rect 350 492 366 509
rect 384 492 400 509
rect 350 468 400 492
rect 350 451 366 468
rect 384 451 400 468
rect 350 440 400 451
rect 418 509 468 530
rect 418 492 434 509
rect 452 492 468 509
rect 418 468 468 492
rect 418 451 434 468
rect 452 451 468 468
rect 418 440 468 451
rect 486 509 536 530
rect 486 492 502 509
rect 520 492 536 509
rect 486 468 536 492
rect 486 451 502 468
rect 520 451 536 468
rect 486 440 536 451
<< ndiffc >>
rect 106 172 124 189
rect 154 172 172 189
rect 202 172 220 189
rect 306 172 324 189
rect 354 172 372 189
rect 402 172 420 189
rect 450 172 468 189
<< pdiffc >>
rect 86 492 104 509
rect 86 451 104 468
rect 154 492 172 509
rect 154 451 172 468
rect 222 492 240 509
rect 222 451 240 468
rect 298 492 316 509
rect 298 451 316 468
rect 366 492 384 509
rect 366 451 384 468
rect 434 492 452 509
rect 434 451 452 468
rect 502 492 520 509
rect 502 451 520 468
<< psubdiff >>
rect 40 70 640 80
rect 40 50 110 70
rect 130 50 170 70
rect 190 50 230 70
rect 250 50 290 70
rect 310 50 350 70
rect 370 50 410 70
rect 430 50 470 70
rect 490 50 530 70
rect 550 50 640 70
rect 40 40 640 50
<< nsubdiff >>
rect 40 630 640 640
rect 40 610 110 630
rect 130 610 170 630
rect 190 610 230 630
rect 250 610 290 630
rect 310 610 350 630
rect 370 610 410 630
rect 430 610 470 630
rect 490 610 530 630
rect 550 610 640 630
rect 40 600 640 610
<< psubdiffcont >>
rect 110 50 130 70
rect 170 50 190 70
rect 230 50 250 70
rect 290 50 310 70
rect 350 50 370 70
rect 410 50 430 70
rect 470 50 490 70
rect 530 50 550 70
<< nsubdiffcont >>
rect 110 610 130 630
rect 170 610 190 630
rect 230 610 250 630
rect 290 610 310 630
rect 350 610 370 630
rect 410 610 430 630
rect 470 610 490 630
rect 530 610 550 630
<< poly >>
rect 105 578 145 583
rect 105 554 113 578
rect 137 554 145 578
rect 105 549 145 554
rect 400 580 649 590
rect 400 572 617 580
rect 120 530 138 549
rect 188 530 206 543
rect 332 530 350 543
rect 400 530 418 572
rect 609 556 617 572
rect 641 556 649 580
rect 609 551 649 556
rect 468 530 486 543
rect 120 293 138 440
rect 188 389 206 440
rect 188 383 246 389
rect 188 359 214 383
rect 238 359 246 383
rect 188 354 246 359
rect 332 363 350 440
rect 400 427 418 440
rect 188 293 206 354
rect 332 345 396 363
rect 120 275 148 293
rect 130 202 148 275
rect 178 275 206 293
rect 308 318 348 323
rect 308 294 316 318
rect 340 294 348 318
rect 308 288 348 294
rect 178 202 196 275
rect 330 202 348 288
rect 378 288 396 345
rect 468 323 486 440
rect 468 317 508 323
rect 468 293 476 317
rect 500 293 508 317
rect 468 288 508 293
rect 378 283 418 288
rect 378 259 386 283
rect 410 259 418 283
rect 378 253 418 259
rect 378 202 396 253
rect 426 202 444 218
rect 130 147 148 160
rect 178 147 196 160
rect 330 147 348 160
rect 378 147 396 160
rect 426 147 444 160
rect 609 159 649 165
rect 609 147 617 159
rect 426 135 617 147
rect 641 135 649 159
rect 426 129 649 135
<< polycont >>
rect 113 554 137 578
rect 617 556 641 580
rect 214 359 238 383
rect 316 294 340 318
rect 476 293 500 317
rect 386 259 410 283
rect 617 135 641 159
<< locali >>
rect 34 517 67 680
rect 101 630 139 638
rect 101 610 110 630
rect 130 610 139 630
rect 101 601 139 610
rect 161 630 199 638
rect 161 610 170 630
rect 190 610 199 630
rect 161 601 199 610
rect 221 630 259 638
rect 221 610 230 630
rect 250 610 259 630
rect 221 601 259 610
rect 281 630 319 638
rect 281 610 290 630
rect 310 610 319 630
rect 281 601 319 610
rect 341 630 379 638
rect 341 610 350 630
rect 370 610 379 630
rect 341 601 379 610
rect 401 637 439 638
rect 461 637 499 638
rect 401 630 499 637
rect 401 610 410 630
rect 430 610 470 630
rect 490 610 499 630
rect 401 601 499 610
rect 521 630 559 638
rect 521 610 530 630
rect 550 610 559 630
rect 521 601 559 610
rect 419 600 481 601
rect 105 578 145 583
rect 105 554 113 578
rect 137 554 145 578
rect 105 549 145 554
rect 34 509 105 517
rect 34 492 86 509
rect 104 492 105 509
rect 34 468 105 492
rect 34 451 86 468
rect 104 451 105 468
rect 34 443 105 451
rect 153 509 173 517
rect 153 492 154 509
rect 172 492 173 509
rect 153 468 173 492
rect 153 451 154 468
rect 172 451 173 468
rect 34 127 67 443
rect 84 233 125 239
rect 84 209 92 233
rect 116 209 125 233
rect 84 203 125 209
rect 106 189 125 203
rect 124 172 125 189
rect 106 164 125 172
rect 153 189 173 451
rect 221 513 317 517
rect 221 509 285 513
rect 309 509 317 513
rect 221 492 222 509
rect 240 492 285 509
rect 316 492 317 509
rect 221 489 285 492
rect 309 489 317 492
rect 221 470 317 489
rect 221 468 286 470
rect 310 468 317 470
rect 221 451 222 468
rect 240 451 286 468
rect 316 451 317 468
rect 221 446 286 451
rect 310 446 317 451
rect 221 443 317 446
rect 365 509 385 542
rect 365 492 366 509
rect 384 492 385 509
rect 365 468 385 492
rect 365 451 366 468
rect 384 451 385 468
rect 365 443 385 451
rect 433 509 453 600
rect 616 590 649 680
rect 609 580 649 590
rect 609 556 617 580
rect 641 556 649 580
rect 609 551 649 556
rect 433 492 434 509
rect 452 492 453 509
rect 433 468 453 492
rect 433 451 434 468
rect 452 451 453 468
rect 433 443 453 451
rect 501 514 541 517
rect 501 509 510 514
rect 501 492 502 509
rect 501 490 510 492
rect 534 490 541 514
rect 501 471 541 490
rect 501 468 510 471
rect 501 451 502 468
rect 501 447 510 451
rect 534 447 541 471
rect 501 443 541 447
rect 206 383 246 389
rect 206 359 214 383
rect 238 359 246 383
rect 206 354 246 359
rect 263 239 282 443
rect 308 318 348 323
rect 308 294 316 318
rect 340 294 348 318
rect 308 288 348 294
rect 468 317 508 323
rect 468 293 476 317
rect 500 293 508 317
rect 468 288 508 293
rect 378 283 418 288
rect 378 259 386 283
rect 410 259 418 283
rect 378 253 418 259
rect 263 233 324 239
rect 263 209 290 233
rect 314 209 324 233
rect 263 203 324 209
rect 153 172 154 189
rect 172 172 173 189
rect 153 164 173 172
rect 202 189 220 197
rect 34 108 41 127
rect 60 108 67 127
rect 34 0 67 108
rect 202 135 220 172
rect 306 189 324 203
rect 306 164 324 172
rect 354 214 468 231
rect 354 189 372 214
rect 354 164 372 172
rect 402 189 420 197
rect 202 128 243 135
rect 202 104 211 128
rect 235 104 243 128
rect 202 99 243 104
rect 402 78 420 172
rect 450 189 468 214
rect 450 164 468 172
rect 616 165 649 551
rect 609 159 649 165
rect 609 135 617 159
rect 641 135 649 159
rect 609 129 649 135
rect 101 70 139 78
rect 101 50 110 70
rect 130 50 139 70
rect 101 41 139 50
rect 161 70 199 78
rect 161 50 170 70
rect 190 50 199 70
rect 161 41 199 50
rect 221 70 259 78
rect 221 50 230 70
rect 250 50 259 70
rect 221 41 259 50
rect 281 70 319 78
rect 281 50 290 70
rect 310 50 319 70
rect 281 41 319 50
rect 341 70 439 78
rect 341 50 350 70
rect 370 50 410 70
rect 430 50 439 70
rect 341 41 439 50
rect 461 70 499 78
rect 461 50 470 70
rect 490 50 499 70
rect 461 41 499 50
rect 521 70 559 78
rect 521 50 530 70
rect 550 50 559 70
rect 521 41 559 50
rect 616 0 649 129
<< viali >>
rect 110 610 130 630
rect 170 610 190 630
rect 230 610 250 630
rect 290 610 310 630
rect 350 610 370 630
rect 410 610 430 630
rect 470 610 490 630
rect 530 610 550 630
rect 113 554 137 578
rect 154 492 172 509
rect 154 451 172 468
rect 92 209 116 233
rect 285 509 309 513
rect 285 492 298 509
rect 298 492 309 509
rect 285 489 309 492
rect 286 468 310 470
rect 286 451 298 468
rect 298 451 310 468
rect 286 446 310 451
rect 510 509 534 514
rect 510 492 520 509
rect 520 492 534 509
rect 510 490 534 492
rect 510 468 534 471
rect 510 451 520 468
rect 520 451 534 468
rect 510 447 534 451
rect 214 359 238 383
rect 316 294 340 318
rect 476 293 500 317
rect 386 259 410 283
rect 290 209 314 233
rect 41 108 60 127
rect 211 104 235 128
rect 110 50 130 70
rect 170 50 190 70
rect 230 50 250 70
rect 290 50 310 70
rect 350 50 370 70
rect 410 50 430 70
rect 470 50 490 70
rect 530 50 550 70
<< metal1 >>
rect 0 630 680 660
rect 0 610 110 630
rect 130 610 170 630
rect 190 610 230 630
rect 250 610 290 630
rect 310 610 350 630
rect 370 610 410 630
rect 430 610 470 630
rect 490 610 530 630
rect 550 610 680 630
rect 0 600 680 610
rect 105 578 145 583
rect 105 572 113 578
rect 0 554 113 572
rect 137 572 145 578
rect 137 554 680 572
rect 0 551 680 554
rect 150 518 176 521
rect 150 468 176 492
rect 277 513 317 517
rect 277 489 285 513
rect 309 489 317 513
rect 277 484 317 489
rect 501 514 541 517
rect 501 490 510 514
rect 534 490 541 514
rect 501 484 541 490
rect 277 471 541 484
rect 277 470 510 471
rect 277 446 286 470
rect 310 446 317 470
rect 277 443 317 446
rect 501 447 510 470
rect 534 447 541 471
rect 501 443 541 447
rect 150 439 176 442
rect 0 383 680 389
rect 0 368 214 383
rect 206 359 214 368
rect 238 368 680 383
rect 238 359 246 368
rect 206 354 246 359
rect 0 318 680 327
rect 0 305 316 318
rect 308 294 316 305
rect 340 317 680 318
rect 340 305 476 317
rect 340 294 348 305
rect 308 288 348 294
rect 468 293 476 305
rect 500 305 680 317
rect 500 293 508 305
rect 468 288 508 293
rect 378 283 418 288
rect 378 274 386 283
rect 0 259 386 274
rect 410 274 418 283
rect 410 259 680 274
rect 0 253 680 259
rect 84 233 324 239
rect 84 209 92 233
rect 116 218 290 233
rect 116 209 125 218
rect 84 203 125 209
rect 282 209 290 218
rect 314 209 324 233
rect 282 203 324 209
rect 34 128 67 131
rect 202 128 243 135
rect 0 127 211 128
rect 0 108 41 127
rect 60 108 211 127
rect 0 107 211 108
rect 34 104 67 107
rect 202 104 211 107
rect 235 107 680 128
rect 235 104 243 107
rect 202 99 243 104
rect 0 70 680 80
rect 0 50 110 70
rect 130 50 170 70
rect 190 50 230 70
rect 250 50 290 70
rect 310 50 350 70
rect 370 50 410 70
rect 430 50 470 70
rect 490 50 530 70
rect 550 50 680 70
rect 0 17 680 50
<< via1 >>
rect 150 509 176 518
rect 150 492 154 509
rect 154 492 172 509
rect 172 492 176 509
rect 150 451 154 468
rect 154 451 172 468
rect 172 451 176 468
rect 150 442 176 451
<< metal2 >>
rect 147 518 179 535
rect 147 492 150 518
rect 176 492 179 518
rect 147 468 179 492
rect 147 442 150 468
rect 176 442 179 468
rect 147 439 179 442
<< labels >>
rlabel metal1 0 634 0 634 7 VDD
port 1 w
rlabel metal1 0 48 0 48 7 VSS
port 6 w
rlabel locali 634 0 634 0 5 ROW_N
port 7 s
rlabel metal1 0 561 0 561 7 SAMPLE_N
port 2 w
rlabel locali 375 542 375 542 1 VINT
port 10 n
rlabel metal1 0 378 0 378 7 SAMPLE
port 3 w
rlabel metal1 0 262 0 262 7 COL_N
port 5 w
rlabel metal1 0 116 0 116 7 VCOM
port 8 w
rlabel metal2 163 535 163 535 1 CBOT
port 9 n
rlabel metal1 0 316 0 316 7 COLON_N
port 4 w
rlabel locali 282 345 282 345 3 VDRV
port 12 e
rlabel locali 409 231 409 231 1 VINT2
port 11 n
<< end >>
