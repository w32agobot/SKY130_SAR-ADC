magic
tech sky130A
timestamp 1662910862
<< nwell >>
rect 117 474 521 661
<< nmos >>
rect 186 347 201 389
rect 234 347 249 389
rect 378 348 393 390
rect 426 348 441 390
<< pmos >>
rect 186 492 201 572
rect 234 492 249 572
rect 378 493 393 573
rect 426 493 441 573
<< ndiff >>
rect 155 383 186 389
rect 155 353 161 383
rect 178 353 186 383
rect 155 347 186 353
rect 201 383 234 389
rect 201 353 209 383
rect 226 353 234 383
rect 201 347 234 353
rect 249 383 280 389
rect 249 353 257 383
rect 274 353 280 383
rect 249 347 280 353
rect 347 384 378 390
rect 347 354 353 384
rect 370 354 378 384
rect 347 348 378 354
rect 393 384 426 390
rect 393 354 401 384
rect 418 354 426 384
rect 393 348 426 354
rect 441 384 472 390
rect 441 354 449 384
rect 466 354 472 384
rect 441 348 472 354
<< pdiff >>
rect 155 566 186 572
rect 155 498 161 566
rect 178 498 186 566
rect 155 492 186 498
rect 201 566 234 572
rect 201 498 209 566
rect 226 498 234 566
rect 201 492 234 498
rect 249 566 280 572
rect 249 498 257 566
rect 274 498 280 566
rect 249 492 280 498
rect 347 567 378 573
rect 347 499 353 567
rect 370 499 378 567
rect 347 493 378 499
rect 393 567 426 573
rect 393 499 401 567
rect 418 499 426 567
rect 393 493 426 499
rect 441 567 472 573
rect 441 499 449 567
rect 466 499 472 567
rect 441 493 472 499
<< ndiffc >>
rect 161 353 178 383
rect 209 353 226 383
rect 257 353 274 383
rect 353 354 370 384
rect 401 354 418 384
rect 449 354 466 384
<< pdiffc >>
rect 161 498 178 566
rect 209 498 226 566
rect 257 498 274 566
rect 353 499 370 567
rect 401 499 418 567
rect 449 499 466 567
<< psubdiff >>
rect 161 295 185 312
rect 202 295 233 312
rect 250 295 285 312
rect 302 295 337 312
rect 354 295 384 312
rect 401 295 433 312
rect 450 295 466 312
<< nsubdiff >>
rect 221 640 473 643
rect 221 623 233 640
rect 250 623 285 640
rect 302 623 337 640
rect 354 623 385 640
rect 402 623 432 640
rect 449 623 473 640
rect 221 620 473 623
<< psubdiffcont >>
rect 185 295 202 312
rect 233 295 250 312
rect 285 295 302 312
rect 337 295 354 312
rect 384 295 401 312
rect 433 295 450 312
<< nsubdiffcont >>
rect 233 623 250 640
rect 285 623 302 640
rect 337 623 354 640
rect 385 623 402 640
rect 432 623 449 640
<< poly >>
rect 176 630 210 635
rect 176 612 184 630
rect 202 612 210 630
rect 176 595 210 612
rect 176 580 249 595
rect 186 572 201 580
rect 234 572 249 580
rect 378 573 393 586
rect 426 573 441 586
rect 186 389 201 492
rect 234 389 249 492
rect 378 436 393 493
rect 275 435 393 436
rect 426 435 441 493
rect 275 430 441 435
rect 275 413 283 430
rect 300 421 441 430
rect 300 413 319 421
rect 275 408 319 413
rect 378 408 441 421
rect 378 390 393 408
rect 426 390 441 408
rect 186 334 201 347
rect 234 334 249 347
rect 378 335 393 348
rect 426 335 441 348
rect 487 331 514 339
rect 487 314 492 331
rect 509 314 514 331
rect 487 306 514 314
<< polycont >>
rect 184 612 202 630
rect 283 413 300 430
rect 492 314 509 331
<< locali >>
rect 127 354 144 664
rect 221 640 473 643
rect 184 630 202 638
rect 221 623 233 640
rect 250 623 285 640
rect 302 623 337 640
rect 354 623 385 640
rect 402 623 432 640
rect 449 623 473 640
rect 221 620 473 623
rect 184 607 202 612
rect 184 590 185 607
rect 161 566 178 574
rect 161 490 178 498
rect 209 566 226 574
rect 127 285 144 337
rect 161 383 178 391
rect 161 312 178 353
rect 209 385 226 498
rect 257 566 274 620
rect 257 490 274 498
rect 353 567 370 620
rect 353 491 370 499
rect 401 567 418 575
rect 248 430 308 431
rect 248 425 283 430
rect 267 413 283 425
rect 300 413 308 430
rect 267 408 308 413
rect 209 345 226 353
rect 257 383 274 391
rect 257 312 274 353
rect 353 384 370 392
rect 353 312 370 354
rect 401 384 418 499
rect 449 567 466 620
rect 449 491 466 499
rect 401 346 418 354
rect 449 384 466 392
rect 449 312 466 354
rect 497 339 514 664
rect 161 295 185 312
rect 202 295 233 312
rect 250 295 285 312
rect 302 295 337 312
rect 354 295 384 312
rect 401 295 433 312
rect 450 295 466 312
rect 490 331 514 339
rect 490 314 492 331
rect 509 314 514 331
rect 490 306 514 314
rect 497 285 514 306
<< viali >>
rect 233 623 250 640
rect 285 623 302 640
rect 337 623 354 640
rect 385 623 402 640
rect 432 623 449 640
rect 185 590 202 607
rect 161 519 178 542
rect 127 337 144 354
rect 257 521 274 544
rect 401 521 418 556
rect 248 408 267 425
rect 209 383 226 385
rect 209 365 226 383
rect 185 295 202 312
rect 233 295 250 312
rect 285 295 302 312
rect 337 295 354 312
rect 384 295 401 312
rect 433 295 450 312
<< metal1 >>
rect 117 640 521 648
rect 117 624 233 640
rect 117 620 168 624
rect 219 623 233 624
rect 250 623 285 640
rect 302 623 337 640
rect 354 623 385 640
rect 402 623 432 640
rect 449 623 521 640
rect 219 620 521 623
rect 179 607 208 610
rect 179 606 185 607
rect 117 591 185 606
rect 179 590 185 591
rect 202 590 208 607
rect 179 587 208 590
rect 401 591 521 606
rect 401 563 418 591
rect 397 556 421 563
rect 155 544 280 548
rect 155 542 257 544
rect 155 519 161 542
rect 178 521 257 542
rect 274 521 280 544
rect 178 519 280 521
rect 155 516 280 519
rect 397 521 401 556
rect 418 521 421 556
rect 397 508 421 521
rect 117 477 521 491
rect 148 450 491 463
rect 117 449 521 450
rect 117 436 167 449
rect 474 436 521 449
rect 242 425 273 429
rect 242 422 248 425
rect 117 408 248 422
rect 267 408 273 425
rect 242 403 273 408
rect 314 408 521 422
rect 205 385 229 393
rect 205 365 209 385
rect 226 377 229 385
rect 314 377 329 408
rect 226 365 329 377
rect 205 361 329 365
rect 124 354 147 360
rect 205 359 229 361
rect 124 345 127 354
rect 117 337 127 345
rect 144 345 147 354
rect 144 337 521 345
rect 117 331 521 337
rect 117 312 521 317
rect 117 295 185 312
rect 202 295 233 312
rect 250 295 285 312
rect 302 295 337 312
rect 354 295 384 312
rect 401 295 433 312
rect 450 295 521 312
rect 117 289 521 295
<< labels >>
rlabel metal1 117 436 117 450 7 col_n
port 6 w
rlabel metal1 117 477 117 491 7 colon_n
port 7 w
rlabel metal1 117 331 117 345 7 vcom
port 3 w
rlabel metal1 117 289 117 317 7 VSS
port 2 w
rlabel metal1 117 620 117 648 7 VDD
port 1 w
rlabel locali 497 285 514 285 5 row_n
port 8 s
rlabel metal1 117 591 117 606 3 sample_n_in
port 9 e
rlabel metal1 117 408 117 422 3 sample_in
port 10 e
rlabel metal1 521 408 521 422 7 sample_out
port 11 w
rlabel metal1 521 591 521 606 7 sample_n_out
port 12 w
<< end >>
