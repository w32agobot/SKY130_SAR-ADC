* SPICE3 file created from adc_array_wafflecap_16(4)x296aF_28um2.ext - technology: sky130A

.subckt adc_array_wafflecap_16(4)x296aF_28um2 cbot ctop
C0 cfloating cbot 3.51fF
C1 ctop cbot 1.18fF
C2 cfloating ctop 0.43fF
C3 cbot VSUBS 2.16fF
C4 cfloating VSUBS 0.56fF
.ends
