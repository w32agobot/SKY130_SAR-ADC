magic
tech sky130A
timestamp 1667056780
<< nwell >>
rect 3065 6600 3124 6804
rect 1446 6361 1628 6406
rect 1423 6349 1628 6361
rect 1423 6220 1451 6349
rect 1506 6294 1628 6349
rect 1500 6275 1628 6294
rect 1506 6220 1628 6275
rect 1423 6207 1628 6220
rect 3064 6028 3204 6230
<< poly >>
rect 3119 6556 3135 6570
rect 3119 6474 3134 6556
rect 3119 6465 3156 6474
rect 3119 6448 3134 6465
rect 3151 6448 3156 6465
rect 3119 6440 3156 6448
rect 2318 6062 2357 6067
rect 2318 6045 2326 6062
rect 2343 6045 2357 6062
rect 2318 6040 2357 6045
<< polycont >>
rect 3134 6448 3151 6465
rect 1418 6187 1435 6204
rect 2326 6045 2343 6062
<< locali >>
rect 1570 6740 1678 6743
rect 1570 6722 1576 6740
rect 1593 6722 1615 6740
rect 1632 6722 1651 6740
rect 1668 6722 1678 6740
rect 1570 6719 1678 6722
rect 1570 6406 1613 6719
rect 3550 6570 3617 6573
rect 3550 6552 3556 6570
rect 3574 6552 3593 6570
rect 3611 6552 3617 6570
rect 3550 6549 3617 6552
rect 1454 6386 1613 6406
rect 3130 6465 3154 6473
rect 3130 6448 3134 6465
rect 3151 6448 3154 6465
rect 3183 6448 3733 6474
rect 1523 6294 1545 6386
rect 1523 6275 1569 6294
rect 3130 6282 3154 6448
rect 3130 6264 3133 6282
rect 3151 6264 3154 6282
rect 1410 6204 1437 6212
rect 1410 6187 1418 6204
rect 1435 6187 1437 6204
rect 1410 6179 1437 6187
rect 1527 6204 1554 6212
rect 1527 6187 1535 6204
rect 1552 6187 1554 6204
rect 1527 6179 1554 6187
rect 3130 6106 3154 6264
rect 3171 6420 3195 6426
rect 3171 6402 3174 6420
rect 3192 6402 3195 6420
rect 3171 6252 3195 6402
rect 3264 6365 3307 6448
rect 3437 6275 3537 6278
rect 3437 6259 3475 6275
rect 3469 6257 3475 6259
rect 3493 6257 3513 6275
rect 3531 6257 3537 6275
rect 3469 6254 3537 6257
rect 3171 6234 3174 6252
rect 3192 6234 3195 6252
rect 3171 6228 3195 6234
rect 3130 6080 3259 6106
rect 2318 6062 2357 6067
rect 2318 6045 2326 6062
rect 2343 6045 2357 6062
rect 3081 6046 3249 6063
rect 2318 6040 2357 6045
<< viali >>
rect 1576 6722 1593 6740
rect 1615 6722 1632 6740
rect 1651 6722 1668 6740
rect 3556 6552 3574 6570
rect 3593 6552 3611 6570
rect 3133 6264 3151 6282
rect 1418 6187 1435 6204
rect 1535 6187 1552 6204
rect 3174 6402 3192 6420
rect 3475 6257 3493 6275
rect 3513 6257 3531 6275
rect 3174 6234 3192 6252
rect 2326 6045 2343 6062
rect 2365 6045 2382 6062
<< metal1 >>
rect 1000 6770 1014 6885
rect 1570 6740 1678 6770
rect 1570 6722 1576 6740
rect 1593 6722 1615 6740
rect 1632 6722 1651 6740
rect 1668 6722 1678 6740
rect 1570 6719 1678 6722
rect 3060 6738 3121 6755
rect 1000 6541 1007 6555
rect 1000 6513 1007 6527
rect 3060 6426 3078 6738
rect 3607 6588 4005 6602
rect 3550 6570 3617 6573
rect 3550 6552 3556 6570
rect 3574 6552 3593 6570
rect 3611 6568 3617 6570
rect 3611 6554 4005 6568
rect 3611 6552 3617 6554
rect 3550 6549 3617 6552
rect 3060 6420 3195 6426
rect 3060 6407 3174 6420
rect 3171 6402 3174 6407
rect 3192 6402 3195 6420
rect 3171 6396 3195 6402
rect 3130 6282 3154 6288
rect 3130 6277 3133 6282
rect 3032 6264 3133 6277
rect 3151 6264 3154 6282
rect 3032 6258 3154 6264
rect 3469 6275 3537 6278
rect 3171 6252 3195 6258
rect 3469 6257 3475 6275
rect 3493 6257 3513 6275
rect 3531 6273 3537 6275
rect 3531 6259 4005 6273
rect 3531 6257 3537 6259
rect 3469 6254 3537 6257
rect 3171 6234 3174 6252
rect 3192 6245 3195 6252
rect 3192 6234 3220 6245
rect 3171 6226 3220 6234
rect 1407 6204 1438 6212
rect 1407 6203 1418 6204
rect 1000 6189 1418 6203
rect 1407 6187 1418 6189
rect 1435 6187 1438 6204
rect 1407 6179 1438 6187
rect 1527 6204 1555 6212
rect 1527 6187 1535 6204
rect 1552 6195 1555 6204
rect 1552 6187 1657 6195
rect 1527 6179 1657 6187
rect 1000 5910 1011 6026
rect 1393 6025 1621 6078
rect 1636 6067 1657 6179
rect 1636 6062 2390 6067
rect 1636 6045 2326 6062
rect 2343 6045 2365 6062
rect 2382 6045 2390 6062
rect 1636 6040 2390 6045
use adc_comp_circuit  adc_comp_circuit_0
timestamp 1665574574
transform 1 0 1637 0 1 6689
box -637 -1689 2355 1109
use adc_inverter  adc_inverter_0
timestamp 1664803391
transform 1 0 1423 0 1 6118
box -13 -65 104 291
use adc_inverter  adc_inverter_1
timestamp 1664803391
transform 1 0 1540 0 1 6118
box -13 -65 104 291
use adc_nor  adc_nor_0
timestamp 1661513809
transform 1 0 3208 0 -1 6258
box -4 -118 253 230
use adc_nor_latch  adc_nor_latch_0
timestamp 1661515501
transform 1 0 3124 0 1 6456
box -3 0 505 348
<< labels >>
flabel metal1 s 3924 6259 4005 6273 3 FreeSans 80 0 0 0 comp_trig
port 6 e signal output
flabel metal1 s 1000 6189 1007 6203 7 FreeSans 80 0 0 0 clk
port 3 w signal input
flabel metal1 s 3924 6554 4005 6568 3 FreeSans 80 0 0 0 latch_qn
port 7 e signal output
flabel metal1 s 3924 6588 4005 6602 3 FreeSans 80 0 0 0 latch_q
port 8 e signal output
flabel metal1 s 1000 5910 1011 6026 7 FreeSans 80 0 0 0 VGND
port 2 w ground bidirectional
flabel metal1 s 1000 6770 1014 6885 7 FreeSans 80 0 0 0 VPWR
port 1 w power bidirectional
flabel metal1 s 1000 6541 1007 6555 7 FreeSans 80 0 0 0 inp
port 4 w signal input
flabel metal1 s 1000 6513 1007 6527 7 FreeSans 80 0 0 0 inn
port 5 w signal input
<< properties >>
string FIXED_BBOX 0 0 4200 12900
string LEFclass BLOCK
string LEForigin 0 0
string LEFsource USER
<< end >>
