magic
tech sky130A
magscale 1 2
timestamp 1664545144
<< nwell >>
rect -224 -36 223 138
<< pmos >>
rect -129 0 -29 100
rect 29 0 129 100
<< pdiff >>
rect -187 88 -129 100
rect -187 12 -175 88
rect -141 12 -129 88
rect -187 0 -129 12
rect -29 88 29 100
rect -29 12 -17 88
rect 17 12 29 88
rect -29 0 29 12
rect 129 88 187 100
rect 129 12 141 88
rect 175 12 187 88
rect 129 0 187 12
<< pdiffc >>
rect -175 12 -141 88
rect -17 12 17 88
rect 141 12 175 88
<< poly >>
rect -129 100 -29 126
rect 29 100 129 126
rect -129 -26 -29 0
rect 29 -26 129 0
<< locali >>
rect -175 88 -141 104
rect -175 -4 -141 12
rect -17 88 17 104
rect -17 -4 17 12
rect 141 88 175 104
rect 141 -4 175 12
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 1 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
