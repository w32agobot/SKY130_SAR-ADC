VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO adc_vcm_generator
  CLASS BLOCK ;
  FOREIGN adc_vcm_generator ;
  ORIGIN 0.000 0.000 ;
  SIZE 131.850 BY 340.000 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 6.910 174.150 7.750 174.155 ;
        RECT 12.155 174.150 14.705 174.155 ;
        RECT 6.395 172.925 23.795 174.150 ;
        RECT 6.395 171.320 24.255 172.925 ;
        RECT 6.395 167.105 24.255 168.710 ;
        RECT 7.315 165.885 23.795 167.105 ;
        RECT 7.315 165.880 9.625 165.885 ;
        RECT 14.675 165.880 23.795 165.885 ;
      LAYER li1 ;
        RECT 43.835 174.260 47.835 174.460 ;
        RECT 7.185 172.825 7.475 173.990 ;
        RECT 7.100 172.655 7.560 172.825 ;
        RECT 14.950 172.820 15.240 173.985 ;
        RECT 15.560 172.820 15.890 173.970 ;
        RECT 16.400 172.820 16.730 173.620 ;
        RECT 17.250 172.820 17.490 173.620 ;
        RECT 18.320 172.820 18.650 173.970 ;
        RECT 19.160 172.820 19.490 173.620 ;
        RECT 20.010 172.820 20.250 173.620 ;
        RECT 21.675 172.820 21.885 173.960 ;
        RECT 23.055 172.820 23.265 173.960 ;
        RECT 43.835 173.660 44.235 174.260 ;
        RECT 43.835 173.460 47.835 173.660 ;
        RECT 43.835 172.860 44.235 173.460 ;
        RECT 7.965 172.650 24.065 172.820 ;
        RECT 43.835 172.660 47.835 172.860 ;
        RECT 8.050 171.485 8.340 172.650 ;
        RECT 8.510 171.510 8.770 172.650 ;
        RECT 9.440 171.510 9.720 172.650 ;
        RECT 10.500 172.225 10.885 172.650 ;
        RECT 11.915 172.225 12.300 172.650 ;
        RECT 13.330 172.225 13.715 172.650 ;
        RECT 15.100 172.225 15.485 172.650 ;
        RECT 16.515 172.225 16.900 172.650 ;
        RECT 17.930 172.225 18.315 172.650 ;
        RECT 19.700 172.225 20.085 172.650 ;
        RECT 21.115 172.225 21.500 172.650 ;
        RECT 22.530 172.225 22.915 172.650 ;
        RECT 23.690 171.485 23.980 172.650 ;
        RECT 43.835 172.060 44.235 172.660 ;
        RECT 43.835 171.860 47.835 172.060 ;
        RECT 43.835 171.260 44.235 171.860 ;
        RECT 43.835 171.060 47.835 171.260 ;
        RECT 43.835 170.460 44.235 171.060 ;
        RECT 43.835 170.260 47.835 170.460 ;
        RECT 43.835 169.660 44.235 170.260 ;
        RECT 43.835 169.460 47.835 169.660 ;
        RECT 43.835 168.860 44.235 169.460 ;
        RECT 43.835 168.660 47.835 168.860 ;
        RECT 6.670 167.380 6.960 168.545 ;
        RECT 7.385 167.380 7.595 168.520 ;
        RECT 8.510 167.380 8.790 168.520 ;
        RECT 9.460 167.380 9.720 168.520 ;
        RECT 10.500 167.380 10.885 167.805 ;
        RECT 11.915 167.380 12.300 167.805 ;
        RECT 13.330 167.380 13.715 167.805 ;
        RECT 15.100 167.380 15.485 167.805 ;
        RECT 16.515 167.380 16.900 167.805 ;
        RECT 17.930 167.380 18.315 167.805 ;
        RECT 19.700 167.380 20.085 167.805 ;
        RECT 21.115 167.380 21.500 167.805 ;
        RECT 22.530 167.380 22.915 167.805 ;
        RECT 23.690 167.380 23.980 168.545 ;
        RECT 43.835 168.060 44.235 168.660 ;
        RECT 43.835 167.860 47.835 168.060 ;
        RECT 6.585 167.210 24.065 167.380 ;
        RECT 43.835 167.260 44.235 167.860 ;
        RECT 7.590 166.045 7.880 167.210 ;
        RECT 10.570 166.560 10.745 167.210 ;
        RECT 10.575 164.605 10.745 166.560 ;
        RECT 14.950 166.045 15.240 167.210 ;
        RECT 15.560 166.060 15.890 167.210 ;
        RECT 16.400 166.410 16.730 167.210 ;
        RECT 17.250 166.410 17.490 167.210 ;
        RECT 18.320 166.060 18.650 167.210 ;
        RECT 19.160 166.410 19.490 167.210 ;
        RECT 20.010 166.410 20.250 167.210 ;
        RECT 21.675 166.070 21.885 167.210 ;
        RECT 23.055 166.070 23.265 167.210 ;
        RECT 43.835 167.060 47.835 167.260 ;
        RECT 43.835 166.860 44.235 167.060 ;
        RECT 48.585 166.860 48.785 174.460 ;
        RECT 49.385 166.860 49.585 174.460 ;
        RECT 50.185 166.860 50.385 174.460 ;
        RECT 50.985 166.860 51.185 174.460 ;
        RECT 51.785 166.860 51.985 174.460 ;
        RECT 43.835 166.460 51.985 166.860 ;
        RECT 43.835 166.260 44.235 166.460 ;
        RECT 43.835 166.060 47.835 166.260 ;
        RECT 43.835 165.460 44.235 166.060 ;
        RECT 43.835 165.260 47.835 165.460 ;
        RECT 43.835 164.660 44.235 165.260 ;
        RECT 43.835 164.460 47.835 164.660 ;
        RECT 43.835 163.860 44.235 164.460 ;
        RECT 43.835 163.660 47.835 163.860 ;
        RECT 43.835 163.060 44.235 163.660 ;
        RECT 43.835 162.860 47.835 163.060 ;
        RECT 43.835 162.260 44.235 162.860 ;
        RECT 43.835 162.060 47.835 162.260 ;
        RECT 43.835 161.460 44.235 162.060 ;
        RECT 43.835 161.260 47.835 161.460 ;
        RECT 43.835 160.660 44.235 161.260 ;
        RECT 43.835 160.460 47.835 160.660 ;
        RECT 43.835 159.860 44.235 160.460 ;
        RECT 43.835 159.660 47.835 159.860 ;
        RECT 43.835 159.060 44.235 159.660 ;
        RECT 43.835 158.860 47.835 159.060 ;
        RECT 48.585 158.860 48.785 166.460 ;
        RECT 49.385 158.860 49.585 166.460 ;
        RECT 50.185 158.860 50.385 166.460 ;
        RECT 50.985 158.860 51.185 166.460 ;
        RECT 51.785 158.860 51.985 166.460 ;
        RECT 53.285 166.860 53.485 174.460 ;
        RECT 54.085 166.860 54.285 174.460 ;
        RECT 54.885 166.860 55.085 174.460 ;
        RECT 55.685 166.860 55.885 174.460 ;
        RECT 56.485 166.860 56.685 174.460 ;
        RECT 57.435 174.260 61.435 174.460 ;
        RECT 61.035 173.660 61.435 174.260 ;
        RECT 57.435 173.460 61.435 173.660 ;
        RECT 61.035 172.860 61.435 173.460 ;
        RECT 57.435 172.660 61.435 172.860 ;
        RECT 61.035 172.060 61.435 172.660 ;
        RECT 57.435 171.860 61.435 172.060 ;
        RECT 61.035 171.260 61.435 171.860 ;
        RECT 57.435 171.060 61.435 171.260 ;
        RECT 61.035 170.460 61.435 171.060 ;
        RECT 57.435 170.260 61.435 170.460 ;
        RECT 61.035 169.660 61.435 170.260 ;
        RECT 57.435 169.460 61.435 169.660 ;
        RECT 61.035 168.860 61.435 169.460 ;
        RECT 57.435 168.660 61.435 168.860 ;
        RECT 61.035 168.060 61.435 168.660 ;
        RECT 57.435 167.860 61.435 168.060 ;
        RECT 61.035 167.260 61.435 167.860 ;
        RECT 57.435 167.060 61.435 167.260 ;
        RECT 61.035 166.860 61.435 167.060 ;
        RECT 53.285 166.460 61.435 166.860 ;
        RECT 53.285 158.860 53.485 166.460 ;
        RECT 54.085 158.860 54.285 166.460 ;
        RECT 54.885 158.860 55.085 166.460 ;
        RECT 55.685 158.860 55.885 166.460 ;
        RECT 56.485 158.860 56.685 166.460 ;
        RECT 61.035 166.260 61.435 166.460 ;
        RECT 57.435 166.060 61.435 166.260 ;
        RECT 61.035 165.460 61.435 166.060 ;
        RECT 57.435 165.260 61.435 165.460 ;
        RECT 61.035 164.660 61.435 165.260 ;
        RECT 57.435 164.460 61.435 164.660 ;
        RECT 61.035 163.860 61.435 164.460 ;
        RECT 57.435 163.660 61.435 163.860 ;
        RECT 61.035 163.060 61.435 163.660 ;
        RECT 57.435 162.860 61.435 163.060 ;
        RECT 61.035 162.260 61.435 162.860 ;
        RECT 57.435 162.060 61.435 162.260 ;
        RECT 61.035 161.460 61.435 162.060 ;
        RECT 57.435 161.260 61.435 161.460 ;
        RECT 61.035 160.660 61.435 161.260 ;
        RECT 57.435 160.460 61.435 160.660 ;
        RECT 61.035 159.860 61.435 160.460 ;
        RECT 57.435 159.660 61.435 159.860 ;
        RECT 61.035 159.060 61.435 159.660 ;
        RECT 57.435 158.860 61.435 159.060 ;
        RECT 63.835 174.260 67.835 174.460 ;
        RECT 63.835 173.660 64.235 174.260 ;
        RECT 63.835 173.460 67.835 173.660 ;
        RECT 63.835 172.860 64.235 173.460 ;
        RECT 63.835 172.660 67.835 172.860 ;
        RECT 63.835 172.060 64.235 172.660 ;
        RECT 63.835 171.860 67.835 172.060 ;
        RECT 63.835 171.260 64.235 171.860 ;
        RECT 63.835 171.060 67.835 171.260 ;
        RECT 63.835 170.460 64.235 171.060 ;
        RECT 63.835 170.260 67.835 170.460 ;
        RECT 63.835 169.660 64.235 170.260 ;
        RECT 63.835 169.460 67.835 169.660 ;
        RECT 63.835 168.860 64.235 169.460 ;
        RECT 63.835 168.660 67.835 168.860 ;
        RECT 63.835 168.060 64.235 168.660 ;
        RECT 63.835 167.860 67.835 168.060 ;
        RECT 63.835 167.260 64.235 167.860 ;
        RECT 63.835 167.060 67.835 167.260 ;
        RECT 63.835 166.860 64.235 167.060 ;
        RECT 68.585 166.860 68.785 174.460 ;
        RECT 69.385 166.860 69.585 174.460 ;
        RECT 70.185 166.860 70.385 174.460 ;
        RECT 70.985 166.860 71.185 174.460 ;
        RECT 71.785 166.860 71.985 174.460 ;
        RECT 63.835 166.460 71.985 166.860 ;
        RECT 63.835 166.260 64.235 166.460 ;
        RECT 63.835 166.060 67.835 166.260 ;
        RECT 63.835 165.460 64.235 166.060 ;
        RECT 63.835 165.260 67.835 165.460 ;
        RECT 63.835 164.660 64.235 165.260 ;
        RECT 63.835 164.460 67.835 164.660 ;
        RECT 63.835 163.860 64.235 164.460 ;
        RECT 63.835 163.660 67.835 163.860 ;
        RECT 63.835 163.060 64.235 163.660 ;
        RECT 63.835 162.860 67.835 163.060 ;
        RECT 63.835 162.260 64.235 162.860 ;
        RECT 63.835 162.060 67.835 162.260 ;
        RECT 63.835 161.460 64.235 162.060 ;
        RECT 63.835 161.260 67.835 161.460 ;
        RECT 63.835 160.660 64.235 161.260 ;
        RECT 63.835 160.460 67.835 160.660 ;
        RECT 63.835 159.860 64.235 160.460 ;
        RECT 63.835 159.660 67.835 159.860 ;
        RECT 63.835 159.060 64.235 159.660 ;
        RECT 63.835 158.860 67.835 159.060 ;
        RECT 68.585 158.860 68.785 166.460 ;
        RECT 69.385 158.860 69.585 166.460 ;
        RECT 70.185 158.860 70.385 166.460 ;
        RECT 70.985 158.860 71.185 166.460 ;
        RECT 71.785 158.860 71.985 166.460 ;
        RECT 73.285 166.860 73.485 174.460 ;
        RECT 74.085 166.860 74.285 174.460 ;
        RECT 74.885 166.860 75.085 174.460 ;
        RECT 75.685 166.860 75.885 174.460 ;
        RECT 76.485 166.860 76.685 174.460 ;
        RECT 77.435 174.260 81.435 174.460 ;
        RECT 81.035 173.660 81.435 174.260 ;
        RECT 77.435 173.460 81.435 173.660 ;
        RECT 81.035 172.860 81.435 173.460 ;
        RECT 77.435 172.660 81.435 172.860 ;
        RECT 81.035 172.060 81.435 172.660 ;
        RECT 77.435 171.860 81.435 172.060 ;
        RECT 81.035 171.260 81.435 171.860 ;
        RECT 77.435 171.060 81.435 171.260 ;
        RECT 81.035 170.460 81.435 171.060 ;
        RECT 77.435 170.260 81.435 170.460 ;
        RECT 81.035 169.660 81.435 170.260 ;
        RECT 77.435 169.460 81.435 169.660 ;
        RECT 81.035 168.860 81.435 169.460 ;
        RECT 77.435 168.660 81.435 168.860 ;
        RECT 81.035 168.060 81.435 168.660 ;
        RECT 77.435 167.860 81.435 168.060 ;
        RECT 81.035 167.260 81.435 167.860 ;
        RECT 77.435 167.060 81.435 167.260 ;
        RECT 81.035 166.860 81.435 167.060 ;
        RECT 73.285 166.460 81.435 166.860 ;
        RECT 73.285 158.860 73.485 166.460 ;
        RECT 74.085 158.860 74.285 166.460 ;
        RECT 74.885 158.860 75.085 166.460 ;
        RECT 75.685 158.860 75.885 166.460 ;
        RECT 76.485 158.860 76.685 166.460 ;
        RECT 81.035 166.260 81.435 166.460 ;
        RECT 77.435 166.060 81.435 166.260 ;
        RECT 81.035 165.460 81.435 166.060 ;
        RECT 77.435 165.260 81.435 165.460 ;
        RECT 81.035 164.660 81.435 165.260 ;
        RECT 77.435 164.460 81.435 164.660 ;
        RECT 81.035 163.860 81.435 164.460 ;
        RECT 77.435 163.660 81.435 163.860 ;
        RECT 81.035 163.060 81.435 163.660 ;
        RECT 77.435 162.860 81.435 163.060 ;
        RECT 81.035 162.260 81.435 162.860 ;
        RECT 77.435 162.060 81.435 162.260 ;
        RECT 81.035 161.460 81.435 162.060 ;
        RECT 77.435 161.260 81.435 161.460 ;
        RECT 81.035 160.660 81.435 161.260 ;
        RECT 77.435 160.460 81.435 160.660 ;
        RECT 81.035 159.860 81.435 160.460 ;
        RECT 77.435 159.660 81.435 159.860 ;
        RECT 81.035 159.060 81.435 159.660 ;
        RECT 77.435 158.860 81.435 159.060 ;
        RECT 83.835 174.260 87.835 174.460 ;
        RECT 83.835 173.660 84.235 174.260 ;
        RECT 83.835 173.460 87.835 173.660 ;
        RECT 83.835 172.860 84.235 173.460 ;
        RECT 83.835 172.660 87.835 172.860 ;
        RECT 83.835 172.060 84.235 172.660 ;
        RECT 83.835 171.860 87.835 172.060 ;
        RECT 83.835 171.260 84.235 171.860 ;
        RECT 83.835 171.060 87.835 171.260 ;
        RECT 83.835 170.460 84.235 171.060 ;
        RECT 83.835 170.260 87.835 170.460 ;
        RECT 83.835 169.660 84.235 170.260 ;
        RECT 83.835 169.460 87.835 169.660 ;
        RECT 83.835 168.860 84.235 169.460 ;
        RECT 83.835 168.660 87.835 168.860 ;
        RECT 83.835 168.060 84.235 168.660 ;
        RECT 83.835 167.860 87.835 168.060 ;
        RECT 83.835 167.260 84.235 167.860 ;
        RECT 83.835 167.060 87.835 167.260 ;
        RECT 83.835 166.860 84.235 167.060 ;
        RECT 88.585 166.860 88.785 174.460 ;
        RECT 89.385 166.860 89.585 174.460 ;
        RECT 90.185 166.860 90.385 174.460 ;
        RECT 90.985 166.860 91.185 174.460 ;
        RECT 91.785 166.860 91.985 174.460 ;
        RECT 83.835 166.460 91.985 166.860 ;
        RECT 83.835 166.260 84.235 166.460 ;
        RECT 83.835 166.060 87.835 166.260 ;
        RECT 83.835 165.460 84.235 166.060 ;
        RECT 83.835 165.260 87.835 165.460 ;
        RECT 83.835 164.660 84.235 165.260 ;
        RECT 83.835 164.460 87.835 164.660 ;
        RECT 83.835 163.860 84.235 164.460 ;
        RECT 83.835 163.660 87.835 163.860 ;
        RECT 83.835 163.060 84.235 163.660 ;
        RECT 83.835 162.860 87.835 163.060 ;
        RECT 83.835 162.260 84.235 162.860 ;
        RECT 83.835 162.060 87.835 162.260 ;
        RECT 83.835 161.460 84.235 162.060 ;
        RECT 83.835 161.260 87.835 161.460 ;
        RECT 83.835 160.660 84.235 161.260 ;
        RECT 83.835 160.460 87.835 160.660 ;
        RECT 83.835 159.860 84.235 160.460 ;
        RECT 83.835 159.660 87.835 159.860 ;
        RECT 83.835 159.060 84.235 159.660 ;
        RECT 83.835 158.860 87.835 159.060 ;
        RECT 88.585 158.860 88.785 166.460 ;
        RECT 89.385 158.860 89.585 166.460 ;
        RECT 90.185 158.860 90.385 166.460 ;
        RECT 90.985 158.860 91.185 166.460 ;
        RECT 91.785 158.860 91.985 166.460 ;
        RECT 93.285 166.860 93.485 174.460 ;
        RECT 94.085 166.860 94.285 174.460 ;
        RECT 94.885 166.860 95.085 174.460 ;
        RECT 95.685 166.860 95.885 174.460 ;
        RECT 96.485 166.860 96.685 174.460 ;
        RECT 97.435 174.260 101.435 174.460 ;
        RECT 101.035 173.660 101.435 174.260 ;
        RECT 97.435 173.460 101.435 173.660 ;
        RECT 101.035 172.860 101.435 173.460 ;
        RECT 97.435 172.660 101.435 172.860 ;
        RECT 101.035 172.060 101.435 172.660 ;
        RECT 97.435 171.860 101.435 172.060 ;
        RECT 101.035 171.260 101.435 171.860 ;
        RECT 97.435 171.060 101.435 171.260 ;
        RECT 101.035 170.460 101.435 171.060 ;
        RECT 97.435 170.260 101.435 170.460 ;
        RECT 101.035 169.660 101.435 170.260 ;
        RECT 97.435 169.460 101.435 169.660 ;
        RECT 101.035 168.860 101.435 169.460 ;
        RECT 97.435 168.660 101.435 168.860 ;
        RECT 101.035 168.060 101.435 168.660 ;
        RECT 97.435 167.860 101.435 168.060 ;
        RECT 101.035 167.260 101.435 167.860 ;
        RECT 97.435 167.060 101.435 167.260 ;
        RECT 101.035 166.860 101.435 167.060 ;
        RECT 93.285 166.460 101.435 166.860 ;
        RECT 93.285 158.860 93.485 166.460 ;
        RECT 94.085 158.860 94.285 166.460 ;
        RECT 94.885 158.860 95.085 166.460 ;
        RECT 95.685 158.860 95.885 166.460 ;
        RECT 96.485 158.860 96.685 166.460 ;
        RECT 101.035 166.260 101.435 166.460 ;
        RECT 97.435 166.060 101.435 166.260 ;
        RECT 101.035 165.460 101.435 166.060 ;
        RECT 97.435 165.260 101.435 165.460 ;
        RECT 101.035 164.660 101.435 165.260 ;
        RECT 97.435 164.460 101.435 164.660 ;
        RECT 101.035 163.860 101.435 164.460 ;
        RECT 97.435 163.660 101.435 163.860 ;
        RECT 101.035 163.060 101.435 163.660 ;
        RECT 97.435 162.860 101.435 163.060 ;
        RECT 101.035 162.260 101.435 162.860 ;
        RECT 97.435 162.060 101.435 162.260 ;
        RECT 101.035 161.460 101.435 162.060 ;
        RECT 97.435 161.260 101.435 161.460 ;
        RECT 101.035 160.660 101.435 161.260 ;
        RECT 97.435 160.460 101.435 160.660 ;
        RECT 101.035 159.860 101.435 160.460 ;
        RECT 97.435 159.660 101.435 159.860 ;
        RECT 101.035 159.060 101.435 159.660 ;
        RECT 97.435 158.860 101.435 159.060 ;
        RECT 103.835 174.260 107.835 174.460 ;
        RECT 103.835 173.660 104.235 174.260 ;
        RECT 103.835 173.460 107.835 173.660 ;
        RECT 103.835 172.860 104.235 173.460 ;
        RECT 103.835 172.660 107.835 172.860 ;
        RECT 103.835 172.060 104.235 172.660 ;
        RECT 103.835 171.860 107.835 172.060 ;
        RECT 103.835 171.260 104.235 171.860 ;
        RECT 103.835 171.060 107.835 171.260 ;
        RECT 103.835 170.460 104.235 171.060 ;
        RECT 103.835 170.260 107.835 170.460 ;
        RECT 103.835 169.660 104.235 170.260 ;
        RECT 103.835 169.460 107.835 169.660 ;
        RECT 103.835 168.860 104.235 169.460 ;
        RECT 103.835 168.660 107.835 168.860 ;
        RECT 103.835 168.060 104.235 168.660 ;
        RECT 103.835 167.860 107.835 168.060 ;
        RECT 103.835 167.260 104.235 167.860 ;
        RECT 103.835 167.060 107.835 167.260 ;
        RECT 103.835 166.860 104.235 167.060 ;
        RECT 108.585 166.860 108.785 174.460 ;
        RECT 109.385 166.860 109.585 174.460 ;
        RECT 110.185 166.860 110.385 174.460 ;
        RECT 110.985 166.860 111.185 174.460 ;
        RECT 111.785 166.860 111.985 174.460 ;
        RECT 103.835 166.460 111.985 166.860 ;
        RECT 103.835 166.260 104.235 166.460 ;
        RECT 103.835 166.060 107.835 166.260 ;
        RECT 103.835 165.460 104.235 166.060 ;
        RECT 103.835 165.260 107.835 165.460 ;
        RECT 103.835 164.660 104.235 165.260 ;
        RECT 103.835 164.460 107.835 164.660 ;
        RECT 103.835 163.860 104.235 164.460 ;
        RECT 103.835 163.660 107.835 163.860 ;
        RECT 103.835 163.060 104.235 163.660 ;
        RECT 103.835 162.860 107.835 163.060 ;
        RECT 103.835 162.260 104.235 162.860 ;
        RECT 103.835 162.060 107.835 162.260 ;
        RECT 103.835 161.460 104.235 162.060 ;
        RECT 103.835 161.260 107.835 161.460 ;
        RECT 103.835 160.660 104.235 161.260 ;
        RECT 103.835 160.460 107.835 160.660 ;
        RECT 103.835 159.860 104.235 160.460 ;
        RECT 103.835 159.660 107.835 159.860 ;
        RECT 103.835 159.060 104.235 159.660 ;
        RECT 103.835 158.860 107.835 159.060 ;
        RECT 108.585 158.860 108.785 166.460 ;
        RECT 109.385 158.860 109.585 166.460 ;
        RECT 110.185 158.860 110.385 166.460 ;
        RECT 110.985 158.860 111.185 166.460 ;
        RECT 111.785 158.860 111.985 166.460 ;
        RECT 113.285 166.860 113.485 174.460 ;
        RECT 114.085 166.860 114.285 174.460 ;
        RECT 114.885 166.860 115.085 174.460 ;
        RECT 115.685 166.860 115.885 174.460 ;
        RECT 116.485 166.860 116.685 174.460 ;
        RECT 117.435 174.260 121.435 174.460 ;
        RECT 121.035 173.660 121.435 174.260 ;
        RECT 117.435 173.460 121.435 173.660 ;
        RECT 121.035 172.860 121.435 173.460 ;
        RECT 117.435 172.660 121.435 172.860 ;
        RECT 121.035 172.060 121.435 172.660 ;
        RECT 117.435 171.860 121.435 172.060 ;
        RECT 121.035 171.260 121.435 171.860 ;
        RECT 117.435 171.060 121.435 171.260 ;
        RECT 121.035 170.460 121.435 171.060 ;
        RECT 117.435 170.260 121.435 170.460 ;
        RECT 121.035 169.660 121.435 170.260 ;
        RECT 117.435 169.460 121.435 169.660 ;
        RECT 121.035 168.860 121.435 169.460 ;
        RECT 117.435 168.660 121.435 168.860 ;
        RECT 121.035 168.060 121.435 168.660 ;
        RECT 117.435 167.860 121.435 168.060 ;
        RECT 121.035 167.260 121.435 167.860 ;
        RECT 117.435 167.060 121.435 167.260 ;
        RECT 121.035 166.860 121.435 167.060 ;
        RECT 113.285 166.460 121.435 166.860 ;
        RECT 113.285 158.860 113.485 166.460 ;
        RECT 114.085 158.860 114.285 166.460 ;
        RECT 114.885 158.860 115.085 166.460 ;
        RECT 115.685 158.860 115.885 166.460 ;
        RECT 116.485 158.860 116.685 166.460 ;
        RECT 121.035 166.260 121.435 166.460 ;
        RECT 117.435 166.060 121.435 166.260 ;
        RECT 121.035 165.460 121.435 166.060 ;
        RECT 117.435 165.260 121.435 165.460 ;
        RECT 121.035 164.660 121.435 165.260 ;
        RECT 117.435 164.460 121.435 164.660 ;
        RECT 121.035 163.860 121.435 164.460 ;
        RECT 117.435 163.660 121.435 163.860 ;
        RECT 121.035 163.060 121.435 163.660 ;
        RECT 117.435 162.860 121.435 163.060 ;
        RECT 121.035 162.260 121.435 162.860 ;
        RECT 117.435 162.060 121.435 162.260 ;
        RECT 121.035 161.460 121.435 162.060 ;
        RECT 117.435 161.260 121.435 161.460 ;
        RECT 121.035 160.660 121.435 161.260 ;
        RECT 117.435 160.460 121.435 160.660 ;
        RECT 121.035 159.860 121.435 160.460 ;
        RECT 117.435 159.660 121.435 159.860 ;
        RECT 121.035 159.060 121.435 159.660 ;
        RECT 117.435 158.860 121.435 159.060 ;
      LAYER mcon ;
        RECT 7.245 172.655 7.415 172.825 ;
        RECT 8.110 172.650 8.280 172.820 ;
        RECT 8.570 172.650 8.740 172.820 ;
        RECT 9.030 172.650 9.200 172.820 ;
        RECT 9.490 172.650 9.660 172.820 ;
        RECT 9.950 172.650 10.120 172.820 ;
        RECT 10.410 172.650 10.580 172.820 ;
        RECT 10.870 172.650 11.040 172.820 ;
        RECT 11.330 172.650 11.500 172.820 ;
        RECT 11.790 172.650 11.960 172.820 ;
        RECT 12.250 172.650 12.420 172.820 ;
        RECT 12.710 172.650 12.880 172.820 ;
        RECT 13.170 172.650 13.340 172.820 ;
        RECT 13.630 172.650 13.800 172.820 ;
        RECT 14.090 172.650 14.260 172.820 ;
        RECT 14.550 172.650 14.720 172.820 ;
        RECT 15.010 172.650 15.180 172.820 ;
        RECT 15.470 172.650 15.640 172.820 ;
        RECT 15.930 172.650 16.100 172.820 ;
        RECT 16.390 172.650 16.560 172.820 ;
        RECT 16.850 172.650 17.020 172.820 ;
        RECT 17.310 172.650 17.480 172.820 ;
        RECT 17.770 172.650 17.940 172.820 ;
        RECT 18.230 172.650 18.400 172.820 ;
        RECT 18.690 172.650 18.860 172.820 ;
        RECT 19.150 172.650 19.320 172.820 ;
        RECT 19.610 172.650 19.780 172.820 ;
        RECT 20.070 172.650 20.240 172.820 ;
        RECT 20.530 172.650 20.700 172.820 ;
        RECT 20.990 172.650 21.160 172.820 ;
        RECT 21.450 172.650 21.620 172.820 ;
        RECT 21.910 172.650 22.080 172.820 ;
        RECT 22.370 172.650 22.540 172.820 ;
        RECT 22.830 172.650 23.000 172.820 ;
        RECT 23.290 172.650 23.460 172.820 ;
        RECT 23.750 172.650 23.920 172.820 ;
        RECT 43.885 170.960 44.185 171.410 ;
        RECT 43.885 170.210 44.185 170.660 ;
        RECT 43.885 169.460 44.185 169.910 ;
        RECT 43.885 168.710 44.185 169.160 ;
        RECT 43.885 167.960 44.185 168.410 ;
        RECT 6.730 167.210 6.900 167.380 ;
        RECT 7.190 167.210 7.360 167.380 ;
        RECT 7.650 167.210 7.820 167.380 ;
        RECT 8.110 167.210 8.280 167.380 ;
        RECT 8.570 167.210 8.740 167.380 ;
        RECT 9.030 167.210 9.200 167.380 ;
        RECT 9.490 167.210 9.660 167.380 ;
        RECT 9.950 167.210 10.120 167.380 ;
        RECT 10.410 167.210 10.580 167.380 ;
        RECT 10.870 167.210 11.040 167.380 ;
        RECT 11.330 167.210 11.500 167.380 ;
        RECT 11.790 167.210 11.960 167.380 ;
        RECT 12.250 167.210 12.420 167.380 ;
        RECT 12.710 167.210 12.880 167.380 ;
        RECT 13.170 167.210 13.340 167.380 ;
        RECT 13.630 167.210 13.800 167.380 ;
        RECT 14.090 167.210 14.260 167.380 ;
        RECT 14.550 167.210 14.720 167.380 ;
        RECT 15.010 167.210 15.180 167.380 ;
        RECT 15.470 167.210 15.640 167.380 ;
        RECT 15.930 167.210 16.100 167.380 ;
        RECT 16.390 167.210 16.560 167.380 ;
        RECT 16.850 167.210 17.020 167.380 ;
        RECT 17.310 167.210 17.480 167.380 ;
        RECT 17.770 167.210 17.940 167.380 ;
        RECT 18.230 167.210 18.400 167.380 ;
        RECT 18.690 167.210 18.860 167.380 ;
        RECT 19.150 167.210 19.320 167.380 ;
        RECT 19.610 167.210 19.780 167.380 ;
        RECT 20.070 167.210 20.240 167.380 ;
        RECT 20.530 167.210 20.700 167.380 ;
        RECT 20.990 167.210 21.160 167.380 ;
        RECT 21.450 167.210 21.620 167.380 ;
        RECT 21.910 167.210 22.080 167.380 ;
        RECT 22.370 167.210 22.540 167.380 ;
        RECT 22.830 167.210 23.000 167.380 ;
        RECT 23.290 167.210 23.460 167.380 ;
        RECT 23.750 167.210 23.920 167.380 ;
        RECT 43.885 167.210 44.185 167.660 ;
        RECT 43.885 166.460 44.185 166.910 ;
        RECT 43.885 165.710 44.185 166.160 ;
        RECT 43.885 164.960 44.185 165.410 ;
        RECT 43.885 164.210 44.185 164.660 ;
        RECT 43.885 163.460 44.185 163.910 ;
        RECT 43.885 162.710 44.185 163.160 ;
        RECT 43.885 161.960 44.185 162.410 ;
        RECT 61.085 170.960 61.385 171.410 ;
        RECT 61.085 170.210 61.385 170.660 ;
        RECT 61.085 169.460 61.385 169.910 ;
        RECT 61.085 168.710 61.385 169.160 ;
        RECT 61.085 167.960 61.385 168.410 ;
        RECT 61.085 167.210 61.385 167.660 ;
        RECT 61.085 166.460 61.385 166.910 ;
        RECT 61.085 165.710 61.385 166.160 ;
        RECT 61.085 164.960 61.385 165.410 ;
        RECT 61.085 164.210 61.385 164.660 ;
        RECT 61.085 163.460 61.385 163.910 ;
        RECT 61.085 162.710 61.385 163.160 ;
        RECT 61.085 161.960 61.385 162.410 ;
        RECT 63.885 170.960 64.185 171.410 ;
        RECT 63.885 170.210 64.185 170.660 ;
        RECT 63.885 169.460 64.185 169.910 ;
        RECT 63.885 168.710 64.185 169.160 ;
        RECT 63.885 167.960 64.185 168.410 ;
        RECT 63.885 167.210 64.185 167.660 ;
        RECT 63.885 166.460 64.185 166.910 ;
        RECT 63.885 165.710 64.185 166.160 ;
        RECT 63.885 164.960 64.185 165.410 ;
        RECT 63.885 164.210 64.185 164.660 ;
        RECT 63.885 163.460 64.185 163.910 ;
        RECT 63.885 162.710 64.185 163.160 ;
        RECT 63.885 161.960 64.185 162.410 ;
        RECT 81.085 170.960 81.385 171.410 ;
        RECT 81.085 170.210 81.385 170.660 ;
        RECT 81.085 169.460 81.385 169.910 ;
        RECT 81.085 168.710 81.385 169.160 ;
        RECT 81.085 167.960 81.385 168.410 ;
        RECT 81.085 167.210 81.385 167.660 ;
        RECT 81.085 166.460 81.385 166.910 ;
        RECT 81.085 165.710 81.385 166.160 ;
        RECT 81.085 164.960 81.385 165.410 ;
        RECT 81.085 164.210 81.385 164.660 ;
        RECT 81.085 163.460 81.385 163.910 ;
        RECT 81.085 162.710 81.385 163.160 ;
        RECT 81.085 161.960 81.385 162.410 ;
        RECT 83.885 170.960 84.185 171.410 ;
        RECT 83.885 170.210 84.185 170.660 ;
        RECT 83.885 169.460 84.185 169.910 ;
        RECT 83.885 168.710 84.185 169.160 ;
        RECT 83.885 167.960 84.185 168.410 ;
        RECT 83.885 167.210 84.185 167.660 ;
        RECT 83.885 166.460 84.185 166.910 ;
        RECT 83.885 165.710 84.185 166.160 ;
        RECT 83.885 164.960 84.185 165.410 ;
        RECT 83.885 164.210 84.185 164.660 ;
        RECT 83.885 163.460 84.185 163.910 ;
        RECT 83.885 162.710 84.185 163.160 ;
        RECT 83.885 161.960 84.185 162.410 ;
        RECT 101.085 170.960 101.385 171.410 ;
        RECT 101.085 170.210 101.385 170.660 ;
        RECT 101.085 169.460 101.385 169.910 ;
        RECT 101.085 168.710 101.385 169.160 ;
        RECT 101.085 167.960 101.385 168.410 ;
        RECT 101.085 167.210 101.385 167.660 ;
        RECT 101.085 166.460 101.385 166.910 ;
        RECT 101.085 165.710 101.385 166.160 ;
        RECT 101.085 164.960 101.385 165.410 ;
        RECT 101.085 164.210 101.385 164.660 ;
        RECT 101.085 163.460 101.385 163.910 ;
        RECT 101.085 162.710 101.385 163.160 ;
        RECT 101.085 161.960 101.385 162.410 ;
        RECT 103.885 170.960 104.185 171.410 ;
        RECT 103.885 170.210 104.185 170.660 ;
        RECT 103.885 169.460 104.185 169.910 ;
        RECT 103.885 168.710 104.185 169.160 ;
        RECT 103.885 167.960 104.185 168.410 ;
        RECT 103.885 167.210 104.185 167.660 ;
        RECT 103.885 166.460 104.185 166.910 ;
        RECT 103.885 165.710 104.185 166.160 ;
        RECT 103.885 164.960 104.185 165.410 ;
        RECT 103.885 164.210 104.185 164.660 ;
        RECT 103.885 163.460 104.185 163.910 ;
        RECT 103.885 162.710 104.185 163.160 ;
        RECT 103.885 161.960 104.185 162.410 ;
        RECT 121.085 170.960 121.385 171.410 ;
        RECT 121.085 170.210 121.385 170.660 ;
        RECT 121.085 169.460 121.385 169.910 ;
        RECT 121.085 168.710 121.385 169.160 ;
        RECT 121.085 167.960 121.385 168.410 ;
        RECT 121.085 167.210 121.385 167.660 ;
        RECT 121.085 166.460 121.385 166.910 ;
        RECT 121.085 165.710 121.385 166.160 ;
        RECT 121.085 164.960 121.385 165.410 ;
        RECT 121.085 164.210 121.385 164.660 ;
        RECT 121.085 163.460 121.385 163.910 ;
        RECT 121.085 162.710 121.385 163.160 ;
        RECT 121.085 161.960 121.385 162.410 ;
      LAYER met1 ;
        RECT 16.435 178.760 22.105 178.765 ;
        RECT 0.000 177.485 129.510 178.760 ;
        RECT 49.435 175.460 55.835 176.660 ;
        RECT 69.435 175.460 75.835 176.660 ;
        RECT 89.435 175.460 95.835 176.660 ;
        RECT 109.435 175.460 115.835 176.660 ;
        RECT 52.135 174.810 53.135 175.460 ;
        RECT 72.135 174.810 73.135 175.460 ;
        RECT 92.135 174.810 93.135 175.460 ;
        RECT 112.135 174.810 113.135 175.460 ;
        RECT 48.785 174.660 56.485 174.810 ;
        RECT 68.785 174.660 76.485 174.810 ;
        RECT 88.785 174.660 96.485 174.810 ;
        RECT 108.785 174.660 116.485 174.810 ;
        RECT 7.100 172.975 7.560 172.980 ;
        RECT 0.000 172.495 24.065 172.975 ;
        RECT 43.835 169.860 44.585 171.660 ;
        RECT 0.000 167.055 24.065 167.535 ;
        RECT 42.635 167.110 44.585 169.860 ;
        RECT 42.635 166.210 42.785 167.110 ;
        RECT 43.435 166.960 44.585 167.110 ;
        RECT 44.735 166.960 44.885 174.510 ;
        RECT 45.335 166.960 45.485 174.510 ;
        RECT 45.935 166.960 46.085 174.510 ;
        RECT 46.535 166.960 46.685 174.510 ;
        RECT 47.135 166.960 47.285 174.510 ;
        RECT 47.735 166.960 47.885 174.510 ;
        RECT 52.135 174.210 53.135 174.660 ;
        RECT 48.785 174.060 56.485 174.210 ;
        RECT 52.135 173.610 53.135 174.060 ;
        RECT 48.785 173.460 56.485 173.610 ;
        RECT 52.135 173.010 53.135 173.460 ;
        RECT 48.785 172.860 56.485 173.010 ;
        RECT 52.135 172.410 53.135 172.860 ;
        RECT 48.785 172.260 56.485 172.410 ;
        RECT 52.135 171.810 53.135 172.260 ;
        RECT 48.785 171.660 56.485 171.810 ;
        RECT 52.135 171.210 53.135 171.660 ;
        RECT 48.785 171.060 56.485 171.210 ;
        RECT 52.135 170.610 53.135 171.060 ;
        RECT 48.785 170.460 56.485 170.610 ;
        RECT 52.135 170.010 53.135 170.460 ;
        RECT 48.785 169.860 56.485 170.010 ;
        RECT 52.135 169.410 53.135 169.860 ;
        RECT 48.785 169.260 56.485 169.410 ;
        RECT 52.135 168.810 53.135 169.260 ;
        RECT 48.785 168.660 56.485 168.810 ;
        RECT 52.135 168.210 53.135 168.660 ;
        RECT 48.785 168.060 56.485 168.210 ;
        RECT 52.135 167.610 53.135 168.060 ;
        RECT 48.785 167.460 56.485 167.610 ;
        RECT 52.135 166.960 53.135 167.460 ;
        RECT 57.385 166.960 57.535 174.510 ;
        RECT 57.985 166.960 58.135 174.510 ;
        RECT 58.585 166.960 58.735 174.510 ;
        RECT 59.185 166.960 59.335 174.510 ;
        RECT 59.785 166.960 59.935 174.510 ;
        RECT 60.385 166.960 60.535 174.510 ;
        RECT 60.685 169.860 61.435 171.660 ;
        RECT 63.835 169.860 64.585 171.660 ;
        RECT 60.685 167.110 64.585 169.860 ;
        RECT 60.685 166.960 61.835 167.110 ;
        RECT 43.435 166.360 61.835 166.960 ;
        RECT 43.435 166.210 44.585 166.360 ;
        RECT 42.635 163.460 44.585 166.210 ;
        RECT 43.835 161.710 44.585 163.460 ;
        RECT 44.735 158.810 44.885 166.360 ;
        RECT 45.335 158.810 45.485 166.360 ;
        RECT 45.935 158.810 46.085 166.360 ;
        RECT 46.535 158.810 46.685 166.360 ;
        RECT 47.135 158.810 47.285 166.360 ;
        RECT 47.735 158.810 47.885 166.360 ;
        RECT 52.135 165.860 53.135 166.360 ;
        RECT 48.785 165.710 56.485 165.860 ;
        RECT 52.135 165.260 53.135 165.710 ;
        RECT 48.785 165.110 56.485 165.260 ;
        RECT 52.135 164.660 53.135 165.110 ;
        RECT 48.785 164.510 56.485 164.660 ;
        RECT 52.135 164.060 53.135 164.510 ;
        RECT 48.785 163.910 56.485 164.060 ;
        RECT 52.135 163.460 53.135 163.910 ;
        RECT 48.785 163.310 56.485 163.460 ;
        RECT 52.135 162.860 53.135 163.310 ;
        RECT 48.785 162.710 56.485 162.860 ;
        RECT 52.135 162.260 53.135 162.710 ;
        RECT 48.785 162.110 56.485 162.260 ;
        RECT 52.135 161.660 53.135 162.110 ;
        RECT 48.785 161.510 56.485 161.660 ;
        RECT 52.135 161.060 53.135 161.510 ;
        RECT 48.785 160.910 56.485 161.060 ;
        RECT 52.135 160.460 53.135 160.910 ;
        RECT 48.785 160.310 56.485 160.460 ;
        RECT 52.135 159.860 53.135 160.310 ;
        RECT 48.785 159.710 56.485 159.860 ;
        RECT 52.135 159.260 53.135 159.710 ;
        RECT 48.785 159.110 56.485 159.260 ;
        RECT 52.135 158.660 53.135 159.110 ;
        RECT 57.385 158.810 57.535 166.360 ;
        RECT 57.985 158.810 58.135 166.360 ;
        RECT 58.585 158.810 58.735 166.360 ;
        RECT 59.185 158.810 59.335 166.360 ;
        RECT 59.785 158.810 59.935 166.360 ;
        RECT 60.385 158.810 60.535 166.360 ;
        RECT 60.685 166.210 61.835 166.360 ;
        RECT 62.485 166.210 62.785 167.110 ;
        RECT 63.435 166.960 64.585 167.110 ;
        RECT 64.735 166.960 64.885 174.510 ;
        RECT 65.335 166.960 65.485 174.510 ;
        RECT 65.935 166.960 66.085 174.510 ;
        RECT 66.535 166.960 66.685 174.510 ;
        RECT 67.135 166.960 67.285 174.510 ;
        RECT 67.735 166.960 67.885 174.510 ;
        RECT 72.135 174.210 73.135 174.660 ;
        RECT 68.785 174.060 76.485 174.210 ;
        RECT 72.135 173.610 73.135 174.060 ;
        RECT 68.785 173.460 76.485 173.610 ;
        RECT 72.135 173.010 73.135 173.460 ;
        RECT 68.785 172.860 76.485 173.010 ;
        RECT 72.135 172.410 73.135 172.860 ;
        RECT 68.785 172.260 76.485 172.410 ;
        RECT 72.135 171.810 73.135 172.260 ;
        RECT 68.785 171.660 76.485 171.810 ;
        RECT 72.135 171.210 73.135 171.660 ;
        RECT 68.785 171.060 76.485 171.210 ;
        RECT 72.135 170.610 73.135 171.060 ;
        RECT 68.785 170.460 76.485 170.610 ;
        RECT 72.135 170.010 73.135 170.460 ;
        RECT 68.785 169.860 76.485 170.010 ;
        RECT 72.135 169.410 73.135 169.860 ;
        RECT 68.785 169.260 76.485 169.410 ;
        RECT 72.135 168.810 73.135 169.260 ;
        RECT 68.785 168.660 76.485 168.810 ;
        RECT 72.135 168.210 73.135 168.660 ;
        RECT 68.785 168.060 76.485 168.210 ;
        RECT 72.135 167.610 73.135 168.060 ;
        RECT 68.785 167.460 76.485 167.610 ;
        RECT 72.135 166.960 73.135 167.460 ;
        RECT 77.385 166.960 77.535 174.510 ;
        RECT 77.985 166.960 78.135 174.510 ;
        RECT 78.585 166.960 78.735 174.510 ;
        RECT 79.185 166.960 79.335 174.510 ;
        RECT 79.785 166.960 79.935 174.510 ;
        RECT 80.385 166.960 80.535 174.510 ;
        RECT 80.685 169.860 81.435 171.660 ;
        RECT 83.835 169.860 84.585 171.660 ;
        RECT 80.685 167.110 84.585 169.860 ;
        RECT 80.685 166.960 81.835 167.110 ;
        RECT 63.435 166.360 81.835 166.960 ;
        RECT 63.435 166.210 64.585 166.360 ;
        RECT 60.685 163.460 64.585 166.210 ;
        RECT 60.685 161.710 61.435 163.460 ;
        RECT 63.835 161.710 64.585 163.460 ;
        RECT 64.735 158.810 64.885 166.360 ;
        RECT 65.335 158.810 65.485 166.360 ;
        RECT 65.935 158.810 66.085 166.360 ;
        RECT 66.535 158.810 66.685 166.360 ;
        RECT 67.135 158.810 67.285 166.360 ;
        RECT 67.735 158.810 67.885 166.360 ;
        RECT 72.135 165.860 73.135 166.360 ;
        RECT 68.785 165.710 76.485 165.860 ;
        RECT 72.135 165.260 73.135 165.710 ;
        RECT 68.785 165.110 76.485 165.260 ;
        RECT 72.135 164.660 73.135 165.110 ;
        RECT 68.785 164.510 76.485 164.660 ;
        RECT 72.135 164.060 73.135 164.510 ;
        RECT 68.785 163.910 76.485 164.060 ;
        RECT 72.135 163.460 73.135 163.910 ;
        RECT 68.785 163.310 76.485 163.460 ;
        RECT 72.135 162.860 73.135 163.310 ;
        RECT 68.785 162.710 76.485 162.860 ;
        RECT 72.135 162.260 73.135 162.710 ;
        RECT 68.785 162.110 76.485 162.260 ;
        RECT 72.135 161.660 73.135 162.110 ;
        RECT 68.785 161.510 76.485 161.660 ;
        RECT 72.135 161.060 73.135 161.510 ;
        RECT 68.785 160.910 76.485 161.060 ;
        RECT 72.135 160.460 73.135 160.910 ;
        RECT 68.785 160.310 76.485 160.460 ;
        RECT 72.135 159.860 73.135 160.310 ;
        RECT 68.785 159.710 76.485 159.860 ;
        RECT 72.135 159.260 73.135 159.710 ;
        RECT 68.785 159.110 76.485 159.260 ;
        RECT 72.135 158.660 73.135 159.110 ;
        RECT 77.385 158.810 77.535 166.360 ;
        RECT 77.985 158.810 78.135 166.360 ;
        RECT 78.585 158.810 78.735 166.360 ;
        RECT 79.185 158.810 79.335 166.360 ;
        RECT 79.785 158.810 79.935 166.360 ;
        RECT 80.385 158.810 80.535 166.360 ;
        RECT 80.685 166.210 81.835 166.360 ;
        RECT 82.485 166.210 82.785 167.110 ;
        RECT 83.435 166.960 84.585 167.110 ;
        RECT 84.735 166.960 84.885 174.510 ;
        RECT 85.335 166.960 85.485 174.510 ;
        RECT 85.935 166.960 86.085 174.510 ;
        RECT 86.535 166.960 86.685 174.510 ;
        RECT 87.135 166.960 87.285 174.510 ;
        RECT 87.735 166.960 87.885 174.510 ;
        RECT 92.135 174.210 93.135 174.660 ;
        RECT 88.785 174.060 96.485 174.210 ;
        RECT 92.135 173.610 93.135 174.060 ;
        RECT 88.785 173.460 96.485 173.610 ;
        RECT 92.135 173.010 93.135 173.460 ;
        RECT 88.785 172.860 96.485 173.010 ;
        RECT 92.135 172.410 93.135 172.860 ;
        RECT 88.785 172.260 96.485 172.410 ;
        RECT 92.135 171.810 93.135 172.260 ;
        RECT 88.785 171.660 96.485 171.810 ;
        RECT 92.135 171.210 93.135 171.660 ;
        RECT 88.785 171.060 96.485 171.210 ;
        RECT 92.135 170.610 93.135 171.060 ;
        RECT 88.785 170.460 96.485 170.610 ;
        RECT 92.135 170.010 93.135 170.460 ;
        RECT 88.785 169.860 96.485 170.010 ;
        RECT 92.135 169.410 93.135 169.860 ;
        RECT 88.785 169.260 96.485 169.410 ;
        RECT 92.135 168.810 93.135 169.260 ;
        RECT 88.785 168.660 96.485 168.810 ;
        RECT 92.135 168.210 93.135 168.660 ;
        RECT 88.785 168.060 96.485 168.210 ;
        RECT 92.135 167.610 93.135 168.060 ;
        RECT 88.785 167.460 96.485 167.610 ;
        RECT 92.135 166.960 93.135 167.460 ;
        RECT 97.385 166.960 97.535 174.510 ;
        RECT 97.985 166.960 98.135 174.510 ;
        RECT 98.585 166.960 98.735 174.510 ;
        RECT 99.185 166.960 99.335 174.510 ;
        RECT 99.785 166.960 99.935 174.510 ;
        RECT 100.385 166.960 100.535 174.510 ;
        RECT 100.685 169.860 101.435 171.660 ;
        RECT 103.835 169.860 104.585 171.660 ;
        RECT 100.685 167.110 104.585 169.860 ;
        RECT 100.685 166.960 101.835 167.110 ;
        RECT 83.435 166.360 101.835 166.960 ;
        RECT 83.435 166.210 84.585 166.360 ;
        RECT 80.685 163.460 84.585 166.210 ;
        RECT 80.685 161.710 81.435 163.460 ;
        RECT 83.835 161.710 84.585 163.460 ;
        RECT 84.735 158.810 84.885 166.360 ;
        RECT 85.335 158.810 85.485 166.360 ;
        RECT 85.935 158.810 86.085 166.360 ;
        RECT 86.535 158.810 86.685 166.360 ;
        RECT 87.135 158.810 87.285 166.360 ;
        RECT 87.735 158.810 87.885 166.360 ;
        RECT 92.135 165.860 93.135 166.360 ;
        RECT 88.785 165.710 96.485 165.860 ;
        RECT 92.135 165.260 93.135 165.710 ;
        RECT 88.785 165.110 96.485 165.260 ;
        RECT 92.135 164.660 93.135 165.110 ;
        RECT 88.785 164.510 96.485 164.660 ;
        RECT 92.135 164.060 93.135 164.510 ;
        RECT 88.785 163.910 96.485 164.060 ;
        RECT 92.135 163.460 93.135 163.910 ;
        RECT 88.785 163.310 96.485 163.460 ;
        RECT 92.135 162.860 93.135 163.310 ;
        RECT 88.785 162.710 96.485 162.860 ;
        RECT 92.135 162.260 93.135 162.710 ;
        RECT 88.785 162.110 96.485 162.260 ;
        RECT 92.135 161.660 93.135 162.110 ;
        RECT 88.785 161.510 96.485 161.660 ;
        RECT 92.135 161.060 93.135 161.510 ;
        RECT 88.785 160.910 96.485 161.060 ;
        RECT 92.135 160.460 93.135 160.910 ;
        RECT 88.785 160.310 96.485 160.460 ;
        RECT 92.135 159.860 93.135 160.310 ;
        RECT 88.785 159.710 96.485 159.860 ;
        RECT 92.135 159.260 93.135 159.710 ;
        RECT 88.785 159.110 96.485 159.260 ;
        RECT 92.135 158.660 93.135 159.110 ;
        RECT 97.385 158.810 97.535 166.360 ;
        RECT 97.985 158.810 98.135 166.360 ;
        RECT 98.585 158.810 98.735 166.360 ;
        RECT 99.185 158.810 99.335 166.360 ;
        RECT 99.785 158.810 99.935 166.360 ;
        RECT 100.385 158.810 100.535 166.360 ;
        RECT 100.685 166.210 101.835 166.360 ;
        RECT 102.485 166.210 102.785 167.110 ;
        RECT 103.435 166.960 104.585 167.110 ;
        RECT 104.735 166.960 104.885 174.510 ;
        RECT 105.335 166.960 105.485 174.510 ;
        RECT 105.935 166.960 106.085 174.510 ;
        RECT 106.535 166.960 106.685 174.510 ;
        RECT 107.135 166.960 107.285 174.510 ;
        RECT 107.735 166.960 107.885 174.510 ;
        RECT 112.135 174.210 113.135 174.660 ;
        RECT 108.785 174.060 116.485 174.210 ;
        RECT 112.135 173.610 113.135 174.060 ;
        RECT 108.785 173.460 116.485 173.610 ;
        RECT 112.135 173.010 113.135 173.460 ;
        RECT 108.785 172.860 116.485 173.010 ;
        RECT 112.135 172.410 113.135 172.860 ;
        RECT 108.785 172.260 116.485 172.410 ;
        RECT 112.135 171.810 113.135 172.260 ;
        RECT 108.785 171.660 116.485 171.810 ;
        RECT 112.135 171.210 113.135 171.660 ;
        RECT 108.785 171.060 116.485 171.210 ;
        RECT 112.135 170.610 113.135 171.060 ;
        RECT 108.785 170.460 116.485 170.610 ;
        RECT 112.135 170.010 113.135 170.460 ;
        RECT 108.785 169.860 116.485 170.010 ;
        RECT 112.135 169.410 113.135 169.860 ;
        RECT 108.785 169.260 116.485 169.410 ;
        RECT 112.135 168.810 113.135 169.260 ;
        RECT 108.785 168.660 116.485 168.810 ;
        RECT 112.135 168.210 113.135 168.660 ;
        RECT 108.785 168.060 116.485 168.210 ;
        RECT 112.135 167.610 113.135 168.060 ;
        RECT 108.785 167.460 116.485 167.610 ;
        RECT 112.135 166.960 113.135 167.460 ;
        RECT 117.385 166.960 117.535 174.510 ;
        RECT 117.985 166.960 118.135 174.510 ;
        RECT 118.585 166.960 118.735 174.510 ;
        RECT 119.185 166.960 119.335 174.510 ;
        RECT 119.785 166.960 119.935 174.510 ;
        RECT 120.385 166.960 120.535 174.510 ;
        RECT 120.685 169.860 121.435 171.660 ;
        RECT 120.685 167.510 122.635 169.860 ;
        RECT 120.685 167.110 129.510 167.510 ;
        RECT 120.685 166.960 121.835 167.110 ;
        RECT 103.435 166.360 121.835 166.960 ;
        RECT 103.435 166.210 104.585 166.360 ;
        RECT 100.685 163.460 104.585 166.210 ;
        RECT 100.685 161.710 101.435 163.460 ;
        RECT 103.835 161.710 104.585 163.460 ;
        RECT 104.735 158.810 104.885 166.360 ;
        RECT 105.335 158.810 105.485 166.360 ;
        RECT 105.935 158.810 106.085 166.360 ;
        RECT 106.535 158.810 106.685 166.360 ;
        RECT 107.135 158.810 107.285 166.360 ;
        RECT 107.735 158.810 107.885 166.360 ;
        RECT 112.135 165.860 113.135 166.360 ;
        RECT 108.785 165.710 116.485 165.860 ;
        RECT 112.135 165.260 113.135 165.710 ;
        RECT 108.785 165.110 116.485 165.260 ;
        RECT 112.135 164.660 113.135 165.110 ;
        RECT 108.785 164.510 116.485 164.660 ;
        RECT 112.135 164.060 113.135 164.510 ;
        RECT 108.785 163.910 116.485 164.060 ;
        RECT 112.135 163.460 113.135 163.910 ;
        RECT 108.785 163.310 116.485 163.460 ;
        RECT 112.135 162.860 113.135 163.310 ;
        RECT 108.785 162.710 116.485 162.860 ;
        RECT 112.135 162.260 113.135 162.710 ;
        RECT 108.785 162.110 116.485 162.260 ;
        RECT 112.135 161.660 113.135 162.110 ;
        RECT 108.785 161.510 116.485 161.660 ;
        RECT 112.135 161.060 113.135 161.510 ;
        RECT 108.785 160.910 116.485 161.060 ;
        RECT 112.135 160.460 113.135 160.910 ;
        RECT 108.785 160.310 116.485 160.460 ;
        RECT 112.135 159.860 113.135 160.310 ;
        RECT 108.785 159.710 116.485 159.860 ;
        RECT 112.135 159.260 113.135 159.710 ;
        RECT 108.785 159.110 116.485 159.260 ;
        RECT 112.135 158.660 113.135 159.110 ;
        RECT 117.385 158.810 117.535 166.360 ;
        RECT 117.985 158.810 118.135 166.360 ;
        RECT 118.585 158.810 118.735 166.360 ;
        RECT 119.185 158.810 119.335 166.360 ;
        RECT 119.785 158.810 119.935 166.360 ;
        RECT 120.385 158.810 120.535 166.360 ;
        RECT 120.685 166.210 121.835 166.360 ;
        RECT 122.485 166.235 129.510 167.110 ;
        RECT 122.485 166.210 122.635 166.235 ;
        RECT 120.685 163.460 122.635 166.210 ;
        RECT 120.685 161.710 121.435 163.460 ;
        RECT 48.785 158.510 56.485 158.660 ;
        RECT 68.785 158.510 76.485 158.660 ;
        RECT 88.785 158.510 96.485 158.660 ;
        RECT 108.785 158.510 116.485 158.660 ;
        RECT 52.135 157.860 53.135 158.510 ;
        RECT 72.135 157.860 73.135 158.510 ;
        RECT 92.135 157.860 93.135 158.510 ;
        RECT 112.135 157.860 113.135 158.510 ;
        RECT 49.435 156.660 55.835 157.860 ;
        RECT 69.435 156.660 75.835 157.860 ;
        RECT 89.435 156.660 95.835 157.860 ;
        RECT 109.435 156.660 115.835 157.860 ;
      LAYER via ;
        RECT 0.160 178.305 0.560 178.705 ;
        RECT 0.785 178.305 1.185 178.705 ;
        RECT 1.410 178.305 1.810 178.705 ;
        RECT 127.675 178.230 128.075 178.630 ;
        RECT 128.300 178.230 128.700 178.630 ;
        RECT 128.925 178.230 129.325 178.630 ;
        RECT 0.160 177.775 0.560 178.175 ;
        RECT 0.785 177.775 1.185 178.175 ;
        RECT 1.410 177.775 1.810 178.175 ;
        RECT 127.670 177.630 128.070 178.030 ;
        RECT 128.295 177.630 128.695 178.030 ;
        RECT 128.920 177.630 129.320 178.030 ;
        RECT 49.535 175.560 50.535 176.560 ;
        RECT 50.685 175.560 51.685 176.560 ;
        RECT 51.835 175.560 53.435 176.560 ;
        RECT 53.585 175.560 54.585 176.560 ;
        RECT 54.735 175.560 55.735 176.560 ;
        RECT 69.535 175.560 70.535 176.560 ;
        RECT 70.685 175.560 71.685 176.560 ;
        RECT 71.835 175.560 73.435 176.560 ;
        RECT 73.585 175.560 74.585 176.560 ;
        RECT 74.735 175.560 75.735 176.560 ;
        RECT 89.535 175.560 90.535 176.560 ;
        RECT 90.685 175.560 91.685 176.560 ;
        RECT 91.835 175.560 93.435 176.560 ;
        RECT 93.585 175.560 94.585 176.560 ;
        RECT 94.735 175.560 95.735 176.560 ;
        RECT 109.535 175.560 110.535 176.560 ;
        RECT 110.685 175.560 111.685 176.560 ;
        RECT 111.835 175.560 113.435 176.560 ;
        RECT 113.585 175.560 114.585 176.560 ;
        RECT 114.735 175.560 115.735 176.560 ;
        RECT 0.080 172.540 0.490 172.930 ;
        RECT 0.650 172.540 1.060 172.930 ;
        RECT 1.220 172.540 1.630 172.930 ;
        RECT 42.735 169.060 43.435 169.760 ;
        RECT 42.735 168.210 43.435 168.910 ;
        RECT 0.080 167.100 0.490 167.490 ;
        RECT 0.650 167.100 1.060 167.490 ;
        RECT 1.220 167.100 1.630 167.490 ;
        RECT 42.735 167.360 43.435 168.060 ;
        RECT 61.835 169.060 62.535 169.760 ;
        RECT 62.735 169.060 63.435 169.760 ;
        RECT 61.835 168.210 62.535 168.910 ;
        RECT 62.735 168.210 63.435 168.910 ;
        RECT 61.835 167.360 62.535 168.060 ;
        RECT 62.735 167.360 63.435 168.060 ;
        RECT 42.735 165.260 43.435 165.960 ;
        RECT 42.735 164.410 43.435 165.110 ;
        RECT 42.735 163.560 43.435 164.260 ;
        RECT 81.835 169.060 82.535 169.760 ;
        RECT 82.735 169.060 83.435 169.760 ;
        RECT 81.835 168.210 82.535 168.910 ;
        RECT 82.735 168.210 83.435 168.910 ;
        RECT 81.835 167.360 82.535 168.060 ;
        RECT 82.735 167.360 83.435 168.060 ;
        RECT 61.835 165.260 62.535 165.960 ;
        RECT 62.735 165.260 63.435 165.960 ;
        RECT 61.835 164.410 62.535 165.110 ;
        RECT 62.735 164.410 63.435 165.110 ;
        RECT 61.835 163.560 62.535 164.260 ;
        RECT 62.735 163.560 63.435 164.260 ;
        RECT 101.835 169.060 102.535 169.760 ;
        RECT 102.735 169.060 103.435 169.760 ;
        RECT 101.835 168.210 102.535 168.910 ;
        RECT 102.735 168.210 103.435 168.910 ;
        RECT 101.835 167.360 102.535 168.060 ;
        RECT 102.735 167.360 103.435 168.060 ;
        RECT 81.835 165.260 82.535 165.960 ;
        RECT 82.735 165.260 83.435 165.960 ;
        RECT 81.835 164.410 82.535 165.110 ;
        RECT 82.735 164.410 83.435 165.110 ;
        RECT 81.835 163.560 82.535 164.260 ;
        RECT 82.735 163.560 83.435 164.260 ;
        RECT 121.835 169.060 122.535 169.760 ;
        RECT 121.835 168.210 122.535 168.910 ;
        RECT 121.835 167.360 122.535 168.060 ;
        RECT 101.835 165.260 102.535 165.960 ;
        RECT 102.735 165.260 103.435 165.960 ;
        RECT 101.835 164.410 102.535 165.110 ;
        RECT 102.735 164.410 103.435 165.110 ;
        RECT 101.835 163.560 102.535 164.260 ;
        RECT 102.735 163.560 103.435 164.260 ;
        RECT 122.800 166.980 123.200 167.380 ;
        RECT 123.425 166.980 123.825 167.380 ;
        RECT 124.050 166.980 124.450 167.380 ;
        RECT 127.675 166.980 128.075 167.380 ;
        RECT 128.300 166.980 128.700 167.380 ;
        RECT 128.925 166.980 129.325 167.380 ;
        RECT 122.795 166.380 123.195 166.780 ;
        RECT 123.420 166.380 123.820 166.780 ;
        RECT 124.045 166.380 124.445 166.780 ;
        RECT 127.670 166.380 128.070 166.780 ;
        RECT 128.295 166.380 128.695 166.780 ;
        RECT 128.920 166.380 129.320 166.780 ;
        RECT 121.835 165.260 122.535 165.960 ;
        RECT 121.835 164.410 122.535 165.110 ;
        RECT 121.835 163.560 122.535 164.260 ;
        RECT 49.535 156.760 50.535 157.760 ;
        RECT 50.635 156.760 51.635 157.760 ;
        RECT 51.785 156.760 53.385 157.760 ;
        RECT 53.585 156.760 54.585 157.760 ;
        RECT 54.735 156.760 55.735 157.760 ;
        RECT 69.535 156.760 70.535 157.760 ;
        RECT 70.635 156.760 71.635 157.760 ;
        RECT 71.785 156.760 73.385 157.760 ;
        RECT 73.585 156.760 74.585 157.760 ;
        RECT 74.735 156.760 75.735 157.760 ;
        RECT 89.535 156.760 90.535 157.760 ;
        RECT 90.635 156.760 91.635 157.760 ;
        RECT 91.785 156.760 93.385 157.760 ;
        RECT 93.585 156.760 94.585 157.760 ;
        RECT 94.735 156.760 95.735 157.760 ;
        RECT 109.535 156.760 110.535 157.760 ;
        RECT 110.635 156.760 111.635 157.760 ;
        RECT 111.785 156.760 113.385 157.760 ;
        RECT 113.585 156.760 114.585 157.760 ;
        RECT 114.735 156.760 115.735 157.760 ;
      LAYER met2 ;
        RECT 0.000 177.640 2.000 178.760 ;
        RECT 127.510 177.485 129.510 178.760 ;
        RECT 49.435 175.760 55.835 176.660 ;
        RECT 69.435 175.760 75.835 176.660 ;
        RECT 89.435 175.760 95.835 176.660 ;
        RECT 109.435 175.760 115.835 176.660 ;
        RECT 47.535 175.260 57.735 175.760 ;
        RECT 67.535 175.260 77.735 175.760 ;
        RECT 87.535 175.260 97.735 175.760 ;
        RECT 107.535 175.260 117.735 175.760 ;
        RECT 44.435 175.210 60.835 175.260 ;
        RECT 44.435 174.660 48.235 175.210 ;
        RECT 47.935 174.210 48.235 174.660 ;
        RECT 44.385 174.060 48.235 174.210 ;
        RECT 47.935 173.610 48.235 174.060 ;
        RECT 44.385 173.460 48.235 173.610 ;
        RECT 47.935 173.010 48.235 173.460 ;
        RECT 0.000 172.495 1.710 172.975 ;
        RECT 44.385 172.860 48.235 173.010 ;
        RECT 47.935 172.410 48.235 172.860 ;
        RECT 44.385 172.260 48.235 172.410 ;
        RECT 47.935 171.810 48.235 172.260 ;
        RECT 44.385 171.660 48.235 171.810 ;
        RECT 47.935 171.210 48.235 171.660 ;
        RECT 44.385 171.060 48.235 171.210 ;
        RECT 47.935 170.610 48.235 171.060 ;
        RECT 44.385 170.460 48.235 170.610 ;
        RECT 47.935 170.010 48.235 170.460 ;
        RECT 44.385 169.860 48.235 170.010 ;
        RECT 0.000 167.055 1.710 167.535 ;
        RECT 42.635 163.460 43.535 169.860 ;
        RECT 47.935 169.410 48.235 169.860 ;
        RECT 44.385 169.260 48.235 169.410 ;
        RECT 47.935 168.810 48.235 169.260 ;
        RECT 44.385 168.660 48.235 168.810 ;
        RECT 47.935 168.210 48.235 168.660 ;
        RECT 44.385 168.060 48.235 168.210 ;
        RECT 47.935 167.610 48.235 168.060 ;
        RECT 44.385 167.460 48.235 167.610 ;
        RECT 47.935 167.010 48.235 167.460 ;
        RECT 48.685 167.010 48.835 175.210 ;
        RECT 49.285 167.010 49.435 175.210 ;
        RECT 49.885 167.010 50.035 175.210 ;
        RECT 50.485 167.010 50.635 175.210 ;
        RECT 51.085 167.010 51.235 175.210 ;
        RECT 51.685 167.010 51.835 175.210 ;
        RECT 47.935 165.860 48.235 166.310 ;
        RECT 44.385 165.710 48.235 165.860 ;
        RECT 47.935 165.260 48.235 165.710 ;
        RECT 44.385 165.110 48.235 165.260 ;
        RECT 47.935 164.660 48.235 165.110 ;
        RECT 44.385 164.510 48.235 164.660 ;
        RECT 47.935 164.060 48.235 164.510 ;
        RECT 44.385 163.910 48.235 164.060 ;
        RECT 47.935 163.460 48.235 163.910 ;
        RECT 44.385 163.310 48.235 163.460 ;
        RECT 47.935 162.860 48.235 163.310 ;
        RECT 44.385 162.710 48.235 162.860 ;
        RECT 47.935 162.260 48.235 162.710 ;
        RECT 44.385 162.110 48.235 162.260 ;
        RECT 47.935 161.660 48.235 162.110 ;
        RECT 44.385 161.510 48.235 161.660 ;
        RECT 47.935 161.060 48.235 161.510 ;
        RECT 44.385 160.910 48.235 161.060 ;
        RECT 47.935 160.460 48.235 160.910 ;
        RECT 44.385 160.310 48.235 160.460 ;
        RECT 47.935 159.860 48.235 160.310 ;
        RECT 44.385 159.710 48.235 159.860 ;
        RECT 47.935 159.260 48.235 159.710 ;
        RECT 44.385 159.110 48.235 159.260 ;
        RECT 47.935 158.660 48.235 159.110 ;
        RECT 44.435 158.110 48.235 158.660 ;
        RECT 48.685 158.110 48.835 166.310 ;
        RECT 49.285 158.110 49.435 166.310 ;
        RECT 49.885 158.110 50.035 166.310 ;
        RECT 50.485 158.110 50.635 166.310 ;
        RECT 51.085 158.110 51.235 166.310 ;
        RECT 51.685 158.110 51.835 166.310 ;
        RECT 52.285 158.110 52.985 175.210 ;
        RECT 53.435 167.010 53.585 175.210 ;
        RECT 54.035 167.010 54.185 175.210 ;
        RECT 54.635 167.010 54.785 175.210 ;
        RECT 55.235 167.010 55.385 175.210 ;
        RECT 55.835 167.010 55.985 175.210 ;
        RECT 56.435 167.010 56.585 175.210 ;
        RECT 57.035 174.660 60.835 175.210 ;
        RECT 64.435 175.210 80.835 175.260 ;
        RECT 64.435 174.660 68.235 175.210 ;
        RECT 57.035 174.210 57.335 174.660 ;
        RECT 67.935 174.210 68.235 174.660 ;
        RECT 57.035 174.060 60.885 174.210 ;
        RECT 64.385 174.060 68.235 174.210 ;
        RECT 57.035 173.610 57.335 174.060 ;
        RECT 67.935 173.610 68.235 174.060 ;
        RECT 57.035 173.460 60.885 173.610 ;
        RECT 64.385 173.460 68.235 173.610 ;
        RECT 57.035 173.010 57.335 173.460 ;
        RECT 67.935 173.010 68.235 173.460 ;
        RECT 57.035 172.860 60.885 173.010 ;
        RECT 64.385 172.860 68.235 173.010 ;
        RECT 57.035 172.410 57.335 172.860 ;
        RECT 67.935 172.410 68.235 172.860 ;
        RECT 57.035 172.260 60.885 172.410 ;
        RECT 64.385 172.260 68.235 172.410 ;
        RECT 57.035 171.810 57.335 172.260 ;
        RECT 67.935 171.810 68.235 172.260 ;
        RECT 57.035 171.660 60.885 171.810 ;
        RECT 64.385 171.660 68.235 171.810 ;
        RECT 57.035 171.210 57.335 171.660 ;
        RECT 67.935 171.210 68.235 171.660 ;
        RECT 57.035 171.060 60.885 171.210 ;
        RECT 64.385 171.060 68.235 171.210 ;
        RECT 57.035 170.610 57.335 171.060 ;
        RECT 67.935 170.610 68.235 171.060 ;
        RECT 57.035 170.460 60.885 170.610 ;
        RECT 64.385 170.460 68.235 170.610 ;
        RECT 57.035 170.010 57.335 170.460 ;
        RECT 67.935 170.010 68.235 170.460 ;
        RECT 57.035 169.860 60.885 170.010 ;
        RECT 64.385 169.860 68.235 170.010 ;
        RECT 57.035 169.410 57.335 169.860 ;
        RECT 57.035 169.260 60.885 169.410 ;
        RECT 57.035 168.810 57.335 169.260 ;
        RECT 57.035 168.660 60.885 168.810 ;
        RECT 57.035 168.210 57.335 168.660 ;
        RECT 57.035 168.060 60.885 168.210 ;
        RECT 57.035 167.610 57.335 168.060 ;
        RECT 57.035 167.460 60.885 167.610 ;
        RECT 57.035 167.010 57.335 167.460 ;
        RECT 53.435 158.110 53.585 166.310 ;
        RECT 54.035 158.110 54.185 166.310 ;
        RECT 54.635 158.110 54.785 166.310 ;
        RECT 55.235 158.110 55.385 166.310 ;
        RECT 55.835 158.110 55.985 166.310 ;
        RECT 56.435 158.110 56.585 166.310 ;
        RECT 57.035 165.860 57.335 166.310 ;
        RECT 57.035 165.710 60.885 165.860 ;
        RECT 57.035 165.260 57.335 165.710 ;
        RECT 57.035 165.110 60.885 165.260 ;
        RECT 57.035 164.660 57.335 165.110 ;
        RECT 57.035 164.510 60.885 164.660 ;
        RECT 57.035 164.060 57.335 164.510 ;
        RECT 57.035 163.910 60.885 164.060 ;
        RECT 57.035 163.460 57.335 163.910 ;
        RECT 61.735 163.460 63.535 169.860 ;
        RECT 67.935 169.410 68.235 169.860 ;
        RECT 64.385 169.260 68.235 169.410 ;
        RECT 67.935 168.810 68.235 169.260 ;
        RECT 64.385 168.660 68.235 168.810 ;
        RECT 67.935 168.210 68.235 168.660 ;
        RECT 64.385 168.060 68.235 168.210 ;
        RECT 67.935 167.610 68.235 168.060 ;
        RECT 64.385 167.460 68.235 167.610 ;
        RECT 67.935 167.010 68.235 167.460 ;
        RECT 68.685 167.010 68.835 175.210 ;
        RECT 69.285 167.010 69.435 175.210 ;
        RECT 69.885 167.010 70.035 175.210 ;
        RECT 70.485 167.010 70.635 175.210 ;
        RECT 71.085 167.010 71.235 175.210 ;
        RECT 71.685 167.010 71.835 175.210 ;
        RECT 67.935 165.860 68.235 166.310 ;
        RECT 64.385 165.710 68.235 165.860 ;
        RECT 67.935 165.260 68.235 165.710 ;
        RECT 64.385 165.110 68.235 165.260 ;
        RECT 67.935 164.660 68.235 165.110 ;
        RECT 64.385 164.510 68.235 164.660 ;
        RECT 67.935 164.060 68.235 164.510 ;
        RECT 64.385 163.910 68.235 164.060 ;
        RECT 67.935 163.460 68.235 163.910 ;
        RECT 57.035 163.310 60.885 163.460 ;
        RECT 64.385 163.310 68.235 163.460 ;
        RECT 57.035 162.860 57.335 163.310 ;
        RECT 67.935 162.860 68.235 163.310 ;
        RECT 57.035 162.710 60.885 162.860 ;
        RECT 64.385 162.710 68.235 162.860 ;
        RECT 57.035 162.260 57.335 162.710 ;
        RECT 67.935 162.260 68.235 162.710 ;
        RECT 57.035 162.110 60.885 162.260 ;
        RECT 64.385 162.110 68.235 162.260 ;
        RECT 57.035 161.660 57.335 162.110 ;
        RECT 67.935 161.660 68.235 162.110 ;
        RECT 57.035 161.510 60.885 161.660 ;
        RECT 64.385 161.510 68.235 161.660 ;
        RECT 57.035 161.060 57.335 161.510 ;
        RECT 67.935 161.060 68.235 161.510 ;
        RECT 57.035 160.910 60.885 161.060 ;
        RECT 64.385 160.910 68.235 161.060 ;
        RECT 57.035 160.460 57.335 160.910 ;
        RECT 67.935 160.460 68.235 160.910 ;
        RECT 57.035 160.310 60.885 160.460 ;
        RECT 64.385 160.310 68.235 160.460 ;
        RECT 57.035 159.860 57.335 160.310 ;
        RECT 67.935 159.860 68.235 160.310 ;
        RECT 57.035 159.710 60.885 159.860 ;
        RECT 64.385 159.710 68.235 159.860 ;
        RECT 57.035 159.260 57.335 159.710 ;
        RECT 67.935 159.260 68.235 159.710 ;
        RECT 57.035 159.110 60.885 159.260 ;
        RECT 64.385 159.110 68.235 159.260 ;
        RECT 57.035 158.660 57.335 159.110 ;
        RECT 67.935 158.660 68.235 159.110 ;
        RECT 57.035 158.110 60.835 158.660 ;
        RECT 44.435 158.060 60.835 158.110 ;
        RECT 64.435 158.110 68.235 158.660 ;
        RECT 68.685 158.110 68.835 166.310 ;
        RECT 69.285 158.110 69.435 166.310 ;
        RECT 69.885 158.110 70.035 166.310 ;
        RECT 70.485 158.110 70.635 166.310 ;
        RECT 71.085 158.110 71.235 166.310 ;
        RECT 71.685 158.110 71.835 166.310 ;
        RECT 72.285 158.110 72.985 175.210 ;
        RECT 73.435 167.010 73.585 175.210 ;
        RECT 74.035 167.010 74.185 175.210 ;
        RECT 74.635 167.010 74.785 175.210 ;
        RECT 75.235 167.010 75.385 175.210 ;
        RECT 75.835 167.010 75.985 175.210 ;
        RECT 76.435 167.010 76.585 175.210 ;
        RECT 77.035 174.660 80.835 175.210 ;
        RECT 84.435 175.210 100.835 175.260 ;
        RECT 84.435 174.660 88.235 175.210 ;
        RECT 77.035 174.210 77.335 174.660 ;
        RECT 87.935 174.210 88.235 174.660 ;
        RECT 77.035 174.060 80.885 174.210 ;
        RECT 84.385 174.060 88.235 174.210 ;
        RECT 77.035 173.610 77.335 174.060 ;
        RECT 87.935 173.610 88.235 174.060 ;
        RECT 77.035 173.460 80.885 173.610 ;
        RECT 84.385 173.460 88.235 173.610 ;
        RECT 77.035 173.010 77.335 173.460 ;
        RECT 87.935 173.010 88.235 173.460 ;
        RECT 77.035 172.860 80.885 173.010 ;
        RECT 84.385 172.860 88.235 173.010 ;
        RECT 77.035 172.410 77.335 172.860 ;
        RECT 87.935 172.410 88.235 172.860 ;
        RECT 77.035 172.260 80.885 172.410 ;
        RECT 84.385 172.260 88.235 172.410 ;
        RECT 77.035 171.810 77.335 172.260 ;
        RECT 87.935 171.810 88.235 172.260 ;
        RECT 77.035 171.660 80.885 171.810 ;
        RECT 84.385 171.660 88.235 171.810 ;
        RECT 77.035 171.210 77.335 171.660 ;
        RECT 87.935 171.210 88.235 171.660 ;
        RECT 77.035 171.060 80.885 171.210 ;
        RECT 84.385 171.060 88.235 171.210 ;
        RECT 77.035 170.610 77.335 171.060 ;
        RECT 87.935 170.610 88.235 171.060 ;
        RECT 77.035 170.460 80.885 170.610 ;
        RECT 84.385 170.460 88.235 170.610 ;
        RECT 77.035 170.010 77.335 170.460 ;
        RECT 87.935 170.010 88.235 170.460 ;
        RECT 77.035 169.860 80.885 170.010 ;
        RECT 84.385 169.860 88.235 170.010 ;
        RECT 77.035 169.410 77.335 169.860 ;
        RECT 77.035 169.260 80.885 169.410 ;
        RECT 77.035 168.810 77.335 169.260 ;
        RECT 77.035 168.660 80.885 168.810 ;
        RECT 77.035 168.210 77.335 168.660 ;
        RECT 77.035 168.060 80.885 168.210 ;
        RECT 77.035 167.610 77.335 168.060 ;
        RECT 77.035 167.460 80.885 167.610 ;
        RECT 77.035 167.010 77.335 167.460 ;
        RECT 73.435 158.110 73.585 166.310 ;
        RECT 74.035 158.110 74.185 166.310 ;
        RECT 74.635 158.110 74.785 166.310 ;
        RECT 75.235 158.110 75.385 166.310 ;
        RECT 75.835 158.110 75.985 166.310 ;
        RECT 76.435 158.110 76.585 166.310 ;
        RECT 77.035 165.860 77.335 166.310 ;
        RECT 77.035 165.710 80.885 165.860 ;
        RECT 77.035 165.260 77.335 165.710 ;
        RECT 77.035 165.110 80.885 165.260 ;
        RECT 77.035 164.660 77.335 165.110 ;
        RECT 77.035 164.510 80.885 164.660 ;
        RECT 77.035 164.060 77.335 164.510 ;
        RECT 77.035 163.910 80.885 164.060 ;
        RECT 77.035 163.460 77.335 163.910 ;
        RECT 81.735 163.460 83.535 169.860 ;
        RECT 87.935 169.410 88.235 169.860 ;
        RECT 84.385 169.260 88.235 169.410 ;
        RECT 87.935 168.810 88.235 169.260 ;
        RECT 84.385 168.660 88.235 168.810 ;
        RECT 87.935 168.210 88.235 168.660 ;
        RECT 84.385 168.060 88.235 168.210 ;
        RECT 87.935 167.610 88.235 168.060 ;
        RECT 84.385 167.460 88.235 167.610 ;
        RECT 87.935 167.010 88.235 167.460 ;
        RECT 88.685 167.010 88.835 175.210 ;
        RECT 89.285 167.010 89.435 175.210 ;
        RECT 89.885 167.010 90.035 175.210 ;
        RECT 90.485 167.010 90.635 175.210 ;
        RECT 91.085 167.010 91.235 175.210 ;
        RECT 91.685 167.010 91.835 175.210 ;
        RECT 87.935 165.860 88.235 166.310 ;
        RECT 84.385 165.710 88.235 165.860 ;
        RECT 87.935 165.260 88.235 165.710 ;
        RECT 84.385 165.110 88.235 165.260 ;
        RECT 87.935 164.660 88.235 165.110 ;
        RECT 84.385 164.510 88.235 164.660 ;
        RECT 87.935 164.060 88.235 164.510 ;
        RECT 84.385 163.910 88.235 164.060 ;
        RECT 87.935 163.460 88.235 163.910 ;
        RECT 77.035 163.310 80.885 163.460 ;
        RECT 84.385 163.310 88.235 163.460 ;
        RECT 77.035 162.860 77.335 163.310 ;
        RECT 87.935 162.860 88.235 163.310 ;
        RECT 77.035 162.710 80.885 162.860 ;
        RECT 84.385 162.710 88.235 162.860 ;
        RECT 77.035 162.260 77.335 162.710 ;
        RECT 87.935 162.260 88.235 162.710 ;
        RECT 77.035 162.110 80.885 162.260 ;
        RECT 84.385 162.110 88.235 162.260 ;
        RECT 77.035 161.660 77.335 162.110 ;
        RECT 87.935 161.660 88.235 162.110 ;
        RECT 77.035 161.510 80.885 161.660 ;
        RECT 84.385 161.510 88.235 161.660 ;
        RECT 77.035 161.060 77.335 161.510 ;
        RECT 87.935 161.060 88.235 161.510 ;
        RECT 77.035 160.910 80.885 161.060 ;
        RECT 84.385 160.910 88.235 161.060 ;
        RECT 77.035 160.460 77.335 160.910 ;
        RECT 87.935 160.460 88.235 160.910 ;
        RECT 77.035 160.310 80.885 160.460 ;
        RECT 84.385 160.310 88.235 160.460 ;
        RECT 77.035 159.860 77.335 160.310 ;
        RECT 87.935 159.860 88.235 160.310 ;
        RECT 77.035 159.710 80.885 159.860 ;
        RECT 84.385 159.710 88.235 159.860 ;
        RECT 77.035 159.260 77.335 159.710 ;
        RECT 87.935 159.260 88.235 159.710 ;
        RECT 77.035 159.110 80.885 159.260 ;
        RECT 84.385 159.110 88.235 159.260 ;
        RECT 77.035 158.660 77.335 159.110 ;
        RECT 87.935 158.660 88.235 159.110 ;
        RECT 77.035 158.110 80.835 158.660 ;
        RECT 64.435 158.060 80.835 158.110 ;
        RECT 84.435 158.110 88.235 158.660 ;
        RECT 88.685 158.110 88.835 166.310 ;
        RECT 89.285 158.110 89.435 166.310 ;
        RECT 89.885 158.110 90.035 166.310 ;
        RECT 90.485 158.110 90.635 166.310 ;
        RECT 91.085 158.110 91.235 166.310 ;
        RECT 91.685 158.110 91.835 166.310 ;
        RECT 92.285 158.110 92.985 175.210 ;
        RECT 93.435 167.010 93.585 175.210 ;
        RECT 94.035 167.010 94.185 175.210 ;
        RECT 94.635 167.010 94.785 175.210 ;
        RECT 95.235 167.010 95.385 175.210 ;
        RECT 95.835 167.010 95.985 175.210 ;
        RECT 96.435 167.010 96.585 175.210 ;
        RECT 97.035 174.660 100.835 175.210 ;
        RECT 104.435 175.210 120.835 175.260 ;
        RECT 104.435 174.660 108.235 175.210 ;
        RECT 97.035 174.210 97.335 174.660 ;
        RECT 107.935 174.210 108.235 174.660 ;
        RECT 97.035 174.060 100.885 174.210 ;
        RECT 104.385 174.060 108.235 174.210 ;
        RECT 97.035 173.610 97.335 174.060 ;
        RECT 107.935 173.610 108.235 174.060 ;
        RECT 97.035 173.460 100.885 173.610 ;
        RECT 104.385 173.460 108.235 173.610 ;
        RECT 97.035 173.010 97.335 173.460 ;
        RECT 107.935 173.010 108.235 173.460 ;
        RECT 97.035 172.860 100.885 173.010 ;
        RECT 104.385 172.860 108.235 173.010 ;
        RECT 97.035 172.410 97.335 172.860 ;
        RECT 107.935 172.410 108.235 172.860 ;
        RECT 97.035 172.260 100.885 172.410 ;
        RECT 104.385 172.260 108.235 172.410 ;
        RECT 97.035 171.810 97.335 172.260 ;
        RECT 107.935 171.810 108.235 172.260 ;
        RECT 97.035 171.660 100.885 171.810 ;
        RECT 104.385 171.660 108.235 171.810 ;
        RECT 97.035 171.210 97.335 171.660 ;
        RECT 107.935 171.210 108.235 171.660 ;
        RECT 97.035 171.060 100.885 171.210 ;
        RECT 104.385 171.060 108.235 171.210 ;
        RECT 97.035 170.610 97.335 171.060 ;
        RECT 107.935 170.610 108.235 171.060 ;
        RECT 97.035 170.460 100.885 170.610 ;
        RECT 104.385 170.460 108.235 170.610 ;
        RECT 97.035 170.010 97.335 170.460 ;
        RECT 107.935 170.010 108.235 170.460 ;
        RECT 97.035 169.860 100.885 170.010 ;
        RECT 104.385 169.860 108.235 170.010 ;
        RECT 97.035 169.410 97.335 169.860 ;
        RECT 97.035 169.260 100.885 169.410 ;
        RECT 97.035 168.810 97.335 169.260 ;
        RECT 97.035 168.660 100.885 168.810 ;
        RECT 97.035 168.210 97.335 168.660 ;
        RECT 97.035 168.060 100.885 168.210 ;
        RECT 97.035 167.610 97.335 168.060 ;
        RECT 97.035 167.460 100.885 167.610 ;
        RECT 97.035 167.010 97.335 167.460 ;
        RECT 93.435 158.110 93.585 166.310 ;
        RECT 94.035 158.110 94.185 166.310 ;
        RECT 94.635 158.110 94.785 166.310 ;
        RECT 95.235 158.110 95.385 166.310 ;
        RECT 95.835 158.110 95.985 166.310 ;
        RECT 96.435 158.110 96.585 166.310 ;
        RECT 97.035 165.860 97.335 166.310 ;
        RECT 97.035 165.710 100.885 165.860 ;
        RECT 97.035 165.260 97.335 165.710 ;
        RECT 97.035 165.110 100.885 165.260 ;
        RECT 97.035 164.660 97.335 165.110 ;
        RECT 97.035 164.510 100.885 164.660 ;
        RECT 97.035 164.060 97.335 164.510 ;
        RECT 97.035 163.910 100.885 164.060 ;
        RECT 97.035 163.460 97.335 163.910 ;
        RECT 101.735 163.460 103.535 169.860 ;
        RECT 107.935 169.410 108.235 169.860 ;
        RECT 104.385 169.260 108.235 169.410 ;
        RECT 107.935 168.810 108.235 169.260 ;
        RECT 104.385 168.660 108.235 168.810 ;
        RECT 107.935 168.210 108.235 168.660 ;
        RECT 104.385 168.060 108.235 168.210 ;
        RECT 107.935 167.610 108.235 168.060 ;
        RECT 104.385 167.460 108.235 167.610 ;
        RECT 107.935 167.010 108.235 167.460 ;
        RECT 108.685 167.010 108.835 175.210 ;
        RECT 109.285 167.010 109.435 175.210 ;
        RECT 109.885 167.010 110.035 175.210 ;
        RECT 110.485 167.010 110.635 175.210 ;
        RECT 111.085 167.010 111.235 175.210 ;
        RECT 111.685 167.010 111.835 175.210 ;
        RECT 107.935 165.860 108.235 166.310 ;
        RECT 104.385 165.710 108.235 165.860 ;
        RECT 107.935 165.260 108.235 165.710 ;
        RECT 104.385 165.110 108.235 165.260 ;
        RECT 107.935 164.660 108.235 165.110 ;
        RECT 104.385 164.510 108.235 164.660 ;
        RECT 107.935 164.060 108.235 164.510 ;
        RECT 104.385 163.910 108.235 164.060 ;
        RECT 107.935 163.460 108.235 163.910 ;
        RECT 97.035 163.310 100.885 163.460 ;
        RECT 104.385 163.310 108.235 163.460 ;
        RECT 97.035 162.860 97.335 163.310 ;
        RECT 107.935 162.860 108.235 163.310 ;
        RECT 97.035 162.710 100.885 162.860 ;
        RECT 104.385 162.710 108.235 162.860 ;
        RECT 97.035 162.260 97.335 162.710 ;
        RECT 107.935 162.260 108.235 162.710 ;
        RECT 97.035 162.110 100.885 162.260 ;
        RECT 104.385 162.110 108.235 162.260 ;
        RECT 97.035 161.660 97.335 162.110 ;
        RECT 107.935 161.660 108.235 162.110 ;
        RECT 97.035 161.510 100.885 161.660 ;
        RECT 104.385 161.510 108.235 161.660 ;
        RECT 97.035 161.060 97.335 161.510 ;
        RECT 107.935 161.060 108.235 161.510 ;
        RECT 97.035 160.910 100.885 161.060 ;
        RECT 104.385 160.910 108.235 161.060 ;
        RECT 97.035 160.460 97.335 160.910 ;
        RECT 107.935 160.460 108.235 160.910 ;
        RECT 97.035 160.310 100.885 160.460 ;
        RECT 104.385 160.310 108.235 160.460 ;
        RECT 97.035 159.860 97.335 160.310 ;
        RECT 107.935 159.860 108.235 160.310 ;
        RECT 97.035 159.710 100.885 159.860 ;
        RECT 104.385 159.710 108.235 159.860 ;
        RECT 97.035 159.260 97.335 159.710 ;
        RECT 107.935 159.260 108.235 159.710 ;
        RECT 97.035 159.110 100.885 159.260 ;
        RECT 104.385 159.110 108.235 159.260 ;
        RECT 97.035 158.660 97.335 159.110 ;
        RECT 107.935 158.660 108.235 159.110 ;
        RECT 97.035 158.110 100.835 158.660 ;
        RECT 84.435 158.060 100.835 158.110 ;
        RECT 104.435 158.110 108.235 158.660 ;
        RECT 108.685 158.110 108.835 166.310 ;
        RECT 109.285 158.110 109.435 166.310 ;
        RECT 109.885 158.110 110.035 166.310 ;
        RECT 110.485 158.110 110.635 166.310 ;
        RECT 111.085 158.110 111.235 166.310 ;
        RECT 111.685 158.110 111.835 166.310 ;
        RECT 112.285 158.110 112.985 175.210 ;
        RECT 113.435 167.010 113.585 175.210 ;
        RECT 114.035 167.010 114.185 175.210 ;
        RECT 114.635 167.010 114.785 175.210 ;
        RECT 115.235 167.010 115.385 175.210 ;
        RECT 115.835 167.010 115.985 175.210 ;
        RECT 116.435 167.010 116.585 175.210 ;
        RECT 117.035 174.660 120.835 175.210 ;
        RECT 117.035 174.210 117.335 174.660 ;
        RECT 117.035 174.060 120.885 174.210 ;
        RECT 117.035 173.610 117.335 174.060 ;
        RECT 117.035 173.460 120.885 173.610 ;
        RECT 117.035 173.010 117.335 173.460 ;
        RECT 117.035 172.860 120.885 173.010 ;
        RECT 117.035 172.410 117.335 172.860 ;
        RECT 117.035 172.260 120.885 172.410 ;
        RECT 117.035 171.810 117.335 172.260 ;
        RECT 117.035 171.660 120.885 171.810 ;
        RECT 117.035 171.210 117.335 171.660 ;
        RECT 117.035 171.060 120.885 171.210 ;
        RECT 117.035 170.610 117.335 171.060 ;
        RECT 117.035 170.460 120.885 170.610 ;
        RECT 117.035 170.010 117.335 170.460 ;
        RECT 117.035 169.860 120.885 170.010 ;
        RECT 117.035 169.410 117.335 169.860 ;
        RECT 117.035 169.260 120.885 169.410 ;
        RECT 117.035 168.810 117.335 169.260 ;
        RECT 117.035 168.660 120.885 168.810 ;
        RECT 117.035 168.210 117.335 168.660 ;
        RECT 117.035 168.060 120.885 168.210 ;
        RECT 117.035 167.610 117.335 168.060 ;
        RECT 117.035 167.460 120.885 167.610 ;
        RECT 121.735 167.510 122.635 169.860 ;
        RECT 117.035 167.010 117.335 167.460 ;
        RECT 113.435 158.110 113.585 166.310 ;
        RECT 114.035 158.110 114.185 166.310 ;
        RECT 114.635 158.110 114.785 166.310 ;
        RECT 115.235 158.110 115.385 166.310 ;
        RECT 115.835 158.110 115.985 166.310 ;
        RECT 116.435 158.110 116.585 166.310 ;
        RECT 117.035 165.860 117.335 166.310 ;
        RECT 121.735 166.235 124.635 167.510 ;
        RECT 127.510 166.235 129.510 167.510 ;
        RECT 117.035 165.710 120.885 165.860 ;
        RECT 117.035 165.260 117.335 165.710 ;
        RECT 117.035 165.110 120.885 165.260 ;
        RECT 117.035 164.660 117.335 165.110 ;
        RECT 117.035 164.510 120.885 164.660 ;
        RECT 117.035 164.060 117.335 164.510 ;
        RECT 117.035 163.910 120.885 164.060 ;
        RECT 117.035 163.460 117.335 163.910 ;
        RECT 121.735 163.460 122.635 166.235 ;
        RECT 117.035 163.310 120.885 163.460 ;
        RECT 117.035 162.860 117.335 163.310 ;
        RECT 117.035 162.710 120.885 162.860 ;
        RECT 117.035 162.260 117.335 162.710 ;
        RECT 117.035 162.110 120.885 162.260 ;
        RECT 117.035 161.660 117.335 162.110 ;
        RECT 117.035 161.510 120.885 161.660 ;
        RECT 117.035 161.060 117.335 161.510 ;
        RECT 117.035 160.910 120.885 161.060 ;
        RECT 117.035 160.460 117.335 160.910 ;
        RECT 117.035 160.310 120.885 160.460 ;
        RECT 117.035 159.860 117.335 160.310 ;
        RECT 117.035 159.710 120.885 159.860 ;
        RECT 117.035 159.260 117.335 159.710 ;
        RECT 117.035 159.110 120.885 159.260 ;
        RECT 117.035 158.660 117.335 159.110 ;
        RECT 117.035 158.110 120.835 158.660 ;
        RECT 104.435 158.060 120.835 158.110 ;
        RECT 47.535 157.560 57.735 158.060 ;
        RECT 67.535 157.560 77.735 158.060 ;
        RECT 87.535 157.560 97.735 158.060 ;
        RECT 107.535 157.560 117.735 158.060 ;
        RECT 49.435 156.660 55.835 157.560 ;
        RECT 69.435 156.660 75.835 157.560 ;
        RECT 89.435 156.660 95.835 157.560 ;
        RECT 109.435 156.660 115.835 157.560 ;
      LAYER via2 ;
        RECT 0.160 178.305 0.560 178.705 ;
        RECT 0.785 178.305 1.185 178.705 ;
        RECT 1.410 178.305 1.810 178.705 ;
        RECT 0.160 177.775 0.560 178.175 ;
        RECT 0.785 177.775 1.185 178.175 ;
        RECT 1.410 177.775 1.810 178.175 ;
        RECT 127.675 178.230 128.075 178.630 ;
        RECT 128.300 178.230 128.700 178.630 ;
        RECT 128.925 178.230 129.325 178.630 ;
        RECT 127.670 177.630 128.070 178.030 ;
        RECT 128.295 177.630 128.695 178.030 ;
        RECT 128.920 177.630 129.320 178.030 ;
        RECT 0.080 172.540 0.490 172.930 ;
        RECT 0.650 172.540 1.060 172.930 ;
        RECT 1.220 172.540 1.630 172.930 ;
        RECT 0.080 167.100 0.490 167.490 ;
        RECT 0.650 167.100 1.060 167.490 ;
        RECT 1.220 167.100 1.630 167.490 ;
        RECT 122.800 166.980 123.200 167.380 ;
        RECT 123.425 166.980 123.825 167.380 ;
        RECT 124.050 166.980 124.450 167.380 ;
        RECT 122.795 166.380 123.195 166.780 ;
        RECT 123.420 166.380 123.820 166.780 ;
        RECT 124.045 166.380 124.445 166.780 ;
        RECT 127.675 166.980 128.075 167.380 ;
        RECT 128.300 166.980 128.700 167.380 ;
        RECT 128.925 166.980 129.325 167.380 ;
        RECT 127.670 166.380 128.070 166.780 ;
        RECT 128.295 166.380 128.695 166.780 ;
        RECT 128.920 166.380 129.320 166.780 ;
      LAYER met3 ;
        RECT 0.000 177.640 2.000 178.760 ;
        RECT 127.510 177.485 129.510 178.760 ;
        RECT 49.435 175.810 55.835 176.660 ;
        RECT 69.435 175.810 75.835 176.660 ;
        RECT 89.435 175.810 95.835 176.660 ;
        RECT 109.435 175.810 115.835 176.660 ;
        RECT 0.000 172.495 1.710 172.975 ;
        RECT 0.000 167.055 1.710 167.535 ;
        RECT 42.635 163.460 43.485 169.860 ;
        RECT 61.785 163.460 63.485 169.860 ;
        RECT 81.785 163.460 83.485 169.860 ;
        RECT 101.785 163.460 103.485 169.860 ;
        RECT 121.785 167.510 122.635 169.860 ;
        RECT 121.785 166.235 124.635 167.510 ;
        RECT 127.510 166.235 129.510 167.510 ;
        RECT 121.785 163.460 122.635 166.235 ;
        RECT 49.435 156.660 55.835 157.510 ;
        RECT 69.435 156.660 75.835 157.510 ;
        RECT 89.435 156.660 95.835 157.510 ;
        RECT 109.435 156.660 115.835 157.510 ;
      LAYER via3 ;
        RECT 0.160 178.305 0.555 178.705 ;
        RECT 0.780 178.305 1.180 178.705 ;
        RECT 1.410 178.305 1.810 178.705 ;
        RECT 0.160 177.775 0.555 178.175 ;
        RECT 0.780 177.775 1.180 178.175 ;
        RECT 1.410 177.775 1.810 178.175 ;
        RECT 127.675 178.230 128.075 178.630 ;
        RECT 128.300 178.230 128.700 178.630 ;
        RECT 128.925 178.230 129.325 178.630 ;
        RECT 127.670 177.630 128.070 178.030 ;
        RECT 128.295 177.630 128.695 178.030 ;
        RECT 128.920 177.630 129.320 178.030 ;
        RECT 49.535 175.910 50.185 176.560 ;
        RECT 50.335 175.910 50.985 176.560 ;
        RECT 51.135 175.910 51.785 176.560 ;
        RECT 53.485 175.910 54.135 176.560 ;
        RECT 54.285 175.910 54.935 176.560 ;
        RECT 55.085 175.910 55.735 176.560 ;
        RECT 69.535 175.910 70.185 176.560 ;
        RECT 70.335 175.910 70.985 176.560 ;
        RECT 71.135 175.910 71.785 176.560 ;
        RECT 73.485 175.910 74.135 176.560 ;
        RECT 74.285 175.910 74.935 176.560 ;
        RECT 75.085 175.910 75.735 176.560 ;
        RECT 89.535 175.910 90.185 176.560 ;
        RECT 90.335 175.910 90.985 176.560 ;
        RECT 91.135 175.910 91.785 176.560 ;
        RECT 93.485 175.910 94.135 176.560 ;
        RECT 94.285 175.910 94.935 176.560 ;
        RECT 95.085 175.910 95.735 176.560 ;
        RECT 109.535 175.910 110.185 176.560 ;
        RECT 110.335 175.910 110.985 176.560 ;
        RECT 111.135 175.910 111.785 176.560 ;
        RECT 113.485 175.910 114.135 176.560 ;
        RECT 114.285 175.910 114.935 176.560 ;
        RECT 115.085 175.910 115.735 176.560 ;
        RECT 0.075 172.535 0.495 172.935 ;
        RECT 0.645 172.535 1.065 172.935 ;
        RECT 1.215 172.535 1.635 172.935 ;
        RECT 42.735 169.110 43.385 169.760 ;
        RECT 42.735 168.310 43.385 168.960 ;
        RECT 0.075 167.095 0.495 167.495 ;
        RECT 0.645 167.095 1.065 167.495 ;
        RECT 1.215 167.095 1.635 167.495 ;
        RECT 42.735 167.510 43.385 168.160 ;
        RECT 42.735 165.160 43.385 165.810 ;
        RECT 42.735 164.360 43.385 165.010 ;
        RECT 42.735 163.560 43.385 164.210 ;
        RECT 61.885 169.110 62.535 169.760 ;
        RECT 62.735 169.110 63.385 169.760 ;
        RECT 61.885 168.310 62.535 168.960 ;
        RECT 62.735 168.310 63.385 168.960 ;
        RECT 61.885 167.510 62.535 168.160 ;
        RECT 62.735 167.510 63.385 168.160 ;
        RECT 61.885 165.160 62.535 165.810 ;
        RECT 62.735 165.160 63.385 165.810 ;
        RECT 61.885 164.360 62.535 165.010 ;
        RECT 62.735 164.360 63.385 165.010 ;
        RECT 61.885 163.560 62.535 164.210 ;
        RECT 62.735 163.560 63.385 164.210 ;
        RECT 81.885 169.110 82.535 169.760 ;
        RECT 82.735 169.110 83.385 169.760 ;
        RECT 81.885 168.310 82.535 168.960 ;
        RECT 82.735 168.310 83.385 168.960 ;
        RECT 81.885 167.510 82.535 168.160 ;
        RECT 82.735 167.510 83.385 168.160 ;
        RECT 81.885 165.160 82.535 165.810 ;
        RECT 82.735 165.160 83.385 165.810 ;
        RECT 81.885 164.360 82.535 165.010 ;
        RECT 82.735 164.360 83.385 165.010 ;
        RECT 81.885 163.560 82.535 164.210 ;
        RECT 82.735 163.560 83.385 164.210 ;
        RECT 101.885 169.110 102.535 169.760 ;
        RECT 102.735 169.110 103.385 169.760 ;
        RECT 101.885 168.310 102.535 168.960 ;
        RECT 102.735 168.310 103.385 168.960 ;
        RECT 101.885 167.510 102.535 168.160 ;
        RECT 102.735 167.510 103.385 168.160 ;
        RECT 101.885 165.160 102.535 165.810 ;
        RECT 102.735 165.160 103.385 165.810 ;
        RECT 101.885 164.360 102.535 165.010 ;
        RECT 102.735 164.360 103.385 165.010 ;
        RECT 101.885 163.560 102.535 164.210 ;
        RECT 102.735 163.560 103.385 164.210 ;
        RECT 121.885 169.110 122.535 169.760 ;
        RECT 121.885 168.310 122.535 168.960 ;
        RECT 121.885 167.510 122.535 168.160 ;
        RECT 122.800 166.980 123.200 167.380 ;
        RECT 123.425 166.980 123.825 167.380 ;
        RECT 124.050 166.980 124.450 167.380 ;
        RECT 122.795 166.380 123.195 166.780 ;
        RECT 123.420 166.380 123.820 166.780 ;
        RECT 124.045 166.380 124.445 166.780 ;
        RECT 127.675 166.980 128.075 167.380 ;
        RECT 128.300 166.980 128.700 167.380 ;
        RECT 128.925 166.980 129.325 167.380 ;
        RECT 127.670 166.380 128.070 166.780 ;
        RECT 128.295 166.380 128.695 166.780 ;
        RECT 128.920 166.380 129.320 166.780 ;
        RECT 121.885 165.160 122.535 165.810 ;
        RECT 121.885 164.360 122.535 165.010 ;
        RECT 121.885 163.560 122.535 164.210 ;
        RECT 49.535 156.760 50.185 157.410 ;
        RECT 50.335 156.760 50.985 157.410 ;
        RECT 51.135 156.760 51.785 157.410 ;
        RECT 53.485 156.760 54.135 157.410 ;
        RECT 54.285 156.760 54.935 157.410 ;
        RECT 55.085 156.760 55.735 157.410 ;
        RECT 69.535 156.760 70.185 157.410 ;
        RECT 70.335 156.760 70.985 157.410 ;
        RECT 71.135 156.760 71.785 157.410 ;
        RECT 73.485 156.760 74.135 157.410 ;
        RECT 74.285 156.760 74.935 157.410 ;
        RECT 75.085 156.760 75.735 157.410 ;
        RECT 89.535 156.760 90.185 157.410 ;
        RECT 90.335 156.760 90.985 157.410 ;
        RECT 91.135 156.760 91.785 157.410 ;
        RECT 93.485 156.760 94.135 157.410 ;
        RECT 94.285 156.760 94.935 157.410 ;
        RECT 95.085 156.760 95.735 157.410 ;
        RECT 109.535 156.760 110.185 157.410 ;
        RECT 110.335 156.760 110.985 157.410 ;
        RECT 111.135 156.760 111.785 157.410 ;
        RECT 113.485 156.760 114.135 157.410 ;
        RECT 114.285 156.760 114.935 157.410 ;
        RECT 115.085 156.760 115.735 157.410 ;
      LAYER met4 ;
        RECT 0.000 0.000 2.000 340.000 ;
        RECT 49.435 175.210 55.835 176.660 ;
        RECT 69.435 175.210 75.835 176.660 ;
        RECT 89.435 175.210 95.835 176.660 ;
        RECT 109.435 175.210 115.835 176.660 ;
        RECT 44.085 169.860 61.185 175.210 ;
        RECT 64.085 169.860 81.185 175.210 ;
        RECT 84.085 169.860 101.185 175.210 ;
        RECT 104.085 169.860 121.185 175.210 ;
        RECT 42.635 167.510 122.635 169.860 ;
        RECT 42.635 166.235 124.635 167.510 ;
        RECT 42.635 163.460 122.635 166.235 ;
        RECT 44.085 158.110 61.185 163.460 ;
        RECT 64.085 158.110 81.185 163.460 ;
        RECT 84.085 158.110 101.185 163.460 ;
        RECT 104.085 158.110 121.185 163.460 ;
        RECT 49.435 156.660 55.835 158.110 ;
        RECT 69.435 156.660 75.835 158.110 ;
        RECT 89.435 156.660 95.835 158.110 ;
        RECT 109.435 156.660 115.835 158.110 ;
        RECT 127.510 0.000 129.510 340.000 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER pwell ;
        RECT 9.130 339.100 11.530 340.000 ;
        RECT 17.930 339.100 20.330 340.000 ;
        RECT 29.130 339.100 31.530 340.000 ;
        RECT 37.930 339.100 40.330 340.000 ;
        RECT 49.130 339.100 51.530 340.000 ;
        RECT 57.930 339.100 60.330 340.000 ;
        RECT 69.130 339.100 71.530 340.000 ;
        RECT 77.930 339.100 80.330 340.000 ;
        RECT 89.130 339.100 91.530 340.000 ;
        RECT 97.930 339.100 100.330 340.000 ;
        RECT 109.130 339.100 111.530 340.000 ;
        RECT 117.930 339.100 120.330 340.000 ;
        RECT 5.880 338.900 23.830 339.100 ;
        RECT 25.880 338.900 43.830 339.100 ;
        RECT 45.880 338.900 63.830 339.100 ;
        RECT 65.880 338.900 83.830 339.100 ;
        RECT 85.880 338.900 103.830 339.100 ;
        RECT 105.880 338.900 123.830 339.100 ;
        RECT 5.830 338.800 23.830 338.900 ;
        RECT 25.830 338.800 43.830 338.900 ;
        RECT 45.830 338.800 63.830 338.900 ;
        RECT 65.830 338.800 83.830 338.900 ;
        RECT 85.830 338.800 103.830 338.900 ;
        RECT 105.830 338.800 123.830 338.900 ;
        RECT 5.680 335.600 23.830 338.800 ;
        RECT 25.680 335.600 43.830 338.800 ;
        RECT 45.680 335.600 63.830 338.800 ;
        RECT 65.680 335.600 83.830 338.800 ;
        RECT 85.680 335.600 103.830 338.800 ;
        RECT 105.680 335.600 123.830 338.800 ;
        RECT 4.730 333.200 124.730 335.600 ;
        RECT 5.630 326.800 23.830 333.200 ;
        RECT 25.630 326.800 43.830 333.200 ;
        RECT 45.630 326.800 63.830 333.200 ;
        RECT 65.630 326.800 83.830 333.200 ;
        RECT 85.630 326.800 103.830 333.200 ;
        RECT 105.630 326.800 123.830 333.200 ;
        RECT 4.730 324.400 124.730 326.800 ;
        RECT 5.630 320.900 23.830 324.400 ;
        RECT 25.630 320.900 43.830 324.400 ;
        RECT 45.630 320.900 63.830 324.400 ;
        RECT 65.630 320.900 83.830 324.400 ;
        RECT 85.630 320.900 103.830 324.400 ;
        RECT 105.630 320.900 123.830 324.400 ;
        RECT 9.130 319.100 11.530 320.900 ;
        RECT 17.930 319.100 20.330 320.900 ;
        RECT 29.130 319.100 31.530 320.900 ;
        RECT 37.930 319.100 40.330 320.900 ;
        RECT 49.130 319.100 51.530 320.900 ;
        RECT 57.930 319.100 60.330 320.900 ;
        RECT 69.130 319.100 71.530 320.900 ;
        RECT 77.930 319.100 80.330 320.900 ;
        RECT 89.130 319.100 91.530 320.900 ;
        RECT 97.930 319.100 100.330 320.900 ;
        RECT 109.130 319.100 111.530 320.900 ;
        RECT 117.930 319.100 120.330 320.900 ;
        RECT 5.880 318.900 23.830 319.100 ;
        RECT 25.880 318.900 43.830 319.100 ;
        RECT 45.880 318.900 63.830 319.100 ;
        RECT 65.880 318.900 83.830 319.100 ;
        RECT 85.880 318.900 103.830 319.100 ;
        RECT 105.880 318.900 123.830 319.100 ;
        RECT 5.830 318.800 23.830 318.900 ;
        RECT 25.830 318.800 43.830 318.900 ;
        RECT 45.830 318.800 63.830 318.900 ;
        RECT 65.830 318.800 83.830 318.900 ;
        RECT 85.830 318.800 103.830 318.900 ;
        RECT 105.830 318.800 123.830 318.900 ;
        RECT 5.680 315.600 23.830 318.800 ;
        RECT 25.680 315.600 43.830 318.800 ;
        RECT 45.680 315.600 63.830 318.800 ;
        RECT 65.680 315.600 83.830 318.800 ;
        RECT 85.680 315.600 103.830 318.800 ;
        RECT 105.680 315.600 123.830 318.800 ;
        RECT 4.730 313.200 124.730 315.600 ;
        RECT 5.630 306.800 23.830 313.200 ;
        RECT 25.630 306.800 43.830 313.200 ;
        RECT 45.630 306.800 63.830 313.200 ;
        RECT 65.630 306.800 83.830 313.200 ;
        RECT 85.630 306.800 103.830 313.200 ;
        RECT 105.630 306.800 123.830 313.200 ;
        RECT 4.730 304.400 124.730 306.800 ;
        RECT 5.630 300.900 23.830 304.400 ;
        RECT 25.630 300.900 43.830 304.400 ;
        RECT 45.630 300.900 63.830 304.400 ;
        RECT 65.630 300.900 83.830 304.400 ;
        RECT 85.630 300.900 103.830 304.400 ;
        RECT 105.630 300.900 123.830 304.400 ;
        RECT 9.130 299.100 11.530 300.900 ;
        RECT 17.930 299.100 20.330 300.900 ;
        RECT 29.130 299.100 31.530 300.900 ;
        RECT 37.930 299.100 40.330 300.900 ;
        RECT 49.130 299.100 51.530 300.900 ;
        RECT 57.930 299.100 60.330 300.900 ;
        RECT 69.130 299.100 71.530 300.900 ;
        RECT 77.930 299.100 80.330 300.900 ;
        RECT 89.130 299.100 91.530 300.900 ;
        RECT 97.930 299.100 100.330 300.900 ;
        RECT 109.130 299.100 111.530 300.900 ;
        RECT 117.930 299.100 120.330 300.900 ;
        RECT 5.880 298.900 23.830 299.100 ;
        RECT 25.880 298.900 43.830 299.100 ;
        RECT 45.880 298.900 63.830 299.100 ;
        RECT 65.880 298.900 83.830 299.100 ;
        RECT 85.880 298.900 103.830 299.100 ;
        RECT 105.880 298.900 123.830 299.100 ;
        RECT 5.830 298.800 23.830 298.900 ;
        RECT 25.830 298.800 43.830 298.900 ;
        RECT 45.830 298.800 63.830 298.900 ;
        RECT 65.830 298.800 83.830 298.900 ;
        RECT 85.830 298.800 103.830 298.900 ;
        RECT 105.830 298.800 123.830 298.900 ;
        RECT 5.680 295.600 23.830 298.800 ;
        RECT 25.680 295.600 43.830 298.800 ;
        RECT 45.680 295.600 63.830 298.800 ;
        RECT 65.680 295.600 83.830 298.800 ;
        RECT 85.680 295.600 103.830 298.800 ;
        RECT 105.680 295.600 123.830 298.800 ;
        RECT 4.730 293.200 124.730 295.600 ;
        RECT 5.630 286.800 23.830 293.200 ;
        RECT 25.630 286.800 43.830 293.200 ;
        RECT 45.630 286.800 63.830 293.200 ;
        RECT 65.630 286.800 83.830 293.200 ;
        RECT 85.630 286.800 103.830 293.200 ;
        RECT 105.630 286.800 123.830 293.200 ;
        RECT 4.730 284.400 124.730 286.800 ;
        RECT 5.630 280.900 23.830 284.400 ;
        RECT 25.630 280.900 43.830 284.400 ;
        RECT 45.630 280.900 63.830 284.400 ;
        RECT 65.630 280.900 83.830 284.400 ;
        RECT 85.630 280.900 103.830 284.400 ;
        RECT 105.630 280.900 123.830 284.400 ;
        RECT 9.130 279.100 11.530 280.900 ;
        RECT 17.930 279.100 20.330 280.900 ;
        RECT 29.130 279.100 31.530 280.900 ;
        RECT 37.930 279.100 40.330 280.900 ;
        RECT 49.130 279.100 51.530 280.900 ;
        RECT 57.930 279.100 60.330 280.900 ;
        RECT 69.130 279.100 71.530 280.900 ;
        RECT 77.930 279.100 80.330 280.900 ;
        RECT 89.130 279.100 91.530 280.900 ;
        RECT 97.930 279.100 100.330 280.900 ;
        RECT 109.130 279.100 111.530 280.900 ;
        RECT 117.930 279.100 120.330 280.900 ;
        RECT 5.880 278.900 23.830 279.100 ;
        RECT 25.880 278.900 43.830 279.100 ;
        RECT 45.880 278.900 63.830 279.100 ;
        RECT 65.880 278.900 83.830 279.100 ;
        RECT 85.880 278.900 103.830 279.100 ;
        RECT 105.880 278.900 123.830 279.100 ;
        RECT 5.830 278.800 23.830 278.900 ;
        RECT 25.830 278.800 43.830 278.900 ;
        RECT 45.830 278.800 63.830 278.900 ;
        RECT 65.830 278.800 83.830 278.900 ;
        RECT 85.830 278.800 103.830 278.900 ;
        RECT 105.830 278.800 123.830 278.900 ;
        RECT 5.680 275.600 23.830 278.800 ;
        RECT 25.680 275.600 43.830 278.800 ;
        RECT 45.680 275.600 63.830 278.800 ;
        RECT 65.680 275.600 83.830 278.800 ;
        RECT 85.680 275.600 103.830 278.800 ;
        RECT 105.680 275.600 123.830 278.800 ;
        RECT 4.730 273.200 124.730 275.600 ;
        RECT 5.630 266.800 23.830 273.200 ;
        RECT 25.630 266.800 43.830 273.200 ;
        RECT 45.630 266.800 63.830 273.200 ;
        RECT 65.630 266.800 83.830 273.200 ;
        RECT 85.630 266.800 103.830 273.200 ;
        RECT 105.630 266.800 123.830 273.200 ;
        RECT 4.730 264.400 124.730 266.800 ;
        RECT 5.630 260.900 23.830 264.400 ;
        RECT 25.630 260.900 43.830 264.400 ;
        RECT 45.630 260.900 63.830 264.400 ;
        RECT 65.630 260.900 83.830 264.400 ;
        RECT 85.630 260.900 103.830 264.400 ;
        RECT 105.630 260.900 123.830 264.400 ;
        RECT 9.130 259.100 11.530 260.900 ;
        RECT 17.930 259.100 20.330 260.900 ;
        RECT 29.130 259.100 31.530 260.900 ;
        RECT 37.930 259.100 40.330 260.900 ;
        RECT 49.130 259.100 51.530 260.900 ;
        RECT 57.930 259.100 60.330 260.900 ;
        RECT 69.130 259.100 71.530 260.900 ;
        RECT 77.930 259.100 80.330 260.900 ;
        RECT 89.130 259.100 91.530 260.900 ;
        RECT 97.930 259.100 100.330 260.900 ;
        RECT 109.130 259.100 111.530 260.900 ;
        RECT 117.930 259.100 120.330 260.900 ;
        RECT 5.880 258.900 23.830 259.100 ;
        RECT 25.880 258.900 43.830 259.100 ;
        RECT 45.880 258.900 63.830 259.100 ;
        RECT 65.880 258.900 83.830 259.100 ;
        RECT 85.880 258.900 103.830 259.100 ;
        RECT 105.880 258.900 123.830 259.100 ;
        RECT 5.830 258.800 23.830 258.900 ;
        RECT 25.830 258.800 43.830 258.900 ;
        RECT 45.830 258.800 63.830 258.900 ;
        RECT 65.830 258.800 83.830 258.900 ;
        RECT 85.830 258.800 103.830 258.900 ;
        RECT 105.830 258.800 123.830 258.900 ;
        RECT 5.680 255.600 23.830 258.800 ;
        RECT 25.680 255.600 43.830 258.800 ;
        RECT 45.680 255.600 63.830 258.800 ;
        RECT 65.680 255.600 83.830 258.800 ;
        RECT 85.680 255.600 103.830 258.800 ;
        RECT 105.680 255.600 123.830 258.800 ;
        RECT 4.730 253.200 124.730 255.600 ;
        RECT 5.630 246.800 23.830 253.200 ;
        RECT 25.630 246.800 43.830 253.200 ;
        RECT 45.630 246.800 63.830 253.200 ;
        RECT 65.630 246.800 83.830 253.200 ;
        RECT 85.630 246.800 103.830 253.200 ;
        RECT 105.630 246.800 123.830 253.200 ;
        RECT 4.730 244.400 124.730 246.800 ;
        RECT 5.630 240.900 23.830 244.400 ;
        RECT 25.630 240.900 43.830 244.400 ;
        RECT 45.630 240.900 63.830 244.400 ;
        RECT 65.630 240.900 83.830 244.400 ;
        RECT 85.630 240.900 103.830 244.400 ;
        RECT 105.630 240.900 123.830 244.400 ;
        RECT 9.130 239.100 11.530 240.900 ;
        RECT 17.930 239.100 20.330 240.900 ;
        RECT 29.130 239.100 31.530 240.900 ;
        RECT 37.930 239.100 40.330 240.900 ;
        RECT 49.130 239.100 51.530 240.900 ;
        RECT 57.930 239.100 60.330 240.900 ;
        RECT 69.130 239.100 71.530 240.900 ;
        RECT 77.930 239.100 80.330 240.900 ;
        RECT 89.130 239.100 91.530 240.900 ;
        RECT 97.930 239.100 100.330 240.900 ;
        RECT 109.130 239.100 111.530 240.900 ;
        RECT 117.930 239.100 120.330 240.900 ;
        RECT 5.880 238.900 23.830 239.100 ;
        RECT 25.880 238.900 43.830 239.100 ;
        RECT 45.880 238.900 63.830 239.100 ;
        RECT 65.880 238.900 83.830 239.100 ;
        RECT 85.880 238.900 103.830 239.100 ;
        RECT 105.880 238.900 123.830 239.100 ;
        RECT 5.830 238.800 23.830 238.900 ;
        RECT 25.830 238.800 43.830 238.900 ;
        RECT 45.830 238.800 63.830 238.900 ;
        RECT 65.830 238.800 83.830 238.900 ;
        RECT 85.830 238.800 103.830 238.900 ;
        RECT 105.830 238.800 123.830 238.900 ;
        RECT 5.680 235.600 23.830 238.800 ;
        RECT 25.680 235.600 43.830 238.800 ;
        RECT 45.680 235.600 63.830 238.800 ;
        RECT 65.680 235.600 83.830 238.800 ;
        RECT 85.680 235.600 103.830 238.800 ;
        RECT 105.680 235.600 123.830 238.800 ;
        RECT 4.730 233.200 124.730 235.600 ;
        RECT 5.630 226.800 23.830 233.200 ;
        RECT 25.630 226.800 43.830 233.200 ;
        RECT 45.630 226.800 63.830 233.200 ;
        RECT 65.630 226.800 83.830 233.200 ;
        RECT 85.630 226.800 103.830 233.200 ;
        RECT 105.630 226.800 123.830 233.200 ;
        RECT 4.730 224.400 124.730 226.800 ;
        RECT 5.630 220.900 23.830 224.400 ;
        RECT 25.630 220.900 43.830 224.400 ;
        RECT 45.630 220.900 63.830 224.400 ;
        RECT 65.630 220.900 83.830 224.400 ;
        RECT 85.630 220.900 103.830 224.400 ;
        RECT 105.630 220.900 123.830 224.400 ;
        RECT 9.130 219.100 11.530 220.900 ;
        RECT 17.930 219.100 20.330 220.900 ;
        RECT 29.130 219.100 31.530 220.900 ;
        RECT 37.930 219.100 40.330 220.900 ;
        RECT 49.130 219.100 51.530 220.900 ;
        RECT 57.930 219.100 60.330 220.900 ;
        RECT 69.130 219.100 71.530 220.900 ;
        RECT 77.930 219.100 80.330 220.900 ;
        RECT 89.130 219.100 91.530 220.900 ;
        RECT 97.930 219.100 100.330 220.900 ;
        RECT 109.130 219.100 111.530 220.900 ;
        RECT 117.930 219.100 120.330 220.900 ;
        RECT 5.880 218.900 23.830 219.100 ;
        RECT 25.880 218.900 43.830 219.100 ;
        RECT 45.880 218.900 63.830 219.100 ;
        RECT 65.880 218.900 83.830 219.100 ;
        RECT 85.880 218.900 103.830 219.100 ;
        RECT 105.880 218.900 123.830 219.100 ;
        RECT 5.830 218.800 23.830 218.900 ;
        RECT 25.830 218.800 43.830 218.900 ;
        RECT 45.830 218.800 63.830 218.900 ;
        RECT 65.830 218.800 83.830 218.900 ;
        RECT 85.830 218.800 103.830 218.900 ;
        RECT 105.830 218.800 123.830 218.900 ;
        RECT 5.680 215.600 23.830 218.800 ;
        RECT 25.680 215.600 43.830 218.800 ;
        RECT 45.680 215.600 63.830 218.800 ;
        RECT 65.680 215.600 83.830 218.800 ;
        RECT 85.680 215.600 103.830 218.800 ;
        RECT 105.680 215.600 123.830 218.800 ;
        RECT 4.730 213.200 124.730 215.600 ;
        RECT 5.630 206.800 23.830 213.200 ;
        RECT 25.630 206.800 43.830 213.200 ;
        RECT 45.630 206.800 63.830 213.200 ;
        RECT 65.630 206.800 83.830 213.200 ;
        RECT 85.630 206.800 103.830 213.200 ;
        RECT 105.630 206.800 123.830 213.200 ;
        RECT 4.730 204.400 124.730 206.800 ;
        RECT 5.630 200.900 23.830 204.400 ;
        RECT 25.630 200.900 43.830 204.400 ;
        RECT 45.630 200.900 63.830 204.400 ;
        RECT 65.630 200.900 83.830 204.400 ;
        RECT 85.630 200.900 103.830 204.400 ;
        RECT 105.630 200.900 123.830 204.400 ;
        RECT 9.130 200.000 11.530 200.900 ;
        RECT 17.930 200.000 20.330 200.900 ;
        RECT 29.130 200.000 31.530 200.900 ;
        RECT 37.930 200.000 40.330 200.900 ;
        RECT 49.130 200.000 51.530 200.900 ;
        RECT 57.930 200.000 60.330 200.900 ;
        RECT 69.130 200.000 71.530 200.900 ;
        RECT 77.930 200.000 80.330 200.900 ;
        RECT 89.130 200.000 91.530 200.900 ;
        RECT 97.930 200.000 100.330 200.900 ;
        RECT 109.130 200.000 111.530 200.900 ;
        RECT 117.930 200.000 120.330 200.900 ;
        RECT 47.035 175.760 49.435 176.660 ;
        RECT 55.835 175.760 58.235 176.660 ;
        RECT 67.035 175.760 69.435 176.660 ;
        RECT 75.835 175.760 78.235 176.660 ;
        RECT 87.035 175.760 89.435 176.660 ;
        RECT 95.835 175.760 98.235 176.660 ;
        RECT 107.035 175.760 109.435 176.660 ;
        RECT 115.835 175.760 118.235 176.660 ;
        RECT 43.785 175.560 61.735 175.760 ;
        RECT 63.785 175.560 81.735 175.760 ;
        RECT 83.785 175.560 101.735 175.760 ;
        RECT 103.785 175.560 121.735 175.760 ;
        RECT 43.735 175.460 61.735 175.560 ;
        RECT 63.735 175.460 81.735 175.560 ;
        RECT 83.735 175.460 101.735 175.560 ;
        RECT 103.735 175.460 121.735 175.560 ;
        RECT 7.115 174.485 7.545 175.270 ;
        RECT 14.880 174.480 15.310 175.265 ;
        RECT 43.585 172.260 61.735 175.460 ;
        RECT 63.585 172.260 81.735 175.460 ;
        RECT 83.585 172.260 101.735 175.460 ;
        RECT 103.585 172.260 121.735 175.460 ;
        RECT 7.980 170.205 8.410 170.990 ;
        RECT 23.620 170.205 24.050 170.990 ;
        RECT 42.635 169.860 122.635 172.260 ;
        RECT 6.600 169.040 7.030 169.825 ;
        RECT 23.620 169.040 24.050 169.825 ;
        RECT 7.520 164.765 7.950 165.550 ;
        RECT 14.880 164.765 15.310 165.550 ;
        RECT 43.535 163.460 61.735 169.860 ;
        RECT 63.535 163.460 81.735 169.860 ;
        RECT 83.535 163.460 101.735 169.860 ;
        RECT 103.535 163.460 121.735 169.860 ;
        RECT 42.635 161.060 122.635 163.460 ;
        RECT 43.535 157.560 61.735 161.060 ;
        RECT 63.535 157.560 81.735 161.060 ;
        RECT 83.535 157.560 101.735 161.060 ;
        RECT 103.535 157.560 121.735 161.060 ;
        RECT 47.035 156.660 49.435 157.560 ;
        RECT 55.835 156.660 58.235 157.560 ;
        RECT 67.035 156.660 69.435 157.560 ;
        RECT 75.835 156.660 78.235 157.560 ;
        RECT 87.035 156.660 89.435 157.560 ;
        RECT 95.835 156.660 98.235 157.560 ;
        RECT 107.035 156.660 109.435 157.560 ;
        RECT 115.835 156.660 118.235 157.560 ;
        RECT 9.130 139.100 11.530 140.000 ;
        RECT 17.930 139.100 20.330 140.000 ;
        RECT 29.130 139.100 31.530 140.000 ;
        RECT 37.930 139.100 40.330 140.000 ;
        RECT 49.130 139.100 51.530 140.000 ;
        RECT 57.930 139.100 60.330 140.000 ;
        RECT 69.130 139.100 71.530 140.000 ;
        RECT 77.930 139.100 80.330 140.000 ;
        RECT 89.130 139.100 91.530 140.000 ;
        RECT 97.930 139.100 100.330 140.000 ;
        RECT 109.130 139.100 111.530 140.000 ;
        RECT 117.930 139.100 120.330 140.000 ;
        RECT 5.880 138.900 23.830 139.100 ;
        RECT 25.880 138.900 43.830 139.100 ;
        RECT 45.880 138.900 63.830 139.100 ;
        RECT 65.880 138.900 83.830 139.100 ;
        RECT 85.880 138.900 103.830 139.100 ;
        RECT 105.880 138.900 123.830 139.100 ;
        RECT 5.830 138.800 23.830 138.900 ;
        RECT 25.830 138.800 43.830 138.900 ;
        RECT 45.830 138.800 63.830 138.900 ;
        RECT 65.830 138.800 83.830 138.900 ;
        RECT 85.830 138.800 103.830 138.900 ;
        RECT 105.830 138.800 123.830 138.900 ;
        RECT 5.680 135.600 23.830 138.800 ;
        RECT 25.680 135.600 43.830 138.800 ;
        RECT 45.680 135.600 63.830 138.800 ;
        RECT 65.680 135.600 83.830 138.800 ;
        RECT 85.680 135.600 103.830 138.800 ;
        RECT 105.680 135.600 123.830 138.800 ;
        RECT 4.730 133.200 124.730 135.600 ;
        RECT 5.630 126.800 23.830 133.200 ;
        RECT 25.630 126.800 43.830 133.200 ;
        RECT 45.630 126.800 63.830 133.200 ;
        RECT 65.630 126.800 83.830 133.200 ;
        RECT 85.630 126.800 103.830 133.200 ;
        RECT 105.630 126.800 123.830 133.200 ;
        RECT 4.730 124.400 124.730 126.800 ;
        RECT 5.630 120.900 23.830 124.400 ;
        RECT 25.630 120.900 43.830 124.400 ;
        RECT 45.630 120.900 63.830 124.400 ;
        RECT 65.630 120.900 83.830 124.400 ;
        RECT 85.630 120.900 103.830 124.400 ;
        RECT 105.630 120.900 123.830 124.400 ;
        RECT 9.130 119.100 11.530 120.900 ;
        RECT 17.930 119.100 20.330 120.900 ;
        RECT 29.130 119.100 31.530 120.900 ;
        RECT 37.930 119.100 40.330 120.900 ;
        RECT 49.130 119.100 51.530 120.900 ;
        RECT 57.930 119.100 60.330 120.900 ;
        RECT 69.130 119.100 71.530 120.900 ;
        RECT 77.930 119.100 80.330 120.900 ;
        RECT 89.130 119.100 91.530 120.900 ;
        RECT 97.930 119.100 100.330 120.900 ;
        RECT 109.130 119.100 111.530 120.900 ;
        RECT 117.930 119.100 120.330 120.900 ;
        RECT 5.880 118.900 23.830 119.100 ;
        RECT 25.880 118.900 43.830 119.100 ;
        RECT 45.880 118.900 63.830 119.100 ;
        RECT 65.880 118.900 83.830 119.100 ;
        RECT 85.880 118.900 103.830 119.100 ;
        RECT 105.880 118.900 123.830 119.100 ;
        RECT 5.830 118.800 23.830 118.900 ;
        RECT 25.830 118.800 43.830 118.900 ;
        RECT 45.830 118.800 63.830 118.900 ;
        RECT 65.830 118.800 83.830 118.900 ;
        RECT 85.830 118.800 103.830 118.900 ;
        RECT 105.830 118.800 123.830 118.900 ;
        RECT 5.680 115.600 23.830 118.800 ;
        RECT 25.680 115.600 43.830 118.800 ;
        RECT 45.680 115.600 63.830 118.800 ;
        RECT 65.680 115.600 83.830 118.800 ;
        RECT 85.680 115.600 103.830 118.800 ;
        RECT 105.680 115.600 123.830 118.800 ;
        RECT 4.730 113.200 124.730 115.600 ;
        RECT 5.630 106.800 23.830 113.200 ;
        RECT 25.630 106.800 43.830 113.200 ;
        RECT 45.630 106.800 63.830 113.200 ;
        RECT 65.630 106.800 83.830 113.200 ;
        RECT 85.630 106.800 103.830 113.200 ;
        RECT 105.630 106.800 123.830 113.200 ;
        RECT 4.730 104.400 124.730 106.800 ;
        RECT 5.630 100.900 23.830 104.400 ;
        RECT 25.630 100.900 43.830 104.400 ;
        RECT 45.630 100.900 63.830 104.400 ;
        RECT 65.630 100.900 83.830 104.400 ;
        RECT 85.630 100.900 103.830 104.400 ;
        RECT 105.630 100.900 123.830 104.400 ;
        RECT 9.130 99.100 11.530 100.900 ;
        RECT 17.930 99.100 20.330 100.900 ;
        RECT 29.130 99.100 31.530 100.900 ;
        RECT 37.930 99.100 40.330 100.900 ;
        RECT 49.130 99.100 51.530 100.900 ;
        RECT 57.930 99.100 60.330 100.900 ;
        RECT 69.130 99.100 71.530 100.900 ;
        RECT 77.930 99.100 80.330 100.900 ;
        RECT 89.130 99.100 91.530 100.900 ;
        RECT 97.930 99.100 100.330 100.900 ;
        RECT 109.130 99.100 111.530 100.900 ;
        RECT 117.930 99.100 120.330 100.900 ;
        RECT 5.880 98.900 23.830 99.100 ;
        RECT 25.880 98.900 43.830 99.100 ;
        RECT 45.880 98.900 63.830 99.100 ;
        RECT 65.880 98.900 83.830 99.100 ;
        RECT 85.880 98.900 103.830 99.100 ;
        RECT 105.880 98.900 123.830 99.100 ;
        RECT 5.830 98.800 23.830 98.900 ;
        RECT 25.830 98.800 43.830 98.900 ;
        RECT 45.830 98.800 63.830 98.900 ;
        RECT 65.830 98.800 83.830 98.900 ;
        RECT 85.830 98.800 103.830 98.900 ;
        RECT 105.830 98.800 123.830 98.900 ;
        RECT 5.680 95.600 23.830 98.800 ;
        RECT 25.680 95.600 43.830 98.800 ;
        RECT 45.680 95.600 63.830 98.800 ;
        RECT 65.680 95.600 83.830 98.800 ;
        RECT 85.680 95.600 103.830 98.800 ;
        RECT 105.680 95.600 123.830 98.800 ;
        RECT 4.730 93.200 124.730 95.600 ;
        RECT 5.630 86.800 23.830 93.200 ;
        RECT 25.630 86.800 43.830 93.200 ;
        RECT 45.630 86.800 63.830 93.200 ;
        RECT 65.630 86.800 83.830 93.200 ;
        RECT 85.630 86.800 103.830 93.200 ;
        RECT 105.630 86.800 123.830 93.200 ;
        RECT 4.730 84.400 124.730 86.800 ;
        RECT 5.630 80.900 23.830 84.400 ;
        RECT 25.630 80.900 43.830 84.400 ;
        RECT 45.630 80.900 63.830 84.400 ;
        RECT 65.630 80.900 83.830 84.400 ;
        RECT 85.630 80.900 103.830 84.400 ;
        RECT 105.630 80.900 123.830 84.400 ;
        RECT 9.130 79.100 11.530 80.900 ;
        RECT 17.930 79.100 20.330 80.900 ;
        RECT 29.130 79.100 31.530 80.900 ;
        RECT 37.930 79.100 40.330 80.900 ;
        RECT 49.130 79.100 51.530 80.900 ;
        RECT 57.930 79.100 60.330 80.900 ;
        RECT 69.130 79.100 71.530 80.900 ;
        RECT 77.930 79.100 80.330 80.900 ;
        RECT 89.130 79.100 91.530 80.900 ;
        RECT 97.930 79.100 100.330 80.900 ;
        RECT 109.130 79.100 111.530 80.900 ;
        RECT 117.930 79.100 120.330 80.900 ;
        RECT 5.880 78.900 23.830 79.100 ;
        RECT 25.880 78.900 43.830 79.100 ;
        RECT 45.880 78.900 63.830 79.100 ;
        RECT 65.880 78.900 83.830 79.100 ;
        RECT 85.880 78.900 103.830 79.100 ;
        RECT 105.880 78.900 123.830 79.100 ;
        RECT 5.830 78.800 23.830 78.900 ;
        RECT 25.830 78.800 43.830 78.900 ;
        RECT 45.830 78.800 63.830 78.900 ;
        RECT 65.830 78.800 83.830 78.900 ;
        RECT 85.830 78.800 103.830 78.900 ;
        RECT 105.830 78.800 123.830 78.900 ;
        RECT 5.680 75.600 23.830 78.800 ;
        RECT 25.680 75.600 43.830 78.800 ;
        RECT 45.680 75.600 63.830 78.800 ;
        RECT 65.680 75.600 83.830 78.800 ;
        RECT 85.680 75.600 103.830 78.800 ;
        RECT 105.680 75.600 123.830 78.800 ;
        RECT 4.730 73.200 124.730 75.600 ;
        RECT 5.630 66.800 23.830 73.200 ;
        RECT 25.630 66.800 43.830 73.200 ;
        RECT 45.630 66.800 63.830 73.200 ;
        RECT 65.630 66.800 83.830 73.200 ;
        RECT 85.630 66.800 103.830 73.200 ;
        RECT 105.630 66.800 123.830 73.200 ;
        RECT 4.730 64.400 124.730 66.800 ;
        RECT 5.630 60.900 23.830 64.400 ;
        RECT 25.630 60.900 43.830 64.400 ;
        RECT 45.630 60.900 63.830 64.400 ;
        RECT 65.630 60.900 83.830 64.400 ;
        RECT 85.630 60.900 103.830 64.400 ;
        RECT 105.630 60.900 123.830 64.400 ;
        RECT 9.130 59.100 11.530 60.900 ;
        RECT 17.930 59.100 20.330 60.900 ;
        RECT 29.130 59.100 31.530 60.900 ;
        RECT 37.930 59.100 40.330 60.900 ;
        RECT 49.130 59.100 51.530 60.900 ;
        RECT 57.930 59.100 60.330 60.900 ;
        RECT 69.130 59.100 71.530 60.900 ;
        RECT 77.930 59.100 80.330 60.900 ;
        RECT 89.130 59.100 91.530 60.900 ;
        RECT 97.930 59.100 100.330 60.900 ;
        RECT 109.130 59.100 111.530 60.900 ;
        RECT 117.930 59.100 120.330 60.900 ;
        RECT 5.880 58.900 23.830 59.100 ;
        RECT 25.880 58.900 43.830 59.100 ;
        RECT 45.880 58.900 63.830 59.100 ;
        RECT 65.880 58.900 83.830 59.100 ;
        RECT 85.880 58.900 103.830 59.100 ;
        RECT 105.880 58.900 123.830 59.100 ;
        RECT 5.830 58.800 23.830 58.900 ;
        RECT 25.830 58.800 43.830 58.900 ;
        RECT 45.830 58.800 63.830 58.900 ;
        RECT 65.830 58.800 83.830 58.900 ;
        RECT 85.830 58.800 103.830 58.900 ;
        RECT 105.830 58.800 123.830 58.900 ;
        RECT 5.680 55.600 23.830 58.800 ;
        RECT 25.680 55.600 43.830 58.800 ;
        RECT 45.680 55.600 63.830 58.800 ;
        RECT 65.680 55.600 83.830 58.800 ;
        RECT 85.680 55.600 103.830 58.800 ;
        RECT 105.680 55.600 123.830 58.800 ;
        RECT 4.730 53.200 124.730 55.600 ;
        RECT 5.630 46.800 23.830 53.200 ;
        RECT 25.630 46.800 43.830 53.200 ;
        RECT 45.630 46.800 63.830 53.200 ;
        RECT 65.630 46.800 83.830 53.200 ;
        RECT 85.630 46.800 103.830 53.200 ;
        RECT 105.630 46.800 123.830 53.200 ;
        RECT 4.730 44.400 124.730 46.800 ;
        RECT 5.630 40.900 23.830 44.400 ;
        RECT 25.630 40.900 43.830 44.400 ;
        RECT 45.630 40.900 63.830 44.400 ;
        RECT 65.630 40.900 83.830 44.400 ;
        RECT 85.630 40.900 103.830 44.400 ;
        RECT 105.630 40.900 123.830 44.400 ;
        RECT 9.130 39.100 11.530 40.900 ;
        RECT 17.930 39.100 20.330 40.900 ;
        RECT 29.130 39.100 31.530 40.900 ;
        RECT 37.930 39.100 40.330 40.900 ;
        RECT 49.130 39.100 51.530 40.900 ;
        RECT 57.930 39.100 60.330 40.900 ;
        RECT 69.130 39.100 71.530 40.900 ;
        RECT 77.930 39.100 80.330 40.900 ;
        RECT 89.130 39.100 91.530 40.900 ;
        RECT 97.930 39.100 100.330 40.900 ;
        RECT 109.130 39.100 111.530 40.900 ;
        RECT 117.930 39.100 120.330 40.900 ;
        RECT 5.880 38.900 23.830 39.100 ;
        RECT 25.880 38.900 43.830 39.100 ;
        RECT 45.880 38.900 63.830 39.100 ;
        RECT 65.880 38.900 83.830 39.100 ;
        RECT 85.880 38.900 103.830 39.100 ;
        RECT 105.880 38.900 123.830 39.100 ;
        RECT 5.830 38.800 23.830 38.900 ;
        RECT 25.830 38.800 43.830 38.900 ;
        RECT 45.830 38.800 63.830 38.900 ;
        RECT 65.830 38.800 83.830 38.900 ;
        RECT 85.830 38.800 103.830 38.900 ;
        RECT 105.830 38.800 123.830 38.900 ;
        RECT 5.680 35.600 23.830 38.800 ;
        RECT 25.680 35.600 43.830 38.800 ;
        RECT 45.680 35.600 63.830 38.800 ;
        RECT 65.680 35.600 83.830 38.800 ;
        RECT 85.680 35.600 103.830 38.800 ;
        RECT 105.680 35.600 123.830 38.800 ;
        RECT 4.730 33.200 124.730 35.600 ;
        RECT 5.630 26.800 23.830 33.200 ;
        RECT 25.630 26.800 43.830 33.200 ;
        RECT 45.630 26.800 63.830 33.200 ;
        RECT 65.630 26.800 83.830 33.200 ;
        RECT 85.630 26.800 103.830 33.200 ;
        RECT 105.630 26.800 123.830 33.200 ;
        RECT 4.730 24.400 124.730 26.800 ;
        RECT 5.630 20.900 23.830 24.400 ;
        RECT 25.630 20.900 43.830 24.400 ;
        RECT 45.630 20.900 63.830 24.400 ;
        RECT 65.630 20.900 83.830 24.400 ;
        RECT 85.630 20.900 103.830 24.400 ;
        RECT 105.630 20.900 123.830 24.400 ;
        RECT 9.130 19.100 11.530 20.900 ;
        RECT 17.930 19.100 20.330 20.900 ;
        RECT 29.130 19.100 31.530 20.900 ;
        RECT 37.930 19.100 40.330 20.900 ;
        RECT 49.130 19.100 51.530 20.900 ;
        RECT 57.930 19.100 60.330 20.900 ;
        RECT 69.130 19.100 71.530 20.900 ;
        RECT 77.930 19.100 80.330 20.900 ;
        RECT 89.130 19.100 91.530 20.900 ;
        RECT 97.930 19.100 100.330 20.900 ;
        RECT 109.130 19.100 111.530 20.900 ;
        RECT 117.930 19.100 120.330 20.900 ;
        RECT 5.880 18.900 23.830 19.100 ;
        RECT 25.880 18.900 43.830 19.100 ;
        RECT 45.880 18.900 63.830 19.100 ;
        RECT 65.880 18.900 83.830 19.100 ;
        RECT 85.880 18.900 103.830 19.100 ;
        RECT 105.880 18.900 123.830 19.100 ;
        RECT 5.830 18.800 23.830 18.900 ;
        RECT 25.830 18.800 43.830 18.900 ;
        RECT 45.830 18.800 63.830 18.900 ;
        RECT 65.830 18.800 83.830 18.900 ;
        RECT 85.830 18.800 103.830 18.900 ;
        RECT 105.830 18.800 123.830 18.900 ;
        RECT 5.680 15.600 23.830 18.800 ;
        RECT 25.680 15.600 43.830 18.800 ;
        RECT 45.680 15.600 63.830 18.800 ;
        RECT 65.680 15.600 83.830 18.800 ;
        RECT 85.680 15.600 103.830 18.800 ;
        RECT 105.680 15.600 123.830 18.800 ;
        RECT 4.730 13.200 124.730 15.600 ;
        RECT 5.630 6.800 23.830 13.200 ;
        RECT 25.630 6.800 43.830 13.200 ;
        RECT 45.630 6.800 63.830 13.200 ;
        RECT 65.630 6.800 83.830 13.200 ;
        RECT 85.630 6.800 103.830 13.200 ;
        RECT 105.630 6.800 123.830 13.200 ;
        RECT 4.730 4.400 124.730 6.800 ;
        RECT 5.630 0.900 23.830 4.400 ;
        RECT 25.630 0.900 43.830 4.400 ;
        RECT 45.630 0.900 63.830 4.400 ;
        RECT 65.630 0.900 83.830 4.400 ;
        RECT 85.630 0.900 103.830 4.400 ;
        RECT 105.630 0.900 123.830 4.400 ;
        RECT 9.130 0.000 11.530 0.900 ;
        RECT 17.930 0.000 20.330 0.900 ;
        RECT 29.130 0.000 31.530 0.900 ;
        RECT 37.930 0.000 40.330 0.900 ;
        RECT 49.130 0.000 51.530 0.900 ;
        RECT 57.930 0.000 60.330 0.900 ;
        RECT 69.130 0.000 71.530 0.900 ;
        RECT 77.930 0.000 80.330 0.900 ;
        RECT 89.130 0.000 91.530 0.900 ;
        RECT 97.930 0.000 100.330 0.900 ;
        RECT 109.130 0.000 111.530 0.900 ;
        RECT 117.930 0.000 120.330 0.900 ;
      LAYER li1 ;
        RECT 9.180 339.600 11.480 340.000 ;
        RECT 17.980 339.600 20.280 340.000 ;
        RECT 29.180 339.600 31.480 340.000 ;
        RECT 37.980 339.600 40.280 340.000 ;
        RECT 49.180 339.600 51.480 340.000 ;
        RECT 57.980 339.600 60.280 340.000 ;
        RECT 69.180 339.600 71.480 340.000 ;
        RECT 77.980 339.600 80.280 340.000 ;
        RECT 89.180 339.600 91.480 340.000 ;
        RECT 97.980 339.600 100.280 340.000 ;
        RECT 109.180 339.600 111.480 340.000 ;
        RECT 117.980 339.600 120.280 340.000 ;
        RECT 5.130 339.200 24.330 339.600 ;
        RECT 2.515 336.880 2.875 337.260 ;
        RECT 3.145 336.880 3.505 337.260 ;
        RECT 3.745 336.880 4.105 337.260 ;
        RECT 2.515 336.290 2.875 336.670 ;
        RECT 3.145 336.290 3.505 336.670 ;
        RECT 3.745 336.290 4.105 336.670 ;
        RECT 5.130 335.550 5.530 339.200 ;
        RECT 9.180 339.150 11.480 339.200 ;
        RECT 17.980 339.150 20.280 339.200 ;
        RECT 6.530 338.000 22.930 338.600 ;
        RECT 10.130 337.400 10.480 338.000 ;
        RECT 6.530 337.200 10.480 337.400 ;
        RECT 10.130 336.600 10.480 337.200 ;
        RECT 6.530 336.400 10.480 336.600 ;
        RECT 10.130 335.800 10.480 336.400 ;
        RECT 6.530 335.600 10.480 335.800 ;
        RECT 4.730 335.545 5.580 335.550 ;
        RECT 2.315 333.250 5.580 335.545 ;
        RECT 10.130 335.000 10.480 335.600 ;
        RECT 6.530 334.800 10.480 335.000 ;
        RECT 10.130 334.200 10.480 334.800 ;
        RECT 6.530 334.000 10.480 334.200 ;
        RECT 10.130 333.400 10.480 334.000 ;
        RECT 5.130 326.750 5.530 333.250 ;
        RECT 6.530 333.200 10.480 333.400 ;
        RECT 10.130 332.600 10.480 333.200 ;
        RECT 6.530 332.400 10.480 332.600 ;
        RECT 10.130 331.800 10.480 332.400 ;
        RECT 6.530 331.600 10.480 331.800 ;
        RECT 10.130 331.000 10.480 331.600 ;
        RECT 6.530 330.800 10.480 331.000 ;
        RECT 10.130 330.400 10.480 330.800 ;
        RECT 11.080 330.400 11.280 338.000 ;
        RECT 11.880 330.400 12.080 338.000 ;
        RECT 12.680 330.400 12.880 338.000 ;
        RECT 13.480 330.400 13.680 338.000 ;
        RECT 10.130 329.200 10.480 329.600 ;
        RECT 6.530 329.000 10.480 329.200 ;
        RECT 10.130 328.400 10.480 329.000 ;
        RECT 6.530 328.200 10.480 328.400 ;
        RECT 10.130 327.600 10.480 328.200 ;
        RECT 6.530 327.400 10.480 327.600 ;
        RECT 10.130 326.800 10.480 327.400 ;
        RECT 4.730 326.745 5.580 326.750 ;
        RECT 2.315 324.450 5.580 326.745 ;
        RECT 6.530 326.600 10.480 326.800 ;
        RECT 10.130 326.000 10.480 326.600 ;
        RECT 6.530 325.800 10.480 326.000 ;
        RECT 10.130 325.200 10.480 325.800 ;
        RECT 6.530 325.000 10.480 325.200 ;
        RECT 2.515 323.515 2.875 323.895 ;
        RECT 3.145 323.515 3.505 323.895 ;
        RECT 3.745 323.515 4.105 323.895 ;
        RECT 2.515 322.925 2.875 323.305 ;
        RECT 3.145 322.925 3.505 323.305 ;
        RECT 3.745 322.925 4.105 323.305 ;
        RECT 5.130 320.800 5.530 324.450 ;
        RECT 10.130 324.400 10.480 325.000 ;
        RECT 6.530 324.200 10.480 324.400 ;
        RECT 10.130 323.600 10.480 324.200 ;
        RECT 6.530 323.400 10.480 323.600 ;
        RECT 10.130 322.800 10.480 323.400 ;
        RECT 6.530 322.600 10.480 322.800 ;
        RECT 10.130 322.000 10.480 322.600 ;
        RECT 11.080 322.000 11.280 329.600 ;
        RECT 11.880 322.000 12.080 329.600 ;
        RECT 12.680 322.000 12.880 329.600 ;
        RECT 13.480 322.000 13.680 329.600 ;
        RECT 14.280 322.000 15.180 338.000 ;
        RECT 15.780 330.400 15.980 338.000 ;
        RECT 16.580 330.400 16.780 338.000 ;
        RECT 17.380 330.400 17.580 338.000 ;
        RECT 18.180 330.400 18.380 338.000 ;
        RECT 18.980 337.400 19.330 338.000 ;
        RECT 18.980 337.200 22.930 337.400 ;
        RECT 18.980 336.600 19.330 337.200 ;
        RECT 18.980 336.400 22.930 336.600 ;
        RECT 18.980 335.800 19.330 336.400 ;
        RECT 18.980 335.600 22.930 335.800 ;
        RECT 18.980 335.000 19.330 335.600 ;
        RECT 23.930 335.550 24.330 339.200 ;
        RECT 25.130 339.200 44.330 339.600 ;
        RECT 25.130 335.550 25.530 339.200 ;
        RECT 29.180 339.150 31.480 339.200 ;
        RECT 37.980 339.150 40.280 339.200 ;
        RECT 26.530 338.000 42.930 338.600 ;
        RECT 30.130 337.400 30.480 338.000 ;
        RECT 26.530 337.200 30.480 337.400 ;
        RECT 30.130 336.600 30.480 337.200 ;
        RECT 26.530 336.400 30.480 336.600 ;
        RECT 30.130 335.800 30.480 336.400 ;
        RECT 26.530 335.600 30.480 335.800 ;
        RECT 18.980 334.800 22.930 335.000 ;
        RECT 18.980 334.200 19.330 334.800 ;
        RECT 18.980 334.000 22.930 334.200 ;
        RECT 18.980 333.400 19.330 334.000 ;
        RECT 18.980 333.200 22.930 333.400 ;
        RECT 23.880 333.250 25.580 335.550 ;
        RECT 30.130 335.000 30.480 335.600 ;
        RECT 26.530 334.800 30.480 335.000 ;
        RECT 30.130 334.200 30.480 334.800 ;
        RECT 26.530 334.000 30.480 334.200 ;
        RECT 30.130 333.400 30.480 334.000 ;
        RECT 18.980 332.600 19.330 333.200 ;
        RECT 18.980 332.400 22.930 332.600 ;
        RECT 18.980 331.800 19.330 332.400 ;
        RECT 18.980 331.600 22.930 331.800 ;
        RECT 18.980 331.000 19.330 331.600 ;
        RECT 18.980 330.800 22.930 331.000 ;
        RECT 18.980 330.400 19.330 330.800 ;
        RECT 15.780 322.000 15.980 329.600 ;
        RECT 16.580 322.000 16.780 329.600 ;
        RECT 17.380 322.000 17.580 329.600 ;
        RECT 18.180 322.000 18.380 329.600 ;
        RECT 18.980 329.200 19.330 329.600 ;
        RECT 18.980 329.000 22.930 329.200 ;
        RECT 18.980 328.400 19.330 329.000 ;
        RECT 18.980 328.200 22.930 328.400 ;
        RECT 18.980 327.600 19.330 328.200 ;
        RECT 18.980 327.400 22.930 327.600 ;
        RECT 18.980 326.800 19.330 327.400 ;
        RECT 18.980 326.600 22.930 326.800 ;
        RECT 23.930 326.750 24.330 333.250 ;
        RECT 25.130 326.750 25.530 333.250 ;
        RECT 26.530 333.200 30.480 333.400 ;
        RECT 30.130 332.600 30.480 333.200 ;
        RECT 26.530 332.400 30.480 332.600 ;
        RECT 30.130 331.800 30.480 332.400 ;
        RECT 26.530 331.600 30.480 331.800 ;
        RECT 30.130 331.000 30.480 331.600 ;
        RECT 26.530 330.800 30.480 331.000 ;
        RECT 30.130 330.400 30.480 330.800 ;
        RECT 31.080 330.400 31.280 338.000 ;
        RECT 31.880 330.400 32.080 338.000 ;
        RECT 32.680 330.400 32.880 338.000 ;
        RECT 33.480 330.400 33.680 338.000 ;
        RECT 30.130 329.200 30.480 329.600 ;
        RECT 26.530 329.000 30.480 329.200 ;
        RECT 30.130 328.400 30.480 329.000 ;
        RECT 26.530 328.200 30.480 328.400 ;
        RECT 30.130 327.600 30.480 328.200 ;
        RECT 26.530 327.400 30.480 327.600 ;
        RECT 30.130 326.800 30.480 327.400 ;
        RECT 18.980 326.000 19.330 326.600 ;
        RECT 18.980 325.800 22.930 326.000 ;
        RECT 18.980 325.200 19.330 325.800 ;
        RECT 18.980 325.000 22.930 325.200 ;
        RECT 18.980 324.400 19.330 325.000 ;
        RECT 23.880 324.450 25.580 326.750 ;
        RECT 26.530 326.600 30.480 326.800 ;
        RECT 30.130 326.000 30.480 326.600 ;
        RECT 26.530 325.800 30.480 326.000 ;
        RECT 30.130 325.200 30.480 325.800 ;
        RECT 26.530 325.000 30.480 325.200 ;
        RECT 18.980 324.200 22.930 324.400 ;
        RECT 18.980 323.600 19.330 324.200 ;
        RECT 18.980 323.400 22.930 323.600 ;
        RECT 18.980 322.800 19.330 323.400 ;
        RECT 18.980 322.600 22.930 322.800 ;
        RECT 18.980 322.000 19.330 322.600 ;
        RECT 6.530 321.400 22.930 322.000 ;
        RECT 9.180 320.800 11.480 320.850 ;
        RECT 17.980 320.800 20.280 320.850 ;
        RECT 23.930 320.800 24.330 324.450 ;
        RECT 5.130 320.400 24.330 320.800 ;
        RECT 25.130 320.800 25.530 324.450 ;
        RECT 30.130 324.400 30.480 325.000 ;
        RECT 26.530 324.200 30.480 324.400 ;
        RECT 30.130 323.600 30.480 324.200 ;
        RECT 26.530 323.400 30.480 323.600 ;
        RECT 30.130 322.800 30.480 323.400 ;
        RECT 26.530 322.600 30.480 322.800 ;
        RECT 30.130 322.000 30.480 322.600 ;
        RECT 31.080 322.000 31.280 329.600 ;
        RECT 31.880 322.000 32.080 329.600 ;
        RECT 32.680 322.000 32.880 329.600 ;
        RECT 33.480 322.000 33.680 329.600 ;
        RECT 34.280 322.000 35.180 338.000 ;
        RECT 35.780 330.400 35.980 338.000 ;
        RECT 36.580 330.400 36.780 338.000 ;
        RECT 37.380 330.400 37.580 338.000 ;
        RECT 38.180 330.400 38.380 338.000 ;
        RECT 38.980 337.400 39.330 338.000 ;
        RECT 38.980 337.200 42.930 337.400 ;
        RECT 38.980 336.600 39.330 337.200 ;
        RECT 38.980 336.400 42.930 336.600 ;
        RECT 38.980 335.800 39.330 336.400 ;
        RECT 38.980 335.600 42.930 335.800 ;
        RECT 38.980 335.000 39.330 335.600 ;
        RECT 43.930 335.550 44.330 339.200 ;
        RECT 45.130 339.200 64.330 339.600 ;
        RECT 45.130 335.550 45.530 339.200 ;
        RECT 49.180 339.150 51.480 339.200 ;
        RECT 57.980 339.150 60.280 339.200 ;
        RECT 46.530 338.000 62.930 338.600 ;
        RECT 50.130 337.400 50.480 338.000 ;
        RECT 46.530 337.200 50.480 337.400 ;
        RECT 50.130 336.600 50.480 337.200 ;
        RECT 46.530 336.400 50.480 336.600 ;
        RECT 50.130 335.800 50.480 336.400 ;
        RECT 46.530 335.600 50.480 335.800 ;
        RECT 38.980 334.800 42.930 335.000 ;
        RECT 38.980 334.200 39.330 334.800 ;
        RECT 38.980 334.000 42.930 334.200 ;
        RECT 38.980 333.400 39.330 334.000 ;
        RECT 38.980 333.200 42.930 333.400 ;
        RECT 43.880 333.250 45.580 335.550 ;
        RECT 50.130 335.000 50.480 335.600 ;
        RECT 46.530 334.800 50.480 335.000 ;
        RECT 50.130 334.200 50.480 334.800 ;
        RECT 46.530 334.000 50.480 334.200 ;
        RECT 50.130 333.400 50.480 334.000 ;
        RECT 38.980 332.600 39.330 333.200 ;
        RECT 38.980 332.400 42.930 332.600 ;
        RECT 38.980 331.800 39.330 332.400 ;
        RECT 38.980 331.600 42.930 331.800 ;
        RECT 38.980 331.000 39.330 331.600 ;
        RECT 38.980 330.800 42.930 331.000 ;
        RECT 38.980 330.400 39.330 330.800 ;
        RECT 35.780 322.000 35.980 329.600 ;
        RECT 36.580 322.000 36.780 329.600 ;
        RECT 37.380 322.000 37.580 329.600 ;
        RECT 38.180 322.000 38.380 329.600 ;
        RECT 38.980 329.200 39.330 329.600 ;
        RECT 38.980 329.000 42.930 329.200 ;
        RECT 38.980 328.400 39.330 329.000 ;
        RECT 38.980 328.200 42.930 328.400 ;
        RECT 38.980 327.600 39.330 328.200 ;
        RECT 38.980 327.400 42.930 327.600 ;
        RECT 38.980 326.800 39.330 327.400 ;
        RECT 38.980 326.600 42.930 326.800 ;
        RECT 43.930 326.750 44.330 333.250 ;
        RECT 45.130 326.750 45.530 333.250 ;
        RECT 46.530 333.200 50.480 333.400 ;
        RECT 50.130 332.600 50.480 333.200 ;
        RECT 46.530 332.400 50.480 332.600 ;
        RECT 50.130 331.800 50.480 332.400 ;
        RECT 46.530 331.600 50.480 331.800 ;
        RECT 50.130 331.000 50.480 331.600 ;
        RECT 46.530 330.800 50.480 331.000 ;
        RECT 50.130 330.400 50.480 330.800 ;
        RECT 51.080 330.400 51.280 338.000 ;
        RECT 51.880 330.400 52.080 338.000 ;
        RECT 52.680 330.400 52.880 338.000 ;
        RECT 53.480 330.400 53.680 338.000 ;
        RECT 50.130 329.200 50.480 329.600 ;
        RECT 46.530 329.000 50.480 329.200 ;
        RECT 50.130 328.400 50.480 329.000 ;
        RECT 46.530 328.200 50.480 328.400 ;
        RECT 50.130 327.600 50.480 328.200 ;
        RECT 46.530 327.400 50.480 327.600 ;
        RECT 50.130 326.800 50.480 327.400 ;
        RECT 38.980 326.000 39.330 326.600 ;
        RECT 38.980 325.800 42.930 326.000 ;
        RECT 38.980 325.200 39.330 325.800 ;
        RECT 38.980 325.000 42.930 325.200 ;
        RECT 38.980 324.400 39.330 325.000 ;
        RECT 43.880 324.450 45.580 326.750 ;
        RECT 46.530 326.600 50.480 326.800 ;
        RECT 50.130 326.000 50.480 326.600 ;
        RECT 46.530 325.800 50.480 326.000 ;
        RECT 50.130 325.200 50.480 325.800 ;
        RECT 46.530 325.000 50.480 325.200 ;
        RECT 38.980 324.200 42.930 324.400 ;
        RECT 38.980 323.600 39.330 324.200 ;
        RECT 38.980 323.400 42.930 323.600 ;
        RECT 38.980 322.800 39.330 323.400 ;
        RECT 38.980 322.600 42.930 322.800 ;
        RECT 38.980 322.000 39.330 322.600 ;
        RECT 26.530 321.400 42.930 322.000 ;
        RECT 29.180 320.800 31.480 320.850 ;
        RECT 37.980 320.800 40.280 320.850 ;
        RECT 43.930 320.800 44.330 324.450 ;
        RECT 25.130 320.400 44.330 320.800 ;
        RECT 45.130 320.800 45.530 324.450 ;
        RECT 50.130 324.400 50.480 325.000 ;
        RECT 46.530 324.200 50.480 324.400 ;
        RECT 50.130 323.600 50.480 324.200 ;
        RECT 46.530 323.400 50.480 323.600 ;
        RECT 50.130 322.800 50.480 323.400 ;
        RECT 46.530 322.600 50.480 322.800 ;
        RECT 50.130 322.000 50.480 322.600 ;
        RECT 51.080 322.000 51.280 329.600 ;
        RECT 51.880 322.000 52.080 329.600 ;
        RECT 52.680 322.000 52.880 329.600 ;
        RECT 53.480 322.000 53.680 329.600 ;
        RECT 54.280 322.000 55.180 338.000 ;
        RECT 55.780 330.400 55.980 338.000 ;
        RECT 56.580 330.400 56.780 338.000 ;
        RECT 57.380 330.400 57.580 338.000 ;
        RECT 58.180 330.400 58.380 338.000 ;
        RECT 58.980 337.400 59.330 338.000 ;
        RECT 58.980 337.200 62.930 337.400 ;
        RECT 58.980 336.600 59.330 337.200 ;
        RECT 58.980 336.400 62.930 336.600 ;
        RECT 58.980 335.800 59.330 336.400 ;
        RECT 58.980 335.600 62.930 335.800 ;
        RECT 58.980 335.000 59.330 335.600 ;
        RECT 63.930 335.550 64.330 339.200 ;
        RECT 65.130 339.200 84.330 339.600 ;
        RECT 65.130 335.550 65.530 339.200 ;
        RECT 69.180 339.150 71.480 339.200 ;
        RECT 77.980 339.150 80.280 339.200 ;
        RECT 66.530 338.000 82.930 338.600 ;
        RECT 70.130 337.400 70.480 338.000 ;
        RECT 66.530 337.200 70.480 337.400 ;
        RECT 70.130 336.600 70.480 337.200 ;
        RECT 66.530 336.400 70.480 336.600 ;
        RECT 70.130 335.800 70.480 336.400 ;
        RECT 66.530 335.600 70.480 335.800 ;
        RECT 58.980 334.800 62.930 335.000 ;
        RECT 58.980 334.200 59.330 334.800 ;
        RECT 58.980 334.000 62.930 334.200 ;
        RECT 58.980 333.400 59.330 334.000 ;
        RECT 58.980 333.200 62.930 333.400 ;
        RECT 63.880 333.250 65.580 335.550 ;
        RECT 70.130 335.000 70.480 335.600 ;
        RECT 66.530 334.800 70.480 335.000 ;
        RECT 70.130 334.200 70.480 334.800 ;
        RECT 66.530 334.000 70.480 334.200 ;
        RECT 70.130 333.400 70.480 334.000 ;
        RECT 58.980 332.600 59.330 333.200 ;
        RECT 58.980 332.400 62.930 332.600 ;
        RECT 58.980 331.800 59.330 332.400 ;
        RECT 58.980 331.600 62.930 331.800 ;
        RECT 58.980 331.000 59.330 331.600 ;
        RECT 58.980 330.800 62.930 331.000 ;
        RECT 58.980 330.400 59.330 330.800 ;
        RECT 55.780 322.000 55.980 329.600 ;
        RECT 56.580 322.000 56.780 329.600 ;
        RECT 57.380 322.000 57.580 329.600 ;
        RECT 58.180 322.000 58.380 329.600 ;
        RECT 58.980 329.200 59.330 329.600 ;
        RECT 58.980 329.000 62.930 329.200 ;
        RECT 58.980 328.400 59.330 329.000 ;
        RECT 58.980 328.200 62.930 328.400 ;
        RECT 58.980 327.600 59.330 328.200 ;
        RECT 58.980 327.400 62.930 327.600 ;
        RECT 58.980 326.800 59.330 327.400 ;
        RECT 58.980 326.600 62.930 326.800 ;
        RECT 63.930 326.750 64.330 333.250 ;
        RECT 65.130 326.750 65.530 333.250 ;
        RECT 66.530 333.200 70.480 333.400 ;
        RECT 70.130 332.600 70.480 333.200 ;
        RECT 66.530 332.400 70.480 332.600 ;
        RECT 70.130 331.800 70.480 332.400 ;
        RECT 66.530 331.600 70.480 331.800 ;
        RECT 70.130 331.000 70.480 331.600 ;
        RECT 66.530 330.800 70.480 331.000 ;
        RECT 70.130 330.400 70.480 330.800 ;
        RECT 71.080 330.400 71.280 338.000 ;
        RECT 71.880 330.400 72.080 338.000 ;
        RECT 72.680 330.400 72.880 338.000 ;
        RECT 73.480 330.400 73.680 338.000 ;
        RECT 70.130 329.200 70.480 329.600 ;
        RECT 66.530 329.000 70.480 329.200 ;
        RECT 70.130 328.400 70.480 329.000 ;
        RECT 66.530 328.200 70.480 328.400 ;
        RECT 70.130 327.600 70.480 328.200 ;
        RECT 66.530 327.400 70.480 327.600 ;
        RECT 70.130 326.800 70.480 327.400 ;
        RECT 58.980 326.000 59.330 326.600 ;
        RECT 58.980 325.800 62.930 326.000 ;
        RECT 58.980 325.200 59.330 325.800 ;
        RECT 58.980 325.000 62.930 325.200 ;
        RECT 58.980 324.400 59.330 325.000 ;
        RECT 63.880 324.450 65.580 326.750 ;
        RECT 66.530 326.600 70.480 326.800 ;
        RECT 70.130 326.000 70.480 326.600 ;
        RECT 66.530 325.800 70.480 326.000 ;
        RECT 70.130 325.200 70.480 325.800 ;
        RECT 66.530 325.000 70.480 325.200 ;
        RECT 58.980 324.200 62.930 324.400 ;
        RECT 58.980 323.600 59.330 324.200 ;
        RECT 58.980 323.400 62.930 323.600 ;
        RECT 58.980 322.800 59.330 323.400 ;
        RECT 58.980 322.600 62.930 322.800 ;
        RECT 58.980 322.000 59.330 322.600 ;
        RECT 46.530 321.400 62.930 322.000 ;
        RECT 49.180 320.800 51.480 320.850 ;
        RECT 57.980 320.800 60.280 320.850 ;
        RECT 63.930 320.800 64.330 324.450 ;
        RECT 45.130 320.400 64.330 320.800 ;
        RECT 65.130 320.800 65.530 324.450 ;
        RECT 70.130 324.400 70.480 325.000 ;
        RECT 66.530 324.200 70.480 324.400 ;
        RECT 70.130 323.600 70.480 324.200 ;
        RECT 66.530 323.400 70.480 323.600 ;
        RECT 70.130 322.800 70.480 323.400 ;
        RECT 66.530 322.600 70.480 322.800 ;
        RECT 70.130 322.000 70.480 322.600 ;
        RECT 71.080 322.000 71.280 329.600 ;
        RECT 71.880 322.000 72.080 329.600 ;
        RECT 72.680 322.000 72.880 329.600 ;
        RECT 73.480 322.000 73.680 329.600 ;
        RECT 74.280 322.000 75.180 338.000 ;
        RECT 75.780 330.400 75.980 338.000 ;
        RECT 76.580 330.400 76.780 338.000 ;
        RECT 77.380 330.400 77.580 338.000 ;
        RECT 78.180 330.400 78.380 338.000 ;
        RECT 78.980 337.400 79.330 338.000 ;
        RECT 78.980 337.200 82.930 337.400 ;
        RECT 78.980 336.600 79.330 337.200 ;
        RECT 78.980 336.400 82.930 336.600 ;
        RECT 78.980 335.800 79.330 336.400 ;
        RECT 78.980 335.600 82.930 335.800 ;
        RECT 78.980 335.000 79.330 335.600 ;
        RECT 83.930 335.550 84.330 339.200 ;
        RECT 85.130 339.200 104.330 339.600 ;
        RECT 85.130 335.550 85.530 339.200 ;
        RECT 89.180 339.150 91.480 339.200 ;
        RECT 97.980 339.150 100.280 339.200 ;
        RECT 86.530 338.000 102.930 338.600 ;
        RECT 90.130 337.400 90.480 338.000 ;
        RECT 86.530 337.200 90.480 337.400 ;
        RECT 90.130 336.600 90.480 337.200 ;
        RECT 86.530 336.400 90.480 336.600 ;
        RECT 90.130 335.800 90.480 336.400 ;
        RECT 86.530 335.600 90.480 335.800 ;
        RECT 78.980 334.800 82.930 335.000 ;
        RECT 78.980 334.200 79.330 334.800 ;
        RECT 78.980 334.000 82.930 334.200 ;
        RECT 78.980 333.400 79.330 334.000 ;
        RECT 78.980 333.200 82.930 333.400 ;
        RECT 83.880 333.250 85.580 335.550 ;
        RECT 90.130 335.000 90.480 335.600 ;
        RECT 86.530 334.800 90.480 335.000 ;
        RECT 90.130 334.200 90.480 334.800 ;
        RECT 86.530 334.000 90.480 334.200 ;
        RECT 90.130 333.400 90.480 334.000 ;
        RECT 78.980 332.600 79.330 333.200 ;
        RECT 78.980 332.400 82.930 332.600 ;
        RECT 78.980 331.800 79.330 332.400 ;
        RECT 78.980 331.600 82.930 331.800 ;
        RECT 78.980 331.000 79.330 331.600 ;
        RECT 78.980 330.800 82.930 331.000 ;
        RECT 78.980 330.400 79.330 330.800 ;
        RECT 75.780 322.000 75.980 329.600 ;
        RECT 76.580 322.000 76.780 329.600 ;
        RECT 77.380 322.000 77.580 329.600 ;
        RECT 78.180 322.000 78.380 329.600 ;
        RECT 78.980 329.200 79.330 329.600 ;
        RECT 78.980 329.000 82.930 329.200 ;
        RECT 78.980 328.400 79.330 329.000 ;
        RECT 78.980 328.200 82.930 328.400 ;
        RECT 78.980 327.600 79.330 328.200 ;
        RECT 78.980 327.400 82.930 327.600 ;
        RECT 78.980 326.800 79.330 327.400 ;
        RECT 78.980 326.600 82.930 326.800 ;
        RECT 83.930 326.750 84.330 333.250 ;
        RECT 85.130 326.750 85.530 333.250 ;
        RECT 86.530 333.200 90.480 333.400 ;
        RECT 90.130 332.600 90.480 333.200 ;
        RECT 86.530 332.400 90.480 332.600 ;
        RECT 90.130 331.800 90.480 332.400 ;
        RECT 86.530 331.600 90.480 331.800 ;
        RECT 90.130 331.000 90.480 331.600 ;
        RECT 86.530 330.800 90.480 331.000 ;
        RECT 90.130 330.400 90.480 330.800 ;
        RECT 91.080 330.400 91.280 338.000 ;
        RECT 91.880 330.400 92.080 338.000 ;
        RECT 92.680 330.400 92.880 338.000 ;
        RECT 93.480 330.400 93.680 338.000 ;
        RECT 90.130 329.200 90.480 329.600 ;
        RECT 86.530 329.000 90.480 329.200 ;
        RECT 90.130 328.400 90.480 329.000 ;
        RECT 86.530 328.200 90.480 328.400 ;
        RECT 90.130 327.600 90.480 328.200 ;
        RECT 86.530 327.400 90.480 327.600 ;
        RECT 90.130 326.800 90.480 327.400 ;
        RECT 78.980 326.000 79.330 326.600 ;
        RECT 78.980 325.800 82.930 326.000 ;
        RECT 78.980 325.200 79.330 325.800 ;
        RECT 78.980 325.000 82.930 325.200 ;
        RECT 78.980 324.400 79.330 325.000 ;
        RECT 83.880 324.450 85.580 326.750 ;
        RECT 86.530 326.600 90.480 326.800 ;
        RECT 90.130 326.000 90.480 326.600 ;
        RECT 86.530 325.800 90.480 326.000 ;
        RECT 90.130 325.200 90.480 325.800 ;
        RECT 86.530 325.000 90.480 325.200 ;
        RECT 78.980 324.200 82.930 324.400 ;
        RECT 78.980 323.600 79.330 324.200 ;
        RECT 78.980 323.400 82.930 323.600 ;
        RECT 78.980 322.800 79.330 323.400 ;
        RECT 78.980 322.600 82.930 322.800 ;
        RECT 78.980 322.000 79.330 322.600 ;
        RECT 66.530 321.400 82.930 322.000 ;
        RECT 69.180 320.800 71.480 320.850 ;
        RECT 77.980 320.800 80.280 320.850 ;
        RECT 83.930 320.800 84.330 324.450 ;
        RECT 65.130 320.400 84.330 320.800 ;
        RECT 85.130 320.800 85.530 324.450 ;
        RECT 90.130 324.400 90.480 325.000 ;
        RECT 86.530 324.200 90.480 324.400 ;
        RECT 90.130 323.600 90.480 324.200 ;
        RECT 86.530 323.400 90.480 323.600 ;
        RECT 90.130 322.800 90.480 323.400 ;
        RECT 86.530 322.600 90.480 322.800 ;
        RECT 90.130 322.000 90.480 322.600 ;
        RECT 91.080 322.000 91.280 329.600 ;
        RECT 91.880 322.000 92.080 329.600 ;
        RECT 92.680 322.000 92.880 329.600 ;
        RECT 93.480 322.000 93.680 329.600 ;
        RECT 94.280 322.000 95.180 338.000 ;
        RECT 95.780 330.400 95.980 338.000 ;
        RECT 96.580 330.400 96.780 338.000 ;
        RECT 97.380 330.400 97.580 338.000 ;
        RECT 98.180 330.400 98.380 338.000 ;
        RECT 98.980 337.400 99.330 338.000 ;
        RECT 98.980 337.200 102.930 337.400 ;
        RECT 98.980 336.600 99.330 337.200 ;
        RECT 98.980 336.400 102.930 336.600 ;
        RECT 98.980 335.800 99.330 336.400 ;
        RECT 98.980 335.600 102.930 335.800 ;
        RECT 98.980 335.000 99.330 335.600 ;
        RECT 103.930 335.550 104.330 339.200 ;
        RECT 105.130 339.200 124.330 339.600 ;
        RECT 105.130 335.550 105.530 339.200 ;
        RECT 109.180 339.150 111.480 339.200 ;
        RECT 117.980 339.150 120.280 339.200 ;
        RECT 106.530 338.000 122.930 338.600 ;
        RECT 110.130 337.400 110.480 338.000 ;
        RECT 106.530 337.200 110.480 337.400 ;
        RECT 110.130 336.600 110.480 337.200 ;
        RECT 106.530 336.400 110.480 336.600 ;
        RECT 110.130 335.800 110.480 336.400 ;
        RECT 106.530 335.600 110.480 335.800 ;
        RECT 98.980 334.800 102.930 335.000 ;
        RECT 98.980 334.200 99.330 334.800 ;
        RECT 98.980 334.000 102.930 334.200 ;
        RECT 98.980 333.400 99.330 334.000 ;
        RECT 98.980 333.200 102.930 333.400 ;
        RECT 103.880 333.250 105.580 335.550 ;
        RECT 110.130 335.000 110.480 335.600 ;
        RECT 106.530 334.800 110.480 335.000 ;
        RECT 110.130 334.200 110.480 334.800 ;
        RECT 106.530 334.000 110.480 334.200 ;
        RECT 110.130 333.400 110.480 334.000 ;
        RECT 98.980 332.600 99.330 333.200 ;
        RECT 98.980 332.400 102.930 332.600 ;
        RECT 98.980 331.800 99.330 332.400 ;
        RECT 98.980 331.600 102.930 331.800 ;
        RECT 98.980 331.000 99.330 331.600 ;
        RECT 98.980 330.800 102.930 331.000 ;
        RECT 98.980 330.400 99.330 330.800 ;
        RECT 95.780 322.000 95.980 329.600 ;
        RECT 96.580 322.000 96.780 329.600 ;
        RECT 97.380 322.000 97.580 329.600 ;
        RECT 98.180 322.000 98.380 329.600 ;
        RECT 98.980 329.200 99.330 329.600 ;
        RECT 98.980 329.000 102.930 329.200 ;
        RECT 98.980 328.400 99.330 329.000 ;
        RECT 98.980 328.200 102.930 328.400 ;
        RECT 98.980 327.600 99.330 328.200 ;
        RECT 98.980 327.400 102.930 327.600 ;
        RECT 98.980 326.800 99.330 327.400 ;
        RECT 98.980 326.600 102.930 326.800 ;
        RECT 103.930 326.750 104.330 333.250 ;
        RECT 105.130 326.750 105.530 333.250 ;
        RECT 106.530 333.200 110.480 333.400 ;
        RECT 110.130 332.600 110.480 333.200 ;
        RECT 106.530 332.400 110.480 332.600 ;
        RECT 110.130 331.800 110.480 332.400 ;
        RECT 106.530 331.600 110.480 331.800 ;
        RECT 110.130 331.000 110.480 331.600 ;
        RECT 106.530 330.800 110.480 331.000 ;
        RECT 110.130 330.400 110.480 330.800 ;
        RECT 111.080 330.400 111.280 338.000 ;
        RECT 111.880 330.400 112.080 338.000 ;
        RECT 112.680 330.400 112.880 338.000 ;
        RECT 113.480 330.400 113.680 338.000 ;
        RECT 110.130 329.200 110.480 329.600 ;
        RECT 106.530 329.000 110.480 329.200 ;
        RECT 110.130 328.400 110.480 329.000 ;
        RECT 106.530 328.200 110.480 328.400 ;
        RECT 110.130 327.600 110.480 328.200 ;
        RECT 106.530 327.400 110.480 327.600 ;
        RECT 110.130 326.800 110.480 327.400 ;
        RECT 98.980 326.000 99.330 326.600 ;
        RECT 98.980 325.800 102.930 326.000 ;
        RECT 98.980 325.200 99.330 325.800 ;
        RECT 98.980 325.000 102.930 325.200 ;
        RECT 98.980 324.400 99.330 325.000 ;
        RECT 103.880 324.450 105.580 326.750 ;
        RECT 106.530 326.600 110.480 326.800 ;
        RECT 110.130 326.000 110.480 326.600 ;
        RECT 106.530 325.800 110.480 326.000 ;
        RECT 110.130 325.200 110.480 325.800 ;
        RECT 106.530 325.000 110.480 325.200 ;
        RECT 98.980 324.200 102.930 324.400 ;
        RECT 98.980 323.600 99.330 324.200 ;
        RECT 98.980 323.400 102.930 323.600 ;
        RECT 98.980 322.800 99.330 323.400 ;
        RECT 98.980 322.600 102.930 322.800 ;
        RECT 98.980 322.000 99.330 322.600 ;
        RECT 86.530 321.400 102.930 322.000 ;
        RECT 89.180 320.800 91.480 320.850 ;
        RECT 97.980 320.800 100.280 320.850 ;
        RECT 103.930 320.800 104.330 324.450 ;
        RECT 85.130 320.400 104.330 320.800 ;
        RECT 105.130 320.800 105.530 324.450 ;
        RECT 110.130 324.400 110.480 325.000 ;
        RECT 106.530 324.200 110.480 324.400 ;
        RECT 110.130 323.600 110.480 324.200 ;
        RECT 106.530 323.400 110.480 323.600 ;
        RECT 110.130 322.800 110.480 323.400 ;
        RECT 106.530 322.600 110.480 322.800 ;
        RECT 110.130 322.000 110.480 322.600 ;
        RECT 111.080 322.000 111.280 329.600 ;
        RECT 111.880 322.000 112.080 329.600 ;
        RECT 112.680 322.000 112.880 329.600 ;
        RECT 113.480 322.000 113.680 329.600 ;
        RECT 114.280 322.000 115.180 338.000 ;
        RECT 115.780 330.400 115.980 338.000 ;
        RECT 116.580 330.400 116.780 338.000 ;
        RECT 117.380 330.400 117.580 338.000 ;
        RECT 118.180 330.400 118.380 338.000 ;
        RECT 118.980 337.400 119.330 338.000 ;
        RECT 118.980 337.200 122.930 337.400 ;
        RECT 118.980 336.600 119.330 337.200 ;
        RECT 118.980 336.400 122.930 336.600 ;
        RECT 118.980 335.800 119.330 336.400 ;
        RECT 118.980 335.600 122.930 335.800 ;
        RECT 118.980 335.000 119.330 335.600 ;
        RECT 123.930 335.550 124.330 339.200 ;
        RECT 125.340 337.080 125.700 337.460 ;
        RECT 125.970 337.080 126.330 337.460 ;
        RECT 126.570 337.080 126.930 337.460 ;
        RECT 125.340 336.490 125.700 336.870 ;
        RECT 125.970 336.490 126.330 336.870 ;
        RECT 126.570 336.490 126.930 336.870 ;
        RECT 118.980 334.800 122.930 335.000 ;
        RECT 118.980 334.200 119.330 334.800 ;
        RECT 118.980 334.000 122.930 334.200 ;
        RECT 118.980 333.400 119.330 334.000 ;
        RECT 118.980 333.200 122.930 333.400 ;
        RECT 123.880 333.250 124.730 335.550 ;
        RECT 118.980 332.600 119.330 333.200 ;
        RECT 118.980 332.400 122.930 332.600 ;
        RECT 118.980 331.800 119.330 332.400 ;
        RECT 118.980 331.600 122.930 331.800 ;
        RECT 118.980 331.000 119.330 331.600 ;
        RECT 118.980 330.800 122.930 331.000 ;
        RECT 118.980 330.400 119.330 330.800 ;
        RECT 115.780 322.000 115.980 329.600 ;
        RECT 116.580 322.000 116.780 329.600 ;
        RECT 117.380 322.000 117.580 329.600 ;
        RECT 118.180 322.000 118.380 329.600 ;
        RECT 118.980 329.200 119.330 329.600 ;
        RECT 118.980 329.000 122.930 329.200 ;
        RECT 118.980 328.400 119.330 329.000 ;
        RECT 118.980 328.200 122.930 328.400 ;
        RECT 118.980 327.600 119.330 328.200 ;
        RECT 118.980 327.400 122.930 327.600 ;
        RECT 118.980 326.800 119.330 327.400 ;
        RECT 118.980 326.600 122.930 326.800 ;
        RECT 123.930 326.750 124.330 333.250 ;
        RECT 118.980 326.000 119.330 326.600 ;
        RECT 118.980 325.800 122.930 326.000 ;
        RECT 118.980 325.200 119.330 325.800 ;
        RECT 118.980 325.000 122.930 325.200 ;
        RECT 118.980 324.400 119.330 325.000 ;
        RECT 123.880 324.450 124.730 326.750 ;
        RECT 118.980 324.200 122.930 324.400 ;
        RECT 118.980 323.600 119.330 324.200 ;
        RECT 118.980 323.400 122.930 323.600 ;
        RECT 118.980 322.800 119.330 323.400 ;
        RECT 118.980 322.600 122.930 322.800 ;
        RECT 118.980 322.000 119.330 322.600 ;
        RECT 106.530 321.400 122.930 322.000 ;
        RECT 109.180 320.800 111.480 320.850 ;
        RECT 117.980 320.800 120.280 320.850 ;
        RECT 123.930 320.800 124.330 324.450 ;
        RECT 125.340 323.095 125.700 323.475 ;
        RECT 125.970 323.095 126.330 323.475 ;
        RECT 126.570 323.095 126.930 323.475 ;
        RECT 125.340 322.505 125.700 322.885 ;
        RECT 125.970 322.505 126.330 322.885 ;
        RECT 126.570 322.505 126.930 322.885 ;
        RECT 105.130 320.400 124.330 320.800 ;
        RECT 9.180 319.600 11.480 320.400 ;
        RECT 17.980 319.600 20.280 320.400 ;
        RECT 29.180 319.600 31.480 320.400 ;
        RECT 37.980 319.600 40.280 320.400 ;
        RECT 49.180 319.600 51.480 320.400 ;
        RECT 57.980 319.600 60.280 320.400 ;
        RECT 69.180 319.600 71.480 320.400 ;
        RECT 77.980 319.600 80.280 320.400 ;
        RECT 89.180 319.600 91.480 320.400 ;
        RECT 97.980 319.600 100.280 320.400 ;
        RECT 109.180 319.600 111.480 320.400 ;
        RECT 117.980 319.600 120.280 320.400 ;
        RECT 5.130 319.200 24.330 319.600 ;
        RECT 2.515 316.870 2.875 317.250 ;
        RECT 3.145 316.870 3.505 317.250 ;
        RECT 3.745 316.870 4.105 317.250 ;
        RECT 2.515 316.280 2.875 316.660 ;
        RECT 3.145 316.280 3.505 316.660 ;
        RECT 3.745 316.280 4.105 316.660 ;
        RECT 5.130 315.550 5.530 319.200 ;
        RECT 9.180 319.150 11.480 319.200 ;
        RECT 17.980 319.150 20.280 319.200 ;
        RECT 6.530 318.000 22.930 318.600 ;
        RECT 10.130 317.400 10.480 318.000 ;
        RECT 6.530 317.200 10.480 317.400 ;
        RECT 10.130 316.600 10.480 317.200 ;
        RECT 6.530 316.400 10.480 316.600 ;
        RECT 10.130 315.800 10.480 316.400 ;
        RECT 6.530 315.600 10.480 315.800 ;
        RECT 4.730 315.545 5.580 315.550 ;
        RECT 2.315 313.250 5.580 315.545 ;
        RECT 10.130 315.000 10.480 315.600 ;
        RECT 6.530 314.800 10.480 315.000 ;
        RECT 10.130 314.200 10.480 314.800 ;
        RECT 6.530 314.000 10.480 314.200 ;
        RECT 10.130 313.400 10.480 314.000 ;
        RECT 5.130 306.750 5.530 313.250 ;
        RECT 6.530 313.200 10.480 313.400 ;
        RECT 10.130 312.600 10.480 313.200 ;
        RECT 6.530 312.400 10.480 312.600 ;
        RECT 10.130 311.800 10.480 312.400 ;
        RECT 6.530 311.600 10.480 311.800 ;
        RECT 10.130 311.000 10.480 311.600 ;
        RECT 6.530 310.800 10.480 311.000 ;
        RECT 10.130 310.400 10.480 310.800 ;
        RECT 11.080 310.400 11.280 318.000 ;
        RECT 11.880 310.400 12.080 318.000 ;
        RECT 12.680 310.400 12.880 318.000 ;
        RECT 13.480 310.400 13.680 318.000 ;
        RECT 10.130 309.200 10.480 309.600 ;
        RECT 6.530 309.000 10.480 309.200 ;
        RECT 10.130 308.400 10.480 309.000 ;
        RECT 6.530 308.200 10.480 308.400 ;
        RECT 10.130 307.600 10.480 308.200 ;
        RECT 6.530 307.400 10.480 307.600 ;
        RECT 10.130 306.800 10.480 307.400 ;
        RECT 2.315 304.455 5.580 306.750 ;
        RECT 6.530 306.600 10.480 306.800 ;
        RECT 10.130 306.000 10.480 306.600 ;
        RECT 6.530 305.800 10.480 306.000 ;
        RECT 10.130 305.200 10.480 305.800 ;
        RECT 6.530 305.000 10.480 305.200 ;
        RECT 4.730 304.450 5.580 304.455 ;
        RECT 2.515 303.170 2.875 303.550 ;
        RECT 3.145 303.170 3.505 303.550 ;
        RECT 3.745 303.170 4.105 303.550 ;
        RECT 2.515 302.580 2.875 302.960 ;
        RECT 3.145 302.580 3.505 302.960 ;
        RECT 3.745 302.580 4.105 302.960 ;
        RECT 5.130 300.800 5.530 304.450 ;
        RECT 10.130 304.400 10.480 305.000 ;
        RECT 6.530 304.200 10.480 304.400 ;
        RECT 10.130 303.600 10.480 304.200 ;
        RECT 6.530 303.400 10.480 303.600 ;
        RECT 10.130 302.800 10.480 303.400 ;
        RECT 6.530 302.600 10.480 302.800 ;
        RECT 10.130 302.000 10.480 302.600 ;
        RECT 11.080 302.000 11.280 309.600 ;
        RECT 11.880 302.000 12.080 309.600 ;
        RECT 12.680 302.000 12.880 309.600 ;
        RECT 13.480 302.000 13.680 309.600 ;
        RECT 14.280 302.000 15.180 318.000 ;
        RECT 15.780 310.400 15.980 318.000 ;
        RECT 16.580 310.400 16.780 318.000 ;
        RECT 17.380 310.400 17.580 318.000 ;
        RECT 18.180 310.400 18.380 318.000 ;
        RECT 18.980 317.400 19.330 318.000 ;
        RECT 18.980 317.200 22.930 317.400 ;
        RECT 18.980 316.600 19.330 317.200 ;
        RECT 18.980 316.400 22.930 316.600 ;
        RECT 18.980 315.800 19.330 316.400 ;
        RECT 18.980 315.600 22.930 315.800 ;
        RECT 18.980 315.000 19.330 315.600 ;
        RECT 23.930 315.550 24.330 319.200 ;
        RECT 25.130 319.200 44.330 319.600 ;
        RECT 25.130 315.550 25.530 319.200 ;
        RECT 29.180 319.150 31.480 319.200 ;
        RECT 37.980 319.150 40.280 319.200 ;
        RECT 26.530 318.000 42.930 318.600 ;
        RECT 30.130 317.400 30.480 318.000 ;
        RECT 26.530 317.200 30.480 317.400 ;
        RECT 30.130 316.600 30.480 317.200 ;
        RECT 26.530 316.400 30.480 316.600 ;
        RECT 30.130 315.800 30.480 316.400 ;
        RECT 26.530 315.600 30.480 315.800 ;
        RECT 18.980 314.800 22.930 315.000 ;
        RECT 18.980 314.200 19.330 314.800 ;
        RECT 18.980 314.000 22.930 314.200 ;
        RECT 18.980 313.400 19.330 314.000 ;
        RECT 18.980 313.200 22.930 313.400 ;
        RECT 23.880 313.250 25.580 315.550 ;
        RECT 30.130 315.000 30.480 315.600 ;
        RECT 26.530 314.800 30.480 315.000 ;
        RECT 30.130 314.200 30.480 314.800 ;
        RECT 26.530 314.000 30.480 314.200 ;
        RECT 30.130 313.400 30.480 314.000 ;
        RECT 18.980 312.600 19.330 313.200 ;
        RECT 18.980 312.400 22.930 312.600 ;
        RECT 18.980 311.800 19.330 312.400 ;
        RECT 18.980 311.600 22.930 311.800 ;
        RECT 18.980 311.000 19.330 311.600 ;
        RECT 18.980 310.800 22.930 311.000 ;
        RECT 18.980 310.400 19.330 310.800 ;
        RECT 15.780 302.000 15.980 309.600 ;
        RECT 16.580 302.000 16.780 309.600 ;
        RECT 17.380 302.000 17.580 309.600 ;
        RECT 18.180 302.000 18.380 309.600 ;
        RECT 18.980 309.200 19.330 309.600 ;
        RECT 18.980 309.000 22.930 309.200 ;
        RECT 18.980 308.400 19.330 309.000 ;
        RECT 18.980 308.200 22.930 308.400 ;
        RECT 18.980 307.600 19.330 308.200 ;
        RECT 18.980 307.400 22.930 307.600 ;
        RECT 18.980 306.800 19.330 307.400 ;
        RECT 18.980 306.600 22.930 306.800 ;
        RECT 23.930 306.750 24.330 313.250 ;
        RECT 25.130 306.750 25.530 313.250 ;
        RECT 26.530 313.200 30.480 313.400 ;
        RECT 30.130 312.600 30.480 313.200 ;
        RECT 26.530 312.400 30.480 312.600 ;
        RECT 30.130 311.800 30.480 312.400 ;
        RECT 26.530 311.600 30.480 311.800 ;
        RECT 30.130 311.000 30.480 311.600 ;
        RECT 26.530 310.800 30.480 311.000 ;
        RECT 30.130 310.400 30.480 310.800 ;
        RECT 31.080 310.400 31.280 318.000 ;
        RECT 31.880 310.400 32.080 318.000 ;
        RECT 32.680 310.400 32.880 318.000 ;
        RECT 33.480 310.400 33.680 318.000 ;
        RECT 30.130 309.200 30.480 309.600 ;
        RECT 26.530 309.000 30.480 309.200 ;
        RECT 30.130 308.400 30.480 309.000 ;
        RECT 26.530 308.200 30.480 308.400 ;
        RECT 30.130 307.600 30.480 308.200 ;
        RECT 26.530 307.400 30.480 307.600 ;
        RECT 30.130 306.800 30.480 307.400 ;
        RECT 18.980 306.000 19.330 306.600 ;
        RECT 18.980 305.800 22.930 306.000 ;
        RECT 18.980 305.200 19.330 305.800 ;
        RECT 18.980 305.000 22.930 305.200 ;
        RECT 18.980 304.400 19.330 305.000 ;
        RECT 23.880 304.450 25.580 306.750 ;
        RECT 26.530 306.600 30.480 306.800 ;
        RECT 30.130 306.000 30.480 306.600 ;
        RECT 26.530 305.800 30.480 306.000 ;
        RECT 30.130 305.200 30.480 305.800 ;
        RECT 26.530 305.000 30.480 305.200 ;
        RECT 18.980 304.200 22.930 304.400 ;
        RECT 18.980 303.600 19.330 304.200 ;
        RECT 18.980 303.400 22.930 303.600 ;
        RECT 18.980 302.800 19.330 303.400 ;
        RECT 18.980 302.600 22.930 302.800 ;
        RECT 18.980 302.000 19.330 302.600 ;
        RECT 6.530 301.400 22.930 302.000 ;
        RECT 9.180 300.800 11.480 300.850 ;
        RECT 17.980 300.800 20.280 300.850 ;
        RECT 23.930 300.800 24.330 304.450 ;
        RECT 5.130 300.400 24.330 300.800 ;
        RECT 25.130 300.800 25.530 304.450 ;
        RECT 30.130 304.400 30.480 305.000 ;
        RECT 26.530 304.200 30.480 304.400 ;
        RECT 30.130 303.600 30.480 304.200 ;
        RECT 26.530 303.400 30.480 303.600 ;
        RECT 30.130 302.800 30.480 303.400 ;
        RECT 26.530 302.600 30.480 302.800 ;
        RECT 30.130 302.000 30.480 302.600 ;
        RECT 31.080 302.000 31.280 309.600 ;
        RECT 31.880 302.000 32.080 309.600 ;
        RECT 32.680 302.000 32.880 309.600 ;
        RECT 33.480 302.000 33.680 309.600 ;
        RECT 34.280 302.000 35.180 318.000 ;
        RECT 35.780 310.400 35.980 318.000 ;
        RECT 36.580 310.400 36.780 318.000 ;
        RECT 37.380 310.400 37.580 318.000 ;
        RECT 38.180 310.400 38.380 318.000 ;
        RECT 38.980 317.400 39.330 318.000 ;
        RECT 38.980 317.200 42.930 317.400 ;
        RECT 38.980 316.600 39.330 317.200 ;
        RECT 38.980 316.400 42.930 316.600 ;
        RECT 38.980 315.800 39.330 316.400 ;
        RECT 38.980 315.600 42.930 315.800 ;
        RECT 38.980 315.000 39.330 315.600 ;
        RECT 43.930 315.550 44.330 319.200 ;
        RECT 45.130 319.200 64.330 319.600 ;
        RECT 45.130 315.550 45.530 319.200 ;
        RECT 49.180 319.150 51.480 319.200 ;
        RECT 57.980 319.150 60.280 319.200 ;
        RECT 46.530 318.000 62.930 318.600 ;
        RECT 50.130 317.400 50.480 318.000 ;
        RECT 46.530 317.200 50.480 317.400 ;
        RECT 50.130 316.600 50.480 317.200 ;
        RECT 46.530 316.400 50.480 316.600 ;
        RECT 50.130 315.800 50.480 316.400 ;
        RECT 46.530 315.600 50.480 315.800 ;
        RECT 38.980 314.800 42.930 315.000 ;
        RECT 38.980 314.200 39.330 314.800 ;
        RECT 38.980 314.000 42.930 314.200 ;
        RECT 38.980 313.400 39.330 314.000 ;
        RECT 38.980 313.200 42.930 313.400 ;
        RECT 43.880 313.250 45.580 315.550 ;
        RECT 50.130 315.000 50.480 315.600 ;
        RECT 46.530 314.800 50.480 315.000 ;
        RECT 50.130 314.200 50.480 314.800 ;
        RECT 46.530 314.000 50.480 314.200 ;
        RECT 50.130 313.400 50.480 314.000 ;
        RECT 38.980 312.600 39.330 313.200 ;
        RECT 38.980 312.400 42.930 312.600 ;
        RECT 38.980 311.800 39.330 312.400 ;
        RECT 38.980 311.600 42.930 311.800 ;
        RECT 38.980 311.000 39.330 311.600 ;
        RECT 38.980 310.800 42.930 311.000 ;
        RECT 38.980 310.400 39.330 310.800 ;
        RECT 35.780 302.000 35.980 309.600 ;
        RECT 36.580 302.000 36.780 309.600 ;
        RECT 37.380 302.000 37.580 309.600 ;
        RECT 38.180 302.000 38.380 309.600 ;
        RECT 38.980 309.200 39.330 309.600 ;
        RECT 38.980 309.000 42.930 309.200 ;
        RECT 38.980 308.400 39.330 309.000 ;
        RECT 38.980 308.200 42.930 308.400 ;
        RECT 38.980 307.600 39.330 308.200 ;
        RECT 38.980 307.400 42.930 307.600 ;
        RECT 38.980 306.800 39.330 307.400 ;
        RECT 38.980 306.600 42.930 306.800 ;
        RECT 43.930 306.750 44.330 313.250 ;
        RECT 45.130 306.750 45.530 313.250 ;
        RECT 46.530 313.200 50.480 313.400 ;
        RECT 50.130 312.600 50.480 313.200 ;
        RECT 46.530 312.400 50.480 312.600 ;
        RECT 50.130 311.800 50.480 312.400 ;
        RECT 46.530 311.600 50.480 311.800 ;
        RECT 50.130 311.000 50.480 311.600 ;
        RECT 46.530 310.800 50.480 311.000 ;
        RECT 50.130 310.400 50.480 310.800 ;
        RECT 51.080 310.400 51.280 318.000 ;
        RECT 51.880 310.400 52.080 318.000 ;
        RECT 52.680 310.400 52.880 318.000 ;
        RECT 53.480 310.400 53.680 318.000 ;
        RECT 50.130 309.200 50.480 309.600 ;
        RECT 46.530 309.000 50.480 309.200 ;
        RECT 50.130 308.400 50.480 309.000 ;
        RECT 46.530 308.200 50.480 308.400 ;
        RECT 50.130 307.600 50.480 308.200 ;
        RECT 46.530 307.400 50.480 307.600 ;
        RECT 50.130 306.800 50.480 307.400 ;
        RECT 38.980 306.000 39.330 306.600 ;
        RECT 38.980 305.800 42.930 306.000 ;
        RECT 38.980 305.200 39.330 305.800 ;
        RECT 38.980 305.000 42.930 305.200 ;
        RECT 38.980 304.400 39.330 305.000 ;
        RECT 43.880 304.450 45.580 306.750 ;
        RECT 46.530 306.600 50.480 306.800 ;
        RECT 50.130 306.000 50.480 306.600 ;
        RECT 46.530 305.800 50.480 306.000 ;
        RECT 50.130 305.200 50.480 305.800 ;
        RECT 46.530 305.000 50.480 305.200 ;
        RECT 38.980 304.200 42.930 304.400 ;
        RECT 38.980 303.600 39.330 304.200 ;
        RECT 38.980 303.400 42.930 303.600 ;
        RECT 38.980 302.800 39.330 303.400 ;
        RECT 38.980 302.600 42.930 302.800 ;
        RECT 38.980 302.000 39.330 302.600 ;
        RECT 26.530 301.400 42.930 302.000 ;
        RECT 29.180 300.800 31.480 300.850 ;
        RECT 37.980 300.800 40.280 300.850 ;
        RECT 43.930 300.800 44.330 304.450 ;
        RECT 25.130 300.400 44.330 300.800 ;
        RECT 45.130 300.800 45.530 304.450 ;
        RECT 50.130 304.400 50.480 305.000 ;
        RECT 46.530 304.200 50.480 304.400 ;
        RECT 50.130 303.600 50.480 304.200 ;
        RECT 46.530 303.400 50.480 303.600 ;
        RECT 50.130 302.800 50.480 303.400 ;
        RECT 46.530 302.600 50.480 302.800 ;
        RECT 50.130 302.000 50.480 302.600 ;
        RECT 51.080 302.000 51.280 309.600 ;
        RECT 51.880 302.000 52.080 309.600 ;
        RECT 52.680 302.000 52.880 309.600 ;
        RECT 53.480 302.000 53.680 309.600 ;
        RECT 54.280 302.000 55.180 318.000 ;
        RECT 55.780 310.400 55.980 318.000 ;
        RECT 56.580 310.400 56.780 318.000 ;
        RECT 57.380 310.400 57.580 318.000 ;
        RECT 58.180 310.400 58.380 318.000 ;
        RECT 58.980 317.400 59.330 318.000 ;
        RECT 58.980 317.200 62.930 317.400 ;
        RECT 58.980 316.600 59.330 317.200 ;
        RECT 58.980 316.400 62.930 316.600 ;
        RECT 58.980 315.800 59.330 316.400 ;
        RECT 58.980 315.600 62.930 315.800 ;
        RECT 58.980 315.000 59.330 315.600 ;
        RECT 63.930 315.550 64.330 319.200 ;
        RECT 65.130 319.200 84.330 319.600 ;
        RECT 65.130 315.550 65.530 319.200 ;
        RECT 69.180 319.150 71.480 319.200 ;
        RECT 77.980 319.150 80.280 319.200 ;
        RECT 66.530 318.000 82.930 318.600 ;
        RECT 70.130 317.400 70.480 318.000 ;
        RECT 66.530 317.200 70.480 317.400 ;
        RECT 70.130 316.600 70.480 317.200 ;
        RECT 66.530 316.400 70.480 316.600 ;
        RECT 70.130 315.800 70.480 316.400 ;
        RECT 66.530 315.600 70.480 315.800 ;
        RECT 58.980 314.800 62.930 315.000 ;
        RECT 58.980 314.200 59.330 314.800 ;
        RECT 58.980 314.000 62.930 314.200 ;
        RECT 58.980 313.400 59.330 314.000 ;
        RECT 58.980 313.200 62.930 313.400 ;
        RECT 63.880 313.250 65.580 315.550 ;
        RECT 70.130 315.000 70.480 315.600 ;
        RECT 66.530 314.800 70.480 315.000 ;
        RECT 70.130 314.200 70.480 314.800 ;
        RECT 66.530 314.000 70.480 314.200 ;
        RECT 70.130 313.400 70.480 314.000 ;
        RECT 58.980 312.600 59.330 313.200 ;
        RECT 58.980 312.400 62.930 312.600 ;
        RECT 58.980 311.800 59.330 312.400 ;
        RECT 58.980 311.600 62.930 311.800 ;
        RECT 58.980 311.000 59.330 311.600 ;
        RECT 58.980 310.800 62.930 311.000 ;
        RECT 58.980 310.400 59.330 310.800 ;
        RECT 55.780 302.000 55.980 309.600 ;
        RECT 56.580 302.000 56.780 309.600 ;
        RECT 57.380 302.000 57.580 309.600 ;
        RECT 58.180 302.000 58.380 309.600 ;
        RECT 58.980 309.200 59.330 309.600 ;
        RECT 58.980 309.000 62.930 309.200 ;
        RECT 58.980 308.400 59.330 309.000 ;
        RECT 58.980 308.200 62.930 308.400 ;
        RECT 58.980 307.600 59.330 308.200 ;
        RECT 58.980 307.400 62.930 307.600 ;
        RECT 58.980 306.800 59.330 307.400 ;
        RECT 58.980 306.600 62.930 306.800 ;
        RECT 63.930 306.750 64.330 313.250 ;
        RECT 65.130 306.750 65.530 313.250 ;
        RECT 66.530 313.200 70.480 313.400 ;
        RECT 70.130 312.600 70.480 313.200 ;
        RECT 66.530 312.400 70.480 312.600 ;
        RECT 70.130 311.800 70.480 312.400 ;
        RECT 66.530 311.600 70.480 311.800 ;
        RECT 70.130 311.000 70.480 311.600 ;
        RECT 66.530 310.800 70.480 311.000 ;
        RECT 70.130 310.400 70.480 310.800 ;
        RECT 71.080 310.400 71.280 318.000 ;
        RECT 71.880 310.400 72.080 318.000 ;
        RECT 72.680 310.400 72.880 318.000 ;
        RECT 73.480 310.400 73.680 318.000 ;
        RECT 70.130 309.200 70.480 309.600 ;
        RECT 66.530 309.000 70.480 309.200 ;
        RECT 70.130 308.400 70.480 309.000 ;
        RECT 66.530 308.200 70.480 308.400 ;
        RECT 70.130 307.600 70.480 308.200 ;
        RECT 66.530 307.400 70.480 307.600 ;
        RECT 70.130 306.800 70.480 307.400 ;
        RECT 58.980 306.000 59.330 306.600 ;
        RECT 58.980 305.800 62.930 306.000 ;
        RECT 58.980 305.200 59.330 305.800 ;
        RECT 58.980 305.000 62.930 305.200 ;
        RECT 58.980 304.400 59.330 305.000 ;
        RECT 63.880 304.450 65.580 306.750 ;
        RECT 66.530 306.600 70.480 306.800 ;
        RECT 70.130 306.000 70.480 306.600 ;
        RECT 66.530 305.800 70.480 306.000 ;
        RECT 70.130 305.200 70.480 305.800 ;
        RECT 66.530 305.000 70.480 305.200 ;
        RECT 58.980 304.200 62.930 304.400 ;
        RECT 58.980 303.600 59.330 304.200 ;
        RECT 58.980 303.400 62.930 303.600 ;
        RECT 58.980 302.800 59.330 303.400 ;
        RECT 58.980 302.600 62.930 302.800 ;
        RECT 58.980 302.000 59.330 302.600 ;
        RECT 46.530 301.400 62.930 302.000 ;
        RECT 49.180 300.800 51.480 300.850 ;
        RECT 57.980 300.800 60.280 300.850 ;
        RECT 63.930 300.800 64.330 304.450 ;
        RECT 45.130 300.400 64.330 300.800 ;
        RECT 65.130 300.800 65.530 304.450 ;
        RECT 70.130 304.400 70.480 305.000 ;
        RECT 66.530 304.200 70.480 304.400 ;
        RECT 70.130 303.600 70.480 304.200 ;
        RECT 66.530 303.400 70.480 303.600 ;
        RECT 70.130 302.800 70.480 303.400 ;
        RECT 66.530 302.600 70.480 302.800 ;
        RECT 70.130 302.000 70.480 302.600 ;
        RECT 71.080 302.000 71.280 309.600 ;
        RECT 71.880 302.000 72.080 309.600 ;
        RECT 72.680 302.000 72.880 309.600 ;
        RECT 73.480 302.000 73.680 309.600 ;
        RECT 74.280 302.000 75.180 318.000 ;
        RECT 75.780 310.400 75.980 318.000 ;
        RECT 76.580 310.400 76.780 318.000 ;
        RECT 77.380 310.400 77.580 318.000 ;
        RECT 78.180 310.400 78.380 318.000 ;
        RECT 78.980 317.400 79.330 318.000 ;
        RECT 78.980 317.200 82.930 317.400 ;
        RECT 78.980 316.600 79.330 317.200 ;
        RECT 78.980 316.400 82.930 316.600 ;
        RECT 78.980 315.800 79.330 316.400 ;
        RECT 78.980 315.600 82.930 315.800 ;
        RECT 78.980 315.000 79.330 315.600 ;
        RECT 83.930 315.550 84.330 319.200 ;
        RECT 85.130 319.200 104.330 319.600 ;
        RECT 85.130 315.550 85.530 319.200 ;
        RECT 89.180 319.150 91.480 319.200 ;
        RECT 97.980 319.150 100.280 319.200 ;
        RECT 86.530 318.000 102.930 318.600 ;
        RECT 90.130 317.400 90.480 318.000 ;
        RECT 86.530 317.200 90.480 317.400 ;
        RECT 90.130 316.600 90.480 317.200 ;
        RECT 86.530 316.400 90.480 316.600 ;
        RECT 90.130 315.800 90.480 316.400 ;
        RECT 86.530 315.600 90.480 315.800 ;
        RECT 78.980 314.800 82.930 315.000 ;
        RECT 78.980 314.200 79.330 314.800 ;
        RECT 78.980 314.000 82.930 314.200 ;
        RECT 78.980 313.400 79.330 314.000 ;
        RECT 78.980 313.200 82.930 313.400 ;
        RECT 83.880 313.250 85.580 315.550 ;
        RECT 90.130 315.000 90.480 315.600 ;
        RECT 86.530 314.800 90.480 315.000 ;
        RECT 90.130 314.200 90.480 314.800 ;
        RECT 86.530 314.000 90.480 314.200 ;
        RECT 90.130 313.400 90.480 314.000 ;
        RECT 78.980 312.600 79.330 313.200 ;
        RECT 78.980 312.400 82.930 312.600 ;
        RECT 78.980 311.800 79.330 312.400 ;
        RECT 78.980 311.600 82.930 311.800 ;
        RECT 78.980 311.000 79.330 311.600 ;
        RECT 78.980 310.800 82.930 311.000 ;
        RECT 78.980 310.400 79.330 310.800 ;
        RECT 75.780 302.000 75.980 309.600 ;
        RECT 76.580 302.000 76.780 309.600 ;
        RECT 77.380 302.000 77.580 309.600 ;
        RECT 78.180 302.000 78.380 309.600 ;
        RECT 78.980 309.200 79.330 309.600 ;
        RECT 78.980 309.000 82.930 309.200 ;
        RECT 78.980 308.400 79.330 309.000 ;
        RECT 78.980 308.200 82.930 308.400 ;
        RECT 78.980 307.600 79.330 308.200 ;
        RECT 78.980 307.400 82.930 307.600 ;
        RECT 78.980 306.800 79.330 307.400 ;
        RECT 78.980 306.600 82.930 306.800 ;
        RECT 83.930 306.750 84.330 313.250 ;
        RECT 85.130 306.750 85.530 313.250 ;
        RECT 86.530 313.200 90.480 313.400 ;
        RECT 90.130 312.600 90.480 313.200 ;
        RECT 86.530 312.400 90.480 312.600 ;
        RECT 90.130 311.800 90.480 312.400 ;
        RECT 86.530 311.600 90.480 311.800 ;
        RECT 90.130 311.000 90.480 311.600 ;
        RECT 86.530 310.800 90.480 311.000 ;
        RECT 90.130 310.400 90.480 310.800 ;
        RECT 91.080 310.400 91.280 318.000 ;
        RECT 91.880 310.400 92.080 318.000 ;
        RECT 92.680 310.400 92.880 318.000 ;
        RECT 93.480 310.400 93.680 318.000 ;
        RECT 90.130 309.200 90.480 309.600 ;
        RECT 86.530 309.000 90.480 309.200 ;
        RECT 90.130 308.400 90.480 309.000 ;
        RECT 86.530 308.200 90.480 308.400 ;
        RECT 90.130 307.600 90.480 308.200 ;
        RECT 86.530 307.400 90.480 307.600 ;
        RECT 90.130 306.800 90.480 307.400 ;
        RECT 78.980 306.000 79.330 306.600 ;
        RECT 78.980 305.800 82.930 306.000 ;
        RECT 78.980 305.200 79.330 305.800 ;
        RECT 78.980 305.000 82.930 305.200 ;
        RECT 78.980 304.400 79.330 305.000 ;
        RECT 83.880 304.450 85.580 306.750 ;
        RECT 86.530 306.600 90.480 306.800 ;
        RECT 90.130 306.000 90.480 306.600 ;
        RECT 86.530 305.800 90.480 306.000 ;
        RECT 90.130 305.200 90.480 305.800 ;
        RECT 86.530 305.000 90.480 305.200 ;
        RECT 78.980 304.200 82.930 304.400 ;
        RECT 78.980 303.600 79.330 304.200 ;
        RECT 78.980 303.400 82.930 303.600 ;
        RECT 78.980 302.800 79.330 303.400 ;
        RECT 78.980 302.600 82.930 302.800 ;
        RECT 78.980 302.000 79.330 302.600 ;
        RECT 66.530 301.400 82.930 302.000 ;
        RECT 69.180 300.800 71.480 300.850 ;
        RECT 77.980 300.800 80.280 300.850 ;
        RECT 83.930 300.800 84.330 304.450 ;
        RECT 65.130 300.400 84.330 300.800 ;
        RECT 85.130 300.800 85.530 304.450 ;
        RECT 90.130 304.400 90.480 305.000 ;
        RECT 86.530 304.200 90.480 304.400 ;
        RECT 90.130 303.600 90.480 304.200 ;
        RECT 86.530 303.400 90.480 303.600 ;
        RECT 90.130 302.800 90.480 303.400 ;
        RECT 86.530 302.600 90.480 302.800 ;
        RECT 90.130 302.000 90.480 302.600 ;
        RECT 91.080 302.000 91.280 309.600 ;
        RECT 91.880 302.000 92.080 309.600 ;
        RECT 92.680 302.000 92.880 309.600 ;
        RECT 93.480 302.000 93.680 309.600 ;
        RECT 94.280 302.000 95.180 318.000 ;
        RECT 95.780 310.400 95.980 318.000 ;
        RECT 96.580 310.400 96.780 318.000 ;
        RECT 97.380 310.400 97.580 318.000 ;
        RECT 98.180 310.400 98.380 318.000 ;
        RECT 98.980 317.400 99.330 318.000 ;
        RECT 98.980 317.200 102.930 317.400 ;
        RECT 98.980 316.600 99.330 317.200 ;
        RECT 98.980 316.400 102.930 316.600 ;
        RECT 98.980 315.800 99.330 316.400 ;
        RECT 98.980 315.600 102.930 315.800 ;
        RECT 98.980 315.000 99.330 315.600 ;
        RECT 103.930 315.550 104.330 319.200 ;
        RECT 105.130 319.200 124.330 319.600 ;
        RECT 105.130 315.550 105.530 319.200 ;
        RECT 109.180 319.150 111.480 319.200 ;
        RECT 117.980 319.150 120.280 319.200 ;
        RECT 106.530 318.000 122.930 318.600 ;
        RECT 110.130 317.400 110.480 318.000 ;
        RECT 106.530 317.200 110.480 317.400 ;
        RECT 110.130 316.600 110.480 317.200 ;
        RECT 106.530 316.400 110.480 316.600 ;
        RECT 110.130 315.800 110.480 316.400 ;
        RECT 106.530 315.600 110.480 315.800 ;
        RECT 98.980 314.800 102.930 315.000 ;
        RECT 98.980 314.200 99.330 314.800 ;
        RECT 98.980 314.000 102.930 314.200 ;
        RECT 98.980 313.400 99.330 314.000 ;
        RECT 98.980 313.200 102.930 313.400 ;
        RECT 103.880 313.250 105.580 315.550 ;
        RECT 110.130 315.000 110.480 315.600 ;
        RECT 106.530 314.800 110.480 315.000 ;
        RECT 110.130 314.200 110.480 314.800 ;
        RECT 106.530 314.000 110.480 314.200 ;
        RECT 110.130 313.400 110.480 314.000 ;
        RECT 98.980 312.600 99.330 313.200 ;
        RECT 98.980 312.400 102.930 312.600 ;
        RECT 98.980 311.800 99.330 312.400 ;
        RECT 98.980 311.600 102.930 311.800 ;
        RECT 98.980 311.000 99.330 311.600 ;
        RECT 98.980 310.800 102.930 311.000 ;
        RECT 98.980 310.400 99.330 310.800 ;
        RECT 95.780 302.000 95.980 309.600 ;
        RECT 96.580 302.000 96.780 309.600 ;
        RECT 97.380 302.000 97.580 309.600 ;
        RECT 98.180 302.000 98.380 309.600 ;
        RECT 98.980 309.200 99.330 309.600 ;
        RECT 98.980 309.000 102.930 309.200 ;
        RECT 98.980 308.400 99.330 309.000 ;
        RECT 98.980 308.200 102.930 308.400 ;
        RECT 98.980 307.600 99.330 308.200 ;
        RECT 98.980 307.400 102.930 307.600 ;
        RECT 98.980 306.800 99.330 307.400 ;
        RECT 98.980 306.600 102.930 306.800 ;
        RECT 103.930 306.750 104.330 313.250 ;
        RECT 105.130 306.750 105.530 313.250 ;
        RECT 106.530 313.200 110.480 313.400 ;
        RECT 110.130 312.600 110.480 313.200 ;
        RECT 106.530 312.400 110.480 312.600 ;
        RECT 110.130 311.800 110.480 312.400 ;
        RECT 106.530 311.600 110.480 311.800 ;
        RECT 110.130 311.000 110.480 311.600 ;
        RECT 106.530 310.800 110.480 311.000 ;
        RECT 110.130 310.400 110.480 310.800 ;
        RECT 111.080 310.400 111.280 318.000 ;
        RECT 111.880 310.400 112.080 318.000 ;
        RECT 112.680 310.400 112.880 318.000 ;
        RECT 113.480 310.400 113.680 318.000 ;
        RECT 110.130 309.200 110.480 309.600 ;
        RECT 106.530 309.000 110.480 309.200 ;
        RECT 110.130 308.400 110.480 309.000 ;
        RECT 106.530 308.200 110.480 308.400 ;
        RECT 110.130 307.600 110.480 308.200 ;
        RECT 106.530 307.400 110.480 307.600 ;
        RECT 110.130 306.800 110.480 307.400 ;
        RECT 98.980 306.000 99.330 306.600 ;
        RECT 98.980 305.800 102.930 306.000 ;
        RECT 98.980 305.200 99.330 305.800 ;
        RECT 98.980 305.000 102.930 305.200 ;
        RECT 98.980 304.400 99.330 305.000 ;
        RECT 103.880 304.450 105.580 306.750 ;
        RECT 106.530 306.600 110.480 306.800 ;
        RECT 110.130 306.000 110.480 306.600 ;
        RECT 106.530 305.800 110.480 306.000 ;
        RECT 110.130 305.200 110.480 305.800 ;
        RECT 106.530 305.000 110.480 305.200 ;
        RECT 98.980 304.200 102.930 304.400 ;
        RECT 98.980 303.600 99.330 304.200 ;
        RECT 98.980 303.400 102.930 303.600 ;
        RECT 98.980 302.800 99.330 303.400 ;
        RECT 98.980 302.600 102.930 302.800 ;
        RECT 98.980 302.000 99.330 302.600 ;
        RECT 86.530 301.400 102.930 302.000 ;
        RECT 89.180 300.800 91.480 300.850 ;
        RECT 97.980 300.800 100.280 300.850 ;
        RECT 103.930 300.800 104.330 304.450 ;
        RECT 85.130 300.400 104.330 300.800 ;
        RECT 105.130 300.800 105.530 304.450 ;
        RECT 110.130 304.400 110.480 305.000 ;
        RECT 106.530 304.200 110.480 304.400 ;
        RECT 110.130 303.600 110.480 304.200 ;
        RECT 106.530 303.400 110.480 303.600 ;
        RECT 110.130 302.800 110.480 303.400 ;
        RECT 106.530 302.600 110.480 302.800 ;
        RECT 110.130 302.000 110.480 302.600 ;
        RECT 111.080 302.000 111.280 309.600 ;
        RECT 111.880 302.000 112.080 309.600 ;
        RECT 112.680 302.000 112.880 309.600 ;
        RECT 113.480 302.000 113.680 309.600 ;
        RECT 114.280 302.000 115.180 318.000 ;
        RECT 115.780 310.400 115.980 318.000 ;
        RECT 116.580 310.400 116.780 318.000 ;
        RECT 117.380 310.400 117.580 318.000 ;
        RECT 118.180 310.400 118.380 318.000 ;
        RECT 118.980 317.400 119.330 318.000 ;
        RECT 118.980 317.200 122.930 317.400 ;
        RECT 118.980 316.600 119.330 317.200 ;
        RECT 118.980 316.400 122.930 316.600 ;
        RECT 118.980 315.800 119.330 316.400 ;
        RECT 118.980 315.600 122.930 315.800 ;
        RECT 118.980 315.000 119.330 315.600 ;
        RECT 123.930 315.550 124.330 319.200 ;
        RECT 125.340 317.080 125.700 317.460 ;
        RECT 125.970 317.080 126.330 317.460 ;
        RECT 126.570 317.080 126.930 317.460 ;
        RECT 125.340 316.490 125.700 316.870 ;
        RECT 125.970 316.490 126.330 316.870 ;
        RECT 126.570 316.490 126.930 316.870 ;
        RECT 118.980 314.800 122.930 315.000 ;
        RECT 118.980 314.200 119.330 314.800 ;
        RECT 118.980 314.000 122.930 314.200 ;
        RECT 118.980 313.400 119.330 314.000 ;
        RECT 118.980 313.200 122.930 313.400 ;
        RECT 123.880 313.250 124.730 315.550 ;
        RECT 118.980 312.600 119.330 313.200 ;
        RECT 118.980 312.400 122.930 312.600 ;
        RECT 118.980 311.800 119.330 312.400 ;
        RECT 118.980 311.600 122.930 311.800 ;
        RECT 118.980 311.000 119.330 311.600 ;
        RECT 118.980 310.800 122.930 311.000 ;
        RECT 118.980 310.400 119.330 310.800 ;
        RECT 115.780 302.000 115.980 309.600 ;
        RECT 116.580 302.000 116.780 309.600 ;
        RECT 117.380 302.000 117.580 309.600 ;
        RECT 118.180 302.000 118.380 309.600 ;
        RECT 118.980 309.200 119.330 309.600 ;
        RECT 118.980 309.000 122.930 309.200 ;
        RECT 118.980 308.400 119.330 309.000 ;
        RECT 118.980 308.200 122.930 308.400 ;
        RECT 118.980 307.600 119.330 308.200 ;
        RECT 118.980 307.400 122.930 307.600 ;
        RECT 118.980 306.800 119.330 307.400 ;
        RECT 118.980 306.600 122.930 306.800 ;
        RECT 123.930 306.750 124.330 313.250 ;
        RECT 118.980 306.000 119.330 306.600 ;
        RECT 118.980 305.800 122.930 306.000 ;
        RECT 118.980 305.200 119.330 305.800 ;
        RECT 118.980 305.000 122.930 305.200 ;
        RECT 118.980 304.400 119.330 305.000 ;
        RECT 123.880 304.450 124.730 306.750 ;
        RECT 118.980 304.200 122.930 304.400 ;
        RECT 118.980 303.600 119.330 304.200 ;
        RECT 118.980 303.400 122.930 303.600 ;
        RECT 118.980 302.800 119.330 303.400 ;
        RECT 118.980 302.600 122.930 302.800 ;
        RECT 118.980 302.000 119.330 302.600 ;
        RECT 106.530 301.400 122.930 302.000 ;
        RECT 109.180 300.800 111.480 300.850 ;
        RECT 117.980 300.800 120.280 300.850 ;
        RECT 123.930 300.800 124.330 304.450 ;
        RECT 125.340 303.095 125.700 303.475 ;
        RECT 125.970 303.095 126.330 303.475 ;
        RECT 126.570 303.095 126.930 303.475 ;
        RECT 125.340 302.505 125.700 302.885 ;
        RECT 125.970 302.505 126.330 302.885 ;
        RECT 126.570 302.505 126.930 302.885 ;
        RECT 105.130 300.400 124.330 300.800 ;
        RECT 9.180 299.600 11.480 300.400 ;
        RECT 17.980 299.600 20.280 300.400 ;
        RECT 29.180 299.600 31.480 300.400 ;
        RECT 37.980 299.600 40.280 300.400 ;
        RECT 49.180 299.600 51.480 300.400 ;
        RECT 57.980 299.600 60.280 300.400 ;
        RECT 69.180 299.600 71.480 300.400 ;
        RECT 77.980 299.600 80.280 300.400 ;
        RECT 89.180 299.600 91.480 300.400 ;
        RECT 97.980 299.600 100.280 300.400 ;
        RECT 109.180 299.600 111.480 300.400 ;
        RECT 117.980 299.600 120.280 300.400 ;
        RECT 5.130 299.200 24.330 299.600 ;
        RECT 2.515 297.280 2.875 297.660 ;
        RECT 3.145 297.280 3.505 297.660 ;
        RECT 3.745 297.280 4.105 297.660 ;
        RECT 2.515 296.690 2.875 297.070 ;
        RECT 3.145 296.690 3.505 297.070 ;
        RECT 3.745 296.690 4.105 297.070 ;
        RECT 5.130 295.550 5.530 299.200 ;
        RECT 9.180 299.150 11.480 299.200 ;
        RECT 17.980 299.150 20.280 299.200 ;
        RECT 6.530 298.000 22.930 298.600 ;
        RECT 10.130 297.400 10.480 298.000 ;
        RECT 6.530 297.200 10.480 297.400 ;
        RECT 10.130 296.600 10.480 297.200 ;
        RECT 6.530 296.400 10.480 296.600 ;
        RECT 10.130 295.800 10.480 296.400 ;
        RECT 6.530 295.600 10.480 295.800 ;
        RECT 4.730 295.545 5.580 295.550 ;
        RECT 2.320 295.340 5.580 295.545 ;
        RECT 2.315 293.250 5.580 295.340 ;
        RECT 10.130 295.000 10.480 295.600 ;
        RECT 6.530 294.800 10.480 295.000 ;
        RECT 10.130 294.200 10.480 294.800 ;
        RECT 6.530 294.000 10.480 294.200 ;
        RECT 10.130 293.400 10.480 294.000 ;
        RECT 5.130 286.750 5.530 293.250 ;
        RECT 6.530 293.200 10.480 293.400 ;
        RECT 10.130 292.600 10.480 293.200 ;
        RECT 6.530 292.400 10.480 292.600 ;
        RECT 10.130 291.800 10.480 292.400 ;
        RECT 6.530 291.600 10.480 291.800 ;
        RECT 10.130 291.000 10.480 291.600 ;
        RECT 6.530 290.800 10.480 291.000 ;
        RECT 10.130 290.400 10.480 290.800 ;
        RECT 11.080 290.400 11.280 298.000 ;
        RECT 11.880 290.400 12.080 298.000 ;
        RECT 12.680 290.400 12.880 298.000 ;
        RECT 13.480 290.400 13.680 298.000 ;
        RECT 10.130 289.200 10.480 289.600 ;
        RECT 6.530 289.000 10.480 289.200 ;
        RECT 10.130 288.400 10.480 289.000 ;
        RECT 6.530 288.200 10.480 288.400 ;
        RECT 10.130 287.600 10.480 288.200 ;
        RECT 6.530 287.400 10.480 287.600 ;
        RECT 10.130 286.800 10.480 287.400 ;
        RECT 2.315 284.455 5.580 286.750 ;
        RECT 6.530 286.600 10.480 286.800 ;
        RECT 10.130 286.000 10.480 286.600 ;
        RECT 6.530 285.800 10.480 286.000 ;
        RECT 10.130 285.200 10.480 285.800 ;
        RECT 6.530 285.000 10.480 285.200 ;
        RECT 4.730 284.450 5.580 284.455 ;
        RECT 2.515 283.040 2.875 283.420 ;
        RECT 3.145 283.040 3.505 283.420 ;
        RECT 3.745 283.040 4.105 283.420 ;
        RECT 2.515 282.450 2.875 282.830 ;
        RECT 3.145 282.450 3.505 282.830 ;
        RECT 3.745 282.450 4.105 282.830 ;
        RECT 5.130 280.800 5.530 284.450 ;
        RECT 10.130 284.400 10.480 285.000 ;
        RECT 6.530 284.200 10.480 284.400 ;
        RECT 10.130 283.600 10.480 284.200 ;
        RECT 6.530 283.400 10.480 283.600 ;
        RECT 10.130 282.800 10.480 283.400 ;
        RECT 6.530 282.600 10.480 282.800 ;
        RECT 10.130 282.000 10.480 282.600 ;
        RECT 11.080 282.000 11.280 289.600 ;
        RECT 11.880 282.000 12.080 289.600 ;
        RECT 12.680 282.000 12.880 289.600 ;
        RECT 13.480 282.000 13.680 289.600 ;
        RECT 14.280 282.000 15.180 298.000 ;
        RECT 15.780 290.400 15.980 298.000 ;
        RECT 16.580 290.400 16.780 298.000 ;
        RECT 17.380 290.400 17.580 298.000 ;
        RECT 18.180 290.400 18.380 298.000 ;
        RECT 18.980 297.400 19.330 298.000 ;
        RECT 18.980 297.200 22.930 297.400 ;
        RECT 18.980 296.600 19.330 297.200 ;
        RECT 18.980 296.400 22.930 296.600 ;
        RECT 18.980 295.800 19.330 296.400 ;
        RECT 18.980 295.600 22.930 295.800 ;
        RECT 18.980 295.000 19.330 295.600 ;
        RECT 23.930 295.550 24.330 299.200 ;
        RECT 25.130 299.200 44.330 299.600 ;
        RECT 25.130 295.550 25.530 299.200 ;
        RECT 29.180 299.150 31.480 299.200 ;
        RECT 37.980 299.150 40.280 299.200 ;
        RECT 26.530 298.000 42.930 298.600 ;
        RECT 30.130 297.400 30.480 298.000 ;
        RECT 26.530 297.200 30.480 297.400 ;
        RECT 30.130 296.600 30.480 297.200 ;
        RECT 26.530 296.400 30.480 296.600 ;
        RECT 30.130 295.800 30.480 296.400 ;
        RECT 26.530 295.600 30.480 295.800 ;
        RECT 18.980 294.800 22.930 295.000 ;
        RECT 18.980 294.200 19.330 294.800 ;
        RECT 18.980 294.000 22.930 294.200 ;
        RECT 18.980 293.400 19.330 294.000 ;
        RECT 18.980 293.200 22.930 293.400 ;
        RECT 23.880 293.250 25.580 295.550 ;
        RECT 30.130 295.000 30.480 295.600 ;
        RECT 26.530 294.800 30.480 295.000 ;
        RECT 30.130 294.200 30.480 294.800 ;
        RECT 26.530 294.000 30.480 294.200 ;
        RECT 30.130 293.400 30.480 294.000 ;
        RECT 18.980 292.600 19.330 293.200 ;
        RECT 18.980 292.400 22.930 292.600 ;
        RECT 18.980 291.800 19.330 292.400 ;
        RECT 18.980 291.600 22.930 291.800 ;
        RECT 18.980 291.000 19.330 291.600 ;
        RECT 18.980 290.800 22.930 291.000 ;
        RECT 18.980 290.400 19.330 290.800 ;
        RECT 15.780 282.000 15.980 289.600 ;
        RECT 16.580 282.000 16.780 289.600 ;
        RECT 17.380 282.000 17.580 289.600 ;
        RECT 18.180 282.000 18.380 289.600 ;
        RECT 18.980 289.200 19.330 289.600 ;
        RECT 18.980 289.000 22.930 289.200 ;
        RECT 18.980 288.400 19.330 289.000 ;
        RECT 18.980 288.200 22.930 288.400 ;
        RECT 18.980 287.600 19.330 288.200 ;
        RECT 18.980 287.400 22.930 287.600 ;
        RECT 18.980 286.800 19.330 287.400 ;
        RECT 18.980 286.600 22.930 286.800 ;
        RECT 23.930 286.750 24.330 293.250 ;
        RECT 25.130 286.750 25.530 293.250 ;
        RECT 26.530 293.200 30.480 293.400 ;
        RECT 30.130 292.600 30.480 293.200 ;
        RECT 26.530 292.400 30.480 292.600 ;
        RECT 30.130 291.800 30.480 292.400 ;
        RECT 26.530 291.600 30.480 291.800 ;
        RECT 30.130 291.000 30.480 291.600 ;
        RECT 26.530 290.800 30.480 291.000 ;
        RECT 30.130 290.400 30.480 290.800 ;
        RECT 31.080 290.400 31.280 298.000 ;
        RECT 31.880 290.400 32.080 298.000 ;
        RECT 32.680 290.400 32.880 298.000 ;
        RECT 33.480 290.400 33.680 298.000 ;
        RECT 30.130 289.200 30.480 289.600 ;
        RECT 26.530 289.000 30.480 289.200 ;
        RECT 30.130 288.400 30.480 289.000 ;
        RECT 26.530 288.200 30.480 288.400 ;
        RECT 30.130 287.600 30.480 288.200 ;
        RECT 26.530 287.400 30.480 287.600 ;
        RECT 30.130 286.800 30.480 287.400 ;
        RECT 18.980 286.000 19.330 286.600 ;
        RECT 18.980 285.800 22.930 286.000 ;
        RECT 18.980 285.200 19.330 285.800 ;
        RECT 18.980 285.000 22.930 285.200 ;
        RECT 18.980 284.400 19.330 285.000 ;
        RECT 23.880 284.450 25.580 286.750 ;
        RECT 26.530 286.600 30.480 286.800 ;
        RECT 30.130 286.000 30.480 286.600 ;
        RECT 26.530 285.800 30.480 286.000 ;
        RECT 30.130 285.200 30.480 285.800 ;
        RECT 26.530 285.000 30.480 285.200 ;
        RECT 18.980 284.200 22.930 284.400 ;
        RECT 18.980 283.600 19.330 284.200 ;
        RECT 18.980 283.400 22.930 283.600 ;
        RECT 18.980 282.800 19.330 283.400 ;
        RECT 18.980 282.600 22.930 282.800 ;
        RECT 18.980 282.000 19.330 282.600 ;
        RECT 6.530 281.400 22.930 282.000 ;
        RECT 9.180 280.800 11.480 280.850 ;
        RECT 17.980 280.800 20.280 280.850 ;
        RECT 23.930 280.800 24.330 284.450 ;
        RECT 5.130 280.400 24.330 280.800 ;
        RECT 25.130 280.800 25.530 284.450 ;
        RECT 30.130 284.400 30.480 285.000 ;
        RECT 26.530 284.200 30.480 284.400 ;
        RECT 30.130 283.600 30.480 284.200 ;
        RECT 26.530 283.400 30.480 283.600 ;
        RECT 30.130 282.800 30.480 283.400 ;
        RECT 26.530 282.600 30.480 282.800 ;
        RECT 30.130 282.000 30.480 282.600 ;
        RECT 31.080 282.000 31.280 289.600 ;
        RECT 31.880 282.000 32.080 289.600 ;
        RECT 32.680 282.000 32.880 289.600 ;
        RECT 33.480 282.000 33.680 289.600 ;
        RECT 34.280 282.000 35.180 298.000 ;
        RECT 35.780 290.400 35.980 298.000 ;
        RECT 36.580 290.400 36.780 298.000 ;
        RECT 37.380 290.400 37.580 298.000 ;
        RECT 38.180 290.400 38.380 298.000 ;
        RECT 38.980 297.400 39.330 298.000 ;
        RECT 38.980 297.200 42.930 297.400 ;
        RECT 38.980 296.600 39.330 297.200 ;
        RECT 38.980 296.400 42.930 296.600 ;
        RECT 38.980 295.800 39.330 296.400 ;
        RECT 38.980 295.600 42.930 295.800 ;
        RECT 38.980 295.000 39.330 295.600 ;
        RECT 43.930 295.550 44.330 299.200 ;
        RECT 45.130 299.200 64.330 299.600 ;
        RECT 45.130 295.550 45.530 299.200 ;
        RECT 49.180 299.150 51.480 299.200 ;
        RECT 57.980 299.150 60.280 299.200 ;
        RECT 46.530 298.000 62.930 298.600 ;
        RECT 50.130 297.400 50.480 298.000 ;
        RECT 46.530 297.200 50.480 297.400 ;
        RECT 50.130 296.600 50.480 297.200 ;
        RECT 46.530 296.400 50.480 296.600 ;
        RECT 50.130 295.800 50.480 296.400 ;
        RECT 46.530 295.600 50.480 295.800 ;
        RECT 38.980 294.800 42.930 295.000 ;
        RECT 38.980 294.200 39.330 294.800 ;
        RECT 38.980 294.000 42.930 294.200 ;
        RECT 38.980 293.400 39.330 294.000 ;
        RECT 38.980 293.200 42.930 293.400 ;
        RECT 43.880 293.250 45.580 295.550 ;
        RECT 50.130 295.000 50.480 295.600 ;
        RECT 46.530 294.800 50.480 295.000 ;
        RECT 50.130 294.200 50.480 294.800 ;
        RECT 46.530 294.000 50.480 294.200 ;
        RECT 50.130 293.400 50.480 294.000 ;
        RECT 38.980 292.600 39.330 293.200 ;
        RECT 38.980 292.400 42.930 292.600 ;
        RECT 38.980 291.800 39.330 292.400 ;
        RECT 38.980 291.600 42.930 291.800 ;
        RECT 38.980 291.000 39.330 291.600 ;
        RECT 38.980 290.800 42.930 291.000 ;
        RECT 38.980 290.400 39.330 290.800 ;
        RECT 35.780 282.000 35.980 289.600 ;
        RECT 36.580 282.000 36.780 289.600 ;
        RECT 37.380 282.000 37.580 289.600 ;
        RECT 38.180 282.000 38.380 289.600 ;
        RECT 38.980 289.200 39.330 289.600 ;
        RECT 38.980 289.000 42.930 289.200 ;
        RECT 38.980 288.400 39.330 289.000 ;
        RECT 38.980 288.200 42.930 288.400 ;
        RECT 38.980 287.600 39.330 288.200 ;
        RECT 38.980 287.400 42.930 287.600 ;
        RECT 38.980 286.800 39.330 287.400 ;
        RECT 38.980 286.600 42.930 286.800 ;
        RECT 43.930 286.750 44.330 293.250 ;
        RECT 45.130 286.750 45.530 293.250 ;
        RECT 46.530 293.200 50.480 293.400 ;
        RECT 50.130 292.600 50.480 293.200 ;
        RECT 46.530 292.400 50.480 292.600 ;
        RECT 50.130 291.800 50.480 292.400 ;
        RECT 46.530 291.600 50.480 291.800 ;
        RECT 50.130 291.000 50.480 291.600 ;
        RECT 46.530 290.800 50.480 291.000 ;
        RECT 50.130 290.400 50.480 290.800 ;
        RECT 51.080 290.400 51.280 298.000 ;
        RECT 51.880 290.400 52.080 298.000 ;
        RECT 52.680 290.400 52.880 298.000 ;
        RECT 53.480 290.400 53.680 298.000 ;
        RECT 50.130 289.200 50.480 289.600 ;
        RECT 46.530 289.000 50.480 289.200 ;
        RECT 50.130 288.400 50.480 289.000 ;
        RECT 46.530 288.200 50.480 288.400 ;
        RECT 50.130 287.600 50.480 288.200 ;
        RECT 46.530 287.400 50.480 287.600 ;
        RECT 50.130 286.800 50.480 287.400 ;
        RECT 38.980 286.000 39.330 286.600 ;
        RECT 38.980 285.800 42.930 286.000 ;
        RECT 38.980 285.200 39.330 285.800 ;
        RECT 38.980 285.000 42.930 285.200 ;
        RECT 38.980 284.400 39.330 285.000 ;
        RECT 43.880 284.450 45.580 286.750 ;
        RECT 46.530 286.600 50.480 286.800 ;
        RECT 50.130 286.000 50.480 286.600 ;
        RECT 46.530 285.800 50.480 286.000 ;
        RECT 50.130 285.200 50.480 285.800 ;
        RECT 46.530 285.000 50.480 285.200 ;
        RECT 38.980 284.200 42.930 284.400 ;
        RECT 38.980 283.600 39.330 284.200 ;
        RECT 38.980 283.400 42.930 283.600 ;
        RECT 38.980 282.800 39.330 283.400 ;
        RECT 38.980 282.600 42.930 282.800 ;
        RECT 38.980 282.000 39.330 282.600 ;
        RECT 26.530 281.400 42.930 282.000 ;
        RECT 29.180 280.800 31.480 280.850 ;
        RECT 37.980 280.800 40.280 280.850 ;
        RECT 43.930 280.800 44.330 284.450 ;
        RECT 25.130 280.400 44.330 280.800 ;
        RECT 45.130 280.800 45.530 284.450 ;
        RECT 50.130 284.400 50.480 285.000 ;
        RECT 46.530 284.200 50.480 284.400 ;
        RECT 50.130 283.600 50.480 284.200 ;
        RECT 46.530 283.400 50.480 283.600 ;
        RECT 50.130 282.800 50.480 283.400 ;
        RECT 46.530 282.600 50.480 282.800 ;
        RECT 50.130 282.000 50.480 282.600 ;
        RECT 51.080 282.000 51.280 289.600 ;
        RECT 51.880 282.000 52.080 289.600 ;
        RECT 52.680 282.000 52.880 289.600 ;
        RECT 53.480 282.000 53.680 289.600 ;
        RECT 54.280 282.000 55.180 298.000 ;
        RECT 55.780 290.400 55.980 298.000 ;
        RECT 56.580 290.400 56.780 298.000 ;
        RECT 57.380 290.400 57.580 298.000 ;
        RECT 58.180 290.400 58.380 298.000 ;
        RECT 58.980 297.400 59.330 298.000 ;
        RECT 58.980 297.200 62.930 297.400 ;
        RECT 58.980 296.600 59.330 297.200 ;
        RECT 58.980 296.400 62.930 296.600 ;
        RECT 58.980 295.800 59.330 296.400 ;
        RECT 58.980 295.600 62.930 295.800 ;
        RECT 58.980 295.000 59.330 295.600 ;
        RECT 63.930 295.550 64.330 299.200 ;
        RECT 65.130 299.200 84.330 299.600 ;
        RECT 65.130 295.550 65.530 299.200 ;
        RECT 69.180 299.150 71.480 299.200 ;
        RECT 77.980 299.150 80.280 299.200 ;
        RECT 66.530 298.000 82.930 298.600 ;
        RECT 70.130 297.400 70.480 298.000 ;
        RECT 66.530 297.200 70.480 297.400 ;
        RECT 70.130 296.600 70.480 297.200 ;
        RECT 66.530 296.400 70.480 296.600 ;
        RECT 70.130 295.800 70.480 296.400 ;
        RECT 66.530 295.600 70.480 295.800 ;
        RECT 58.980 294.800 62.930 295.000 ;
        RECT 58.980 294.200 59.330 294.800 ;
        RECT 58.980 294.000 62.930 294.200 ;
        RECT 58.980 293.400 59.330 294.000 ;
        RECT 58.980 293.200 62.930 293.400 ;
        RECT 63.880 293.250 65.580 295.550 ;
        RECT 70.130 295.000 70.480 295.600 ;
        RECT 66.530 294.800 70.480 295.000 ;
        RECT 70.130 294.200 70.480 294.800 ;
        RECT 66.530 294.000 70.480 294.200 ;
        RECT 70.130 293.400 70.480 294.000 ;
        RECT 58.980 292.600 59.330 293.200 ;
        RECT 58.980 292.400 62.930 292.600 ;
        RECT 58.980 291.800 59.330 292.400 ;
        RECT 58.980 291.600 62.930 291.800 ;
        RECT 58.980 291.000 59.330 291.600 ;
        RECT 58.980 290.800 62.930 291.000 ;
        RECT 58.980 290.400 59.330 290.800 ;
        RECT 55.780 282.000 55.980 289.600 ;
        RECT 56.580 282.000 56.780 289.600 ;
        RECT 57.380 282.000 57.580 289.600 ;
        RECT 58.180 282.000 58.380 289.600 ;
        RECT 58.980 289.200 59.330 289.600 ;
        RECT 58.980 289.000 62.930 289.200 ;
        RECT 58.980 288.400 59.330 289.000 ;
        RECT 58.980 288.200 62.930 288.400 ;
        RECT 58.980 287.600 59.330 288.200 ;
        RECT 58.980 287.400 62.930 287.600 ;
        RECT 58.980 286.800 59.330 287.400 ;
        RECT 58.980 286.600 62.930 286.800 ;
        RECT 63.930 286.750 64.330 293.250 ;
        RECT 65.130 286.750 65.530 293.250 ;
        RECT 66.530 293.200 70.480 293.400 ;
        RECT 70.130 292.600 70.480 293.200 ;
        RECT 66.530 292.400 70.480 292.600 ;
        RECT 70.130 291.800 70.480 292.400 ;
        RECT 66.530 291.600 70.480 291.800 ;
        RECT 70.130 291.000 70.480 291.600 ;
        RECT 66.530 290.800 70.480 291.000 ;
        RECT 70.130 290.400 70.480 290.800 ;
        RECT 71.080 290.400 71.280 298.000 ;
        RECT 71.880 290.400 72.080 298.000 ;
        RECT 72.680 290.400 72.880 298.000 ;
        RECT 73.480 290.400 73.680 298.000 ;
        RECT 70.130 289.200 70.480 289.600 ;
        RECT 66.530 289.000 70.480 289.200 ;
        RECT 70.130 288.400 70.480 289.000 ;
        RECT 66.530 288.200 70.480 288.400 ;
        RECT 70.130 287.600 70.480 288.200 ;
        RECT 66.530 287.400 70.480 287.600 ;
        RECT 70.130 286.800 70.480 287.400 ;
        RECT 58.980 286.000 59.330 286.600 ;
        RECT 58.980 285.800 62.930 286.000 ;
        RECT 58.980 285.200 59.330 285.800 ;
        RECT 58.980 285.000 62.930 285.200 ;
        RECT 58.980 284.400 59.330 285.000 ;
        RECT 63.880 284.450 65.580 286.750 ;
        RECT 66.530 286.600 70.480 286.800 ;
        RECT 70.130 286.000 70.480 286.600 ;
        RECT 66.530 285.800 70.480 286.000 ;
        RECT 70.130 285.200 70.480 285.800 ;
        RECT 66.530 285.000 70.480 285.200 ;
        RECT 58.980 284.200 62.930 284.400 ;
        RECT 58.980 283.600 59.330 284.200 ;
        RECT 58.980 283.400 62.930 283.600 ;
        RECT 58.980 282.800 59.330 283.400 ;
        RECT 58.980 282.600 62.930 282.800 ;
        RECT 58.980 282.000 59.330 282.600 ;
        RECT 46.530 281.400 62.930 282.000 ;
        RECT 49.180 280.800 51.480 280.850 ;
        RECT 57.980 280.800 60.280 280.850 ;
        RECT 63.930 280.800 64.330 284.450 ;
        RECT 45.130 280.400 64.330 280.800 ;
        RECT 65.130 280.800 65.530 284.450 ;
        RECT 70.130 284.400 70.480 285.000 ;
        RECT 66.530 284.200 70.480 284.400 ;
        RECT 70.130 283.600 70.480 284.200 ;
        RECT 66.530 283.400 70.480 283.600 ;
        RECT 70.130 282.800 70.480 283.400 ;
        RECT 66.530 282.600 70.480 282.800 ;
        RECT 70.130 282.000 70.480 282.600 ;
        RECT 71.080 282.000 71.280 289.600 ;
        RECT 71.880 282.000 72.080 289.600 ;
        RECT 72.680 282.000 72.880 289.600 ;
        RECT 73.480 282.000 73.680 289.600 ;
        RECT 74.280 282.000 75.180 298.000 ;
        RECT 75.780 290.400 75.980 298.000 ;
        RECT 76.580 290.400 76.780 298.000 ;
        RECT 77.380 290.400 77.580 298.000 ;
        RECT 78.180 290.400 78.380 298.000 ;
        RECT 78.980 297.400 79.330 298.000 ;
        RECT 78.980 297.200 82.930 297.400 ;
        RECT 78.980 296.600 79.330 297.200 ;
        RECT 78.980 296.400 82.930 296.600 ;
        RECT 78.980 295.800 79.330 296.400 ;
        RECT 78.980 295.600 82.930 295.800 ;
        RECT 78.980 295.000 79.330 295.600 ;
        RECT 83.930 295.550 84.330 299.200 ;
        RECT 85.130 299.200 104.330 299.600 ;
        RECT 85.130 295.550 85.530 299.200 ;
        RECT 89.180 299.150 91.480 299.200 ;
        RECT 97.980 299.150 100.280 299.200 ;
        RECT 86.530 298.000 102.930 298.600 ;
        RECT 90.130 297.400 90.480 298.000 ;
        RECT 86.530 297.200 90.480 297.400 ;
        RECT 90.130 296.600 90.480 297.200 ;
        RECT 86.530 296.400 90.480 296.600 ;
        RECT 90.130 295.800 90.480 296.400 ;
        RECT 86.530 295.600 90.480 295.800 ;
        RECT 78.980 294.800 82.930 295.000 ;
        RECT 78.980 294.200 79.330 294.800 ;
        RECT 78.980 294.000 82.930 294.200 ;
        RECT 78.980 293.400 79.330 294.000 ;
        RECT 78.980 293.200 82.930 293.400 ;
        RECT 83.880 293.250 85.580 295.550 ;
        RECT 90.130 295.000 90.480 295.600 ;
        RECT 86.530 294.800 90.480 295.000 ;
        RECT 90.130 294.200 90.480 294.800 ;
        RECT 86.530 294.000 90.480 294.200 ;
        RECT 90.130 293.400 90.480 294.000 ;
        RECT 78.980 292.600 79.330 293.200 ;
        RECT 78.980 292.400 82.930 292.600 ;
        RECT 78.980 291.800 79.330 292.400 ;
        RECT 78.980 291.600 82.930 291.800 ;
        RECT 78.980 291.000 79.330 291.600 ;
        RECT 78.980 290.800 82.930 291.000 ;
        RECT 78.980 290.400 79.330 290.800 ;
        RECT 75.780 282.000 75.980 289.600 ;
        RECT 76.580 282.000 76.780 289.600 ;
        RECT 77.380 282.000 77.580 289.600 ;
        RECT 78.180 282.000 78.380 289.600 ;
        RECT 78.980 289.200 79.330 289.600 ;
        RECT 78.980 289.000 82.930 289.200 ;
        RECT 78.980 288.400 79.330 289.000 ;
        RECT 78.980 288.200 82.930 288.400 ;
        RECT 78.980 287.600 79.330 288.200 ;
        RECT 78.980 287.400 82.930 287.600 ;
        RECT 78.980 286.800 79.330 287.400 ;
        RECT 78.980 286.600 82.930 286.800 ;
        RECT 83.930 286.750 84.330 293.250 ;
        RECT 85.130 286.750 85.530 293.250 ;
        RECT 86.530 293.200 90.480 293.400 ;
        RECT 90.130 292.600 90.480 293.200 ;
        RECT 86.530 292.400 90.480 292.600 ;
        RECT 90.130 291.800 90.480 292.400 ;
        RECT 86.530 291.600 90.480 291.800 ;
        RECT 90.130 291.000 90.480 291.600 ;
        RECT 86.530 290.800 90.480 291.000 ;
        RECT 90.130 290.400 90.480 290.800 ;
        RECT 91.080 290.400 91.280 298.000 ;
        RECT 91.880 290.400 92.080 298.000 ;
        RECT 92.680 290.400 92.880 298.000 ;
        RECT 93.480 290.400 93.680 298.000 ;
        RECT 90.130 289.200 90.480 289.600 ;
        RECT 86.530 289.000 90.480 289.200 ;
        RECT 90.130 288.400 90.480 289.000 ;
        RECT 86.530 288.200 90.480 288.400 ;
        RECT 90.130 287.600 90.480 288.200 ;
        RECT 86.530 287.400 90.480 287.600 ;
        RECT 90.130 286.800 90.480 287.400 ;
        RECT 78.980 286.000 79.330 286.600 ;
        RECT 78.980 285.800 82.930 286.000 ;
        RECT 78.980 285.200 79.330 285.800 ;
        RECT 78.980 285.000 82.930 285.200 ;
        RECT 78.980 284.400 79.330 285.000 ;
        RECT 83.880 284.450 85.580 286.750 ;
        RECT 86.530 286.600 90.480 286.800 ;
        RECT 90.130 286.000 90.480 286.600 ;
        RECT 86.530 285.800 90.480 286.000 ;
        RECT 90.130 285.200 90.480 285.800 ;
        RECT 86.530 285.000 90.480 285.200 ;
        RECT 78.980 284.200 82.930 284.400 ;
        RECT 78.980 283.600 79.330 284.200 ;
        RECT 78.980 283.400 82.930 283.600 ;
        RECT 78.980 282.800 79.330 283.400 ;
        RECT 78.980 282.600 82.930 282.800 ;
        RECT 78.980 282.000 79.330 282.600 ;
        RECT 66.530 281.400 82.930 282.000 ;
        RECT 69.180 280.800 71.480 280.850 ;
        RECT 77.980 280.800 80.280 280.850 ;
        RECT 83.930 280.800 84.330 284.450 ;
        RECT 65.130 280.400 84.330 280.800 ;
        RECT 85.130 280.800 85.530 284.450 ;
        RECT 90.130 284.400 90.480 285.000 ;
        RECT 86.530 284.200 90.480 284.400 ;
        RECT 90.130 283.600 90.480 284.200 ;
        RECT 86.530 283.400 90.480 283.600 ;
        RECT 90.130 282.800 90.480 283.400 ;
        RECT 86.530 282.600 90.480 282.800 ;
        RECT 90.130 282.000 90.480 282.600 ;
        RECT 91.080 282.000 91.280 289.600 ;
        RECT 91.880 282.000 92.080 289.600 ;
        RECT 92.680 282.000 92.880 289.600 ;
        RECT 93.480 282.000 93.680 289.600 ;
        RECT 94.280 282.000 95.180 298.000 ;
        RECT 95.780 290.400 95.980 298.000 ;
        RECT 96.580 290.400 96.780 298.000 ;
        RECT 97.380 290.400 97.580 298.000 ;
        RECT 98.180 290.400 98.380 298.000 ;
        RECT 98.980 297.400 99.330 298.000 ;
        RECT 98.980 297.200 102.930 297.400 ;
        RECT 98.980 296.600 99.330 297.200 ;
        RECT 98.980 296.400 102.930 296.600 ;
        RECT 98.980 295.800 99.330 296.400 ;
        RECT 98.980 295.600 102.930 295.800 ;
        RECT 98.980 295.000 99.330 295.600 ;
        RECT 103.930 295.550 104.330 299.200 ;
        RECT 105.130 299.200 124.330 299.600 ;
        RECT 105.130 295.550 105.530 299.200 ;
        RECT 109.180 299.150 111.480 299.200 ;
        RECT 117.980 299.150 120.280 299.200 ;
        RECT 106.530 298.000 122.930 298.600 ;
        RECT 110.130 297.400 110.480 298.000 ;
        RECT 106.530 297.200 110.480 297.400 ;
        RECT 110.130 296.600 110.480 297.200 ;
        RECT 106.530 296.400 110.480 296.600 ;
        RECT 110.130 295.800 110.480 296.400 ;
        RECT 106.530 295.600 110.480 295.800 ;
        RECT 98.980 294.800 102.930 295.000 ;
        RECT 98.980 294.200 99.330 294.800 ;
        RECT 98.980 294.000 102.930 294.200 ;
        RECT 98.980 293.400 99.330 294.000 ;
        RECT 98.980 293.200 102.930 293.400 ;
        RECT 103.880 293.250 105.580 295.550 ;
        RECT 110.130 295.000 110.480 295.600 ;
        RECT 106.530 294.800 110.480 295.000 ;
        RECT 110.130 294.200 110.480 294.800 ;
        RECT 106.530 294.000 110.480 294.200 ;
        RECT 110.130 293.400 110.480 294.000 ;
        RECT 98.980 292.600 99.330 293.200 ;
        RECT 98.980 292.400 102.930 292.600 ;
        RECT 98.980 291.800 99.330 292.400 ;
        RECT 98.980 291.600 102.930 291.800 ;
        RECT 98.980 291.000 99.330 291.600 ;
        RECT 98.980 290.800 102.930 291.000 ;
        RECT 98.980 290.400 99.330 290.800 ;
        RECT 95.780 282.000 95.980 289.600 ;
        RECT 96.580 282.000 96.780 289.600 ;
        RECT 97.380 282.000 97.580 289.600 ;
        RECT 98.180 282.000 98.380 289.600 ;
        RECT 98.980 289.200 99.330 289.600 ;
        RECT 98.980 289.000 102.930 289.200 ;
        RECT 98.980 288.400 99.330 289.000 ;
        RECT 98.980 288.200 102.930 288.400 ;
        RECT 98.980 287.600 99.330 288.200 ;
        RECT 98.980 287.400 102.930 287.600 ;
        RECT 98.980 286.800 99.330 287.400 ;
        RECT 98.980 286.600 102.930 286.800 ;
        RECT 103.930 286.750 104.330 293.250 ;
        RECT 105.130 286.750 105.530 293.250 ;
        RECT 106.530 293.200 110.480 293.400 ;
        RECT 110.130 292.600 110.480 293.200 ;
        RECT 106.530 292.400 110.480 292.600 ;
        RECT 110.130 291.800 110.480 292.400 ;
        RECT 106.530 291.600 110.480 291.800 ;
        RECT 110.130 291.000 110.480 291.600 ;
        RECT 106.530 290.800 110.480 291.000 ;
        RECT 110.130 290.400 110.480 290.800 ;
        RECT 111.080 290.400 111.280 298.000 ;
        RECT 111.880 290.400 112.080 298.000 ;
        RECT 112.680 290.400 112.880 298.000 ;
        RECT 113.480 290.400 113.680 298.000 ;
        RECT 110.130 289.200 110.480 289.600 ;
        RECT 106.530 289.000 110.480 289.200 ;
        RECT 110.130 288.400 110.480 289.000 ;
        RECT 106.530 288.200 110.480 288.400 ;
        RECT 110.130 287.600 110.480 288.200 ;
        RECT 106.530 287.400 110.480 287.600 ;
        RECT 110.130 286.800 110.480 287.400 ;
        RECT 98.980 286.000 99.330 286.600 ;
        RECT 98.980 285.800 102.930 286.000 ;
        RECT 98.980 285.200 99.330 285.800 ;
        RECT 98.980 285.000 102.930 285.200 ;
        RECT 98.980 284.400 99.330 285.000 ;
        RECT 103.880 284.450 105.580 286.750 ;
        RECT 106.530 286.600 110.480 286.800 ;
        RECT 110.130 286.000 110.480 286.600 ;
        RECT 106.530 285.800 110.480 286.000 ;
        RECT 110.130 285.200 110.480 285.800 ;
        RECT 106.530 285.000 110.480 285.200 ;
        RECT 98.980 284.200 102.930 284.400 ;
        RECT 98.980 283.600 99.330 284.200 ;
        RECT 98.980 283.400 102.930 283.600 ;
        RECT 98.980 282.800 99.330 283.400 ;
        RECT 98.980 282.600 102.930 282.800 ;
        RECT 98.980 282.000 99.330 282.600 ;
        RECT 86.530 281.400 102.930 282.000 ;
        RECT 89.180 280.800 91.480 280.850 ;
        RECT 97.980 280.800 100.280 280.850 ;
        RECT 103.930 280.800 104.330 284.450 ;
        RECT 85.130 280.400 104.330 280.800 ;
        RECT 105.130 280.800 105.530 284.450 ;
        RECT 110.130 284.400 110.480 285.000 ;
        RECT 106.530 284.200 110.480 284.400 ;
        RECT 110.130 283.600 110.480 284.200 ;
        RECT 106.530 283.400 110.480 283.600 ;
        RECT 110.130 282.800 110.480 283.400 ;
        RECT 106.530 282.600 110.480 282.800 ;
        RECT 110.130 282.000 110.480 282.600 ;
        RECT 111.080 282.000 111.280 289.600 ;
        RECT 111.880 282.000 112.080 289.600 ;
        RECT 112.680 282.000 112.880 289.600 ;
        RECT 113.480 282.000 113.680 289.600 ;
        RECT 114.280 282.000 115.180 298.000 ;
        RECT 115.780 290.400 115.980 298.000 ;
        RECT 116.580 290.400 116.780 298.000 ;
        RECT 117.380 290.400 117.580 298.000 ;
        RECT 118.180 290.400 118.380 298.000 ;
        RECT 118.980 297.400 119.330 298.000 ;
        RECT 118.980 297.200 122.930 297.400 ;
        RECT 118.980 296.600 119.330 297.200 ;
        RECT 118.980 296.400 122.930 296.600 ;
        RECT 118.980 295.800 119.330 296.400 ;
        RECT 118.980 295.600 122.930 295.800 ;
        RECT 118.980 295.000 119.330 295.600 ;
        RECT 123.930 295.550 124.330 299.200 ;
        RECT 125.340 297.080 125.700 297.460 ;
        RECT 125.970 297.080 126.330 297.460 ;
        RECT 126.570 297.080 126.930 297.460 ;
        RECT 125.340 296.490 125.700 296.870 ;
        RECT 125.970 296.490 126.330 296.870 ;
        RECT 126.570 296.490 126.930 296.870 ;
        RECT 118.980 294.800 122.930 295.000 ;
        RECT 118.980 294.200 119.330 294.800 ;
        RECT 118.980 294.000 122.930 294.200 ;
        RECT 118.980 293.400 119.330 294.000 ;
        RECT 118.980 293.200 122.930 293.400 ;
        RECT 123.880 293.250 124.730 295.550 ;
        RECT 118.980 292.600 119.330 293.200 ;
        RECT 118.980 292.400 122.930 292.600 ;
        RECT 118.980 291.800 119.330 292.400 ;
        RECT 118.980 291.600 122.930 291.800 ;
        RECT 118.980 291.000 119.330 291.600 ;
        RECT 118.980 290.800 122.930 291.000 ;
        RECT 118.980 290.400 119.330 290.800 ;
        RECT 115.780 282.000 115.980 289.600 ;
        RECT 116.580 282.000 116.780 289.600 ;
        RECT 117.380 282.000 117.580 289.600 ;
        RECT 118.180 282.000 118.380 289.600 ;
        RECT 118.980 289.200 119.330 289.600 ;
        RECT 118.980 289.000 122.930 289.200 ;
        RECT 118.980 288.400 119.330 289.000 ;
        RECT 118.980 288.200 122.930 288.400 ;
        RECT 118.980 287.600 119.330 288.200 ;
        RECT 118.980 287.400 122.930 287.600 ;
        RECT 118.980 286.800 119.330 287.400 ;
        RECT 118.980 286.600 122.930 286.800 ;
        RECT 123.930 286.750 124.330 293.250 ;
        RECT 118.980 286.000 119.330 286.600 ;
        RECT 118.980 285.800 122.930 286.000 ;
        RECT 118.980 285.200 119.330 285.800 ;
        RECT 118.980 285.000 122.930 285.200 ;
        RECT 118.980 284.400 119.330 285.000 ;
        RECT 123.880 284.450 124.730 286.750 ;
        RECT 118.980 284.200 122.930 284.400 ;
        RECT 118.980 283.600 119.330 284.200 ;
        RECT 118.980 283.400 122.930 283.600 ;
        RECT 118.980 282.800 119.330 283.400 ;
        RECT 118.980 282.600 122.930 282.800 ;
        RECT 118.980 282.000 119.330 282.600 ;
        RECT 106.530 281.400 122.930 282.000 ;
        RECT 109.180 280.800 111.480 280.850 ;
        RECT 117.980 280.800 120.280 280.850 ;
        RECT 123.930 280.800 124.330 284.450 ;
        RECT 125.340 283.095 125.700 283.475 ;
        RECT 125.970 283.095 126.330 283.475 ;
        RECT 126.570 283.095 126.930 283.475 ;
        RECT 125.340 282.505 125.700 282.885 ;
        RECT 125.970 282.505 126.330 282.885 ;
        RECT 126.570 282.505 126.930 282.885 ;
        RECT 105.130 280.400 124.330 280.800 ;
        RECT 9.180 279.600 11.480 280.400 ;
        RECT 17.980 279.600 20.280 280.400 ;
        RECT 29.180 279.600 31.480 280.400 ;
        RECT 37.980 279.600 40.280 280.400 ;
        RECT 49.180 279.600 51.480 280.400 ;
        RECT 57.980 279.600 60.280 280.400 ;
        RECT 69.180 279.600 71.480 280.400 ;
        RECT 77.980 279.600 80.280 280.400 ;
        RECT 89.180 279.600 91.480 280.400 ;
        RECT 97.980 279.600 100.280 280.400 ;
        RECT 109.180 279.600 111.480 280.400 ;
        RECT 117.980 279.600 120.280 280.400 ;
        RECT 5.130 279.200 24.330 279.600 ;
        RECT 2.515 277.025 2.875 277.405 ;
        RECT 3.145 277.025 3.505 277.405 ;
        RECT 3.745 277.025 4.105 277.405 ;
        RECT 2.515 276.435 2.875 276.815 ;
        RECT 3.145 276.435 3.505 276.815 ;
        RECT 3.745 276.435 4.105 276.815 ;
        RECT 5.130 275.550 5.530 279.200 ;
        RECT 9.180 279.150 11.480 279.200 ;
        RECT 17.980 279.150 20.280 279.200 ;
        RECT 6.530 278.000 22.930 278.600 ;
        RECT 10.130 277.400 10.480 278.000 ;
        RECT 6.530 277.200 10.480 277.400 ;
        RECT 10.130 276.600 10.480 277.200 ;
        RECT 6.530 276.400 10.480 276.600 ;
        RECT 10.130 275.800 10.480 276.400 ;
        RECT 6.530 275.600 10.480 275.800 ;
        RECT 4.730 275.545 5.580 275.550 ;
        RECT 2.320 275.340 5.580 275.545 ;
        RECT 2.315 273.250 5.580 275.340 ;
        RECT 10.130 275.000 10.480 275.600 ;
        RECT 6.530 274.800 10.480 275.000 ;
        RECT 10.130 274.200 10.480 274.800 ;
        RECT 6.530 274.000 10.480 274.200 ;
        RECT 10.130 273.400 10.480 274.000 ;
        RECT 5.130 266.750 5.530 273.250 ;
        RECT 6.530 273.200 10.480 273.400 ;
        RECT 10.130 272.600 10.480 273.200 ;
        RECT 6.530 272.400 10.480 272.600 ;
        RECT 10.130 271.800 10.480 272.400 ;
        RECT 6.530 271.600 10.480 271.800 ;
        RECT 10.130 271.000 10.480 271.600 ;
        RECT 6.530 270.800 10.480 271.000 ;
        RECT 10.130 270.400 10.480 270.800 ;
        RECT 11.080 270.400 11.280 278.000 ;
        RECT 11.880 270.400 12.080 278.000 ;
        RECT 12.680 270.400 12.880 278.000 ;
        RECT 13.480 270.400 13.680 278.000 ;
        RECT 10.130 269.200 10.480 269.600 ;
        RECT 6.530 269.000 10.480 269.200 ;
        RECT 10.130 268.400 10.480 269.000 ;
        RECT 6.530 268.200 10.480 268.400 ;
        RECT 10.130 267.600 10.480 268.200 ;
        RECT 6.530 267.400 10.480 267.600 ;
        RECT 10.130 266.800 10.480 267.400 ;
        RECT 4.730 266.740 5.580 266.750 ;
        RECT 2.315 264.450 5.580 266.740 ;
        RECT 6.530 266.600 10.480 266.800 ;
        RECT 10.130 266.000 10.480 266.600 ;
        RECT 6.530 265.800 10.480 266.000 ;
        RECT 10.130 265.200 10.480 265.800 ;
        RECT 6.530 265.000 10.480 265.200 ;
        RECT 2.315 264.445 4.730 264.450 ;
        RECT 2.515 263.140 2.875 263.520 ;
        RECT 3.145 263.140 3.505 263.520 ;
        RECT 3.745 263.140 4.105 263.520 ;
        RECT 2.515 262.550 2.875 262.930 ;
        RECT 3.145 262.550 3.505 262.930 ;
        RECT 3.745 262.550 4.105 262.930 ;
        RECT 5.130 260.800 5.530 264.450 ;
        RECT 10.130 264.400 10.480 265.000 ;
        RECT 6.530 264.200 10.480 264.400 ;
        RECT 10.130 263.600 10.480 264.200 ;
        RECT 6.530 263.400 10.480 263.600 ;
        RECT 10.130 262.800 10.480 263.400 ;
        RECT 6.530 262.600 10.480 262.800 ;
        RECT 10.130 262.000 10.480 262.600 ;
        RECT 11.080 262.000 11.280 269.600 ;
        RECT 11.880 262.000 12.080 269.600 ;
        RECT 12.680 262.000 12.880 269.600 ;
        RECT 13.480 262.000 13.680 269.600 ;
        RECT 14.280 262.000 15.180 278.000 ;
        RECT 15.780 270.400 15.980 278.000 ;
        RECT 16.580 270.400 16.780 278.000 ;
        RECT 17.380 270.400 17.580 278.000 ;
        RECT 18.180 270.400 18.380 278.000 ;
        RECT 18.980 277.400 19.330 278.000 ;
        RECT 18.980 277.200 22.930 277.400 ;
        RECT 18.980 276.600 19.330 277.200 ;
        RECT 18.980 276.400 22.930 276.600 ;
        RECT 18.980 275.800 19.330 276.400 ;
        RECT 18.980 275.600 22.930 275.800 ;
        RECT 18.980 275.000 19.330 275.600 ;
        RECT 23.930 275.550 24.330 279.200 ;
        RECT 25.130 279.200 44.330 279.600 ;
        RECT 25.130 275.550 25.530 279.200 ;
        RECT 29.180 279.150 31.480 279.200 ;
        RECT 37.980 279.150 40.280 279.200 ;
        RECT 26.530 278.000 42.930 278.600 ;
        RECT 30.130 277.400 30.480 278.000 ;
        RECT 26.530 277.200 30.480 277.400 ;
        RECT 30.130 276.600 30.480 277.200 ;
        RECT 26.530 276.400 30.480 276.600 ;
        RECT 30.130 275.800 30.480 276.400 ;
        RECT 26.530 275.600 30.480 275.800 ;
        RECT 18.980 274.800 22.930 275.000 ;
        RECT 18.980 274.200 19.330 274.800 ;
        RECT 18.980 274.000 22.930 274.200 ;
        RECT 18.980 273.400 19.330 274.000 ;
        RECT 18.980 273.200 22.930 273.400 ;
        RECT 23.880 273.250 25.580 275.550 ;
        RECT 30.130 275.000 30.480 275.600 ;
        RECT 26.530 274.800 30.480 275.000 ;
        RECT 30.130 274.200 30.480 274.800 ;
        RECT 26.530 274.000 30.480 274.200 ;
        RECT 30.130 273.400 30.480 274.000 ;
        RECT 18.980 272.600 19.330 273.200 ;
        RECT 18.980 272.400 22.930 272.600 ;
        RECT 18.980 271.800 19.330 272.400 ;
        RECT 18.980 271.600 22.930 271.800 ;
        RECT 18.980 271.000 19.330 271.600 ;
        RECT 18.980 270.800 22.930 271.000 ;
        RECT 18.980 270.400 19.330 270.800 ;
        RECT 15.780 262.000 15.980 269.600 ;
        RECT 16.580 262.000 16.780 269.600 ;
        RECT 17.380 262.000 17.580 269.600 ;
        RECT 18.180 262.000 18.380 269.600 ;
        RECT 18.980 269.200 19.330 269.600 ;
        RECT 18.980 269.000 22.930 269.200 ;
        RECT 18.980 268.400 19.330 269.000 ;
        RECT 18.980 268.200 22.930 268.400 ;
        RECT 18.980 267.600 19.330 268.200 ;
        RECT 18.980 267.400 22.930 267.600 ;
        RECT 18.980 266.800 19.330 267.400 ;
        RECT 18.980 266.600 22.930 266.800 ;
        RECT 23.930 266.750 24.330 273.250 ;
        RECT 25.130 266.750 25.530 273.250 ;
        RECT 26.530 273.200 30.480 273.400 ;
        RECT 30.130 272.600 30.480 273.200 ;
        RECT 26.530 272.400 30.480 272.600 ;
        RECT 30.130 271.800 30.480 272.400 ;
        RECT 26.530 271.600 30.480 271.800 ;
        RECT 30.130 271.000 30.480 271.600 ;
        RECT 26.530 270.800 30.480 271.000 ;
        RECT 30.130 270.400 30.480 270.800 ;
        RECT 31.080 270.400 31.280 278.000 ;
        RECT 31.880 270.400 32.080 278.000 ;
        RECT 32.680 270.400 32.880 278.000 ;
        RECT 33.480 270.400 33.680 278.000 ;
        RECT 30.130 269.200 30.480 269.600 ;
        RECT 26.530 269.000 30.480 269.200 ;
        RECT 30.130 268.400 30.480 269.000 ;
        RECT 26.530 268.200 30.480 268.400 ;
        RECT 30.130 267.600 30.480 268.200 ;
        RECT 26.530 267.400 30.480 267.600 ;
        RECT 30.130 266.800 30.480 267.400 ;
        RECT 18.980 266.000 19.330 266.600 ;
        RECT 18.980 265.800 22.930 266.000 ;
        RECT 18.980 265.200 19.330 265.800 ;
        RECT 18.980 265.000 22.930 265.200 ;
        RECT 18.980 264.400 19.330 265.000 ;
        RECT 23.880 264.450 25.580 266.750 ;
        RECT 26.530 266.600 30.480 266.800 ;
        RECT 30.130 266.000 30.480 266.600 ;
        RECT 26.530 265.800 30.480 266.000 ;
        RECT 30.130 265.200 30.480 265.800 ;
        RECT 26.530 265.000 30.480 265.200 ;
        RECT 18.980 264.200 22.930 264.400 ;
        RECT 18.980 263.600 19.330 264.200 ;
        RECT 18.980 263.400 22.930 263.600 ;
        RECT 18.980 262.800 19.330 263.400 ;
        RECT 18.980 262.600 22.930 262.800 ;
        RECT 18.980 262.000 19.330 262.600 ;
        RECT 6.530 261.400 22.930 262.000 ;
        RECT 9.180 260.800 11.480 260.850 ;
        RECT 17.980 260.800 20.280 260.850 ;
        RECT 23.930 260.800 24.330 264.450 ;
        RECT 5.130 260.400 24.330 260.800 ;
        RECT 25.130 260.800 25.530 264.450 ;
        RECT 30.130 264.400 30.480 265.000 ;
        RECT 26.530 264.200 30.480 264.400 ;
        RECT 30.130 263.600 30.480 264.200 ;
        RECT 26.530 263.400 30.480 263.600 ;
        RECT 30.130 262.800 30.480 263.400 ;
        RECT 26.530 262.600 30.480 262.800 ;
        RECT 30.130 262.000 30.480 262.600 ;
        RECT 31.080 262.000 31.280 269.600 ;
        RECT 31.880 262.000 32.080 269.600 ;
        RECT 32.680 262.000 32.880 269.600 ;
        RECT 33.480 262.000 33.680 269.600 ;
        RECT 34.280 262.000 35.180 278.000 ;
        RECT 35.780 270.400 35.980 278.000 ;
        RECT 36.580 270.400 36.780 278.000 ;
        RECT 37.380 270.400 37.580 278.000 ;
        RECT 38.180 270.400 38.380 278.000 ;
        RECT 38.980 277.400 39.330 278.000 ;
        RECT 38.980 277.200 42.930 277.400 ;
        RECT 38.980 276.600 39.330 277.200 ;
        RECT 38.980 276.400 42.930 276.600 ;
        RECT 38.980 275.800 39.330 276.400 ;
        RECT 38.980 275.600 42.930 275.800 ;
        RECT 38.980 275.000 39.330 275.600 ;
        RECT 43.930 275.550 44.330 279.200 ;
        RECT 45.130 279.200 64.330 279.600 ;
        RECT 45.130 275.550 45.530 279.200 ;
        RECT 49.180 279.150 51.480 279.200 ;
        RECT 57.980 279.150 60.280 279.200 ;
        RECT 46.530 278.000 62.930 278.600 ;
        RECT 50.130 277.400 50.480 278.000 ;
        RECT 46.530 277.200 50.480 277.400 ;
        RECT 50.130 276.600 50.480 277.200 ;
        RECT 46.530 276.400 50.480 276.600 ;
        RECT 50.130 275.800 50.480 276.400 ;
        RECT 46.530 275.600 50.480 275.800 ;
        RECT 38.980 274.800 42.930 275.000 ;
        RECT 38.980 274.200 39.330 274.800 ;
        RECT 38.980 274.000 42.930 274.200 ;
        RECT 38.980 273.400 39.330 274.000 ;
        RECT 38.980 273.200 42.930 273.400 ;
        RECT 43.880 273.250 45.580 275.550 ;
        RECT 50.130 275.000 50.480 275.600 ;
        RECT 46.530 274.800 50.480 275.000 ;
        RECT 50.130 274.200 50.480 274.800 ;
        RECT 46.530 274.000 50.480 274.200 ;
        RECT 50.130 273.400 50.480 274.000 ;
        RECT 38.980 272.600 39.330 273.200 ;
        RECT 38.980 272.400 42.930 272.600 ;
        RECT 38.980 271.800 39.330 272.400 ;
        RECT 38.980 271.600 42.930 271.800 ;
        RECT 38.980 271.000 39.330 271.600 ;
        RECT 38.980 270.800 42.930 271.000 ;
        RECT 38.980 270.400 39.330 270.800 ;
        RECT 35.780 262.000 35.980 269.600 ;
        RECT 36.580 262.000 36.780 269.600 ;
        RECT 37.380 262.000 37.580 269.600 ;
        RECT 38.180 262.000 38.380 269.600 ;
        RECT 38.980 269.200 39.330 269.600 ;
        RECT 38.980 269.000 42.930 269.200 ;
        RECT 38.980 268.400 39.330 269.000 ;
        RECT 38.980 268.200 42.930 268.400 ;
        RECT 38.980 267.600 39.330 268.200 ;
        RECT 38.980 267.400 42.930 267.600 ;
        RECT 38.980 266.800 39.330 267.400 ;
        RECT 38.980 266.600 42.930 266.800 ;
        RECT 43.930 266.750 44.330 273.250 ;
        RECT 45.130 266.750 45.530 273.250 ;
        RECT 46.530 273.200 50.480 273.400 ;
        RECT 50.130 272.600 50.480 273.200 ;
        RECT 46.530 272.400 50.480 272.600 ;
        RECT 50.130 271.800 50.480 272.400 ;
        RECT 46.530 271.600 50.480 271.800 ;
        RECT 50.130 271.000 50.480 271.600 ;
        RECT 46.530 270.800 50.480 271.000 ;
        RECT 50.130 270.400 50.480 270.800 ;
        RECT 51.080 270.400 51.280 278.000 ;
        RECT 51.880 270.400 52.080 278.000 ;
        RECT 52.680 270.400 52.880 278.000 ;
        RECT 53.480 270.400 53.680 278.000 ;
        RECT 50.130 269.200 50.480 269.600 ;
        RECT 46.530 269.000 50.480 269.200 ;
        RECT 50.130 268.400 50.480 269.000 ;
        RECT 46.530 268.200 50.480 268.400 ;
        RECT 50.130 267.600 50.480 268.200 ;
        RECT 46.530 267.400 50.480 267.600 ;
        RECT 50.130 266.800 50.480 267.400 ;
        RECT 38.980 266.000 39.330 266.600 ;
        RECT 38.980 265.800 42.930 266.000 ;
        RECT 38.980 265.200 39.330 265.800 ;
        RECT 38.980 265.000 42.930 265.200 ;
        RECT 38.980 264.400 39.330 265.000 ;
        RECT 43.880 264.450 45.580 266.750 ;
        RECT 46.530 266.600 50.480 266.800 ;
        RECT 50.130 266.000 50.480 266.600 ;
        RECT 46.530 265.800 50.480 266.000 ;
        RECT 50.130 265.200 50.480 265.800 ;
        RECT 46.530 265.000 50.480 265.200 ;
        RECT 38.980 264.200 42.930 264.400 ;
        RECT 38.980 263.600 39.330 264.200 ;
        RECT 38.980 263.400 42.930 263.600 ;
        RECT 38.980 262.800 39.330 263.400 ;
        RECT 38.980 262.600 42.930 262.800 ;
        RECT 38.980 262.000 39.330 262.600 ;
        RECT 26.530 261.400 42.930 262.000 ;
        RECT 29.180 260.800 31.480 260.850 ;
        RECT 37.980 260.800 40.280 260.850 ;
        RECT 43.930 260.800 44.330 264.450 ;
        RECT 25.130 260.400 44.330 260.800 ;
        RECT 45.130 260.800 45.530 264.450 ;
        RECT 50.130 264.400 50.480 265.000 ;
        RECT 46.530 264.200 50.480 264.400 ;
        RECT 50.130 263.600 50.480 264.200 ;
        RECT 46.530 263.400 50.480 263.600 ;
        RECT 50.130 262.800 50.480 263.400 ;
        RECT 46.530 262.600 50.480 262.800 ;
        RECT 50.130 262.000 50.480 262.600 ;
        RECT 51.080 262.000 51.280 269.600 ;
        RECT 51.880 262.000 52.080 269.600 ;
        RECT 52.680 262.000 52.880 269.600 ;
        RECT 53.480 262.000 53.680 269.600 ;
        RECT 54.280 262.000 55.180 278.000 ;
        RECT 55.780 270.400 55.980 278.000 ;
        RECT 56.580 270.400 56.780 278.000 ;
        RECT 57.380 270.400 57.580 278.000 ;
        RECT 58.180 270.400 58.380 278.000 ;
        RECT 58.980 277.400 59.330 278.000 ;
        RECT 58.980 277.200 62.930 277.400 ;
        RECT 58.980 276.600 59.330 277.200 ;
        RECT 58.980 276.400 62.930 276.600 ;
        RECT 58.980 275.800 59.330 276.400 ;
        RECT 58.980 275.600 62.930 275.800 ;
        RECT 58.980 275.000 59.330 275.600 ;
        RECT 63.930 275.550 64.330 279.200 ;
        RECT 65.130 279.200 84.330 279.600 ;
        RECT 65.130 275.550 65.530 279.200 ;
        RECT 69.180 279.150 71.480 279.200 ;
        RECT 77.980 279.150 80.280 279.200 ;
        RECT 66.530 278.000 82.930 278.600 ;
        RECT 70.130 277.400 70.480 278.000 ;
        RECT 66.530 277.200 70.480 277.400 ;
        RECT 70.130 276.600 70.480 277.200 ;
        RECT 66.530 276.400 70.480 276.600 ;
        RECT 70.130 275.800 70.480 276.400 ;
        RECT 66.530 275.600 70.480 275.800 ;
        RECT 58.980 274.800 62.930 275.000 ;
        RECT 58.980 274.200 59.330 274.800 ;
        RECT 58.980 274.000 62.930 274.200 ;
        RECT 58.980 273.400 59.330 274.000 ;
        RECT 58.980 273.200 62.930 273.400 ;
        RECT 63.880 273.250 65.580 275.550 ;
        RECT 70.130 275.000 70.480 275.600 ;
        RECT 66.530 274.800 70.480 275.000 ;
        RECT 70.130 274.200 70.480 274.800 ;
        RECT 66.530 274.000 70.480 274.200 ;
        RECT 70.130 273.400 70.480 274.000 ;
        RECT 58.980 272.600 59.330 273.200 ;
        RECT 58.980 272.400 62.930 272.600 ;
        RECT 58.980 271.800 59.330 272.400 ;
        RECT 58.980 271.600 62.930 271.800 ;
        RECT 58.980 271.000 59.330 271.600 ;
        RECT 58.980 270.800 62.930 271.000 ;
        RECT 58.980 270.400 59.330 270.800 ;
        RECT 55.780 262.000 55.980 269.600 ;
        RECT 56.580 262.000 56.780 269.600 ;
        RECT 57.380 262.000 57.580 269.600 ;
        RECT 58.180 262.000 58.380 269.600 ;
        RECT 58.980 269.200 59.330 269.600 ;
        RECT 58.980 269.000 62.930 269.200 ;
        RECT 58.980 268.400 59.330 269.000 ;
        RECT 58.980 268.200 62.930 268.400 ;
        RECT 58.980 267.600 59.330 268.200 ;
        RECT 58.980 267.400 62.930 267.600 ;
        RECT 58.980 266.800 59.330 267.400 ;
        RECT 58.980 266.600 62.930 266.800 ;
        RECT 63.930 266.750 64.330 273.250 ;
        RECT 65.130 266.750 65.530 273.250 ;
        RECT 66.530 273.200 70.480 273.400 ;
        RECT 70.130 272.600 70.480 273.200 ;
        RECT 66.530 272.400 70.480 272.600 ;
        RECT 70.130 271.800 70.480 272.400 ;
        RECT 66.530 271.600 70.480 271.800 ;
        RECT 70.130 271.000 70.480 271.600 ;
        RECT 66.530 270.800 70.480 271.000 ;
        RECT 70.130 270.400 70.480 270.800 ;
        RECT 71.080 270.400 71.280 278.000 ;
        RECT 71.880 270.400 72.080 278.000 ;
        RECT 72.680 270.400 72.880 278.000 ;
        RECT 73.480 270.400 73.680 278.000 ;
        RECT 70.130 269.200 70.480 269.600 ;
        RECT 66.530 269.000 70.480 269.200 ;
        RECT 70.130 268.400 70.480 269.000 ;
        RECT 66.530 268.200 70.480 268.400 ;
        RECT 70.130 267.600 70.480 268.200 ;
        RECT 66.530 267.400 70.480 267.600 ;
        RECT 70.130 266.800 70.480 267.400 ;
        RECT 58.980 266.000 59.330 266.600 ;
        RECT 58.980 265.800 62.930 266.000 ;
        RECT 58.980 265.200 59.330 265.800 ;
        RECT 58.980 265.000 62.930 265.200 ;
        RECT 58.980 264.400 59.330 265.000 ;
        RECT 63.880 264.450 65.580 266.750 ;
        RECT 66.530 266.600 70.480 266.800 ;
        RECT 70.130 266.000 70.480 266.600 ;
        RECT 66.530 265.800 70.480 266.000 ;
        RECT 70.130 265.200 70.480 265.800 ;
        RECT 66.530 265.000 70.480 265.200 ;
        RECT 58.980 264.200 62.930 264.400 ;
        RECT 58.980 263.600 59.330 264.200 ;
        RECT 58.980 263.400 62.930 263.600 ;
        RECT 58.980 262.800 59.330 263.400 ;
        RECT 58.980 262.600 62.930 262.800 ;
        RECT 58.980 262.000 59.330 262.600 ;
        RECT 46.530 261.400 62.930 262.000 ;
        RECT 49.180 260.800 51.480 260.850 ;
        RECT 57.980 260.800 60.280 260.850 ;
        RECT 63.930 260.800 64.330 264.450 ;
        RECT 45.130 260.400 64.330 260.800 ;
        RECT 65.130 260.800 65.530 264.450 ;
        RECT 70.130 264.400 70.480 265.000 ;
        RECT 66.530 264.200 70.480 264.400 ;
        RECT 70.130 263.600 70.480 264.200 ;
        RECT 66.530 263.400 70.480 263.600 ;
        RECT 70.130 262.800 70.480 263.400 ;
        RECT 66.530 262.600 70.480 262.800 ;
        RECT 70.130 262.000 70.480 262.600 ;
        RECT 71.080 262.000 71.280 269.600 ;
        RECT 71.880 262.000 72.080 269.600 ;
        RECT 72.680 262.000 72.880 269.600 ;
        RECT 73.480 262.000 73.680 269.600 ;
        RECT 74.280 262.000 75.180 278.000 ;
        RECT 75.780 270.400 75.980 278.000 ;
        RECT 76.580 270.400 76.780 278.000 ;
        RECT 77.380 270.400 77.580 278.000 ;
        RECT 78.180 270.400 78.380 278.000 ;
        RECT 78.980 277.400 79.330 278.000 ;
        RECT 78.980 277.200 82.930 277.400 ;
        RECT 78.980 276.600 79.330 277.200 ;
        RECT 78.980 276.400 82.930 276.600 ;
        RECT 78.980 275.800 79.330 276.400 ;
        RECT 78.980 275.600 82.930 275.800 ;
        RECT 78.980 275.000 79.330 275.600 ;
        RECT 83.930 275.550 84.330 279.200 ;
        RECT 85.130 279.200 104.330 279.600 ;
        RECT 85.130 275.550 85.530 279.200 ;
        RECT 89.180 279.150 91.480 279.200 ;
        RECT 97.980 279.150 100.280 279.200 ;
        RECT 86.530 278.000 102.930 278.600 ;
        RECT 90.130 277.400 90.480 278.000 ;
        RECT 86.530 277.200 90.480 277.400 ;
        RECT 90.130 276.600 90.480 277.200 ;
        RECT 86.530 276.400 90.480 276.600 ;
        RECT 90.130 275.800 90.480 276.400 ;
        RECT 86.530 275.600 90.480 275.800 ;
        RECT 78.980 274.800 82.930 275.000 ;
        RECT 78.980 274.200 79.330 274.800 ;
        RECT 78.980 274.000 82.930 274.200 ;
        RECT 78.980 273.400 79.330 274.000 ;
        RECT 78.980 273.200 82.930 273.400 ;
        RECT 83.880 273.250 85.580 275.550 ;
        RECT 90.130 275.000 90.480 275.600 ;
        RECT 86.530 274.800 90.480 275.000 ;
        RECT 90.130 274.200 90.480 274.800 ;
        RECT 86.530 274.000 90.480 274.200 ;
        RECT 90.130 273.400 90.480 274.000 ;
        RECT 78.980 272.600 79.330 273.200 ;
        RECT 78.980 272.400 82.930 272.600 ;
        RECT 78.980 271.800 79.330 272.400 ;
        RECT 78.980 271.600 82.930 271.800 ;
        RECT 78.980 271.000 79.330 271.600 ;
        RECT 78.980 270.800 82.930 271.000 ;
        RECT 78.980 270.400 79.330 270.800 ;
        RECT 75.780 262.000 75.980 269.600 ;
        RECT 76.580 262.000 76.780 269.600 ;
        RECT 77.380 262.000 77.580 269.600 ;
        RECT 78.180 262.000 78.380 269.600 ;
        RECT 78.980 269.200 79.330 269.600 ;
        RECT 78.980 269.000 82.930 269.200 ;
        RECT 78.980 268.400 79.330 269.000 ;
        RECT 78.980 268.200 82.930 268.400 ;
        RECT 78.980 267.600 79.330 268.200 ;
        RECT 78.980 267.400 82.930 267.600 ;
        RECT 78.980 266.800 79.330 267.400 ;
        RECT 78.980 266.600 82.930 266.800 ;
        RECT 83.930 266.750 84.330 273.250 ;
        RECT 85.130 266.750 85.530 273.250 ;
        RECT 86.530 273.200 90.480 273.400 ;
        RECT 90.130 272.600 90.480 273.200 ;
        RECT 86.530 272.400 90.480 272.600 ;
        RECT 90.130 271.800 90.480 272.400 ;
        RECT 86.530 271.600 90.480 271.800 ;
        RECT 90.130 271.000 90.480 271.600 ;
        RECT 86.530 270.800 90.480 271.000 ;
        RECT 90.130 270.400 90.480 270.800 ;
        RECT 91.080 270.400 91.280 278.000 ;
        RECT 91.880 270.400 92.080 278.000 ;
        RECT 92.680 270.400 92.880 278.000 ;
        RECT 93.480 270.400 93.680 278.000 ;
        RECT 90.130 269.200 90.480 269.600 ;
        RECT 86.530 269.000 90.480 269.200 ;
        RECT 90.130 268.400 90.480 269.000 ;
        RECT 86.530 268.200 90.480 268.400 ;
        RECT 90.130 267.600 90.480 268.200 ;
        RECT 86.530 267.400 90.480 267.600 ;
        RECT 90.130 266.800 90.480 267.400 ;
        RECT 78.980 266.000 79.330 266.600 ;
        RECT 78.980 265.800 82.930 266.000 ;
        RECT 78.980 265.200 79.330 265.800 ;
        RECT 78.980 265.000 82.930 265.200 ;
        RECT 78.980 264.400 79.330 265.000 ;
        RECT 83.880 264.450 85.580 266.750 ;
        RECT 86.530 266.600 90.480 266.800 ;
        RECT 90.130 266.000 90.480 266.600 ;
        RECT 86.530 265.800 90.480 266.000 ;
        RECT 90.130 265.200 90.480 265.800 ;
        RECT 86.530 265.000 90.480 265.200 ;
        RECT 78.980 264.200 82.930 264.400 ;
        RECT 78.980 263.600 79.330 264.200 ;
        RECT 78.980 263.400 82.930 263.600 ;
        RECT 78.980 262.800 79.330 263.400 ;
        RECT 78.980 262.600 82.930 262.800 ;
        RECT 78.980 262.000 79.330 262.600 ;
        RECT 66.530 261.400 82.930 262.000 ;
        RECT 69.180 260.800 71.480 260.850 ;
        RECT 77.980 260.800 80.280 260.850 ;
        RECT 83.930 260.800 84.330 264.450 ;
        RECT 65.130 260.400 84.330 260.800 ;
        RECT 85.130 260.800 85.530 264.450 ;
        RECT 90.130 264.400 90.480 265.000 ;
        RECT 86.530 264.200 90.480 264.400 ;
        RECT 90.130 263.600 90.480 264.200 ;
        RECT 86.530 263.400 90.480 263.600 ;
        RECT 90.130 262.800 90.480 263.400 ;
        RECT 86.530 262.600 90.480 262.800 ;
        RECT 90.130 262.000 90.480 262.600 ;
        RECT 91.080 262.000 91.280 269.600 ;
        RECT 91.880 262.000 92.080 269.600 ;
        RECT 92.680 262.000 92.880 269.600 ;
        RECT 93.480 262.000 93.680 269.600 ;
        RECT 94.280 262.000 95.180 278.000 ;
        RECT 95.780 270.400 95.980 278.000 ;
        RECT 96.580 270.400 96.780 278.000 ;
        RECT 97.380 270.400 97.580 278.000 ;
        RECT 98.180 270.400 98.380 278.000 ;
        RECT 98.980 277.400 99.330 278.000 ;
        RECT 98.980 277.200 102.930 277.400 ;
        RECT 98.980 276.600 99.330 277.200 ;
        RECT 98.980 276.400 102.930 276.600 ;
        RECT 98.980 275.800 99.330 276.400 ;
        RECT 98.980 275.600 102.930 275.800 ;
        RECT 98.980 275.000 99.330 275.600 ;
        RECT 103.930 275.550 104.330 279.200 ;
        RECT 105.130 279.200 124.330 279.600 ;
        RECT 105.130 275.550 105.530 279.200 ;
        RECT 109.180 279.150 111.480 279.200 ;
        RECT 117.980 279.150 120.280 279.200 ;
        RECT 106.530 278.000 122.930 278.600 ;
        RECT 110.130 277.400 110.480 278.000 ;
        RECT 106.530 277.200 110.480 277.400 ;
        RECT 110.130 276.600 110.480 277.200 ;
        RECT 106.530 276.400 110.480 276.600 ;
        RECT 110.130 275.800 110.480 276.400 ;
        RECT 106.530 275.600 110.480 275.800 ;
        RECT 98.980 274.800 102.930 275.000 ;
        RECT 98.980 274.200 99.330 274.800 ;
        RECT 98.980 274.000 102.930 274.200 ;
        RECT 98.980 273.400 99.330 274.000 ;
        RECT 98.980 273.200 102.930 273.400 ;
        RECT 103.880 273.250 105.580 275.550 ;
        RECT 110.130 275.000 110.480 275.600 ;
        RECT 106.530 274.800 110.480 275.000 ;
        RECT 110.130 274.200 110.480 274.800 ;
        RECT 106.530 274.000 110.480 274.200 ;
        RECT 110.130 273.400 110.480 274.000 ;
        RECT 98.980 272.600 99.330 273.200 ;
        RECT 98.980 272.400 102.930 272.600 ;
        RECT 98.980 271.800 99.330 272.400 ;
        RECT 98.980 271.600 102.930 271.800 ;
        RECT 98.980 271.000 99.330 271.600 ;
        RECT 98.980 270.800 102.930 271.000 ;
        RECT 98.980 270.400 99.330 270.800 ;
        RECT 95.780 262.000 95.980 269.600 ;
        RECT 96.580 262.000 96.780 269.600 ;
        RECT 97.380 262.000 97.580 269.600 ;
        RECT 98.180 262.000 98.380 269.600 ;
        RECT 98.980 269.200 99.330 269.600 ;
        RECT 98.980 269.000 102.930 269.200 ;
        RECT 98.980 268.400 99.330 269.000 ;
        RECT 98.980 268.200 102.930 268.400 ;
        RECT 98.980 267.600 99.330 268.200 ;
        RECT 98.980 267.400 102.930 267.600 ;
        RECT 98.980 266.800 99.330 267.400 ;
        RECT 98.980 266.600 102.930 266.800 ;
        RECT 103.930 266.750 104.330 273.250 ;
        RECT 105.130 266.750 105.530 273.250 ;
        RECT 106.530 273.200 110.480 273.400 ;
        RECT 110.130 272.600 110.480 273.200 ;
        RECT 106.530 272.400 110.480 272.600 ;
        RECT 110.130 271.800 110.480 272.400 ;
        RECT 106.530 271.600 110.480 271.800 ;
        RECT 110.130 271.000 110.480 271.600 ;
        RECT 106.530 270.800 110.480 271.000 ;
        RECT 110.130 270.400 110.480 270.800 ;
        RECT 111.080 270.400 111.280 278.000 ;
        RECT 111.880 270.400 112.080 278.000 ;
        RECT 112.680 270.400 112.880 278.000 ;
        RECT 113.480 270.400 113.680 278.000 ;
        RECT 110.130 269.200 110.480 269.600 ;
        RECT 106.530 269.000 110.480 269.200 ;
        RECT 110.130 268.400 110.480 269.000 ;
        RECT 106.530 268.200 110.480 268.400 ;
        RECT 110.130 267.600 110.480 268.200 ;
        RECT 106.530 267.400 110.480 267.600 ;
        RECT 110.130 266.800 110.480 267.400 ;
        RECT 98.980 266.000 99.330 266.600 ;
        RECT 98.980 265.800 102.930 266.000 ;
        RECT 98.980 265.200 99.330 265.800 ;
        RECT 98.980 265.000 102.930 265.200 ;
        RECT 98.980 264.400 99.330 265.000 ;
        RECT 103.880 264.450 105.580 266.750 ;
        RECT 106.530 266.600 110.480 266.800 ;
        RECT 110.130 266.000 110.480 266.600 ;
        RECT 106.530 265.800 110.480 266.000 ;
        RECT 110.130 265.200 110.480 265.800 ;
        RECT 106.530 265.000 110.480 265.200 ;
        RECT 98.980 264.200 102.930 264.400 ;
        RECT 98.980 263.600 99.330 264.200 ;
        RECT 98.980 263.400 102.930 263.600 ;
        RECT 98.980 262.800 99.330 263.400 ;
        RECT 98.980 262.600 102.930 262.800 ;
        RECT 98.980 262.000 99.330 262.600 ;
        RECT 86.530 261.400 102.930 262.000 ;
        RECT 89.180 260.800 91.480 260.850 ;
        RECT 97.980 260.800 100.280 260.850 ;
        RECT 103.930 260.800 104.330 264.450 ;
        RECT 85.130 260.400 104.330 260.800 ;
        RECT 105.130 260.800 105.530 264.450 ;
        RECT 110.130 264.400 110.480 265.000 ;
        RECT 106.530 264.200 110.480 264.400 ;
        RECT 110.130 263.600 110.480 264.200 ;
        RECT 106.530 263.400 110.480 263.600 ;
        RECT 110.130 262.800 110.480 263.400 ;
        RECT 106.530 262.600 110.480 262.800 ;
        RECT 110.130 262.000 110.480 262.600 ;
        RECT 111.080 262.000 111.280 269.600 ;
        RECT 111.880 262.000 112.080 269.600 ;
        RECT 112.680 262.000 112.880 269.600 ;
        RECT 113.480 262.000 113.680 269.600 ;
        RECT 114.280 262.000 115.180 278.000 ;
        RECT 115.780 270.400 115.980 278.000 ;
        RECT 116.580 270.400 116.780 278.000 ;
        RECT 117.380 270.400 117.580 278.000 ;
        RECT 118.180 270.400 118.380 278.000 ;
        RECT 118.980 277.400 119.330 278.000 ;
        RECT 118.980 277.200 122.930 277.400 ;
        RECT 118.980 276.600 119.330 277.200 ;
        RECT 118.980 276.400 122.930 276.600 ;
        RECT 118.980 275.800 119.330 276.400 ;
        RECT 118.980 275.600 122.930 275.800 ;
        RECT 118.980 275.000 119.330 275.600 ;
        RECT 123.930 275.550 124.330 279.200 ;
        RECT 125.340 277.350 125.700 277.730 ;
        RECT 125.970 277.350 126.330 277.730 ;
        RECT 126.570 277.350 126.930 277.730 ;
        RECT 125.340 276.760 125.700 277.140 ;
        RECT 125.970 276.760 126.330 277.140 ;
        RECT 126.570 276.760 126.930 277.140 ;
        RECT 118.980 274.800 122.930 275.000 ;
        RECT 118.980 274.200 119.330 274.800 ;
        RECT 118.980 274.000 122.930 274.200 ;
        RECT 118.980 273.400 119.330 274.000 ;
        RECT 118.980 273.200 122.930 273.400 ;
        RECT 123.880 273.250 124.730 275.550 ;
        RECT 118.980 272.600 119.330 273.200 ;
        RECT 118.980 272.400 122.930 272.600 ;
        RECT 118.980 271.800 119.330 272.400 ;
        RECT 118.980 271.600 122.930 271.800 ;
        RECT 118.980 271.000 119.330 271.600 ;
        RECT 118.980 270.800 122.930 271.000 ;
        RECT 118.980 270.400 119.330 270.800 ;
        RECT 115.780 262.000 115.980 269.600 ;
        RECT 116.580 262.000 116.780 269.600 ;
        RECT 117.380 262.000 117.580 269.600 ;
        RECT 118.180 262.000 118.380 269.600 ;
        RECT 118.980 269.200 119.330 269.600 ;
        RECT 118.980 269.000 122.930 269.200 ;
        RECT 118.980 268.400 119.330 269.000 ;
        RECT 118.980 268.200 122.930 268.400 ;
        RECT 118.980 267.600 119.330 268.200 ;
        RECT 118.980 267.400 122.930 267.600 ;
        RECT 118.980 266.800 119.330 267.400 ;
        RECT 118.980 266.600 122.930 266.800 ;
        RECT 123.930 266.750 124.330 273.250 ;
        RECT 118.980 266.000 119.330 266.600 ;
        RECT 118.980 265.800 122.930 266.000 ;
        RECT 118.980 265.200 119.330 265.800 ;
        RECT 118.980 265.000 122.930 265.200 ;
        RECT 118.980 264.400 119.330 265.000 ;
        RECT 123.880 264.450 124.730 266.750 ;
        RECT 118.980 264.200 122.930 264.400 ;
        RECT 118.980 263.600 119.330 264.200 ;
        RECT 118.980 263.400 122.930 263.600 ;
        RECT 118.980 262.800 119.330 263.400 ;
        RECT 118.980 262.600 122.930 262.800 ;
        RECT 118.980 262.000 119.330 262.600 ;
        RECT 106.530 261.400 122.930 262.000 ;
        RECT 109.180 260.800 111.480 260.850 ;
        RECT 117.980 260.800 120.280 260.850 ;
        RECT 123.930 260.800 124.330 264.450 ;
        RECT 125.340 262.770 125.700 263.150 ;
        RECT 125.970 262.770 126.330 263.150 ;
        RECT 126.570 262.770 126.930 263.150 ;
        RECT 125.340 262.180 125.700 262.560 ;
        RECT 125.970 262.180 126.330 262.560 ;
        RECT 126.570 262.180 126.930 262.560 ;
        RECT 105.130 260.400 124.330 260.800 ;
        RECT 9.180 259.600 11.480 260.400 ;
        RECT 17.980 259.600 20.280 260.400 ;
        RECT 29.180 259.600 31.480 260.400 ;
        RECT 37.980 259.600 40.280 260.400 ;
        RECT 49.180 259.600 51.480 260.400 ;
        RECT 57.980 259.600 60.280 260.400 ;
        RECT 69.180 259.600 71.480 260.400 ;
        RECT 77.980 259.600 80.280 260.400 ;
        RECT 89.180 259.600 91.480 260.400 ;
        RECT 97.980 259.600 100.280 260.400 ;
        RECT 109.180 259.600 111.480 260.400 ;
        RECT 117.980 259.600 120.280 260.400 ;
        RECT 5.130 259.200 24.330 259.600 ;
        RECT 2.515 257.105 2.875 257.485 ;
        RECT 3.145 257.105 3.505 257.485 ;
        RECT 3.745 257.105 4.105 257.485 ;
        RECT 2.515 256.515 2.875 256.895 ;
        RECT 3.145 256.515 3.505 256.895 ;
        RECT 3.745 256.515 4.105 256.895 ;
        RECT 5.130 255.550 5.530 259.200 ;
        RECT 9.180 259.150 11.480 259.200 ;
        RECT 17.980 259.150 20.280 259.200 ;
        RECT 6.530 258.000 22.930 258.600 ;
        RECT 10.130 257.400 10.480 258.000 ;
        RECT 6.530 257.200 10.480 257.400 ;
        RECT 10.130 256.600 10.480 257.200 ;
        RECT 6.530 256.400 10.480 256.600 ;
        RECT 10.130 255.800 10.480 256.400 ;
        RECT 6.530 255.600 10.480 255.800 ;
        RECT 4.730 255.545 5.580 255.550 ;
        RECT 2.315 253.250 5.580 255.545 ;
        RECT 10.130 255.000 10.480 255.600 ;
        RECT 6.530 254.800 10.480 255.000 ;
        RECT 10.130 254.200 10.480 254.800 ;
        RECT 6.530 254.000 10.480 254.200 ;
        RECT 10.130 253.400 10.480 254.000 ;
        RECT 5.130 246.750 5.530 253.250 ;
        RECT 6.530 253.200 10.480 253.400 ;
        RECT 10.130 252.600 10.480 253.200 ;
        RECT 6.530 252.400 10.480 252.600 ;
        RECT 10.130 251.800 10.480 252.400 ;
        RECT 6.530 251.600 10.480 251.800 ;
        RECT 10.130 251.000 10.480 251.600 ;
        RECT 6.530 250.800 10.480 251.000 ;
        RECT 10.130 250.400 10.480 250.800 ;
        RECT 11.080 250.400 11.280 258.000 ;
        RECT 11.880 250.400 12.080 258.000 ;
        RECT 12.680 250.400 12.880 258.000 ;
        RECT 13.480 250.400 13.680 258.000 ;
        RECT 10.130 249.200 10.480 249.600 ;
        RECT 6.530 249.000 10.480 249.200 ;
        RECT 10.130 248.400 10.480 249.000 ;
        RECT 6.530 248.200 10.480 248.400 ;
        RECT 10.130 247.600 10.480 248.200 ;
        RECT 6.530 247.400 10.480 247.600 ;
        RECT 10.130 246.800 10.480 247.400 ;
        RECT 2.315 244.455 5.580 246.750 ;
        RECT 6.530 246.600 10.480 246.800 ;
        RECT 10.130 246.000 10.480 246.600 ;
        RECT 6.530 245.800 10.480 246.000 ;
        RECT 10.130 245.200 10.480 245.800 ;
        RECT 6.530 245.000 10.480 245.200 ;
        RECT 4.730 244.450 5.580 244.455 ;
        RECT 2.515 243.275 2.875 243.655 ;
        RECT 3.145 243.275 3.505 243.655 ;
        RECT 3.745 243.275 4.105 243.655 ;
        RECT 2.515 242.685 2.875 243.065 ;
        RECT 3.145 242.685 3.505 243.065 ;
        RECT 3.745 242.685 4.105 243.065 ;
        RECT 5.130 240.800 5.530 244.450 ;
        RECT 10.130 244.400 10.480 245.000 ;
        RECT 6.530 244.200 10.480 244.400 ;
        RECT 10.130 243.600 10.480 244.200 ;
        RECT 6.530 243.400 10.480 243.600 ;
        RECT 10.130 242.800 10.480 243.400 ;
        RECT 6.530 242.600 10.480 242.800 ;
        RECT 10.130 242.000 10.480 242.600 ;
        RECT 11.080 242.000 11.280 249.600 ;
        RECT 11.880 242.000 12.080 249.600 ;
        RECT 12.680 242.000 12.880 249.600 ;
        RECT 13.480 242.000 13.680 249.600 ;
        RECT 14.280 242.000 15.180 258.000 ;
        RECT 15.780 250.400 15.980 258.000 ;
        RECT 16.580 250.400 16.780 258.000 ;
        RECT 17.380 250.400 17.580 258.000 ;
        RECT 18.180 250.400 18.380 258.000 ;
        RECT 18.980 257.400 19.330 258.000 ;
        RECT 18.980 257.200 22.930 257.400 ;
        RECT 18.980 256.600 19.330 257.200 ;
        RECT 18.980 256.400 22.930 256.600 ;
        RECT 18.980 255.800 19.330 256.400 ;
        RECT 18.980 255.600 22.930 255.800 ;
        RECT 18.980 255.000 19.330 255.600 ;
        RECT 23.930 255.550 24.330 259.200 ;
        RECT 25.130 259.200 44.330 259.600 ;
        RECT 25.130 255.550 25.530 259.200 ;
        RECT 29.180 259.150 31.480 259.200 ;
        RECT 37.980 259.150 40.280 259.200 ;
        RECT 26.530 258.000 42.930 258.600 ;
        RECT 30.130 257.400 30.480 258.000 ;
        RECT 26.530 257.200 30.480 257.400 ;
        RECT 30.130 256.600 30.480 257.200 ;
        RECT 26.530 256.400 30.480 256.600 ;
        RECT 30.130 255.800 30.480 256.400 ;
        RECT 26.530 255.600 30.480 255.800 ;
        RECT 18.980 254.800 22.930 255.000 ;
        RECT 18.980 254.200 19.330 254.800 ;
        RECT 18.980 254.000 22.930 254.200 ;
        RECT 18.980 253.400 19.330 254.000 ;
        RECT 18.980 253.200 22.930 253.400 ;
        RECT 23.880 253.250 25.580 255.550 ;
        RECT 30.130 255.000 30.480 255.600 ;
        RECT 26.530 254.800 30.480 255.000 ;
        RECT 30.130 254.200 30.480 254.800 ;
        RECT 26.530 254.000 30.480 254.200 ;
        RECT 30.130 253.400 30.480 254.000 ;
        RECT 18.980 252.600 19.330 253.200 ;
        RECT 18.980 252.400 22.930 252.600 ;
        RECT 18.980 251.800 19.330 252.400 ;
        RECT 18.980 251.600 22.930 251.800 ;
        RECT 18.980 251.000 19.330 251.600 ;
        RECT 18.980 250.800 22.930 251.000 ;
        RECT 18.980 250.400 19.330 250.800 ;
        RECT 15.780 242.000 15.980 249.600 ;
        RECT 16.580 242.000 16.780 249.600 ;
        RECT 17.380 242.000 17.580 249.600 ;
        RECT 18.180 242.000 18.380 249.600 ;
        RECT 18.980 249.200 19.330 249.600 ;
        RECT 18.980 249.000 22.930 249.200 ;
        RECT 18.980 248.400 19.330 249.000 ;
        RECT 18.980 248.200 22.930 248.400 ;
        RECT 18.980 247.600 19.330 248.200 ;
        RECT 18.980 247.400 22.930 247.600 ;
        RECT 18.980 246.800 19.330 247.400 ;
        RECT 18.980 246.600 22.930 246.800 ;
        RECT 23.930 246.750 24.330 253.250 ;
        RECT 25.130 246.750 25.530 253.250 ;
        RECT 26.530 253.200 30.480 253.400 ;
        RECT 30.130 252.600 30.480 253.200 ;
        RECT 26.530 252.400 30.480 252.600 ;
        RECT 30.130 251.800 30.480 252.400 ;
        RECT 26.530 251.600 30.480 251.800 ;
        RECT 30.130 251.000 30.480 251.600 ;
        RECT 26.530 250.800 30.480 251.000 ;
        RECT 30.130 250.400 30.480 250.800 ;
        RECT 31.080 250.400 31.280 258.000 ;
        RECT 31.880 250.400 32.080 258.000 ;
        RECT 32.680 250.400 32.880 258.000 ;
        RECT 33.480 250.400 33.680 258.000 ;
        RECT 30.130 249.200 30.480 249.600 ;
        RECT 26.530 249.000 30.480 249.200 ;
        RECT 30.130 248.400 30.480 249.000 ;
        RECT 26.530 248.200 30.480 248.400 ;
        RECT 30.130 247.600 30.480 248.200 ;
        RECT 26.530 247.400 30.480 247.600 ;
        RECT 30.130 246.800 30.480 247.400 ;
        RECT 18.980 246.000 19.330 246.600 ;
        RECT 18.980 245.800 22.930 246.000 ;
        RECT 18.980 245.200 19.330 245.800 ;
        RECT 18.980 245.000 22.930 245.200 ;
        RECT 18.980 244.400 19.330 245.000 ;
        RECT 23.880 244.450 25.580 246.750 ;
        RECT 26.530 246.600 30.480 246.800 ;
        RECT 30.130 246.000 30.480 246.600 ;
        RECT 26.530 245.800 30.480 246.000 ;
        RECT 30.130 245.200 30.480 245.800 ;
        RECT 26.530 245.000 30.480 245.200 ;
        RECT 18.980 244.200 22.930 244.400 ;
        RECT 18.980 243.600 19.330 244.200 ;
        RECT 18.980 243.400 22.930 243.600 ;
        RECT 18.980 242.800 19.330 243.400 ;
        RECT 18.980 242.600 22.930 242.800 ;
        RECT 18.980 242.000 19.330 242.600 ;
        RECT 6.530 241.400 22.930 242.000 ;
        RECT 9.180 240.800 11.480 240.850 ;
        RECT 17.980 240.800 20.280 240.850 ;
        RECT 23.930 240.800 24.330 244.450 ;
        RECT 5.130 240.400 24.330 240.800 ;
        RECT 25.130 240.800 25.530 244.450 ;
        RECT 30.130 244.400 30.480 245.000 ;
        RECT 26.530 244.200 30.480 244.400 ;
        RECT 30.130 243.600 30.480 244.200 ;
        RECT 26.530 243.400 30.480 243.600 ;
        RECT 30.130 242.800 30.480 243.400 ;
        RECT 26.530 242.600 30.480 242.800 ;
        RECT 30.130 242.000 30.480 242.600 ;
        RECT 31.080 242.000 31.280 249.600 ;
        RECT 31.880 242.000 32.080 249.600 ;
        RECT 32.680 242.000 32.880 249.600 ;
        RECT 33.480 242.000 33.680 249.600 ;
        RECT 34.280 242.000 35.180 258.000 ;
        RECT 35.780 250.400 35.980 258.000 ;
        RECT 36.580 250.400 36.780 258.000 ;
        RECT 37.380 250.400 37.580 258.000 ;
        RECT 38.180 250.400 38.380 258.000 ;
        RECT 38.980 257.400 39.330 258.000 ;
        RECT 38.980 257.200 42.930 257.400 ;
        RECT 38.980 256.600 39.330 257.200 ;
        RECT 38.980 256.400 42.930 256.600 ;
        RECT 38.980 255.800 39.330 256.400 ;
        RECT 38.980 255.600 42.930 255.800 ;
        RECT 38.980 255.000 39.330 255.600 ;
        RECT 43.930 255.550 44.330 259.200 ;
        RECT 45.130 259.200 64.330 259.600 ;
        RECT 45.130 255.550 45.530 259.200 ;
        RECT 49.180 259.150 51.480 259.200 ;
        RECT 57.980 259.150 60.280 259.200 ;
        RECT 46.530 258.000 62.930 258.600 ;
        RECT 50.130 257.400 50.480 258.000 ;
        RECT 46.530 257.200 50.480 257.400 ;
        RECT 50.130 256.600 50.480 257.200 ;
        RECT 46.530 256.400 50.480 256.600 ;
        RECT 50.130 255.800 50.480 256.400 ;
        RECT 46.530 255.600 50.480 255.800 ;
        RECT 38.980 254.800 42.930 255.000 ;
        RECT 38.980 254.200 39.330 254.800 ;
        RECT 38.980 254.000 42.930 254.200 ;
        RECT 38.980 253.400 39.330 254.000 ;
        RECT 38.980 253.200 42.930 253.400 ;
        RECT 43.880 253.250 45.580 255.550 ;
        RECT 50.130 255.000 50.480 255.600 ;
        RECT 46.530 254.800 50.480 255.000 ;
        RECT 50.130 254.200 50.480 254.800 ;
        RECT 46.530 254.000 50.480 254.200 ;
        RECT 50.130 253.400 50.480 254.000 ;
        RECT 38.980 252.600 39.330 253.200 ;
        RECT 38.980 252.400 42.930 252.600 ;
        RECT 38.980 251.800 39.330 252.400 ;
        RECT 38.980 251.600 42.930 251.800 ;
        RECT 38.980 251.000 39.330 251.600 ;
        RECT 38.980 250.800 42.930 251.000 ;
        RECT 38.980 250.400 39.330 250.800 ;
        RECT 35.780 242.000 35.980 249.600 ;
        RECT 36.580 242.000 36.780 249.600 ;
        RECT 37.380 242.000 37.580 249.600 ;
        RECT 38.180 242.000 38.380 249.600 ;
        RECT 38.980 249.200 39.330 249.600 ;
        RECT 38.980 249.000 42.930 249.200 ;
        RECT 38.980 248.400 39.330 249.000 ;
        RECT 38.980 248.200 42.930 248.400 ;
        RECT 38.980 247.600 39.330 248.200 ;
        RECT 38.980 247.400 42.930 247.600 ;
        RECT 38.980 246.800 39.330 247.400 ;
        RECT 38.980 246.600 42.930 246.800 ;
        RECT 43.930 246.750 44.330 253.250 ;
        RECT 45.130 246.750 45.530 253.250 ;
        RECT 46.530 253.200 50.480 253.400 ;
        RECT 50.130 252.600 50.480 253.200 ;
        RECT 46.530 252.400 50.480 252.600 ;
        RECT 50.130 251.800 50.480 252.400 ;
        RECT 46.530 251.600 50.480 251.800 ;
        RECT 50.130 251.000 50.480 251.600 ;
        RECT 46.530 250.800 50.480 251.000 ;
        RECT 50.130 250.400 50.480 250.800 ;
        RECT 51.080 250.400 51.280 258.000 ;
        RECT 51.880 250.400 52.080 258.000 ;
        RECT 52.680 250.400 52.880 258.000 ;
        RECT 53.480 250.400 53.680 258.000 ;
        RECT 50.130 249.200 50.480 249.600 ;
        RECT 46.530 249.000 50.480 249.200 ;
        RECT 50.130 248.400 50.480 249.000 ;
        RECT 46.530 248.200 50.480 248.400 ;
        RECT 50.130 247.600 50.480 248.200 ;
        RECT 46.530 247.400 50.480 247.600 ;
        RECT 50.130 246.800 50.480 247.400 ;
        RECT 38.980 246.000 39.330 246.600 ;
        RECT 38.980 245.800 42.930 246.000 ;
        RECT 38.980 245.200 39.330 245.800 ;
        RECT 38.980 245.000 42.930 245.200 ;
        RECT 38.980 244.400 39.330 245.000 ;
        RECT 43.880 244.450 45.580 246.750 ;
        RECT 46.530 246.600 50.480 246.800 ;
        RECT 50.130 246.000 50.480 246.600 ;
        RECT 46.530 245.800 50.480 246.000 ;
        RECT 50.130 245.200 50.480 245.800 ;
        RECT 46.530 245.000 50.480 245.200 ;
        RECT 38.980 244.200 42.930 244.400 ;
        RECT 38.980 243.600 39.330 244.200 ;
        RECT 38.980 243.400 42.930 243.600 ;
        RECT 38.980 242.800 39.330 243.400 ;
        RECT 38.980 242.600 42.930 242.800 ;
        RECT 38.980 242.000 39.330 242.600 ;
        RECT 26.530 241.400 42.930 242.000 ;
        RECT 29.180 240.800 31.480 240.850 ;
        RECT 37.980 240.800 40.280 240.850 ;
        RECT 43.930 240.800 44.330 244.450 ;
        RECT 25.130 240.400 44.330 240.800 ;
        RECT 45.130 240.800 45.530 244.450 ;
        RECT 50.130 244.400 50.480 245.000 ;
        RECT 46.530 244.200 50.480 244.400 ;
        RECT 50.130 243.600 50.480 244.200 ;
        RECT 46.530 243.400 50.480 243.600 ;
        RECT 50.130 242.800 50.480 243.400 ;
        RECT 46.530 242.600 50.480 242.800 ;
        RECT 50.130 242.000 50.480 242.600 ;
        RECT 51.080 242.000 51.280 249.600 ;
        RECT 51.880 242.000 52.080 249.600 ;
        RECT 52.680 242.000 52.880 249.600 ;
        RECT 53.480 242.000 53.680 249.600 ;
        RECT 54.280 242.000 55.180 258.000 ;
        RECT 55.780 250.400 55.980 258.000 ;
        RECT 56.580 250.400 56.780 258.000 ;
        RECT 57.380 250.400 57.580 258.000 ;
        RECT 58.180 250.400 58.380 258.000 ;
        RECT 58.980 257.400 59.330 258.000 ;
        RECT 58.980 257.200 62.930 257.400 ;
        RECT 58.980 256.600 59.330 257.200 ;
        RECT 58.980 256.400 62.930 256.600 ;
        RECT 58.980 255.800 59.330 256.400 ;
        RECT 58.980 255.600 62.930 255.800 ;
        RECT 58.980 255.000 59.330 255.600 ;
        RECT 63.930 255.550 64.330 259.200 ;
        RECT 65.130 259.200 84.330 259.600 ;
        RECT 65.130 255.550 65.530 259.200 ;
        RECT 69.180 259.150 71.480 259.200 ;
        RECT 77.980 259.150 80.280 259.200 ;
        RECT 66.530 258.000 82.930 258.600 ;
        RECT 70.130 257.400 70.480 258.000 ;
        RECT 66.530 257.200 70.480 257.400 ;
        RECT 70.130 256.600 70.480 257.200 ;
        RECT 66.530 256.400 70.480 256.600 ;
        RECT 70.130 255.800 70.480 256.400 ;
        RECT 66.530 255.600 70.480 255.800 ;
        RECT 58.980 254.800 62.930 255.000 ;
        RECT 58.980 254.200 59.330 254.800 ;
        RECT 58.980 254.000 62.930 254.200 ;
        RECT 58.980 253.400 59.330 254.000 ;
        RECT 58.980 253.200 62.930 253.400 ;
        RECT 63.880 253.250 65.580 255.550 ;
        RECT 70.130 255.000 70.480 255.600 ;
        RECT 66.530 254.800 70.480 255.000 ;
        RECT 70.130 254.200 70.480 254.800 ;
        RECT 66.530 254.000 70.480 254.200 ;
        RECT 70.130 253.400 70.480 254.000 ;
        RECT 58.980 252.600 59.330 253.200 ;
        RECT 58.980 252.400 62.930 252.600 ;
        RECT 58.980 251.800 59.330 252.400 ;
        RECT 58.980 251.600 62.930 251.800 ;
        RECT 58.980 251.000 59.330 251.600 ;
        RECT 58.980 250.800 62.930 251.000 ;
        RECT 58.980 250.400 59.330 250.800 ;
        RECT 55.780 242.000 55.980 249.600 ;
        RECT 56.580 242.000 56.780 249.600 ;
        RECT 57.380 242.000 57.580 249.600 ;
        RECT 58.180 242.000 58.380 249.600 ;
        RECT 58.980 249.200 59.330 249.600 ;
        RECT 58.980 249.000 62.930 249.200 ;
        RECT 58.980 248.400 59.330 249.000 ;
        RECT 58.980 248.200 62.930 248.400 ;
        RECT 58.980 247.600 59.330 248.200 ;
        RECT 58.980 247.400 62.930 247.600 ;
        RECT 58.980 246.800 59.330 247.400 ;
        RECT 58.980 246.600 62.930 246.800 ;
        RECT 63.930 246.750 64.330 253.250 ;
        RECT 65.130 246.750 65.530 253.250 ;
        RECT 66.530 253.200 70.480 253.400 ;
        RECT 70.130 252.600 70.480 253.200 ;
        RECT 66.530 252.400 70.480 252.600 ;
        RECT 70.130 251.800 70.480 252.400 ;
        RECT 66.530 251.600 70.480 251.800 ;
        RECT 70.130 251.000 70.480 251.600 ;
        RECT 66.530 250.800 70.480 251.000 ;
        RECT 70.130 250.400 70.480 250.800 ;
        RECT 71.080 250.400 71.280 258.000 ;
        RECT 71.880 250.400 72.080 258.000 ;
        RECT 72.680 250.400 72.880 258.000 ;
        RECT 73.480 250.400 73.680 258.000 ;
        RECT 70.130 249.200 70.480 249.600 ;
        RECT 66.530 249.000 70.480 249.200 ;
        RECT 70.130 248.400 70.480 249.000 ;
        RECT 66.530 248.200 70.480 248.400 ;
        RECT 70.130 247.600 70.480 248.200 ;
        RECT 66.530 247.400 70.480 247.600 ;
        RECT 70.130 246.800 70.480 247.400 ;
        RECT 58.980 246.000 59.330 246.600 ;
        RECT 58.980 245.800 62.930 246.000 ;
        RECT 58.980 245.200 59.330 245.800 ;
        RECT 58.980 245.000 62.930 245.200 ;
        RECT 58.980 244.400 59.330 245.000 ;
        RECT 63.880 244.450 65.580 246.750 ;
        RECT 66.530 246.600 70.480 246.800 ;
        RECT 70.130 246.000 70.480 246.600 ;
        RECT 66.530 245.800 70.480 246.000 ;
        RECT 70.130 245.200 70.480 245.800 ;
        RECT 66.530 245.000 70.480 245.200 ;
        RECT 58.980 244.200 62.930 244.400 ;
        RECT 58.980 243.600 59.330 244.200 ;
        RECT 58.980 243.400 62.930 243.600 ;
        RECT 58.980 242.800 59.330 243.400 ;
        RECT 58.980 242.600 62.930 242.800 ;
        RECT 58.980 242.000 59.330 242.600 ;
        RECT 46.530 241.400 62.930 242.000 ;
        RECT 49.180 240.800 51.480 240.850 ;
        RECT 57.980 240.800 60.280 240.850 ;
        RECT 63.930 240.800 64.330 244.450 ;
        RECT 45.130 240.400 64.330 240.800 ;
        RECT 65.130 240.800 65.530 244.450 ;
        RECT 70.130 244.400 70.480 245.000 ;
        RECT 66.530 244.200 70.480 244.400 ;
        RECT 70.130 243.600 70.480 244.200 ;
        RECT 66.530 243.400 70.480 243.600 ;
        RECT 70.130 242.800 70.480 243.400 ;
        RECT 66.530 242.600 70.480 242.800 ;
        RECT 70.130 242.000 70.480 242.600 ;
        RECT 71.080 242.000 71.280 249.600 ;
        RECT 71.880 242.000 72.080 249.600 ;
        RECT 72.680 242.000 72.880 249.600 ;
        RECT 73.480 242.000 73.680 249.600 ;
        RECT 74.280 242.000 75.180 258.000 ;
        RECT 75.780 250.400 75.980 258.000 ;
        RECT 76.580 250.400 76.780 258.000 ;
        RECT 77.380 250.400 77.580 258.000 ;
        RECT 78.180 250.400 78.380 258.000 ;
        RECT 78.980 257.400 79.330 258.000 ;
        RECT 78.980 257.200 82.930 257.400 ;
        RECT 78.980 256.600 79.330 257.200 ;
        RECT 78.980 256.400 82.930 256.600 ;
        RECT 78.980 255.800 79.330 256.400 ;
        RECT 78.980 255.600 82.930 255.800 ;
        RECT 78.980 255.000 79.330 255.600 ;
        RECT 83.930 255.550 84.330 259.200 ;
        RECT 85.130 259.200 104.330 259.600 ;
        RECT 85.130 255.550 85.530 259.200 ;
        RECT 89.180 259.150 91.480 259.200 ;
        RECT 97.980 259.150 100.280 259.200 ;
        RECT 86.530 258.000 102.930 258.600 ;
        RECT 90.130 257.400 90.480 258.000 ;
        RECT 86.530 257.200 90.480 257.400 ;
        RECT 90.130 256.600 90.480 257.200 ;
        RECT 86.530 256.400 90.480 256.600 ;
        RECT 90.130 255.800 90.480 256.400 ;
        RECT 86.530 255.600 90.480 255.800 ;
        RECT 78.980 254.800 82.930 255.000 ;
        RECT 78.980 254.200 79.330 254.800 ;
        RECT 78.980 254.000 82.930 254.200 ;
        RECT 78.980 253.400 79.330 254.000 ;
        RECT 78.980 253.200 82.930 253.400 ;
        RECT 83.880 253.250 85.580 255.550 ;
        RECT 90.130 255.000 90.480 255.600 ;
        RECT 86.530 254.800 90.480 255.000 ;
        RECT 90.130 254.200 90.480 254.800 ;
        RECT 86.530 254.000 90.480 254.200 ;
        RECT 90.130 253.400 90.480 254.000 ;
        RECT 78.980 252.600 79.330 253.200 ;
        RECT 78.980 252.400 82.930 252.600 ;
        RECT 78.980 251.800 79.330 252.400 ;
        RECT 78.980 251.600 82.930 251.800 ;
        RECT 78.980 251.000 79.330 251.600 ;
        RECT 78.980 250.800 82.930 251.000 ;
        RECT 78.980 250.400 79.330 250.800 ;
        RECT 75.780 242.000 75.980 249.600 ;
        RECT 76.580 242.000 76.780 249.600 ;
        RECT 77.380 242.000 77.580 249.600 ;
        RECT 78.180 242.000 78.380 249.600 ;
        RECT 78.980 249.200 79.330 249.600 ;
        RECT 78.980 249.000 82.930 249.200 ;
        RECT 78.980 248.400 79.330 249.000 ;
        RECT 78.980 248.200 82.930 248.400 ;
        RECT 78.980 247.600 79.330 248.200 ;
        RECT 78.980 247.400 82.930 247.600 ;
        RECT 78.980 246.800 79.330 247.400 ;
        RECT 78.980 246.600 82.930 246.800 ;
        RECT 83.930 246.750 84.330 253.250 ;
        RECT 85.130 246.750 85.530 253.250 ;
        RECT 86.530 253.200 90.480 253.400 ;
        RECT 90.130 252.600 90.480 253.200 ;
        RECT 86.530 252.400 90.480 252.600 ;
        RECT 90.130 251.800 90.480 252.400 ;
        RECT 86.530 251.600 90.480 251.800 ;
        RECT 90.130 251.000 90.480 251.600 ;
        RECT 86.530 250.800 90.480 251.000 ;
        RECT 90.130 250.400 90.480 250.800 ;
        RECT 91.080 250.400 91.280 258.000 ;
        RECT 91.880 250.400 92.080 258.000 ;
        RECT 92.680 250.400 92.880 258.000 ;
        RECT 93.480 250.400 93.680 258.000 ;
        RECT 90.130 249.200 90.480 249.600 ;
        RECT 86.530 249.000 90.480 249.200 ;
        RECT 90.130 248.400 90.480 249.000 ;
        RECT 86.530 248.200 90.480 248.400 ;
        RECT 90.130 247.600 90.480 248.200 ;
        RECT 86.530 247.400 90.480 247.600 ;
        RECT 90.130 246.800 90.480 247.400 ;
        RECT 78.980 246.000 79.330 246.600 ;
        RECT 78.980 245.800 82.930 246.000 ;
        RECT 78.980 245.200 79.330 245.800 ;
        RECT 78.980 245.000 82.930 245.200 ;
        RECT 78.980 244.400 79.330 245.000 ;
        RECT 83.880 244.450 85.580 246.750 ;
        RECT 86.530 246.600 90.480 246.800 ;
        RECT 90.130 246.000 90.480 246.600 ;
        RECT 86.530 245.800 90.480 246.000 ;
        RECT 90.130 245.200 90.480 245.800 ;
        RECT 86.530 245.000 90.480 245.200 ;
        RECT 78.980 244.200 82.930 244.400 ;
        RECT 78.980 243.600 79.330 244.200 ;
        RECT 78.980 243.400 82.930 243.600 ;
        RECT 78.980 242.800 79.330 243.400 ;
        RECT 78.980 242.600 82.930 242.800 ;
        RECT 78.980 242.000 79.330 242.600 ;
        RECT 66.530 241.400 82.930 242.000 ;
        RECT 69.180 240.800 71.480 240.850 ;
        RECT 77.980 240.800 80.280 240.850 ;
        RECT 83.930 240.800 84.330 244.450 ;
        RECT 65.130 240.400 84.330 240.800 ;
        RECT 85.130 240.800 85.530 244.450 ;
        RECT 90.130 244.400 90.480 245.000 ;
        RECT 86.530 244.200 90.480 244.400 ;
        RECT 90.130 243.600 90.480 244.200 ;
        RECT 86.530 243.400 90.480 243.600 ;
        RECT 90.130 242.800 90.480 243.400 ;
        RECT 86.530 242.600 90.480 242.800 ;
        RECT 90.130 242.000 90.480 242.600 ;
        RECT 91.080 242.000 91.280 249.600 ;
        RECT 91.880 242.000 92.080 249.600 ;
        RECT 92.680 242.000 92.880 249.600 ;
        RECT 93.480 242.000 93.680 249.600 ;
        RECT 94.280 242.000 95.180 258.000 ;
        RECT 95.780 250.400 95.980 258.000 ;
        RECT 96.580 250.400 96.780 258.000 ;
        RECT 97.380 250.400 97.580 258.000 ;
        RECT 98.180 250.400 98.380 258.000 ;
        RECT 98.980 257.400 99.330 258.000 ;
        RECT 98.980 257.200 102.930 257.400 ;
        RECT 98.980 256.600 99.330 257.200 ;
        RECT 98.980 256.400 102.930 256.600 ;
        RECT 98.980 255.800 99.330 256.400 ;
        RECT 98.980 255.600 102.930 255.800 ;
        RECT 98.980 255.000 99.330 255.600 ;
        RECT 103.930 255.550 104.330 259.200 ;
        RECT 105.130 259.200 124.330 259.600 ;
        RECT 105.130 255.550 105.530 259.200 ;
        RECT 109.180 259.150 111.480 259.200 ;
        RECT 117.980 259.150 120.280 259.200 ;
        RECT 106.530 258.000 122.930 258.600 ;
        RECT 110.130 257.400 110.480 258.000 ;
        RECT 106.530 257.200 110.480 257.400 ;
        RECT 110.130 256.600 110.480 257.200 ;
        RECT 106.530 256.400 110.480 256.600 ;
        RECT 110.130 255.800 110.480 256.400 ;
        RECT 106.530 255.600 110.480 255.800 ;
        RECT 98.980 254.800 102.930 255.000 ;
        RECT 98.980 254.200 99.330 254.800 ;
        RECT 98.980 254.000 102.930 254.200 ;
        RECT 98.980 253.400 99.330 254.000 ;
        RECT 98.980 253.200 102.930 253.400 ;
        RECT 103.880 253.250 105.580 255.550 ;
        RECT 110.130 255.000 110.480 255.600 ;
        RECT 106.530 254.800 110.480 255.000 ;
        RECT 110.130 254.200 110.480 254.800 ;
        RECT 106.530 254.000 110.480 254.200 ;
        RECT 110.130 253.400 110.480 254.000 ;
        RECT 98.980 252.600 99.330 253.200 ;
        RECT 98.980 252.400 102.930 252.600 ;
        RECT 98.980 251.800 99.330 252.400 ;
        RECT 98.980 251.600 102.930 251.800 ;
        RECT 98.980 251.000 99.330 251.600 ;
        RECT 98.980 250.800 102.930 251.000 ;
        RECT 98.980 250.400 99.330 250.800 ;
        RECT 95.780 242.000 95.980 249.600 ;
        RECT 96.580 242.000 96.780 249.600 ;
        RECT 97.380 242.000 97.580 249.600 ;
        RECT 98.180 242.000 98.380 249.600 ;
        RECT 98.980 249.200 99.330 249.600 ;
        RECT 98.980 249.000 102.930 249.200 ;
        RECT 98.980 248.400 99.330 249.000 ;
        RECT 98.980 248.200 102.930 248.400 ;
        RECT 98.980 247.600 99.330 248.200 ;
        RECT 98.980 247.400 102.930 247.600 ;
        RECT 98.980 246.800 99.330 247.400 ;
        RECT 98.980 246.600 102.930 246.800 ;
        RECT 103.930 246.750 104.330 253.250 ;
        RECT 105.130 246.750 105.530 253.250 ;
        RECT 106.530 253.200 110.480 253.400 ;
        RECT 110.130 252.600 110.480 253.200 ;
        RECT 106.530 252.400 110.480 252.600 ;
        RECT 110.130 251.800 110.480 252.400 ;
        RECT 106.530 251.600 110.480 251.800 ;
        RECT 110.130 251.000 110.480 251.600 ;
        RECT 106.530 250.800 110.480 251.000 ;
        RECT 110.130 250.400 110.480 250.800 ;
        RECT 111.080 250.400 111.280 258.000 ;
        RECT 111.880 250.400 112.080 258.000 ;
        RECT 112.680 250.400 112.880 258.000 ;
        RECT 113.480 250.400 113.680 258.000 ;
        RECT 110.130 249.200 110.480 249.600 ;
        RECT 106.530 249.000 110.480 249.200 ;
        RECT 110.130 248.400 110.480 249.000 ;
        RECT 106.530 248.200 110.480 248.400 ;
        RECT 110.130 247.600 110.480 248.200 ;
        RECT 106.530 247.400 110.480 247.600 ;
        RECT 110.130 246.800 110.480 247.400 ;
        RECT 98.980 246.000 99.330 246.600 ;
        RECT 98.980 245.800 102.930 246.000 ;
        RECT 98.980 245.200 99.330 245.800 ;
        RECT 98.980 245.000 102.930 245.200 ;
        RECT 98.980 244.400 99.330 245.000 ;
        RECT 103.880 244.450 105.580 246.750 ;
        RECT 106.530 246.600 110.480 246.800 ;
        RECT 110.130 246.000 110.480 246.600 ;
        RECT 106.530 245.800 110.480 246.000 ;
        RECT 110.130 245.200 110.480 245.800 ;
        RECT 106.530 245.000 110.480 245.200 ;
        RECT 98.980 244.200 102.930 244.400 ;
        RECT 98.980 243.600 99.330 244.200 ;
        RECT 98.980 243.400 102.930 243.600 ;
        RECT 98.980 242.800 99.330 243.400 ;
        RECT 98.980 242.600 102.930 242.800 ;
        RECT 98.980 242.000 99.330 242.600 ;
        RECT 86.530 241.400 102.930 242.000 ;
        RECT 89.180 240.800 91.480 240.850 ;
        RECT 97.980 240.800 100.280 240.850 ;
        RECT 103.930 240.800 104.330 244.450 ;
        RECT 85.130 240.400 104.330 240.800 ;
        RECT 105.130 240.800 105.530 244.450 ;
        RECT 110.130 244.400 110.480 245.000 ;
        RECT 106.530 244.200 110.480 244.400 ;
        RECT 110.130 243.600 110.480 244.200 ;
        RECT 106.530 243.400 110.480 243.600 ;
        RECT 110.130 242.800 110.480 243.400 ;
        RECT 106.530 242.600 110.480 242.800 ;
        RECT 110.130 242.000 110.480 242.600 ;
        RECT 111.080 242.000 111.280 249.600 ;
        RECT 111.880 242.000 112.080 249.600 ;
        RECT 112.680 242.000 112.880 249.600 ;
        RECT 113.480 242.000 113.680 249.600 ;
        RECT 114.280 242.000 115.180 258.000 ;
        RECT 115.780 250.400 115.980 258.000 ;
        RECT 116.580 250.400 116.780 258.000 ;
        RECT 117.380 250.400 117.580 258.000 ;
        RECT 118.180 250.400 118.380 258.000 ;
        RECT 118.980 257.400 119.330 258.000 ;
        RECT 118.980 257.200 122.930 257.400 ;
        RECT 118.980 256.600 119.330 257.200 ;
        RECT 118.980 256.400 122.930 256.600 ;
        RECT 118.980 255.800 119.330 256.400 ;
        RECT 118.980 255.600 122.930 255.800 ;
        RECT 118.980 255.000 119.330 255.600 ;
        RECT 123.930 255.550 124.330 259.200 ;
        RECT 125.340 256.855 125.700 257.235 ;
        RECT 125.970 256.855 126.330 257.235 ;
        RECT 126.570 256.855 126.930 257.235 ;
        RECT 125.340 256.265 125.700 256.645 ;
        RECT 125.970 256.265 126.330 256.645 ;
        RECT 126.570 256.265 126.930 256.645 ;
        RECT 118.980 254.800 122.930 255.000 ;
        RECT 118.980 254.200 119.330 254.800 ;
        RECT 118.980 254.000 122.930 254.200 ;
        RECT 118.980 253.400 119.330 254.000 ;
        RECT 118.980 253.200 122.930 253.400 ;
        RECT 123.880 253.250 124.730 255.550 ;
        RECT 118.980 252.600 119.330 253.200 ;
        RECT 118.980 252.400 122.930 252.600 ;
        RECT 118.980 251.800 119.330 252.400 ;
        RECT 118.980 251.600 122.930 251.800 ;
        RECT 118.980 251.000 119.330 251.600 ;
        RECT 118.980 250.800 122.930 251.000 ;
        RECT 118.980 250.400 119.330 250.800 ;
        RECT 115.780 242.000 115.980 249.600 ;
        RECT 116.580 242.000 116.780 249.600 ;
        RECT 117.380 242.000 117.580 249.600 ;
        RECT 118.180 242.000 118.380 249.600 ;
        RECT 118.980 249.200 119.330 249.600 ;
        RECT 118.980 249.000 122.930 249.200 ;
        RECT 118.980 248.400 119.330 249.000 ;
        RECT 118.980 248.200 122.930 248.400 ;
        RECT 118.980 247.600 119.330 248.200 ;
        RECT 118.980 247.400 122.930 247.600 ;
        RECT 118.980 246.800 119.330 247.400 ;
        RECT 118.980 246.600 122.930 246.800 ;
        RECT 123.930 246.750 124.330 253.250 ;
        RECT 118.980 246.000 119.330 246.600 ;
        RECT 118.980 245.800 122.930 246.000 ;
        RECT 118.980 245.200 119.330 245.800 ;
        RECT 118.980 245.000 122.930 245.200 ;
        RECT 118.980 244.400 119.330 245.000 ;
        RECT 123.880 244.450 124.730 246.750 ;
        RECT 118.980 244.200 122.930 244.400 ;
        RECT 118.980 243.600 119.330 244.200 ;
        RECT 118.980 243.400 122.930 243.600 ;
        RECT 118.980 242.800 119.330 243.400 ;
        RECT 118.980 242.600 122.930 242.800 ;
        RECT 118.980 242.000 119.330 242.600 ;
        RECT 106.530 241.400 122.930 242.000 ;
        RECT 109.180 240.800 111.480 240.850 ;
        RECT 117.980 240.800 120.280 240.850 ;
        RECT 123.930 240.800 124.330 244.450 ;
        RECT 125.340 242.495 125.700 242.875 ;
        RECT 125.970 242.495 126.330 242.875 ;
        RECT 126.570 242.495 126.930 242.875 ;
        RECT 125.340 241.905 125.700 242.285 ;
        RECT 125.970 241.905 126.330 242.285 ;
        RECT 126.570 241.905 126.930 242.285 ;
        RECT 105.130 240.400 124.330 240.800 ;
        RECT 9.180 239.600 11.480 240.400 ;
        RECT 17.980 239.600 20.280 240.400 ;
        RECT 29.180 239.600 31.480 240.400 ;
        RECT 37.980 239.600 40.280 240.400 ;
        RECT 49.180 239.600 51.480 240.400 ;
        RECT 57.980 239.600 60.280 240.400 ;
        RECT 69.180 239.600 71.480 240.400 ;
        RECT 77.980 239.600 80.280 240.400 ;
        RECT 89.180 239.600 91.480 240.400 ;
        RECT 97.980 239.600 100.280 240.400 ;
        RECT 109.180 239.600 111.480 240.400 ;
        RECT 117.980 239.600 120.280 240.400 ;
        RECT 5.130 239.200 24.330 239.600 ;
        RECT 2.515 237.340 2.875 237.720 ;
        RECT 3.145 237.340 3.505 237.720 ;
        RECT 3.745 237.340 4.105 237.720 ;
        RECT 2.515 236.750 2.875 237.130 ;
        RECT 3.145 236.750 3.505 237.130 ;
        RECT 3.745 236.750 4.105 237.130 ;
        RECT 5.130 235.550 5.530 239.200 ;
        RECT 9.180 239.150 11.480 239.200 ;
        RECT 17.980 239.150 20.280 239.200 ;
        RECT 6.530 238.000 22.930 238.600 ;
        RECT 10.130 237.400 10.480 238.000 ;
        RECT 6.530 237.200 10.480 237.400 ;
        RECT 10.130 236.600 10.480 237.200 ;
        RECT 6.530 236.400 10.480 236.600 ;
        RECT 10.130 235.800 10.480 236.400 ;
        RECT 6.530 235.600 10.480 235.800 ;
        RECT 4.730 235.545 5.580 235.550 ;
        RECT 2.315 233.250 5.580 235.545 ;
        RECT 10.130 235.000 10.480 235.600 ;
        RECT 6.530 234.800 10.480 235.000 ;
        RECT 10.130 234.200 10.480 234.800 ;
        RECT 6.530 234.000 10.480 234.200 ;
        RECT 10.130 233.400 10.480 234.000 ;
        RECT 5.130 226.750 5.530 233.250 ;
        RECT 6.530 233.200 10.480 233.400 ;
        RECT 10.130 232.600 10.480 233.200 ;
        RECT 6.530 232.400 10.480 232.600 ;
        RECT 10.130 231.800 10.480 232.400 ;
        RECT 6.530 231.600 10.480 231.800 ;
        RECT 10.130 231.000 10.480 231.600 ;
        RECT 6.530 230.800 10.480 231.000 ;
        RECT 10.130 230.400 10.480 230.800 ;
        RECT 11.080 230.400 11.280 238.000 ;
        RECT 11.880 230.400 12.080 238.000 ;
        RECT 12.680 230.400 12.880 238.000 ;
        RECT 13.480 230.400 13.680 238.000 ;
        RECT 10.130 229.200 10.480 229.600 ;
        RECT 6.530 229.000 10.480 229.200 ;
        RECT 10.130 228.400 10.480 229.000 ;
        RECT 6.530 228.200 10.480 228.400 ;
        RECT 10.130 227.600 10.480 228.200 ;
        RECT 6.530 227.400 10.480 227.600 ;
        RECT 10.130 226.800 10.480 227.400 ;
        RECT 2.315 224.455 5.580 226.750 ;
        RECT 6.530 226.600 10.480 226.800 ;
        RECT 10.130 226.000 10.480 226.600 ;
        RECT 6.530 225.800 10.480 226.000 ;
        RECT 10.130 225.200 10.480 225.800 ;
        RECT 6.530 225.000 10.480 225.200 ;
        RECT 4.730 224.450 5.580 224.455 ;
        RECT 2.515 223.230 2.875 223.610 ;
        RECT 3.145 223.230 3.505 223.610 ;
        RECT 3.745 223.230 4.105 223.610 ;
        RECT 2.515 222.640 2.875 223.020 ;
        RECT 3.145 222.640 3.505 223.020 ;
        RECT 3.745 222.640 4.105 223.020 ;
        RECT 5.130 220.800 5.530 224.450 ;
        RECT 10.130 224.400 10.480 225.000 ;
        RECT 6.530 224.200 10.480 224.400 ;
        RECT 10.130 223.600 10.480 224.200 ;
        RECT 6.530 223.400 10.480 223.600 ;
        RECT 10.130 222.800 10.480 223.400 ;
        RECT 6.530 222.600 10.480 222.800 ;
        RECT 10.130 222.000 10.480 222.600 ;
        RECT 11.080 222.000 11.280 229.600 ;
        RECT 11.880 222.000 12.080 229.600 ;
        RECT 12.680 222.000 12.880 229.600 ;
        RECT 13.480 222.000 13.680 229.600 ;
        RECT 14.280 222.000 15.180 238.000 ;
        RECT 15.780 230.400 15.980 238.000 ;
        RECT 16.580 230.400 16.780 238.000 ;
        RECT 17.380 230.400 17.580 238.000 ;
        RECT 18.180 230.400 18.380 238.000 ;
        RECT 18.980 237.400 19.330 238.000 ;
        RECT 18.980 237.200 22.930 237.400 ;
        RECT 18.980 236.600 19.330 237.200 ;
        RECT 18.980 236.400 22.930 236.600 ;
        RECT 18.980 235.800 19.330 236.400 ;
        RECT 18.980 235.600 22.930 235.800 ;
        RECT 18.980 235.000 19.330 235.600 ;
        RECT 23.930 235.550 24.330 239.200 ;
        RECT 25.130 239.200 44.330 239.600 ;
        RECT 25.130 235.550 25.530 239.200 ;
        RECT 29.180 239.150 31.480 239.200 ;
        RECT 37.980 239.150 40.280 239.200 ;
        RECT 26.530 238.000 42.930 238.600 ;
        RECT 30.130 237.400 30.480 238.000 ;
        RECT 26.530 237.200 30.480 237.400 ;
        RECT 30.130 236.600 30.480 237.200 ;
        RECT 26.530 236.400 30.480 236.600 ;
        RECT 30.130 235.800 30.480 236.400 ;
        RECT 26.530 235.600 30.480 235.800 ;
        RECT 18.980 234.800 22.930 235.000 ;
        RECT 18.980 234.200 19.330 234.800 ;
        RECT 18.980 234.000 22.930 234.200 ;
        RECT 18.980 233.400 19.330 234.000 ;
        RECT 18.980 233.200 22.930 233.400 ;
        RECT 23.880 233.250 25.580 235.550 ;
        RECT 30.130 235.000 30.480 235.600 ;
        RECT 26.530 234.800 30.480 235.000 ;
        RECT 30.130 234.200 30.480 234.800 ;
        RECT 26.530 234.000 30.480 234.200 ;
        RECT 30.130 233.400 30.480 234.000 ;
        RECT 18.980 232.600 19.330 233.200 ;
        RECT 18.980 232.400 22.930 232.600 ;
        RECT 18.980 231.800 19.330 232.400 ;
        RECT 18.980 231.600 22.930 231.800 ;
        RECT 18.980 231.000 19.330 231.600 ;
        RECT 18.980 230.800 22.930 231.000 ;
        RECT 18.980 230.400 19.330 230.800 ;
        RECT 15.780 222.000 15.980 229.600 ;
        RECT 16.580 222.000 16.780 229.600 ;
        RECT 17.380 222.000 17.580 229.600 ;
        RECT 18.180 222.000 18.380 229.600 ;
        RECT 18.980 229.200 19.330 229.600 ;
        RECT 18.980 229.000 22.930 229.200 ;
        RECT 18.980 228.400 19.330 229.000 ;
        RECT 18.980 228.200 22.930 228.400 ;
        RECT 18.980 227.600 19.330 228.200 ;
        RECT 18.980 227.400 22.930 227.600 ;
        RECT 18.980 226.800 19.330 227.400 ;
        RECT 18.980 226.600 22.930 226.800 ;
        RECT 23.930 226.750 24.330 233.250 ;
        RECT 25.130 226.750 25.530 233.250 ;
        RECT 26.530 233.200 30.480 233.400 ;
        RECT 30.130 232.600 30.480 233.200 ;
        RECT 26.530 232.400 30.480 232.600 ;
        RECT 30.130 231.800 30.480 232.400 ;
        RECT 26.530 231.600 30.480 231.800 ;
        RECT 30.130 231.000 30.480 231.600 ;
        RECT 26.530 230.800 30.480 231.000 ;
        RECT 30.130 230.400 30.480 230.800 ;
        RECT 31.080 230.400 31.280 238.000 ;
        RECT 31.880 230.400 32.080 238.000 ;
        RECT 32.680 230.400 32.880 238.000 ;
        RECT 33.480 230.400 33.680 238.000 ;
        RECT 30.130 229.200 30.480 229.600 ;
        RECT 26.530 229.000 30.480 229.200 ;
        RECT 30.130 228.400 30.480 229.000 ;
        RECT 26.530 228.200 30.480 228.400 ;
        RECT 30.130 227.600 30.480 228.200 ;
        RECT 26.530 227.400 30.480 227.600 ;
        RECT 30.130 226.800 30.480 227.400 ;
        RECT 18.980 226.000 19.330 226.600 ;
        RECT 18.980 225.800 22.930 226.000 ;
        RECT 18.980 225.200 19.330 225.800 ;
        RECT 18.980 225.000 22.930 225.200 ;
        RECT 18.980 224.400 19.330 225.000 ;
        RECT 23.880 224.450 25.580 226.750 ;
        RECT 26.530 226.600 30.480 226.800 ;
        RECT 30.130 226.000 30.480 226.600 ;
        RECT 26.530 225.800 30.480 226.000 ;
        RECT 30.130 225.200 30.480 225.800 ;
        RECT 26.530 225.000 30.480 225.200 ;
        RECT 18.980 224.200 22.930 224.400 ;
        RECT 18.980 223.600 19.330 224.200 ;
        RECT 18.980 223.400 22.930 223.600 ;
        RECT 18.980 222.800 19.330 223.400 ;
        RECT 18.980 222.600 22.930 222.800 ;
        RECT 18.980 222.000 19.330 222.600 ;
        RECT 6.530 221.400 22.930 222.000 ;
        RECT 9.180 220.800 11.480 220.850 ;
        RECT 17.980 220.800 20.280 220.850 ;
        RECT 23.930 220.800 24.330 224.450 ;
        RECT 5.130 220.400 24.330 220.800 ;
        RECT 25.130 220.800 25.530 224.450 ;
        RECT 30.130 224.400 30.480 225.000 ;
        RECT 26.530 224.200 30.480 224.400 ;
        RECT 30.130 223.600 30.480 224.200 ;
        RECT 26.530 223.400 30.480 223.600 ;
        RECT 30.130 222.800 30.480 223.400 ;
        RECT 26.530 222.600 30.480 222.800 ;
        RECT 30.130 222.000 30.480 222.600 ;
        RECT 31.080 222.000 31.280 229.600 ;
        RECT 31.880 222.000 32.080 229.600 ;
        RECT 32.680 222.000 32.880 229.600 ;
        RECT 33.480 222.000 33.680 229.600 ;
        RECT 34.280 222.000 35.180 238.000 ;
        RECT 35.780 230.400 35.980 238.000 ;
        RECT 36.580 230.400 36.780 238.000 ;
        RECT 37.380 230.400 37.580 238.000 ;
        RECT 38.180 230.400 38.380 238.000 ;
        RECT 38.980 237.400 39.330 238.000 ;
        RECT 38.980 237.200 42.930 237.400 ;
        RECT 38.980 236.600 39.330 237.200 ;
        RECT 38.980 236.400 42.930 236.600 ;
        RECT 38.980 235.800 39.330 236.400 ;
        RECT 38.980 235.600 42.930 235.800 ;
        RECT 38.980 235.000 39.330 235.600 ;
        RECT 43.930 235.550 44.330 239.200 ;
        RECT 45.130 239.200 64.330 239.600 ;
        RECT 45.130 235.550 45.530 239.200 ;
        RECT 49.180 239.150 51.480 239.200 ;
        RECT 57.980 239.150 60.280 239.200 ;
        RECT 46.530 238.000 62.930 238.600 ;
        RECT 50.130 237.400 50.480 238.000 ;
        RECT 46.530 237.200 50.480 237.400 ;
        RECT 50.130 236.600 50.480 237.200 ;
        RECT 46.530 236.400 50.480 236.600 ;
        RECT 50.130 235.800 50.480 236.400 ;
        RECT 46.530 235.600 50.480 235.800 ;
        RECT 38.980 234.800 42.930 235.000 ;
        RECT 38.980 234.200 39.330 234.800 ;
        RECT 38.980 234.000 42.930 234.200 ;
        RECT 38.980 233.400 39.330 234.000 ;
        RECT 38.980 233.200 42.930 233.400 ;
        RECT 43.880 233.250 45.580 235.550 ;
        RECT 50.130 235.000 50.480 235.600 ;
        RECT 46.530 234.800 50.480 235.000 ;
        RECT 50.130 234.200 50.480 234.800 ;
        RECT 46.530 234.000 50.480 234.200 ;
        RECT 50.130 233.400 50.480 234.000 ;
        RECT 38.980 232.600 39.330 233.200 ;
        RECT 38.980 232.400 42.930 232.600 ;
        RECT 38.980 231.800 39.330 232.400 ;
        RECT 38.980 231.600 42.930 231.800 ;
        RECT 38.980 231.000 39.330 231.600 ;
        RECT 38.980 230.800 42.930 231.000 ;
        RECT 38.980 230.400 39.330 230.800 ;
        RECT 35.780 222.000 35.980 229.600 ;
        RECT 36.580 222.000 36.780 229.600 ;
        RECT 37.380 222.000 37.580 229.600 ;
        RECT 38.180 222.000 38.380 229.600 ;
        RECT 38.980 229.200 39.330 229.600 ;
        RECT 38.980 229.000 42.930 229.200 ;
        RECT 38.980 228.400 39.330 229.000 ;
        RECT 38.980 228.200 42.930 228.400 ;
        RECT 38.980 227.600 39.330 228.200 ;
        RECT 38.980 227.400 42.930 227.600 ;
        RECT 38.980 226.800 39.330 227.400 ;
        RECT 38.980 226.600 42.930 226.800 ;
        RECT 43.930 226.750 44.330 233.250 ;
        RECT 45.130 226.750 45.530 233.250 ;
        RECT 46.530 233.200 50.480 233.400 ;
        RECT 50.130 232.600 50.480 233.200 ;
        RECT 46.530 232.400 50.480 232.600 ;
        RECT 50.130 231.800 50.480 232.400 ;
        RECT 46.530 231.600 50.480 231.800 ;
        RECT 50.130 231.000 50.480 231.600 ;
        RECT 46.530 230.800 50.480 231.000 ;
        RECT 50.130 230.400 50.480 230.800 ;
        RECT 51.080 230.400 51.280 238.000 ;
        RECT 51.880 230.400 52.080 238.000 ;
        RECT 52.680 230.400 52.880 238.000 ;
        RECT 53.480 230.400 53.680 238.000 ;
        RECT 50.130 229.200 50.480 229.600 ;
        RECT 46.530 229.000 50.480 229.200 ;
        RECT 50.130 228.400 50.480 229.000 ;
        RECT 46.530 228.200 50.480 228.400 ;
        RECT 50.130 227.600 50.480 228.200 ;
        RECT 46.530 227.400 50.480 227.600 ;
        RECT 50.130 226.800 50.480 227.400 ;
        RECT 38.980 226.000 39.330 226.600 ;
        RECT 38.980 225.800 42.930 226.000 ;
        RECT 38.980 225.200 39.330 225.800 ;
        RECT 38.980 225.000 42.930 225.200 ;
        RECT 38.980 224.400 39.330 225.000 ;
        RECT 43.880 224.450 45.580 226.750 ;
        RECT 46.530 226.600 50.480 226.800 ;
        RECT 50.130 226.000 50.480 226.600 ;
        RECT 46.530 225.800 50.480 226.000 ;
        RECT 50.130 225.200 50.480 225.800 ;
        RECT 46.530 225.000 50.480 225.200 ;
        RECT 38.980 224.200 42.930 224.400 ;
        RECT 38.980 223.600 39.330 224.200 ;
        RECT 38.980 223.400 42.930 223.600 ;
        RECT 38.980 222.800 39.330 223.400 ;
        RECT 38.980 222.600 42.930 222.800 ;
        RECT 38.980 222.000 39.330 222.600 ;
        RECT 26.530 221.400 42.930 222.000 ;
        RECT 29.180 220.800 31.480 220.850 ;
        RECT 37.980 220.800 40.280 220.850 ;
        RECT 43.930 220.800 44.330 224.450 ;
        RECT 25.130 220.400 44.330 220.800 ;
        RECT 45.130 220.800 45.530 224.450 ;
        RECT 50.130 224.400 50.480 225.000 ;
        RECT 46.530 224.200 50.480 224.400 ;
        RECT 50.130 223.600 50.480 224.200 ;
        RECT 46.530 223.400 50.480 223.600 ;
        RECT 50.130 222.800 50.480 223.400 ;
        RECT 46.530 222.600 50.480 222.800 ;
        RECT 50.130 222.000 50.480 222.600 ;
        RECT 51.080 222.000 51.280 229.600 ;
        RECT 51.880 222.000 52.080 229.600 ;
        RECT 52.680 222.000 52.880 229.600 ;
        RECT 53.480 222.000 53.680 229.600 ;
        RECT 54.280 222.000 55.180 238.000 ;
        RECT 55.780 230.400 55.980 238.000 ;
        RECT 56.580 230.400 56.780 238.000 ;
        RECT 57.380 230.400 57.580 238.000 ;
        RECT 58.180 230.400 58.380 238.000 ;
        RECT 58.980 237.400 59.330 238.000 ;
        RECT 58.980 237.200 62.930 237.400 ;
        RECT 58.980 236.600 59.330 237.200 ;
        RECT 58.980 236.400 62.930 236.600 ;
        RECT 58.980 235.800 59.330 236.400 ;
        RECT 58.980 235.600 62.930 235.800 ;
        RECT 58.980 235.000 59.330 235.600 ;
        RECT 63.930 235.550 64.330 239.200 ;
        RECT 65.130 239.200 84.330 239.600 ;
        RECT 65.130 235.550 65.530 239.200 ;
        RECT 69.180 239.150 71.480 239.200 ;
        RECT 77.980 239.150 80.280 239.200 ;
        RECT 66.530 238.000 82.930 238.600 ;
        RECT 70.130 237.400 70.480 238.000 ;
        RECT 66.530 237.200 70.480 237.400 ;
        RECT 70.130 236.600 70.480 237.200 ;
        RECT 66.530 236.400 70.480 236.600 ;
        RECT 70.130 235.800 70.480 236.400 ;
        RECT 66.530 235.600 70.480 235.800 ;
        RECT 58.980 234.800 62.930 235.000 ;
        RECT 58.980 234.200 59.330 234.800 ;
        RECT 58.980 234.000 62.930 234.200 ;
        RECT 58.980 233.400 59.330 234.000 ;
        RECT 58.980 233.200 62.930 233.400 ;
        RECT 63.880 233.250 65.580 235.550 ;
        RECT 70.130 235.000 70.480 235.600 ;
        RECT 66.530 234.800 70.480 235.000 ;
        RECT 70.130 234.200 70.480 234.800 ;
        RECT 66.530 234.000 70.480 234.200 ;
        RECT 70.130 233.400 70.480 234.000 ;
        RECT 58.980 232.600 59.330 233.200 ;
        RECT 58.980 232.400 62.930 232.600 ;
        RECT 58.980 231.800 59.330 232.400 ;
        RECT 58.980 231.600 62.930 231.800 ;
        RECT 58.980 231.000 59.330 231.600 ;
        RECT 58.980 230.800 62.930 231.000 ;
        RECT 58.980 230.400 59.330 230.800 ;
        RECT 55.780 222.000 55.980 229.600 ;
        RECT 56.580 222.000 56.780 229.600 ;
        RECT 57.380 222.000 57.580 229.600 ;
        RECT 58.180 222.000 58.380 229.600 ;
        RECT 58.980 229.200 59.330 229.600 ;
        RECT 58.980 229.000 62.930 229.200 ;
        RECT 58.980 228.400 59.330 229.000 ;
        RECT 58.980 228.200 62.930 228.400 ;
        RECT 58.980 227.600 59.330 228.200 ;
        RECT 58.980 227.400 62.930 227.600 ;
        RECT 58.980 226.800 59.330 227.400 ;
        RECT 58.980 226.600 62.930 226.800 ;
        RECT 63.930 226.750 64.330 233.250 ;
        RECT 65.130 226.750 65.530 233.250 ;
        RECT 66.530 233.200 70.480 233.400 ;
        RECT 70.130 232.600 70.480 233.200 ;
        RECT 66.530 232.400 70.480 232.600 ;
        RECT 70.130 231.800 70.480 232.400 ;
        RECT 66.530 231.600 70.480 231.800 ;
        RECT 70.130 231.000 70.480 231.600 ;
        RECT 66.530 230.800 70.480 231.000 ;
        RECT 70.130 230.400 70.480 230.800 ;
        RECT 71.080 230.400 71.280 238.000 ;
        RECT 71.880 230.400 72.080 238.000 ;
        RECT 72.680 230.400 72.880 238.000 ;
        RECT 73.480 230.400 73.680 238.000 ;
        RECT 70.130 229.200 70.480 229.600 ;
        RECT 66.530 229.000 70.480 229.200 ;
        RECT 70.130 228.400 70.480 229.000 ;
        RECT 66.530 228.200 70.480 228.400 ;
        RECT 70.130 227.600 70.480 228.200 ;
        RECT 66.530 227.400 70.480 227.600 ;
        RECT 70.130 226.800 70.480 227.400 ;
        RECT 58.980 226.000 59.330 226.600 ;
        RECT 58.980 225.800 62.930 226.000 ;
        RECT 58.980 225.200 59.330 225.800 ;
        RECT 58.980 225.000 62.930 225.200 ;
        RECT 58.980 224.400 59.330 225.000 ;
        RECT 63.880 224.450 65.580 226.750 ;
        RECT 66.530 226.600 70.480 226.800 ;
        RECT 70.130 226.000 70.480 226.600 ;
        RECT 66.530 225.800 70.480 226.000 ;
        RECT 70.130 225.200 70.480 225.800 ;
        RECT 66.530 225.000 70.480 225.200 ;
        RECT 58.980 224.200 62.930 224.400 ;
        RECT 58.980 223.600 59.330 224.200 ;
        RECT 58.980 223.400 62.930 223.600 ;
        RECT 58.980 222.800 59.330 223.400 ;
        RECT 58.980 222.600 62.930 222.800 ;
        RECT 58.980 222.000 59.330 222.600 ;
        RECT 46.530 221.400 62.930 222.000 ;
        RECT 49.180 220.800 51.480 220.850 ;
        RECT 57.980 220.800 60.280 220.850 ;
        RECT 63.930 220.800 64.330 224.450 ;
        RECT 45.130 220.400 64.330 220.800 ;
        RECT 65.130 220.800 65.530 224.450 ;
        RECT 70.130 224.400 70.480 225.000 ;
        RECT 66.530 224.200 70.480 224.400 ;
        RECT 70.130 223.600 70.480 224.200 ;
        RECT 66.530 223.400 70.480 223.600 ;
        RECT 70.130 222.800 70.480 223.400 ;
        RECT 66.530 222.600 70.480 222.800 ;
        RECT 70.130 222.000 70.480 222.600 ;
        RECT 71.080 222.000 71.280 229.600 ;
        RECT 71.880 222.000 72.080 229.600 ;
        RECT 72.680 222.000 72.880 229.600 ;
        RECT 73.480 222.000 73.680 229.600 ;
        RECT 74.280 222.000 75.180 238.000 ;
        RECT 75.780 230.400 75.980 238.000 ;
        RECT 76.580 230.400 76.780 238.000 ;
        RECT 77.380 230.400 77.580 238.000 ;
        RECT 78.180 230.400 78.380 238.000 ;
        RECT 78.980 237.400 79.330 238.000 ;
        RECT 78.980 237.200 82.930 237.400 ;
        RECT 78.980 236.600 79.330 237.200 ;
        RECT 78.980 236.400 82.930 236.600 ;
        RECT 78.980 235.800 79.330 236.400 ;
        RECT 78.980 235.600 82.930 235.800 ;
        RECT 78.980 235.000 79.330 235.600 ;
        RECT 83.930 235.550 84.330 239.200 ;
        RECT 85.130 239.200 104.330 239.600 ;
        RECT 85.130 235.550 85.530 239.200 ;
        RECT 89.180 239.150 91.480 239.200 ;
        RECT 97.980 239.150 100.280 239.200 ;
        RECT 86.530 238.000 102.930 238.600 ;
        RECT 90.130 237.400 90.480 238.000 ;
        RECT 86.530 237.200 90.480 237.400 ;
        RECT 90.130 236.600 90.480 237.200 ;
        RECT 86.530 236.400 90.480 236.600 ;
        RECT 90.130 235.800 90.480 236.400 ;
        RECT 86.530 235.600 90.480 235.800 ;
        RECT 78.980 234.800 82.930 235.000 ;
        RECT 78.980 234.200 79.330 234.800 ;
        RECT 78.980 234.000 82.930 234.200 ;
        RECT 78.980 233.400 79.330 234.000 ;
        RECT 78.980 233.200 82.930 233.400 ;
        RECT 83.880 233.250 85.580 235.550 ;
        RECT 90.130 235.000 90.480 235.600 ;
        RECT 86.530 234.800 90.480 235.000 ;
        RECT 90.130 234.200 90.480 234.800 ;
        RECT 86.530 234.000 90.480 234.200 ;
        RECT 90.130 233.400 90.480 234.000 ;
        RECT 78.980 232.600 79.330 233.200 ;
        RECT 78.980 232.400 82.930 232.600 ;
        RECT 78.980 231.800 79.330 232.400 ;
        RECT 78.980 231.600 82.930 231.800 ;
        RECT 78.980 231.000 79.330 231.600 ;
        RECT 78.980 230.800 82.930 231.000 ;
        RECT 78.980 230.400 79.330 230.800 ;
        RECT 75.780 222.000 75.980 229.600 ;
        RECT 76.580 222.000 76.780 229.600 ;
        RECT 77.380 222.000 77.580 229.600 ;
        RECT 78.180 222.000 78.380 229.600 ;
        RECT 78.980 229.200 79.330 229.600 ;
        RECT 78.980 229.000 82.930 229.200 ;
        RECT 78.980 228.400 79.330 229.000 ;
        RECT 78.980 228.200 82.930 228.400 ;
        RECT 78.980 227.600 79.330 228.200 ;
        RECT 78.980 227.400 82.930 227.600 ;
        RECT 78.980 226.800 79.330 227.400 ;
        RECT 78.980 226.600 82.930 226.800 ;
        RECT 83.930 226.750 84.330 233.250 ;
        RECT 85.130 226.750 85.530 233.250 ;
        RECT 86.530 233.200 90.480 233.400 ;
        RECT 90.130 232.600 90.480 233.200 ;
        RECT 86.530 232.400 90.480 232.600 ;
        RECT 90.130 231.800 90.480 232.400 ;
        RECT 86.530 231.600 90.480 231.800 ;
        RECT 90.130 231.000 90.480 231.600 ;
        RECT 86.530 230.800 90.480 231.000 ;
        RECT 90.130 230.400 90.480 230.800 ;
        RECT 91.080 230.400 91.280 238.000 ;
        RECT 91.880 230.400 92.080 238.000 ;
        RECT 92.680 230.400 92.880 238.000 ;
        RECT 93.480 230.400 93.680 238.000 ;
        RECT 90.130 229.200 90.480 229.600 ;
        RECT 86.530 229.000 90.480 229.200 ;
        RECT 90.130 228.400 90.480 229.000 ;
        RECT 86.530 228.200 90.480 228.400 ;
        RECT 90.130 227.600 90.480 228.200 ;
        RECT 86.530 227.400 90.480 227.600 ;
        RECT 90.130 226.800 90.480 227.400 ;
        RECT 78.980 226.000 79.330 226.600 ;
        RECT 78.980 225.800 82.930 226.000 ;
        RECT 78.980 225.200 79.330 225.800 ;
        RECT 78.980 225.000 82.930 225.200 ;
        RECT 78.980 224.400 79.330 225.000 ;
        RECT 83.880 224.450 85.580 226.750 ;
        RECT 86.530 226.600 90.480 226.800 ;
        RECT 90.130 226.000 90.480 226.600 ;
        RECT 86.530 225.800 90.480 226.000 ;
        RECT 90.130 225.200 90.480 225.800 ;
        RECT 86.530 225.000 90.480 225.200 ;
        RECT 78.980 224.200 82.930 224.400 ;
        RECT 78.980 223.600 79.330 224.200 ;
        RECT 78.980 223.400 82.930 223.600 ;
        RECT 78.980 222.800 79.330 223.400 ;
        RECT 78.980 222.600 82.930 222.800 ;
        RECT 78.980 222.000 79.330 222.600 ;
        RECT 66.530 221.400 82.930 222.000 ;
        RECT 69.180 220.800 71.480 220.850 ;
        RECT 77.980 220.800 80.280 220.850 ;
        RECT 83.930 220.800 84.330 224.450 ;
        RECT 65.130 220.400 84.330 220.800 ;
        RECT 85.130 220.800 85.530 224.450 ;
        RECT 90.130 224.400 90.480 225.000 ;
        RECT 86.530 224.200 90.480 224.400 ;
        RECT 90.130 223.600 90.480 224.200 ;
        RECT 86.530 223.400 90.480 223.600 ;
        RECT 90.130 222.800 90.480 223.400 ;
        RECT 86.530 222.600 90.480 222.800 ;
        RECT 90.130 222.000 90.480 222.600 ;
        RECT 91.080 222.000 91.280 229.600 ;
        RECT 91.880 222.000 92.080 229.600 ;
        RECT 92.680 222.000 92.880 229.600 ;
        RECT 93.480 222.000 93.680 229.600 ;
        RECT 94.280 222.000 95.180 238.000 ;
        RECT 95.780 230.400 95.980 238.000 ;
        RECT 96.580 230.400 96.780 238.000 ;
        RECT 97.380 230.400 97.580 238.000 ;
        RECT 98.180 230.400 98.380 238.000 ;
        RECT 98.980 237.400 99.330 238.000 ;
        RECT 98.980 237.200 102.930 237.400 ;
        RECT 98.980 236.600 99.330 237.200 ;
        RECT 98.980 236.400 102.930 236.600 ;
        RECT 98.980 235.800 99.330 236.400 ;
        RECT 98.980 235.600 102.930 235.800 ;
        RECT 98.980 235.000 99.330 235.600 ;
        RECT 103.930 235.550 104.330 239.200 ;
        RECT 105.130 239.200 124.330 239.600 ;
        RECT 105.130 235.550 105.530 239.200 ;
        RECT 109.180 239.150 111.480 239.200 ;
        RECT 117.980 239.150 120.280 239.200 ;
        RECT 106.530 238.000 122.930 238.600 ;
        RECT 110.130 237.400 110.480 238.000 ;
        RECT 106.530 237.200 110.480 237.400 ;
        RECT 110.130 236.600 110.480 237.200 ;
        RECT 106.530 236.400 110.480 236.600 ;
        RECT 110.130 235.800 110.480 236.400 ;
        RECT 106.530 235.600 110.480 235.800 ;
        RECT 98.980 234.800 102.930 235.000 ;
        RECT 98.980 234.200 99.330 234.800 ;
        RECT 98.980 234.000 102.930 234.200 ;
        RECT 98.980 233.400 99.330 234.000 ;
        RECT 98.980 233.200 102.930 233.400 ;
        RECT 103.880 233.250 105.580 235.550 ;
        RECT 110.130 235.000 110.480 235.600 ;
        RECT 106.530 234.800 110.480 235.000 ;
        RECT 110.130 234.200 110.480 234.800 ;
        RECT 106.530 234.000 110.480 234.200 ;
        RECT 110.130 233.400 110.480 234.000 ;
        RECT 98.980 232.600 99.330 233.200 ;
        RECT 98.980 232.400 102.930 232.600 ;
        RECT 98.980 231.800 99.330 232.400 ;
        RECT 98.980 231.600 102.930 231.800 ;
        RECT 98.980 231.000 99.330 231.600 ;
        RECT 98.980 230.800 102.930 231.000 ;
        RECT 98.980 230.400 99.330 230.800 ;
        RECT 95.780 222.000 95.980 229.600 ;
        RECT 96.580 222.000 96.780 229.600 ;
        RECT 97.380 222.000 97.580 229.600 ;
        RECT 98.180 222.000 98.380 229.600 ;
        RECT 98.980 229.200 99.330 229.600 ;
        RECT 98.980 229.000 102.930 229.200 ;
        RECT 98.980 228.400 99.330 229.000 ;
        RECT 98.980 228.200 102.930 228.400 ;
        RECT 98.980 227.600 99.330 228.200 ;
        RECT 98.980 227.400 102.930 227.600 ;
        RECT 98.980 226.800 99.330 227.400 ;
        RECT 98.980 226.600 102.930 226.800 ;
        RECT 103.930 226.750 104.330 233.250 ;
        RECT 105.130 226.750 105.530 233.250 ;
        RECT 106.530 233.200 110.480 233.400 ;
        RECT 110.130 232.600 110.480 233.200 ;
        RECT 106.530 232.400 110.480 232.600 ;
        RECT 110.130 231.800 110.480 232.400 ;
        RECT 106.530 231.600 110.480 231.800 ;
        RECT 110.130 231.000 110.480 231.600 ;
        RECT 106.530 230.800 110.480 231.000 ;
        RECT 110.130 230.400 110.480 230.800 ;
        RECT 111.080 230.400 111.280 238.000 ;
        RECT 111.880 230.400 112.080 238.000 ;
        RECT 112.680 230.400 112.880 238.000 ;
        RECT 113.480 230.400 113.680 238.000 ;
        RECT 110.130 229.200 110.480 229.600 ;
        RECT 106.530 229.000 110.480 229.200 ;
        RECT 110.130 228.400 110.480 229.000 ;
        RECT 106.530 228.200 110.480 228.400 ;
        RECT 110.130 227.600 110.480 228.200 ;
        RECT 106.530 227.400 110.480 227.600 ;
        RECT 110.130 226.800 110.480 227.400 ;
        RECT 98.980 226.000 99.330 226.600 ;
        RECT 98.980 225.800 102.930 226.000 ;
        RECT 98.980 225.200 99.330 225.800 ;
        RECT 98.980 225.000 102.930 225.200 ;
        RECT 98.980 224.400 99.330 225.000 ;
        RECT 103.880 224.450 105.580 226.750 ;
        RECT 106.530 226.600 110.480 226.800 ;
        RECT 110.130 226.000 110.480 226.600 ;
        RECT 106.530 225.800 110.480 226.000 ;
        RECT 110.130 225.200 110.480 225.800 ;
        RECT 106.530 225.000 110.480 225.200 ;
        RECT 98.980 224.200 102.930 224.400 ;
        RECT 98.980 223.600 99.330 224.200 ;
        RECT 98.980 223.400 102.930 223.600 ;
        RECT 98.980 222.800 99.330 223.400 ;
        RECT 98.980 222.600 102.930 222.800 ;
        RECT 98.980 222.000 99.330 222.600 ;
        RECT 86.530 221.400 102.930 222.000 ;
        RECT 89.180 220.800 91.480 220.850 ;
        RECT 97.980 220.800 100.280 220.850 ;
        RECT 103.930 220.800 104.330 224.450 ;
        RECT 85.130 220.400 104.330 220.800 ;
        RECT 105.130 220.800 105.530 224.450 ;
        RECT 110.130 224.400 110.480 225.000 ;
        RECT 106.530 224.200 110.480 224.400 ;
        RECT 110.130 223.600 110.480 224.200 ;
        RECT 106.530 223.400 110.480 223.600 ;
        RECT 110.130 222.800 110.480 223.400 ;
        RECT 106.530 222.600 110.480 222.800 ;
        RECT 110.130 222.000 110.480 222.600 ;
        RECT 111.080 222.000 111.280 229.600 ;
        RECT 111.880 222.000 112.080 229.600 ;
        RECT 112.680 222.000 112.880 229.600 ;
        RECT 113.480 222.000 113.680 229.600 ;
        RECT 114.280 222.000 115.180 238.000 ;
        RECT 115.780 230.400 115.980 238.000 ;
        RECT 116.580 230.400 116.780 238.000 ;
        RECT 117.380 230.400 117.580 238.000 ;
        RECT 118.180 230.400 118.380 238.000 ;
        RECT 118.980 237.400 119.330 238.000 ;
        RECT 118.980 237.200 122.930 237.400 ;
        RECT 118.980 236.600 119.330 237.200 ;
        RECT 118.980 236.400 122.930 236.600 ;
        RECT 118.980 235.800 119.330 236.400 ;
        RECT 118.980 235.600 122.930 235.800 ;
        RECT 118.980 235.000 119.330 235.600 ;
        RECT 123.930 235.550 124.330 239.200 ;
        RECT 125.340 236.820 125.700 237.200 ;
        RECT 125.970 236.820 126.330 237.200 ;
        RECT 126.570 236.820 126.930 237.200 ;
        RECT 125.340 236.230 125.700 236.610 ;
        RECT 125.970 236.230 126.330 236.610 ;
        RECT 126.570 236.230 126.930 236.610 ;
        RECT 118.980 234.800 122.930 235.000 ;
        RECT 118.980 234.200 119.330 234.800 ;
        RECT 118.980 234.000 122.930 234.200 ;
        RECT 118.980 233.400 119.330 234.000 ;
        RECT 118.980 233.200 122.930 233.400 ;
        RECT 123.880 233.250 124.730 235.550 ;
        RECT 118.980 232.600 119.330 233.200 ;
        RECT 118.980 232.400 122.930 232.600 ;
        RECT 118.980 231.800 119.330 232.400 ;
        RECT 118.980 231.600 122.930 231.800 ;
        RECT 118.980 231.000 119.330 231.600 ;
        RECT 118.980 230.800 122.930 231.000 ;
        RECT 118.980 230.400 119.330 230.800 ;
        RECT 115.780 222.000 115.980 229.600 ;
        RECT 116.580 222.000 116.780 229.600 ;
        RECT 117.380 222.000 117.580 229.600 ;
        RECT 118.180 222.000 118.380 229.600 ;
        RECT 118.980 229.200 119.330 229.600 ;
        RECT 118.980 229.000 122.930 229.200 ;
        RECT 118.980 228.400 119.330 229.000 ;
        RECT 118.980 228.200 122.930 228.400 ;
        RECT 118.980 227.600 119.330 228.200 ;
        RECT 118.980 227.400 122.930 227.600 ;
        RECT 118.980 226.800 119.330 227.400 ;
        RECT 118.980 226.600 122.930 226.800 ;
        RECT 123.930 226.750 124.330 233.250 ;
        RECT 118.980 226.000 119.330 226.600 ;
        RECT 118.980 225.800 122.930 226.000 ;
        RECT 118.980 225.200 119.330 225.800 ;
        RECT 118.980 225.000 122.930 225.200 ;
        RECT 118.980 224.400 119.330 225.000 ;
        RECT 123.880 224.450 124.730 226.750 ;
        RECT 118.980 224.200 122.930 224.400 ;
        RECT 118.980 223.600 119.330 224.200 ;
        RECT 118.980 223.400 122.930 223.600 ;
        RECT 118.980 222.800 119.330 223.400 ;
        RECT 118.980 222.600 122.930 222.800 ;
        RECT 118.980 222.000 119.330 222.600 ;
        RECT 106.530 221.400 122.930 222.000 ;
        RECT 109.180 220.800 111.480 220.850 ;
        RECT 117.980 220.800 120.280 220.850 ;
        RECT 123.930 220.800 124.330 224.450 ;
        RECT 125.340 223.025 125.700 223.405 ;
        RECT 125.970 223.025 126.330 223.405 ;
        RECT 126.570 223.025 126.930 223.405 ;
        RECT 125.340 222.435 125.700 222.815 ;
        RECT 125.970 222.435 126.330 222.815 ;
        RECT 126.570 222.435 126.930 222.815 ;
        RECT 105.130 220.400 124.330 220.800 ;
        RECT 9.180 219.600 11.480 220.400 ;
        RECT 17.980 219.600 20.280 220.400 ;
        RECT 29.180 219.600 31.480 220.400 ;
        RECT 37.980 219.600 40.280 220.400 ;
        RECT 49.180 219.600 51.480 220.400 ;
        RECT 57.980 219.600 60.280 220.400 ;
        RECT 69.180 219.600 71.480 220.400 ;
        RECT 77.980 219.600 80.280 220.400 ;
        RECT 89.180 219.600 91.480 220.400 ;
        RECT 97.980 219.600 100.280 220.400 ;
        RECT 109.180 219.600 111.480 220.400 ;
        RECT 117.980 219.600 120.280 220.400 ;
        RECT 5.130 219.200 24.330 219.600 ;
        RECT 2.515 217.465 2.875 217.845 ;
        RECT 3.145 217.465 3.505 217.845 ;
        RECT 3.745 217.465 4.105 217.845 ;
        RECT 2.515 216.875 2.875 217.255 ;
        RECT 3.145 216.875 3.505 217.255 ;
        RECT 3.745 216.875 4.105 217.255 ;
        RECT 5.130 215.550 5.530 219.200 ;
        RECT 9.180 219.150 11.480 219.200 ;
        RECT 17.980 219.150 20.280 219.200 ;
        RECT 6.530 218.000 22.930 218.600 ;
        RECT 10.130 217.400 10.480 218.000 ;
        RECT 6.530 217.200 10.480 217.400 ;
        RECT 10.130 216.600 10.480 217.200 ;
        RECT 6.530 216.400 10.480 216.600 ;
        RECT 10.130 215.800 10.480 216.400 ;
        RECT 6.530 215.600 10.480 215.800 ;
        RECT 4.730 215.545 5.580 215.550 ;
        RECT 2.315 213.250 5.580 215.545 ;
        RECT 10.130 215.000 10.480 215.600 ;
        RECT 6.530 214.800 10.480 215.000 ;
        RECT 10.130 214.200 10.480 214.800 ;
        RECT 6.530 214.000 10.480 214.200 ;
        RECT 10.130 213.400 10.480 214.000 ;
        RECT 5.130 206.750 5.530 213.250 ;
        RECT 6.530 213.200 10.480 213.400 ;
        RECT 10.130 212.600 10.480 213.200 ;
        RECT 6.530 212.400 10.480 212.600 ;
        RECT 10.130 211.800 10.480 212.400 ;
        RECT 6.530 211.600 10.480 211.800 ;
        RECT 10.130 211.000 10.480 211.600 ;
        RECT 6.530 210.800 10.480 211.000 ;
        RECT 10.130 210.400 10.480 210.800 ;
        RECT 11.080 210.400 11.280 218.000 ;
        RECT 11.880 210.400 12.080 218.000 ;
        RECT 12.680 210.400 12.880 218.000 ;
        RECT 13.480 210.400 13.680 218.000 ;
        RECT 10.130 209.200 10.480 209.600 ;
        RECT 6.530 209.000 10.480 209.200 ;
        RECT 10.130 208.400 10.480 209.000 ;
        RECT 6.530 208.200 10.480 208.400 ;
        RECT 10.130 207.600 10.480 208.200 ;
        RECT 6.530 207.400 10.480 207.600 ;
        RECT 10.130 206.800 10.480 207.400 ;
        RECT 2.315 204.455 5.580 206.750 ;
        RECT 6.530 206.600 10.480 206.800 ;
        RECT 10.130 206.000 10.480 206.600 ;
        RECT 6.530 205.800 10.480 206.000 ;
        RECT 10.130 205.200 10.480 205.800 ;
        RECT 6.530 205.000 10.480 205.200 ;
        RECT 2.315 204.450 4.180 204.455 ;
        RECT 4.730 204.450 5.580 204.455 ;
        RECT 2.515 202.165 2.875 202.545 ;
        RECT 3.145 202.165 3.505 202.545 ;
        RECT 3.745 202.165 4.105 202.545 ;
        RECT 2.515 201.575 2.875 201.955 ;
        RECT 3.145 201.575 3.505 201.955 ;
        RECT 3.745 201.575 4.105 201.955 ;
        RECT 5.130 200.800 5.530 204.450 ;
        RECT 10.130 204.400 10.480 205.000 ;
        RECT 6.530 204.200 10.480 204.400 ;
        RECT 10.130 203.600 10.480 204.200 ;
        RECT 6.530 203.400 10.480 203.600 ;
        RECT 10.130 202.800 10.480 203.400 ;
        RECT 6.530 202.600 10.480 202.800 ;
        RECT 10.130 202.000 10.480 202.600 ;
        RECT 11.080 202.000 11.280 209.600 ;
        RECT 11.880 202.000 12.080 209.600 ;
        RECT 12.680 202.000 12.880 209.600 ;
        RECT 13.480 202.000 13.680 209.600 ;
        RECT 14.280 202.000 15.180 218.000 ;
        RECT 15.780 210.400 15.980 218.000 ;
        RECT 16.580 210.400 16.780 218.000 ;
        RECT 17.380 210.400 17.580 218.000 ;
        RECT 18.180 210.400 18.380 218.000 ;
        RECT 18.980 217.400 19.330 218.000 ;
        RECT 18.980 217.200 22.930 217.400 ;
        RECT 18.980 216.600 19.330 217.200 ;
        RECT 18.980 216.400 22.930 216.600 ;
        RECT 18.980 215.800 19.330 216.400 ;
        RECT 18.980 215.600 22.930 215.800 ;
        RECT 18.980 215.000 19.330 215.600 ;
        RECT 23.930 215.550 24.330 219.200 ;
        RECT 25.130 219.200 44.330 219.600 ;
        RECT 25.130 215.550 25.530 219.200 ;
        RECT 29.180 219.150 31.480 219.200 ;
        RECT 37.980 219.150 40.280 219.200 ;
        RECT 26.530 218.000 42.930 218.600 ;
        RECT 30.130 217.400 30.480 218.000 ;
        RECT 26.530 217.200 30.480 217.400 ;
        RECT 30.130 216.600 30.480 217.200 ;
        RECT 26.530 216.400 30.480 216.600 ;
        RECT 30.130 215.800 30.480 216.400 ;
        RECT 26.530 215.600 30.480 215.800 ;
        RECT 18.980 214.800 22.930 215.000 ;
        RECT 18.980 214.200 19.330 214.800 ;
        RECT 18.980 214.000 22.930 214.200 ;
        RECT 18.980 213.400 19.330 214.000 ;
        RECT 18.980 213.200 22.930 213.400 ;
        RECT 23.880 213.250 25.580 215.550 ;
        RECT 30.130 215.000 30.480 215.600 ;
        RECT 26.530 214.800 30.480 215.000 ;
        RECT 30.130 214.200 30.480 214.800 ;
        RECT 26.530 214.000 30.480 214.200 ;
        RECT 30.130 213.400 30.480 214.000 ;
        RECT 18.980 212.600 19.330 213.200 ;
        RECT 18.980 212.400 22.930 212.600 ;
        RECT 18.980 211.800 19.330 212.400 ;
        RECT 18.980 211.600 22.930 211.800 ;
        RECT 18.980 211.000 19.330 211.600 ;
        RECT 18.980 210.800 22.930 211.000 ;
        RECT 18.980 210.400 19.330 210.800 ;
        RECT 15.780 202.000 15.980 209.600 ;
        RECT 16.580 202.000 16.780 209.600 ;
        RECT 17.380 202.000 17.580 209.600 ;
        RECT 18.180 202.000 18.380 209.600 ;
        RECT 18.980 209.200 19.330 209.600 ;
        RECT 18.980 209.000 22.930 209.200 ;
        RECT 18.980 208.400 19.330 209.000 ;
        RECT 18.980 208.200 22.930 208.400 ;
        RECT 18.980 207.600 19.330 208.200 ;
        RECT 18.980 207.400 22.930 207.600 ;
        RECT 18.980 206.800 19.330 207.400 ;
        RECT 18.980 206.600 22.930 206.800 ;
        RECT 23.930 206.750 24.330 213.250 ;
        RECT 25.130 206.750 25.530 213.250 ;
        RECT 26.530 213.200 30.480 213.400 ;
        RECT 30.130 212.600 30.480 213.200 ;
        RECT 26.530 212.400 30.480 212.600 ;
        RECT 30.130 211.800 30.480 212.400 ;
        RECT 26.530 211.600 30.480 211.800 ;
        RECT 30.130 211.000 30.480 211.600 ;
        RECT 26.530 210.800 30.480 211.000 ;
        RECT 30.130 210.400 30.480 210.800 ;
        RECT 31.080 210.400 31.280 218.000 ;
        RECT 31.880 210.400 32.080 218.000 ;
        RECT 32.680 210.400 32.880 218.000 ;
        RECT 33.480 210.400 33.680 218.000 ;
        RECT 30.130 209.200 30.480 209.600 ;
        RECT 26.530 209.000 30.480 209.200 ;
        RECT 30.130 208.400 30.480 209.000 ;
        RECT 26.530 208.200 30.480 208.400 ;
        RECT 30.130 207.600 30.480 208.200 ;
        RECT 26.530 207.400 30.480 207.600 ;
        RECT 30.130 206.800 30.480 207.400 ;
        RECT 18.980 206.000 19.330 206.600 ;
        RECT 18.980 205.800 22.930 206.000 ;
        RECT 18.980 205.200 19.330 205.800 ;
        RECT 18.980 205.000 22.930 205.200 ;
        RECT 18.980 204.400 19.330 205.000 ;
        RECT 23.880 204.450 25.580 206.750 ;
        RECT 26.530 206.600 30.480 206.800 ;
        RECT 30.130 206.000 30.480 206.600 ;
        RECT 26.530 205.800 30.480 206.000 ;
        RECT 30.130 205.200 30.480 205.800 ;
        RECT 26.530 205.000 30.480 205.200 ;
        RECT 18.980 204.200 22.930 204.400 ;
        RECT 18.980 203.600 19.330 204.200 ;
        RECT 18.980 203.400 22.930 203.600 ;
        RECT 18.980 202.800 19.330 203.400 ;
        RECT 18.980 202.600 22.930 202.800 ;
        RECT 18.980 202.000 19.330 202.600 ;
        RECT 6.530 201.400 22.930 202.000 ;
        RECT 9.180 200.800 11.480 200.850 ;
        RECT 17.980 200.800 20.280 200.850 ;
        RECT 23.930 200.800 24.330 204.450 ;
        RECT 5.130 200.400 24.330 200.800 ;
        RECT 25.130 200.800 25.530 204.450 ;
        RECT 30.130 204.400 30.480 205.000 ;
        RECT 26.530 204.200 30.480 204.400 ;
        RECT 30.130 203.600 30.480 204.200 ;
        RECT 26.530 203.400 30.480 203.600 ;
        RECT 30.130 202.800 30.480 203.400 ;
        RECT 26.530 202.600 30.480 202.800 ;
        RECT 30.130 202.000 30.480 202.600 ;
        RECT 31.080 202.000 31.280 209.600 ;
        RECT 31.880 202.000 32.080 209.600 ;
        RECT 32.680 202.000 32.880 209.600 ;
        RECT 33.480 202.000 33.680 209.600 ;
        RECT 34.280 202.000 35.180 218.000 ;
        RECT 35.780 210.400 35.980 218.000 ;
        RECT 36.580 210.400 36.780 218.000 ;
        RECT 37.380 210.400 37.580 218.000 ;
        RECT 38.180 210.400 38.380 218.000 ;
        RECT 38.980 217.400 39.330 218.000 ;
        RECT 38.980 217.200 42.930 217.400 ;
        RECT 38.980 216.600 39.330 217.200 ;
        RECT 38.980 216.400 42.930 216.600 ;
        RECT 38.980 215.800 39.330 216.400 ;
        RECT 38.980 215.600 42.930 215.800 ;
        RECT 38.980 215.000 39.330 215.600 ;
        RECT 43.930 215.550 44.330 219.200 ;
        RECT 45.130 219.200 64.330 219.600 ;
        RECT 45.130 215.550 45.530 219.200 ;
        RECT 49.180 219.150 51.480 219.200 ;
        RECT 57.980 219.150 60.280 219.200 ;
        RECT 46.530 218.000 62.930 218.600 ;
        RECT 50.130 217.400 50.480 218.000 ;
        RECT 46.530 217.200 50.480 217.400 ;
        RECT 50.130 216.600 50.480 217.200 ;
        RECT 46.530 216.400 50.480 216.600 ;
        RECT 50.130 215.800 50.480 216.400 ;
        RECT 46.530 215.600 50.480 215.800 ;
        RECT 38.980 214.800 42.930 215.000 ;
        RECT 38.980 214.200 39.330 214.800 ;
        RECT 38.980 214.000 42.930 214.200 ;
        RECT 38.980 213.400 39.330 214.000 ;
        RECT 38.980 213.200 42.930 213.400 ;
        RECT 43.880 213.250 45.580 215.550 ;
        RECT 50.130 215.000 50.480 215.600 ;
        RECT 46.530 214.800 50.480 215.000 ;
        RECT 50.130 214.200 50.480 214.800 ;
        RECT 46.530 214.000 50.480 214.200 ;
        RECT 50.130 213.400 50.480 214.000 ;
        RECT 38.980 212.600 39.330 213.200 ;
        RECT 38.980 212.400 42.930 212.600 ;
        RECT 38.980 211.800 39.330 212.400 ;
        RECT 38.980 211.600 42.930 211.800 ;
        RECT 38.980 211.000 39.330 211.600 ;
        RECT 38.980 210.800 42.930 211.000 ;
        RECT 38.980 210.400 39.330 210.800 ;
        RECT 35.780 202.000 35.980 209.600 ;
        RECT 36.580 202.000 36.780 209.600 ;
        RECT 37.380 202.000 37.580 209.600 ;
        RECT 38.180 202.000 38.380 209.600 ;
        RECT 38.980 209.200 39.330 209.600 ;
        RECT 38.980 209.000 42.930 209.200 ;
        RECT 38.980 208.400 39.330 209.000 ;
        RECT 38.980 208.200 42.930 208.400 ;
        RECT 38.980 207.600 39.330 208.200 ;
        RECT 38.980 207.400 42.930 207.600 ;
        RECT 38.980 206.800 39.330 207.400 ;
        RECT 38.980 206.600 42.930 206.800 ;
        RECT 43.930 206.750 44.330 213.250 ;
        RECT 45.130 206.750 45.530 213.250 ;
        RECT 46.530 213.200 50.480 213.400 ;
        RECT 50.130 212.600 50.480 213.200 ;
        RECT 46.530 212.400 50.480 212.600 ;
        RECT 50.130 211.800 50.480 212.400 ;
        RECT 46.530 211.600 50.480 211.800 ;
        RECT 50.130 211.000 50.480 211.600 ;
        RECT 46.530 210.800 50.480 211.000 ;
        RECT 50.130 210.400 50.480 210.800 ;
        RECT 51.080 210.400 51.280 218.000 ;
        RECT 51.880 210.400 52.080 218.000 ;
        RECT 52.680 210.400 52.880 218.000 ;
        RECT 53.480 210.400 53.680 218.000 ;
        RECT 50.130 209.200 50.480 209.600 ;
        RECT 46.530 209.000 50.480 209.200 ;
        RECT 50.130 208.400 50.480 209.000 ;
        RECT 46.530 208.200 50.480 208.400 ;
        RECT 50.130 207.600 50.480 208.200 ;
        RECT 46.530 207.400 50.480 207.600 ;
        RECT 50.130 206.800 50.480 207.400 ;
        RECT 38.980 206.000 39.330 206.600 ;
        RECT 38.980 205.800 42.930 206.000 ;
        RECT 38.980 205.200 39.330 205.800 ;
        RECT 38.980 205.000 42.930 205.200 ;
        RECT 38.980 204.400 39.330 205.000 ;
        RECT 43.880 204.450 45.580 206.750 ;
        RECT 46.530 206.600 50.480 206.800 ;
        RECT 50.130 206.000 50.480 206.600 ;
        RECT 46.530 205.800 50.480 206.000 ;
        RECT 50.130 205.200 50.480 205.800 ;
        RECT 46.530 205.000 50.480 205.200 ;
        RECT 38.980 204.200 42.930 204.400 ;
        RECT 38.980 203.600 39.330 204.200 ;
        RECT 38.980 203.400 42.930 203.600 ;
        RECT 38.980 202.800 39.330 203.400 ;
        RECT 38.980 202.600 42.930 202.800 ;
        RECT 38.980 202.000 39.330 202.600 ;
        RECT 26.530 201.400 42.930 202.000 ;
        RECT 29.180 200.800 31.480 200.850 ;
        RECT 37.980 200.800 40.280 200.850 ;
        RECT 43.930 200.800 44.330 204.450 ;
        RECT 25.130 200.400 44.330 200.800 ;
        RECT 45.130 200.800 45.530 204.450 ;
        RECT 50.130 204.400 50.480 205.000 ;
        RECT 46.530 204.200 50.480 204.400 ;
        RECT 50.130 203.600 50.480 204.200 ;
        RECT 46.530 203.400 50.480 203.600 ;
        RECT 50.130 202.800 50.480 203.400 ;
        RECT 46.530 202.600 50.480 202.800 ;
        RECT 50.130 202.000 50.480 202.600 ;
        RECT 51.080 202.000 51.280 209.600 ;
        RECT 51.880 202.000 52.080 209.600 ;
        RECT 52.680 202.000 52.880 209.600 ;
        RECT 53.480 202.000 53.680 209.600 ;
        RECT 54.280 202.000 55.180 218.000 ;
        RECT 55.780 210.400 55.980 218.000 ;
        RECT 56.580 210.400 56.780 218.000 ;
        RECT 57.380 210.400 57.580 218.000 ;
        RECT 58.180 210.400 58.380 218.000 ;
        RECT 58.980 217.400 59.330 218.000 ;
        RECT 58.980 217.200 62.930 217.400 ;
        RECT 58.980 216.600 59.330 217.200 ;
        RECT 58.980 216.400 62.930 216.600 ;
        RECT 58.980 215.800 59.330 216.400 ;
        RECT 58.980 215.600 62.930 215.800 ;
        RECT 58.980 215.000 59.330 215.600 ;
        RECT 63.930 215.550 64.330 219.200 ;
        RECT 65.130 219.200 84.330 219.600 ;
        RECT 65.130 215.550 65.530 219.200 ;
        RECT 69.180 219.150 71.480 219.200 ;
        RECT 77.980 219.150 80.280 219.200 ;
        RECT 66.530 218.000 82.930 218.600 ;
        RECT 70.130 217.400 70.480 218.000 ;
        RECT 66.530 217.200 70.480 217.400 ;
        RECT 70.130 216.600 70.480 217.200 ;
        RECT 66.530 216.400 70.480 216.600 ;
        RECT 70.130 215.800 70.480 216.400 ;
        RECT 66.530 215.600 70.480 215.800 ;
        RECT 58.980 214.800 62.930 215.000 ;
        RECT 58.980 214.200 59.330 214.800 ;
        RECT 58.980 214.000 62.930 214.200 ;
        RECT 58.980 213.400 59.330 214.000 ;
        RECT 58.980 213.200 62.930 213.400 ;
        RECT 63.880 213.250 65.580 215.550 ;
        RECT 70.130 215.000 70.480 215.600 ;
        RECT 66.530 214.800 70.480 215.000 ;
        RECT 70.130 214.200 70.480 214.800 ;
        RECT 66.530 214.000 70.480 214.200 ;
        RECT 70.130 213.400 70.480 214.000 ;
        RECT 58.980 212.600 59.330 213.200 ;
        RECT 58.980 212.400 62.930 212.600 ;
        RECT 58.980 211.800 59.330 212.400 ;
        RECT 58.980 211.600 62.930 211.800 ;
        RECT 58.980 211.000 59.330 211.600 ;
        RECT 58.980 210.800 62.930 211.000 ;
        RECT 58.980 210.400 59.330 210.800 ;
        RECT 55.780 202.000 55.980 209.600 ;
        RECT 56.580 202.000 56.780 209.600 ;
        RECT 57.380 202.000 57.580 209.600 ;
        RECT 58.180 202.000 58.380 209.600 ;
        RECT 58.980 209.200 59.330 209.600 ;
        RECT 58.980 209.000 62.930 209.200 ;
        RECT 58.980 208.400 59.330 209.000 ;
        RECT 58.980 208.200 62.930 208.400 ;
        RECT 58.980 207.600 59.330 208.200 ;
        RECT 58.980 207.400 62.930 207.600 ;
        RECT 58.980 206.800 59.330 207.400 ;
        RECT 58.980 206.600 62.930 206.800 ;
        RECT 63.930 206.750 64.330 213.250 ;
        RECT 65.130 206.750 65.530 213.250 ;
        RECT 66.530 213.200 70.480 213.400 ;
        RECT 70.130 212.600 70.480 213.200 ;
        RECT 66.530 212.400 70.480 212.600 ;
        RECT 70.130 211.800 70.480 212.400 ;
        RECT 66.530 211.600 70.480 211.800 ;
        RECT 70.130 211.000 70.480 211.600 ;
        RECT 66.530 210.800 70.480 211.000 ;
        RECT 70.130 210.400 70.480 210.800 ;
        RECT 71.080 210.400 71.280 218.000 ;
        RECT 71.880 210.400 72.080 218.000 ;
        RECT 72.680 210.400 72.880 218.000 ;
        RECT 73.480 210.400 73.680 218.000 ;
        RECT 70.130 209.200 70.480 209.600 ;
        RECT 66.530 209.000 70.480 209.200 ;
        RECT 70.130 208.400 70.480 209.000 ;
        RECT 66.530 208.200 70.480 208.400 ;
        RECT 70.130 207.600 70.480 208.200 ;
        RECT 66.530 207.400 70.480 207.600 ;
        RECT 70.130 206.800 70.480 207.400 ;
        RECT 58.980 206.000 59.330 206.600 ;
        RECT 58.980 205.800 62.930 206.000 ;
        RECT 58.980 205.200 59.330 205.800 ;
        RECT 58.980 205.000 62.930 205.200 ;
        RECT 58.980 204.400 59.330 205.000 ;
        RECT 63.880 204.450 65.580 206.750 ;
        RECT 66.530 206.600 70.480 206.800 ;
        RECT 70.130 206.000 70.480 206.600 ;
        RECT 66.530 205.800 70.480 206.000 ;
        RECT 70.130 205.200 70.480 205.800 ;
        RECT 66.530 205.000 70.480 205.200 ;
        RECT 58.980 204.200 62.930 204.400 ;
        RECT 58.980 203.600 59.330 204.200 ;
        RECT 58.980 203.400 62.930 203.600 ;
        RECT 58.980 202.800 59.330 203.400 ;
        RECT 58.980 202.600 62.930 202.800 ;
        RECT 58.980 202.000 59.330 202.600 ;
        RECT 46.530 201.400 62.930 202.000 ;
        RECT 49.180 200.800 51.480 200.850 ;
        RECT 57.980 200.800 60.280 200.850 ;
        RECT 63.930 200.800 64.330 204.450 ;
        RECT 45.130 200.400 64.330 200.800 ;
        RECT 65.130 200.800 65.530 204.450 ;
        RECT 70.130 204.400 70.480 205.000 ;
        RECT 66.530 204.200 70.480 204.400 ;
        RECT 70.130 203.600 70.480 204.200 ;
        RECT 66.530 203.400 70.480 203.600 ;
        RECT 70.130 202.800 70.480 203.400 ;
        RECT 66.530 202.600 70.480 202.800 ;
        RECT 70.130 202.000 70.480 202.600 ;
        RECT 71.080 202.000 71.280 209.600 ;
        RECT 71.880 202.000 72.080 209.600 ;
        RECT 72.680 202.000 72.880 209.600 ;
        RECT 73.480 202.000 73.680 209.600 ;
        RECT 74.280 202.000 75.180 218.000 ;
        RECT 75.780 210.400 75.980 218.000 ;
        RECT 76.580 210.400 76.780 218.000 ;
        RECT 77.380 210.400 77.580 218.000 ;
        RECT 78.180 210.400 78.380 218.000 ;
        RECT 78.980 217.400 79.330 218.000 ;
        RECT 78.980 217.200 82.930 217.400 ;
        RECT 78.980 216.600 79.330 217.200 ;
        RECT 78.980 216.400 82.930 216.600 ;
        RECT 78.980 215.800 79.330 216.400 ;
        RECT 78.980 215.600 82.930 215.800 ;
        RECT 78.980 215.000 79.330 215.600 ;
        RECT 83.930 215.550 84.330 219.200 ;
        RECT 85.130 219.200 104.330 219.600 ;
        RECT 85.130 215.550 85.530 219.200 ;
        RECT 89.180 219.150 91.480 219.200 ;
        RECT 97.980 219.150 100.280 219.200 ;
        RECT 86.530 218.000 102.930 218.600 ;
        RECT 90.130 217.400 90.480 218.000 ;
        RECT 86.530 217.200 90.480 217.400 ;
        RECT 90.130 216.600 90.480 217.200 ;
        RECT 86.530 216.400 90.480 216.600 ;
        RECT 90.130 215.800 90.480 216.400 ;
        RECT 86.530 215.600 90.480 215.800 ;
        RECT 78.980 214.800 82.930 215.000 ;
        RECT 78.980 214.200 79.330 214.800 ;
        RECT 78.980 214.000 82.930 214.200 ;
        RECT 78.980 213.400 79.330 214.000 ;
        RECT 78.980 213.200 82.930 213.400 ;
        RECT 83.880 213.250 85.580 215.550 ;
        RECT 90.130 215.000 90.480 215.600 ;
        RECT 86.530 214.800 90.480 215.000 ;
        RECT 90.130 214.200 90.480 214.800 ;
        RECT 86.530 214.000 90.480 214.200 ;
        RECT 90.130 213.400 90.480 214.000 ;
        RECT 78.980 212.600 79.330 213.200 ;
        RECT 78.980 212.400 82.930 212.600 ;
        RECT 78.980 211.800 79.330 212.400 ;
        RECT 78.980 211.600 82.930 211.800 ;
        RECT 78.980 211.000 79.330 211.600 ;
        RECT 78.980 210.800 82.930 211.000 ;
        RECT 78.980 210.400 79.330 210.800 ;
        RECT 75.780 202.000 75.980 209.600 ;
        RECT 76.580 202.000 76.780 209.600 ;
        RECT 77.380 202.000 77.580 209.600 ;
        RECT 78.180 202.000 78.380 209.600 ;
        RECT 78.980 209.200 79.330 209.600 ;
        RECT 78.980 209.000 82.930 209.200 ;
        RECT 78.980 208.400 79.330 209.000 ;
        RECT 78.980 208.200 82.930 208.400 ;
        RECT 78.980 207.600 79.330 208.200 ;
        RECT 78.980 207.400 82.930 207.600 ;
        RECT 78.980 206.800 79.330 207.400 ;
        RECT 78.980 206.600 82.930 206.800 ;
        RECT 83.930 206.750 84.330 213.250 ;
        RECT 85.130 206.750 85.530 213.250 ;
        RECT 86.530 213.200 90.480 213.400 ;
        RECT 90.130 212.600 90.480 213.200 ;
        RECT 86.530 212.400 90.480 212.600 ;
        RECT 90.130 211.800 90.480 212.400 ;
        RECT 86.530 211.600 90.480 211.800 ;
        RECT 90.130 211.000 90.480 211.600 ;
        RECT 86.530 210.800 90.480 211.000 ;
        RECT 90.130 210.400 90.480 210.800 ;
        RECT 91.080 210.400 91.280 218.000 ;
        RECT 91.880 210.400 92.080 218.000 ;
        RECT 92.680 210.400 92.880 218.000 ;
        RECT 93.480 210.400 93.680 218.000 ;
        RECT 90.130 209.200 90.480 209.600 ;
        RECT 86.530 209.000 90.480 209.200 ;
        RECT 90.130 208.400 90.480 209.000 ;
        RECT 86.530 208.200 90.480 208.400 ;
        RECT 90.130 207.600 90.480 208.200 ;
        RECT 86.530 207.400 90.480 207.600 ;
        RECT 90.130 206.800 90.480 207.400 ;
        RECT 78.980 206.000 79.330 206.600 ;
        RECT 78.980 205.800 82.930 206.000 ;
        RECT 78.980 205.200 79.330 205.800 ;
        RECT 78.980 205.000 82.930 205.200 ;
        RECT 78.980 204.400 79.330 205.000 ;
        RECT 83.880 204.450 85.580 206.750 ;
        RECT 86.530 206.600 90.480 206.800 ;
        RECT 90.130 206.000 90.480 206.600 ;
        RECT 86.530 205.800 90.480 206.000 ;
        RECT 90.130 205.200 90.480 205.800 ;
        RECT 86.530 205.000 90.480 205.200 ;
        RECT 78.980 204.200 82.930 204.400 ;
        RECT 78.980 203.600 79.330 204.200 ;
        RECT 78.980 203.400 82.930 203.600 ;
        RECT 78.980 202.800 79.330 203.400 ;
        RECT 78.980 202.600 82.930 202.800 ;
        RECT 78.980 202.000 79.330 202.600 ;
        RECT 66.530 201.400 82.930 202.000 ;
        RECT 69.180 200.800 71.480 200.850 ;
        RECT 77.980 200.800 80.280 200.850 ;
        RECT 83.930 200.800 84.330 204.450 ;
        RECT 65.130 200.400 84.330 200.800 ;
        RECT 85.130 200.800 85.530 204.450 ;
        RECT 90.130 204.400 90.480 205.000 ;
        RECT 86.530 204.200 90.480 204.400 ;
        RECT 90.130 203.600 90.480 204.200 ;
        RECT 86.530 203.400 90.480 203.600 ;
        RECT 90.130 202.800 90.480 203.400 ;
        RECT 86.530 202.600 90.480 202.800 ;
        RECT 90.130 202.000 90.480 202.600 ;
        RECT 91.080 202.000 91.280 209.600 ;
        RECT 91.880 202.000 92.080 209.600 ;
        RECT 92.680 202.000 92.880 209.600 ;
        RECT 93.480 202.000 93.680 209.600 ;
        RECT 94.280 202.000 95.180 218.000 ;
        RECT 95.780 210.400 95.980 218.000 ;
        RECT 96.580 210.400 96.780 218.000 ;
        RECT 97.380 210.400 97.580 218.000 ;
        RECT 98.180 210.400 98.380 218.000 ;
        RECT 98.980 217.400 99.330 218.000 ;
        RECT 98.980 217.200 102.930 217.400 ;
        RECT 98.980 216.600 99.330 217.200 ;
        RECT 98.980 216.400 102.930 216.600 ;
        RECT 98.980 215.800 99.330 216.400 ;
        RECT 98.980 215.600 102.930 215.800 ;
        RECT 98.980 215.000 99.330 215.600 ;
        RECT 103.930 215.550 104.330 219.200 ;
        RECT 105.130 219.200 124.330 219.600 ;
        RECT 105.130 215.550 105.530 219.200 ;
        RECT 109.180 219.150 111.480 219.200 ;
        RECT 117.980 219.150 120.280 219.200 ;
        RECT 106.530 218.000 122.930 218.600 ;
        RECT 110.130 217.400 110.480 218.000 ;
        RECT 106.530 217.200 110.480 217.400 ;
        RECT 110.130 216.600 110.480 217.200 ;
        RECT 106.530 216.400 110.480 216.600 ;
        RECT 110.130 215.800 110.480 216.400 ;
        RECT 106.530 215.600 110.480 215.800 ;
        RECT 98.980 214.800 102.930 215.000 ;
        RECT 98.980 214.200 99.330 214.800 ;
        RECT 98.980 214.000 102.930 214.200 ;
        RECT 98.980 213.400 99.330 214.000 ;
        RECT 98.980 213.200 102.930 213.400 ;
        RECT 103.880 213.250 105.580 215.550 ;
        RECT 110.130 215.000 110.480 215.600 ;
        RECT 106.530 214.800 110.480 215.000 ;
        RECT 110.130 214.200 110.480 214.800 ;
        RECT 106.530 214.000 110.480 214.200 ;
        RECT 110.130 213.400 110.480 214.000 ;
        RECT 98.980 212.600 99.330 213.200 ;
        RECT 98.980 212.400 102.930 212.600 ;
        RECT 98.980 211.800 99.330 212.400 ;
        RECT 98.980 211.600 102.930 211.800 ;
        RECT 98.980 211.000 99.330 211.600 ;
        RECT 98.980 210.800 102.930 211.000 ;
        RECT 98.980 210.400 99.330 210.800 ;
        RECT 95.780 202.000 95.980 209.600 ;
        RECT 96.580 202.000 96.780 209.600 ;
        RECT 97.380 202.000 97.580 209.600 ;
        RECT 98.180 202.000 98.380 209.600 ;
        RECT 98.980 209.200 99.330 209.600 ;
        RECT 98.980 209.000 102.930 209.200 ;
        RECT 98.980 208.400 99.330 209.000 ;
        RECT 98.980 208.200 102.930 208.400 ;
        RECT 98.980 207.600 99.330 208.200 ;
        RECT 98.980 207.400 102.930 207.600 ;
        RECT 98.980 206.800 99.330 207.400 ;
        RECT 98.980 206.600 102.930 206.800 ;
        RECT 103.930 206.750 104.330 213.250 ;
        RECT 105.130 206.750 105.530 213.250 ;
        RECT 106.530 213.200 110.480 213.400 ;
        RECT 110.130 212.600 110.480 213.200 ;
        RECT 106.530 212.400 110.480 212.600 ;
        RECT 110.130 211.800 110.480 212.400 ;
        RECT 106.530 211.600 110.480 211.800 ;
        RECT 110.130 211.000 110.480 211.600 ;
        RECT 106.530 210.800 110.480 211.000 ;
        RECT 110.130 210.400 110.480 210.800 ;
        RECT 111.080 210.400 111.280 218.000 ;
        RECT 111.880 210.400 112.080 218.000 ;
        RECT 112.680 210.400 112.880 218.000 ;
        RECT 113.480 210.400 113.680 218.000 ;
        RECT 110.130 209.200 110.480 209.600 ;
        RECT 106.530 209.000 110.480 209.200 ;
        RECT 110.130 208.400 110.480 209.000 ;
        RECT 106.530 208.200 110.480 208.400 ;
        RECT 110.130 207.600 110.480 208.200 ;
        RECT 106.530 207.400 110.480 207.600 ;
        RECT 110.130 206.800 110.480 207.400 ;
        RECT 98.980 206.000 99.330 206.600 ;
        RECT 98.980 205.800 102.930 206.000 ;
        RECT 98.980 205.200 99.330 205.800 ;
        RECT 98.980 205.000 102.930 205.200 ;
        RECT 98.980 204.400 99.330 205.000 ;
        RECT 103.880 204.450 105.580 206.750 ;
        RECT 106.530 206.600 110.480 206.800 ;
        RECT 110.130 206.000 110.480 206.600 ;
        RECT 106.530 205.800 110.480 206.000 ;
        RECT 110.130 205.200 110.480 205.800 ;
        RECT 106.530 205.000 110.480 205.200 ;
        RECT 98.980 204.200 102.930 204.400 ;
        RECT 98.980 203.600 99.330 204.200 ;
        RECT 98.980 203.400 102.930 203.600 ;
        RECT 98.980 202.800 99.330 203.400 ;
        RECT 98.980 202.600 102.930 202.800 ;
        RECT 98.980 202.000 99.330 202.600 ;
        RECT 86.530 201.400 102.930 202.000 ;
        RECT 89.180 200.800 91.480 200.850 ;
        RECT 97.980 200.800 100.280 200.850 ;
        RECT 103.930 200.800 104.330 204.450 ;
        RECT 85.130 200.400 104.330 200.800 ;
        RECT 105.130 200.800 105.530 204.450 ;
        RECT 110.130 204.400 110.480 205.000 ;
        RECT 106.530 204.200 110.480 204.400 ;
        RECT 110.130 203.600 110.480 204.200 ;
        RECT 106.530 203.400 110.480 203.600 ;
        RECT 110.130 202.800 110.480 203.400 ;
        RECT 106.530 202.600 110.480 202.800 ;
        RECT 110.130 202.000 110.480 202.600 ;
        RECT 111.080 202.000 111.280 209.600 ;
        RECT 111.880 202.000 112.080 209.600 ;
        RECT 112.680 202.000 112.880 209.600 ;
        RECT 113.480 202.000 113.680 209.600 ;
        RECT 114.280 202.000 115.180 218.000 ;
        RECT 115.780 210.400 115.980 218.000 ;
        RECT 116.580 210.400 116.780 218.000 ;
        RECT 117.380 210.400 117.580 218.000 ;
        RECT 118.180 210.400 118.380 218.000 ;
        RECT 118.980 217.400 119.330 218.000 ;
        RECT 118.980 217.200 122.930 217.400 ;
        RECT 118.980 216.600 119.330 217.200 ;
        RECT 118.980 216.400 122.930 216.600 ;
        RECT 118.980 215.800 119.330 216.400 ;
        RECT 118.980 215.600 122.930 215.800 ;
        RECT 118.980 215.000 119.330 215.600 ;
        RECT 123.930 215.550 124.330 219.200 ;
        RECT 125.340 217.260 125.700 217.640 ;
        RECT 125.970 217.260 126.330 217.640 ;
        RECT 126.570 217.260 126.930 217.640 ;
        RECT 125.340 216.670 125.700 217.050 ;
        RECT 125.970 216.670 126.330 217.050 ;
        RECT 126.570 216.670 126.930 217.050 ;
        RECT 118.980 214.800 122.930 215.000 ;
        RECT 118.980 214.200 119.330 214.800 ;
        RECT 118.980 214.000 122.930 214.200 ;
        RECT 118.980 213.400 119.330 214.000 ;
        RECT 118.980 213.200 122.930 213.400 ;
        RECT 123.880 213.250 124.730 215.550 ;
        RECT 118.980 212.600 119.330 213.200 ;
        RECT 118.980 212.400 122.930 212.600 ;
        RECT 118.980 211.800 119.330 212.400 ;
        RECT 118.980 211.600 122.930 211.800 ;
        RECT 118.980 211.000 119.330 211.600 ;
        RECT 118.980 210.800 122.930 211.000 ;
        RECT 118.980 210.400 119.330 210.800 ;
        RECT 115.780 202.000 115.980 209.600 ;
        RECT 116.580 202.000 116.780 209.600 ;
        RECT 117.380 202.000 117.580 209.600 ;
        RECT 118.180 202.000 118.380 209.600 ;
        RECT 118.980 209.200 119.330 209.600 ;
        RECT 118.980 209.000 122.930 209.200 ;
        RECT 118.980 208.400 119.330 209.000 ;
        RECT 118.980 208.200 122.930 208.400 ;
        RECT 118.980 207.600 119.330 208.200 ;
        RECT 118.980 207.400 122.930 207.600 ;
        RECT 118.980 206.800 119.330 207.400 ;
        RECT 118.980 206.600 122.930 206.800 ;
        RECT 123.930 206.750 124.330 213.250 ;
        RECT 118.980 206.000 119.330 206.600 ;
        RECT 118.980 205.800 122.930 206.000 ;
        RECT 118.980 205.200 119.330 205.800 ;
        RECT 118.980 205.000 122.930 205.200 ;
        RECT 118.980 204.400 119.330 205.000 ;
        RECT 123.880 204.450 124.730 206.750 ;
        RECT 118.980 204.200 122.930 204.400 ;
        RECT 118.980 203.600 119.330 204.200 ;
        RECT 118.980 203.400 122.930 203.600 ;
        RECT 118.980 202.800 119.330 203.400 ;
        RECT 118.980 202.600 122.930 202.800 ;
        RECT 118.980 202.000 119.330 202.600 ;
        RECT 106.530 201.400 122.930 202.000 ;
        RECT 109.180 200.800 111.480 200.850 ;
        RECT 117.980 200.800 120.280 200.850 ;
        RECT 123.930 200.800 124.330 204.450 ;
        RECT 125.340 201.680 125.700 202.060 ;
        RECT 125.970 201.680 126.330 202.060 ;
        RECT 126.570 201.680 126.930 202.060 ;
        RECT 125.340 201.090 125.700 201.470 ;
        RECT 125.970 201.090 126.330 201.470 ;
        RECT 126.570 201.090 126.930 201.470 ;
        RECT 105.130 200.400 124.330 200.800 ;
        RECT 9.180 200.000 11.480 200.400 ;
        RECT 17.980 200.000 20.280 200.400 ;
        RECT 29.180 200.000 31.480 200.400 ;
        RECT 37.980 200.000 40.280 200.400 ;
        RECT 49.180 200.000 51.480 200.400 ;
        RECT 57.980 200.000 60.280 200.400 ;
        RECT 69.180 200.000 71.480 200.400 ;
        RECT 77.980 200.000 80.280 200.400 ;
        RECT 89.180 200.000 91.480 200.400 ;
        RECT 97.980 200.000 100.280 200.400 ;
        RECT 109.180 200.000 111.480 200.400 ;
        RECT 117.980 200.000 120.280 200.400 ;
        RECT 4.720 177.380 26.020 178.635 ;
        RECT 4.720 163.250 6.190 177.380 ;
        RECT 7.100 175.375 7.560 175.545 ;
        RECT 7.185 174.650 7.475 175.375 ;
        RECT 8.020 173.450 8.190 175.695 ;
        RECT 9.595 175.290 9.770 175.695 ;
        RECT 24.570 175.540 26.020 177.380 ;
        RECT 47.085 176.260 49.385 176.660 ;
        RECT 55.885 176.260 58.185 176.660 ;
        RECT 67.085 176.260 69.385 176.660 ;
        RECT 75.885 176.260 78.185 176.660 ;
        RECT 87.085 176.260 89.385 176.660 ;
        RECT 95.885 176.260 98.185 176.660 ;
        RECT 107.085 176.260 109.385 176.660 ;
        RECT 115.885 176.260 118.185 176.660 ;
        RECT 14.865 175.370 26.020 175.540 ;
        RECT 9.600 173.450 9.770 175.290 ;
        RECT 14.950 174.645 15.240 175.370 ;
        RECT 15.560 174.570 15.890 175.370 ;
        RECT 16.400 174.890 16.730 175.370 ;
        RECT 17.320 174.890 17.560 175.370 ;
        RECT 18.320 174.570 18.650 175.370 ;
        RECT 19.160 174.890 19.490 175.370 ;
        RECT 20.080 174.890 20.320 175.370 ;
        RECT 21.675 174.550 21.905 175.370 ;
        RECT 23.055 174.550 23.285 175.370 ;
        RECT 8.050 170.100 8.340 170.825 ;
        RECT 9.410 170.100 9.720 170.900 ;
        RECT 10.500 170.100 10.885 170.500 ;
        RECT 11.915 170.100 12.300 170.500 ;
        RECT 13.330 170.100 13.715 170.500 ;
        RECT 15.100 170.100 15.485 170.500 ;
        RECT 16.515 170.100 16.900 170.500 ;
        RECT 17.930 170.100 18.315 170.500 ;
        RECT 19.700 170.100 20.085 170.500 ;
        RECT 21.115 170.100 21.500 170.500 ;
        RECT 22.530 170.100 22.915 170.500 ;
        RECT 23.690 170.100 23.980 170.825 ;
        RECT 24.570 170.100 26.020 175.370 ;
        RECT 43.035 175.860 62.235 176.260 ;
        RECT 43.035 172.210 43.435 175.860 ;
        RECT 47.085 175.810 49.385 175.860 ;
        RECT 55.885 175.810 58.185 175.860 ;
        RECT 44.435 174.660 60.835 175.260 ;
        RECT 48.035 174.060 48.385 174.660 ;
        RECT 44.435 173.860 48.385 174.060 ;
        RECT 48.035 173.260 48.385 173.860 ;
        RECT 44.435 173.060 48.385 173.260 ;
        RECT 48.035 172.460 48.385 173.060 ;
        RECT 44.435 172.260 48.385 172.460 ;
        RECT 6.585 169.930 26.020 170.100 ;
        RECT 6.670 169.205 6.960 169.930 ;
        RECT 7.365 169.110 7.595 169.930 ;
        RECT 8.510 169.130 8.820 169.930 ;
        RECT 10.500 169.530 10.885 169.930 ;
        RECT 11.915 169.530 12.300 169.930 ;
        RECT 13.330 169.530 13.715 169.930 ;
        RECT 15.100 169.530 15.485 169.930 ;
        RECT 16.515 169.530 16.900 169.930 ;
        RECT 17.930 169.530 18.315 169.930 ;
        RECT 19.700 169.530 20.085 169.930 ;
        RECT 21.115 169.530 21.500 169.930 ;
        RECT 22.530 169.530 22.915 169.930 ;
        RECT 23.690 169.205 23.980 169.930 ;
        RECT 7.590 164.660 7.880 165.385 ;
        RECT 14.950 164.660 15.240 165.385 ;
        RECT 15.560 164.660 15.890 165.460 ;
        RECT 16.400 164.660 16.730 165.140 ;
        RECT 17.320 164.660 17.560 165.140 ;
        RECT 18.320 164.660 18.650 165.460 ;
        RECT 19.160 164.660 19.490 165.140 ;
        RECT 20.080 164.660 20.320 165.140 ;
        RECT 21.675 164.660 21.905 165.480 ;
        RECT 23.055 164.660 23.285 165.480 ;
        RECT 24.570 164.660 26.020 169.930 ;
        RECT 42.635 169.910 43.485 172.210 ;
        RECT 48.035 171.660 48.385 172.260 ;
        RECT 44.435 171.460 48.385 171.660 ;
        RECT 48.035 170.860 48.385 171.460 ;
        RECT 44.435 170.660 48.385 170.860 ;
        RECT 48.035 170.060 48.385 170.660 ;
        RECT 7.505 164.490 7.965 164.660 ;
        RECT 14.865 164.490 26.020 164.660 ;
        RECT 24.570 163.250 26.020 164.490 ;
        RECT 43.035 163.410 43.435 169.910 ;
        RECT 44.435 169.860 48.385 170.060 ;
        RECT 48.035 169.260 48.385 169.860 ;
        RECT 44.435 169.060 48.385 169.260 ;
        RECT 48.035 168.460 48.385 169.060 ;
        RECT 44.435 168.260 48.385 168.460 ;
        RECT 48.035 167.660 48.385 168.260 ;
        RECT 44.435 167.460 48.385 167.660 ;
        RECT 48.035 167.060 48.385 167.460 ;
        RECT 48.985 167.060 49.185 174.660 ;
        RECT 49.785 167.060 49.985 174.660 ;
        RECT 50.585 167.060 50.785 174.660 ;
        RECT 51.385 167.060 51.585 174.660 ;
        RECT 48.035 165.860 48.385 166.260 ;
        RECT 44.435 165.660 48.385 165.860 ;
        RECT 48.035 165.060 48.385 165.660 ;
        RECT 44.435 164.860 48.385 165.060 ;
        RECT 48.035 164.260 48.385 164.860 ;
        RECT 44.435 164.060 48.385 164.260 ;
        RECT 48.035 163.460 48.385 164.060 ;
        RECT 4.720 162.245 26.020 163.250 ;
        RECT 4.720 162.055 26.015 162.245 ;
        RECT 42.635 161.110 43.485 163.410 ;
        RECT 44.435 163.260 48.385 163.460 ;
        RECT 48.035 162.660 48.385 163.260 ;
        RECT 44.435 162.460 48.385 162.660 ;
        RECT 48.035 161.860 48.385 162.460 ;
        RECT 44.435 161.660 48.385 161.860 ;
        RECT 43.035 157.460 43.435 161.110 ;
        RECT 48.035 161.060 48.385 161.660 ;
        RECT 44.435 160.860 48.385 161.060 ;
        RECT 48.035 160.260 48.385 160.860 ;
        RECT 44.435 160.060 48.385 160.260 ;
        RECT 48.035 159.460 48.385 160.060 ;
        RECT 44.435 159.260 48.385 159.460 ;
        RECT 48.035 158.660 48.385 159.260 ;
        RECT 48.985 158.660 49.185 166.260 ;
        RECT 49.785 158.660 49.985 166.260 ;
        RECT 50.585 158.660 50.785 166.260 ;
        RECT 51.385 158.660 51.585 166.260 ;
        RECT 52.185 158.660 53.085 174.660 ;
        RECT 53.685 167.060 53.885 174.660 ;
        RECT 54.485 167.060 54.685 174.660 ;
        RECT 55.285 167.060 55.485 174.660 ;
        RECT 56.085 167.060 56.285 174.660 ;
        RECT 56.885 174.060 57.235 174.660 ;
        RECT 56.885 173.860 60.835 174.060 ;
        RECT 56.885 173.260 57.235 173.860 ;
        RECT 56.885 173.060 60.835 173.260 ;
        RECT 56.885 172.460 57.235 173.060 ;
        RECT 56.885 172.260 60.835 172.460 ;
        RECT 56.885 171.660 57.235 172.260 ;
        RECT 61.835 172.210 62.235 175.860 ;
        RECT 63.035 175.860 82.235 176.260 ;
        RECT 63.035 172.210 63.435 175.860 ;
        RECT 67.085 175.810 69.385 175.860 ;
        RECT 75.885 175.810 78.185 175.860 ;
        RECT 64.435 174.660 80.835 175.260 ;
        RECT 68.035 174.060 68.385 174.660 ;
        RECT 64.435 173.860 68.385 174.060 ;
        RECT 68.035 173.260 68.385 173.860 ;
        RECT 64.435 173.060 68.385 173.260 ;
        RECT 68.035 172.460 68.385 173.060 ;
        RECT 64.435 172.260 68.385 172.460 ;
        RECT 56.885 171.460 60.835 171.660 ;
        RECT 56.885 170.860 57.235 171.460 ;
        RECT 56.885 170.660 60.835 170.860 ;
        RECT 56.885 170.060 57.235 170.660 ;
        RECT 56.885 169.860 60.835 170.060 ;
        RECT 61.785 169.910 63.485 172.210 ;
        RECT 68.035 171.660 68.385 172.260 ;
        RECT 64.435 171.460 68.385 171.660 ;
        RECT 68.035 170.860 68.385 171.460 ;
        RECT 64.435 170.660 68.385 170.860 ;
        RECT 68.035 170.060 68.385 170.660 ;
        RECT 56.885 169.260 57.235 169.860 ;
        RECT 56.885 169.060 60.835 169.260 ;
        RECT 56.885 168.460 57.235 169.060 ;
        RECT 56.885 168.260 60.835 168.460 ;
        RECT 56.885 167.660 57.235 168.260 ;
        RECT 56.885 167.460 60.835 167.660 ;
        RECT 56.885 167.060 57.235 167.460 ;
        RECT 53.685 158.660 53.885 166.260 ;
        RECT 54.485 158.660 54.685 166.260 ;
        RECT 55.285 158.660 55.485 166.260 ;
        RECT 56.085 158.660 56.285 166.260 ;
        RECT 56.885 165.860 57.235 166.260 ;
        RECT 56.885 165.660 60.835 165.860 ;
        RECT 56.885 165.060 57.235 165.660 ;
        RECT 56.885 164.860 60.835 165.060 ;
        RECT 56.885 164.260 57.235 164.860 ;
        RECT 56.885 164.060 60.835 164.260 ;
        RECT 56.885 163.460 57.235 164.060 ;
        RECT 56.885 163.260 60.835 163.460 ;
        RECT 61.835 163.410 62.235 169.910 ;
        RECT 63.035 163.410 63.435 169.910 ;
        RECT 64.435 169.860 68.385 170.060 ;
        RECT 68.035 169.260 68.385 169.860 ;
        RECT 64.435 169.060 68.385 169.260 ;
        RECT 68.035 168.460 68.385 169.060 ;
        RECT 64.435 168.260 68.385 168.460 ;
        RECT 68.035 167.660 68.385 168.260 ;
        RECT 64.435 167.460 68.385 167.660 ;
        RECT 68.035 167.060 68.385 167.460 ;
        RECT 68.985 167.060 69.185 174.660 ;
        RECT 69.785 167.060 69.985 174.660 ;
        RECT 70.585 167.060 70.785 174.660 ;
        RECT 71.385 167.060 71.585 174.660 ;
        RECT 68.035 165.860 68.385 166.260 ;
        RECT 64.435 165.660 68.385 165.860 ;
        RECT 68.035 165.060 68.385 165.660 ;
        RECT 64.435 164.860 68.385 165.060 ;
        RECT 68.035 164.260 68.385 164.860 ;
        RECT 64.435 164.060 68.385 164.260 ;
        RECT 68.035 163.460 68.385 164.060 ;
        RECT 56.885 162.660 57.235 163.260 ;
        RECT 56.885 162.460 60.835 162.660 ;
        RECT 56.885 161.860 57.235 162.460 ;
        RECT 56.885 161.660 60.835 161.860 ;
        RECT 56.885 161.060 57.235 161.660 ;
        RECT 61.785 161.110 63.485 163.410 ;
        RECT 64.435 163.260 68.385 163.460 ;
        RECT 68.035 162.660 68.385 163.260 ;
        RECT 64.435 162.460 68.385 162.660 ;
        RECT 68.035 161.860 68.385 162.460 ;
        RECT 64.435 161.660 68.385 161.860 ;
        RECT 56.885 160.860 60.835 161.060 ;
        RECT 56.885 160.260 57.235 160.860 ;
        RECT 56.885 160.060 60.835 160.260 ;
        RECT 56.885 159.460 57.235 160.060 ;
        RECT 56.885 159.260 60.835 159.460 ;
        RECT 56.885 158.660 57.235 159.260 ;
        RECT 44.435 158.060 60.835 158.660 ;
        RECT 47.085 157.460 49.385 157.510 ;
        RECT 55.885 157.460 58.185 157.510 ;
        RECT 61.835 157.460 62.235 161.110 ;
        RECT 43.035 157.060 62.235 157.460 ;
        RECT 63.035 157.460 63.435 161.110 ;
        RECT 68.035 161.060 68.385 161.660 ;
        RECT 64.435 160.860 68.385 161.060 ;
        RECT 68.035 160.260 68.385 160.860 ;
        RECT 64.435 160.060 68.385 160.260 ;
        RECT 68.035 159.460 68.385 160.060 ;
        RECT 64.435 159.260 68.385 159.460 ;
        RECT 68.035 158.660 68.385 159.260 ;
        RECT 68.985 158.660 69.185 166.260 ;
        RECT 69.785 158.660 69.985 166.260 ;
        RECT 70.585 158.660 70.785 166.260 ;
        RECT 71.385 158.660 71.585 166.260 ;
        RECT 72.185 158.660 73.085 174.660 ;
        RECT 73.685 167.060 73.885 174.660 ;
        RECT 74.485 167.060 74.685 174.660 ;
        RECT 75.285 167.060 75.485 174.660 ;
        RECT 76.085 167.060 76.285 174.660 ;
        RECT 76.885 174.060 77.235 174.660 ;
        RECT 76.885 173.860 80.835 174.060 ;
        RECT 76.885 173.260 77.235 173.860 ;
        RECT 76.885 173.060 80.835 173.260 ;
        RECT 76.885 172.460 77.235 173.060 ;
        RECT 76.885 172.260 80.835 172.460 ;
        RECT 76.885 171.660 77.235 172.260 ;
        RECT 81.835 172.210 82.235 175.860 ;
        RECT 83.035 175.860 102.235 176.260 ;
        RECT 83.035 172.210 83.435 175.860 ;
        RECT 87.085 175.810 89.385 175.860 ;
        RECT 95.885 175.810 98.185 175.860 ;
        RECT 84.435 174.660 100.835 175.260 ;
        RECT 88.035 174.060 88.385 174.660 ;
        RECT 84.435 173.860 88.385 174.060 ;
        RECT 88.035 173.260 88.385 173.860 ;
        RECT 84.435 173.060 88.385 173.260 ;
        RECT 88.035 172.460 88.385 173.060 ;
        RECT 84.435 172.260 88.385 172.460 ;
        RECT 76.885 171.460 80.835 171.660 ;
        RECT 76.885 170.860 77.235 171.460 ;
        RECT 76.885 170.660 80.835 170.860 ;
        RECT 76.885 170.060 77.235 170.660 ;
        RECT 76.885 169.860 80.835 170.060 ;
        RECT 81.785 169.910 83.485 172.210 ;
        RECT 88.035 171.660 88.385 172.260 ;
        RECT 84.435 171.460 88.385 171.660 ;
        RECT 88.035 170.860 88.385 171.460 ;
        RECT 84.435 170.660 88.385 170.860 ;
        RECT 88.035 170.060 88.385 170.660 ;
        RECT 76.885 169.260 77.235 169.860 ;
        RECT 76.885 169.060 80.835 169.260 ;
        RECT 76.885 168.460 77.235 169.060 ;
        RECT 76.885 168.260 80.835 168.460 ;
        RECT 76.885 167.660 77.235 168.260 ;
        RECT 76.885 167.460 80.835 167.660 ;
        RECT 76.885 167.060 77.235 167.460 ;
        RECT 73.685 158.660 73.885 166.260 ;
        RECT 74.485 158.660 74.685 166.260 ;
        RECT 75.285 158.660 75.485 166.260 ;
        RECT 76.085 158.660 76.285 166.260 ;
        RECT 76.885 165.860 77.235 166.260 ;
        RECT 76.885 165.660 80.835 165.860 ;
        RECT 76.885 165.060 77.235 165.660 ;
        RECT 76.885 164.860 80.835 165.060 ;
        RECT 76.885 164.260 77.235 164.860 ;
        RECT 76.885 164.060 80.835 164.260 ;
        RECT 76.885 163.460 77.235 164.060 ;
        RECT 76.885 163.260 80.835 163.460 ;
        RECT 81.835 163.410 82.235 169.910 ;
        RECT 83.035 163.410 83.435 169.910 ;
        RECT 84.435 169.860 88.385 170.060 ;
        RECT 88.035 169.260 88.385 169.860 ;
        RECT 84.435 169.060 88.385 169.260 ;
        RECT 88.035 168.460 88.385 169.060 ;
        RECT 84.435 168.260 88.385 168.460 ;
        RECT 88.035 167.660 88.385 168.260 ;
        RECT 84.435 167.460 88.385 167.660 ;
        RECT 88.035 167.060 88.385 167.460 ;
        RECT 88.985 167.060 89.185 174.660 ;
        RECT 89.785 167.060 89.985 174.660 ;
        RECT 90.585 167.060 90.785 174.660 ;
        RECT 91.385 167.060 91.585 174.660 ;
        RECT 88.035 165.860 88.385 166.260 ;
        RECT 84.435 165.660 88.385 165.860 ;
        RECT 88.035 165.060 88.385 165.660 ;
        RECT 84.435 164.860 88.385 165.060 ;
        RECT 88.035 164.260 88.385 164.860 ;
        RECT 84.435 164.060 88.385 164.260 ;
        RECT 88.035 163.460 88.385 164.060 ;
        RECT 76.885 162.660 77.235 163.260 ;
        RECT 76.885 162.460 80.835 162.660 ;
        RECT 76.885 161.860 77.235 162.460 ;
        RECT 76.885 161.660 80.835 161.860 ;
        RECT 76.885 161.060 77.235 161.660 ;
        RECT 81.785 161.110 83.485 163.410 ;
        RECT 84.435 163.260 88.385 163.460 ;
        RECT 88.035 162.660 88.385 163.260 ;
        RECT 84.435 162.460 88.385 162.660 ;
        RECT 88.035 161.860 88.385 162.460 ;
        RECT 84.435 161.660 88.385 161.860 ;
        RECT 76.885 160.860 80.835 161.060 ;
        RECT 76.885 160.260 77.235 160.860 ;
        RECT 76.885 160.060 80.835 160.260 ;
        RECT 76.885 159.460 77.235 160.060 ;
        RECT 76.885 159.260 80.835 159.460 ;
        RECT 76.885 158.660 77.235 159.260 ;
        RECT 64.435 158.060 80.835 158.660 ;
        RECT 67.085 157.460 69.385 157.510 ;
        RECT 75.885 157.460 78.185 157.510 ;
        RECT 81.835 157.460 82.235 161.110 ;
        RECT 63.035 157.060 82.235 157.460 ;
        RECT 83.035 157.460 83.435 161.110 ;
        RECT 88.035 161.060 88.385 161.660 ;
        RECT 84.435 160.860 88.385 161.060 ;
        RECT 88.035 160.260 88.385 160.860 ;
        RECT 84.435 160.060 88.385 160.260 ;
        RECT 88.035 159.460 88.385 160.060 ;
        RECT 84.435 159.260 88.385 159.460 ;
        RECT 88.035 158.660 88.385 159.260 ;
        RECT 88.985 158.660 89.185 166.260 ;
        RECT 89.785 158.660 89.985 166.260 ;
        RECT 90.585 158.660 90.785 166.260 ;
        RECT 91.385 158.660 91.585 166.260 ;
        RECT 92.185 158.660 93.085 174.660 ;
        RECT 93.685 167.060 93.885 174.660 ;
        RECT 94.485 167.060 94.685 174.660 ;
        RECT 95.285 167.060 95.485 174.660 ;
        RECT 96.085 167.060 96.285 174.660 ;
        RECT 96.885 174.060 97.235 174.660 ;
        RECT 96.885 173.860 100.835 174.060 ;
        RECT 96.885 173.260 97.235 173.860 ;
        RECT 96.885 173.060 100.835 173.260 ;
        RECT 96.885 172.460 97.235 173.060 ;
        RECT 96.885 172.260 100.835 172.460 ;
        RECT 96.885 171.660 97.235 172.260 ;
        RECT 101.835 172.210 102.235 175.860 ;
        RECT 103.035 175.860 122.235 176.260 ;
        RECT 103.035 172.210 103.435 175.860 ;
        RECT 107.085 175.810 109.385 175.860 ;
        RECT 115.885 175.810 118.185 175.860 ;
        RECT 104.435 174.660 120.835 175.260 ;
        RECT 108.035 174.060 108.385 174.660 ;
        RECT 104.435 173.860 108.385 174.060 ;
        RECT 108.035 173.260 108.385 173.860 ;
        RECT 104.435 173.060 108.385 173.260 ;
        RECT 108.035 172.460 108.385 173.060 ;
        RECT 104.435 172.260 108.385 172.460 ;
        RECT 96.885 171.460 100.835 171.660 ;
        RECT 96.885 170.860 97.235 171.460 ;
        RECT 96.885 170.660 100.835 170.860 ;
        RECT 96.885 170.060 97.235 170.660 ;
        RECT 96.885 169.860 100.835 170.060 ;
        RECT 101.785 169.910 103.485 172.210 ;
        RECT 108.035 171.660 108.385 172.260 ;
        RECT 104.435 171.460 108.385 171.660 ;
        RECT 108.035 170.860 108.385 171.460 ;
        RECT 104.435 170.660 108.385 170.860 ;
        RECT 108.035 170.060 108.385 170.660 ;
        RECT 96.885 169.260 97.235 169.860 ;
        RECT 96.885 169.060 100.835 169.260 ;
        RECT 96.885 168.460 97.235 169.060 ;
        RECT 96.885 168.260 100.835 168.460 ;
        RECT 96.885 167.660 97.235 168.260 ;
        RECT 96.885 167.460 100.835 167.660 ;
        RECT 96.885 167.060 97.235 167.460 ;
        RECT 93.685 158.660 93.885 166.260 ;
        RECT 94.485 158.660 94.685 166.260 ;
        RECT 95.285 158.660 95.485 166.260 ;
        RECT 96.085 158.660 96.285 166.260 ;
        RECT 96.885 165.860 97.235 166.260 ;
        RECT 96.885 165.660 100.835 165.860 ;
        RECT 96.885 165.060 97.235 165.660 ;
        RECT 96.885 164.860 100.835 165.060 ;
        RECT 96.885 164.260 97.235 164.860 ;
        RECT 96.885 164.060 100.835 164.260 ;
        RECT 96.885 163.460 97.235 164.060 ;
        RECT 96.885 163.260 100.835 163.460 ;
        RECT 101.835 163.410 102.235 169.910 ;
        RECT 103.035 163.410 103.435 169.910 ;
        RECT 104.435 169.860 108.385 170.060 ;
        RECT 108.035 169.260 108.385 169.860 ;
        RECT 104.435 169.060 108.385 169.260 ;
        RECT 108.035 168.460 108.385 169.060 ;
        RECT 104.435 168.260 108.385 168.460 ;
        RECT 108.035 167.660 108.385 168.260 ;
        RECT 104.435 167.460 108.385 167.660 ;
        RECT 108.035 167.060 108.385 167.460 ;
        RECT 108.985 167.060 109.185 174.660 ;
        RECT 109.785 167.060 109.985 174.660 ;
        RECT 110.585 167.060 110.785 174.660 ;
        RECT 111.385 167.060 111.585 174.660 ;
        RECT 108.035 165.860 108.385 166.260 ;
        RECT 104.435 165.660 108.385 165.860 ;
        RECT 108.035 165.060 108.385 165.660 ;
        RECT 104.435 164.860 108.385 165.060 ;
        RECT 108.035 164.260 108.385 164.860 ;
        RECT 104.435 164.060 108.385 164.260 ;
        RECT 108.035 163.460 108.385 164.060 ;
        RECT 96.885 162.660 97.235 163.260 ;
        RECT 96.885 162.460 100.835 162.660 ;
        RECT 96.885 161.860 97.235 162.460 ;
        RECT 96.885 161.660 100.835 161.860 ;
        RECT 96.885 161.060 97.235 161.660 ;
        RECT 101.785 161.110 103.485 163.410 ;
        RECT 104.435 163.260 108.385 163.460 ;
        RECT 108.035 162.660 108.385 163.260 ;
        RECT 104.435 162.460 108.385 162.660 ;
        RECT 108.035 161.860 108.385 162.460 ;
        RECT 104.435 161.660 108.385 161.860 ;
        RECT 96.885 160.860 100.835 161.060 ;
        RECT 96.885 160.260 97.235 160.860 ;
        RECT 96.885 160.060 100.835 160.260 ;
        RECT 96.885 159.460 97.235 160.060 ;
        RECT 96.885 159.260 100.835 159.460 ;
        RECT 96.885 158.660 97.235 159.260 ;
        RECT 84.435 158.060 100.835 158.660 ;
        RECT 87.085 157.460 89.385 157.510 ;
        RECT 95.885 157.460 98.185 157.510 ;
        RECT 101.835 157.460 102.235 161.110 ;
        RECT 83.035 157.060 102.235 157.460 ;
        RECT 103.035 157.460 103.435 161.110 ;
        RECT 108.035 161.060 108.385 161.660 ;
        RECT 104.435 160.860 108.385 161.060 ;
        RECT 108.035 160.260 108.385 160.860 ;
        RECT 104.435 160.060 108.385 160.260 ;
        RECT 108.035 159.460 108.385 160.060 ;
        RECT 104.435 159.260 108.385 159.460 ;
        RECT 108.035 158.660 108.385 159.260 ;
        RECT 108.985 158.660 109.185 166.260 ;
        RECT 109.785 158.660 109.985 166.260 ;
        RECT 110.585 158.660 110.785 166.260 ;
        RECT 111.385 158.660 111.585 166.260 ;
        RECT 112.185 158.660 113.085 174.660 ;
        RECT 113.685 167.060 113.885 174.660 ;
        RECT 114.485 167.060 114.685 174.660 ;
        RECT 115.285 167.060 115.485 174.660 ;
        RECT 116.085 167.060 116.285 174.660 ;
        RECT 116.885 174.060 117.235 174.660 ;
        RECT 116.885 173.860 120.835 174.060 ;
        RECT 116.885 173.260 117.235 173.860 ;
        RECT 116.885 173.060 120.835 173.260 ;
        RECT 116.885 172.460 117.235 173.060 ;
        RECT 116.885 172.260 120.835 172.460 ;
        RECT 116.885 171.660 117.235 172.260 ;
        RECT 121.835 172.210 122.235 175.860 ;
        RECT 116.885 171.460 120.835 171.660 ;
        RECT 116.885 170.860 117.235 171.460 ;
        RECT 116.885 170.660 120.835 170.860 ;
        RECT 116.885 170.060 117.235 170.660 ;
        RECT 116.885 169.860 120.835 170.060 ;
        RECT 121.785 169.915 127.140 172.210 ;
        RECT 121.785 169.910 127.005 169.915 ;
        RECT 116.885 169.260 117.235 169.860 ;
        RECT 116.885 169.060 120.835 169.260 ;
        RECT 116.885 168.460 117.235 169.060 ;
        RECT 116.885 168.260 120.835 168.460 ;
        RECT 116.885 167.660 117.235 168.260 ;
        RECT 116.885 167.460 120.835 167.660 ;
        RECT 116.885 167.060 117.235 167.460 ;
        RECT 113.685 158.660 113.885 166.260 ;
        RECT 114.485 158.660 114.685 166.260 ;
        RECT 115.285 158.660 115.485 166.260 ;
        RECT 116.085 158.660 116.285 166.260 ;
        RECT 116.885 165.860 117.235 166.260 ;
        RECT 116.885 165.660 120.835 165.860 ;
        RECT 116.885 165.060 117.235 165.660 ;
        RECT 116.885 164.860 120.835 165.060 ;
        RECT 116.885 164.260 117.235 164.860 ;
        RECT 116.885 164.060 120.835 164.260 ;
        RECT 116.885 163.460 117.235 164.060 ;
        RECT 116.885 163.260 120.835 163.460 ;
        RECT 121.835 163.410 122.235 169.910 ;
        RECT 116.885 162.660 117.235 163.260 ;
        RECT 116.885 162.460 120.835 162.660 ;
        RECT 116.885 161.860 117.235 162.460 ;
        RECT 116.885 161.660 120.835 161.860 ;
        RECT 116.885 161.060 117.235 161.660 ;
        RECT 121.785 161.115 127.140 163.410 ;
        RECT 121.785 161.110 127.005 161.115 ;
        RECT 116.885 160.860 120.835 161.060 ;
        RECT 116.885 160.260 117.235 160.860 ;
        RECT 116.885 160.060 120.835 160.260 ;
        RECT 116.885 159.460 117.235 160.060 ;
        RECT 116.885 159.260 120.835 159.460 ;
        RECT 116.885 158.660 117.235 159.260 ;
        RECT 104.435 158.060 120.835 158.660 ;
        RECT 107.085 157.460 109.385 157.510 ;
        RECT 115.885 157.460 118.185 157.510 ;
        RECT 121.835 157.460 122.235 161.110 ;
        RECT 103.035 157.060 122.235 157.460 ;
        RECT 47.085 156.660 49.385 157.060 ;
        RECT 55.885 156.660 58.185 157.060 ;
        RECT 67.085 156.660 69.385 157.060 ;
        RECT 75.885 156.660 78.185 157.060 ;
        RECT 87.085 156.660 89.385 157.060 ;
        RECT 95.885 156.660 98.185 157.060 ;
        RECT 107.085 156.660 109.385 157.060 ;
        RECT 115.885 156.660 118.185 157.060 ;
        RECT 2.515 141.130 2.875 141.510 ;
        RECT 3.145 141.130 3.505 141.510 ;
        RECT 3.745 141.130 4.105 141.510 ;
        RECT 125.340 141.130 125.700 141.510 ;
        RECT 125.970 141.130 126.330 141.510 ;
        RECT 126.570 141.130 126.930 141.510 ;
        RECT 2.515 140.540 2.875 140.920 ;
        RECT 3.145 140.540 3.505 140.920 ;
        RECT 3.745 140.540 4.105 140.920 ;
        RECT 125.340 140.540 125.700 140.920 ;
        RECT 125.970 140.540 126.330 140.920 ;
        RECT 126.570 140.540 126.930 140.920 ;
        RECT 9.180 139.600 11.480 140.000 ;
        RECT 17.980 139.600 20.280 140.000 ;
        RECT 29.180 139.600 31.480 140.000 ;
        RECT 37.980 139.600 40.280 140.000 ;
        RECT 49.180 139.600 51.480 140.000 ;
        RECT 57.980 139.600 60.280 140.000 ;
        RECT 69.180 139.600 71.480 140.000 ;
        RECT 77.980 139.600 80.280 140.000 ;
        RECT 89.180 139.600 91.480 140.000 ;
        RECT 97.980 139.600 100.280 140.000 ;
        RECT 109.180 139.600 111.480 140.000 ;
        RECT 117.980 139.600 120.280 140.000 ;
        RECT 5.130 139.200 24.330 139.600 ;
        RECT 2.515 137.220 2.875 137.600 ;
        RECT 3.145 137.220 3.505 137.600 ;
        RECT 3.745 137.220 4.105 137.600 ;
        RECT 2.515 136.630 2.875 137.010 ;
        RECT 3.145 136.630 3.505 137.010 ;
        RECT 3.745 136.630 4.105 137.010 ;
        RECT 2.425 135.550 4.235 135.555 ;
        RECT 5.130 135.550 5.530 139.200 ;
        RECT 9.180 139.150 11.480 139.200 ;
        RECT 17.980 139.150 20.280 139.200 ;
        RECT 6.530 138.000 22.930 138.600 ;
        RECT 10.130 137.400 10.480 138.000 ;
        RECT 6.530 137.200 10.480 137.400 ;
        RECT 10.130 136.600 10.480 137.200 ;
        RECT 6.530 136.400 10.480 136.600 ;
        RECT 10.130 135.800 10.480 136.400 ;
        RECT 6.530 135.600 10.480 135.800 ;
        RECT 2.315 133.255 5.580 135.550 ;
        RECT 10.130 135.000 10.480 135.600 ;
        RECT 6.530 134.800 10.480 135.000 ;
        RECT 10.130 134.200 10.480 134.800 ;
        RECT 6.530 134.000 10.480 134.200 ;
        RECT 10.130 133.400 10.480 134.000 ;
        RECT 4.730 133.250 5.580 133.255 ;
        RECT 5.130 126.750 5.530 133.250 ;
        RECT 6.530 133.200 10.480 133.400 ;
        RECT 10.130 132.600 10.480 133.200 ;
        RECT 6.530 132.400 10.480 132.600 ;
        RECT 10.130 131.800 10.480 132.400 ;
        RECT 6.530 131.600 10.480 131.800 ;
        RECT 10.130 131.000 10.480 131.600 ;
        RECT 6.530 130.800 10.480 131.000 ;
        RECT 10.130 130.400 10.480 130.800 ;
        RECT 11.080 130.400 11.280 138.000 ;
        RECT 11.880 130.400 12.080 138.000 ;
        RECT 12.680 130.400 12.880 138.000 ;
        RECT 13.480 130.400 13.680 138.000 ;
        RECT 10.130 129.200 10.480 129.600 ;
        RECT 6.530 129.000 10.480 129.200 ;
        RECT 10.130 128.400 10.480 129.000 ;
        RECT 6.530 128.200 10.480 128.400 ;
        RECT 10.130 127.600 10.480 128.200 ;
        RECT 6.530 127.400 10.480 127.600 ;
        RECT 10.130 126.800 10.480 127.400 ;
        RECT 2.315 124.450 5.580 126.750 ;
        RECT 6.530 126.600 10.480 126.800 ;
        RECT 10.130 126.000 10.480 126.600 ;
        RECT 6.530 125.800 10.480 126.000 ;
        RECT 10.130 125.200 10.480 125.800 ;
        RECT 6.530 125.000 10.480 125.200 ;
        RECT 2.315 124.425 4.315 124.450 ;
        RECT 2.315 124.420 4.310 124.425 ;
        RECT 2.515 122.660 2.875 123.040 ;
        RECT 3.145 122.660 3.505 123.040 ;
        RECT 3.745 122.660 4.105 123.040 ;
        RECT 2.515 122.070 2.875 122.450 ;
        RECT 3.145 122.070 3.505 122.450 ;
        RECT 3.745 122.070 4.105 122.450 ;
        RECT 5.130 120.800 5.530 124.450 ;
        RECT 10.130 124.400 10.480 125.000 ;
        RECT 6.530 124.200 10.480 124.400 ;
        RECT 10.130 123.600 10.480 124.200 ;
        RECT 6.530 123.400 10.480 123.600 ;
        RECT 10.130 122.800 10.480 123.400 ;
        RECT 6.530 122.600 10.480 122.800 ;
        RECT 10.130 122.000 10.480 122.600 ;
        RECT 11.080 122.000 11.280 129.600 ;
        RECT 11.880 122.000 12.080 129.600 ;
        RECT 12.680 122.000 12.880 129.600 ;
        RECT 13.480 122.000 13.680 129.600 ;
        RECT 14.280 122.000 15.180 138.000 ;
        RECT 15.780 130.400 15.980 138.000 ;
        RECT 16.580 130.400 16.780 138.000 ;
        RECT 17.380 130.400 17.580 138.000 ;
        RECT 18.180 130.400 18.380 138.000 ;
        RECT 18.980 137.400 19.330 138.000 ;
        RECT 18.980 137.200 22.930 137.400 ;
        RECT 18.980 136.600 19.330 137.200 ;
        RECT 18.980 136.400 22.930 136.600 ;
        RECT 18.980 135.800 19.330 136.400 ;
        RECT 18.980 135.600 22.930 135.800 ;
        RECT 18.980 135.000 19.330 135.600 ;
        RECT 23.930 135.550 24.330 139.200 ;
        RECT 25.130 139.200 44.330 139.600 ;
        RECT 25.130 135.550 25.530 139.200 ;
        RECT 29.180 139.150 31.480 139.200 ;
        RECT 37.980 139.150 40.280 139.200 ;
        RECT 26.530 138.000 42.930 138.600 ;
        RECT 30.130 137.400 30.480 138.000 ;
        RECT 26.530 137.200 30.480 137.400 ;
        RECT 30.130 136.600 30.480 137.200 ;
        RECT 26.530 136.400 30.480 136.600 ;
        RECT 30.130 135.800 30.480 136.400 ;
        RECT 26.530 135.600 30.480 135.800 ;
        RECT 18.980 134.800 22.930 135.000 ;
        RECT 18.980 134.200 19.330 134.800 ;
        RECT 18.980 134.000 22.930 134.200 ;
        RECT 18.980 133.400 19.330 134.000 ;
        RECT 18.980 133.200 22.930 133.400 ;
        RECT 23.880 133.250 25.580 135.550 ;
        RECT 30.130 135.000 30.480 135.600 ;
        RECT 26.530 134.800 30.480 135.000 ;
        RECT 30.130 134.200 30.480 134.800 ;
        RECT 26.530 134.000 30.480 134.200 ;
        RECT 30.130 133.400 30.480 134.000 ;
        RECT 18.980 132.600 19.330 133.200 ;
        RECT 18.980 132.400 22.930 132.600 ;
        RECT 18.980 131.800 19.330 132.400 ;
        RECT 18.980 131.600 22.930 131.800 ;
        RECT 18.980 131.000 19.330 131.600 ;
        RECT 18.980 130.800 22.930 131.000 ;
        RECT 18.980 130.400 19.330 130.800 ;
        RECT 15.780 122.000 15.980 129.600 ;
        RECT 16.580 122.000 16.780 129.600 ;
        RECT 17.380 122.000 17.580 129.600 ;
        RECT 18.180 122.000 18.380 129.600 ;
        RECT 18.980 129.200 19.330 129.600 ;
        RECT 18.980 129.000 22.930 129.200 ;
        RECT 18.980 128.400 19.330 129.000 ;
        RECT 18.980 128.200 22.930 128.400 ;
        RECT 18.980 127.600 19.330 128.200 ;
        RECT 18.980 127.400 22.930 127.600 ;
        RECT 18.980 126.800 19.330 127.400 ;
        RECT 18.980 126.600 22.930 126.800 ;
        RECT 23.930 126.750 24.330 133.250 ;
        RECT 25.130 126.750 25.530 133.250 ;
        RECT 26.530 133.200 30.480 133.400 ;
        RECT 30.130 132.600 30.480 133.200 ;
        RECT 26.530 132.400 30.480 132.600 ;
        RECT 30.130 131.800 30.480 132.400 ;
        RECT 26.530 131.600 30.480 131.800 ;
        RECT 30.130 131.000 30.480 131.600 ;
        RECT 26.530 130.800 30.480 131.000 ;
        RECT 30.130 130.400 30.480 130.800 ;
        RECT 31.080 130.400 31.280 138.000 ;
        RECT 31.880 130.400 32.080 138.000 ;
        RECT 32.680 130.400 32.880 138.000 ;
        RECT 33.480 130.400 33.680 138.000 ;
        RECT 30.130 129.200 30.480 129.600 ;
        RECT 26.530 129.000 30.480 129.200 ;
        RECT 30.130 128.400 30.480 129.000 ;
        RECT 26.530 128.200 30.480 128.400 ;
        RECT 30.130 127.600 30.480 128.200 ;
        RECT 26.530 127.400 30.480 127.600 ;
        RECT 30.130 126.800 30.480 127.400 ;
        RECT 18.980 126.000 19.330 126.600 ;
        RECT 18.980 125.800 22.930 126.000 ;
        RECT 18.980 125.200 19.330 125.800 ;
        RECT 18.980 125.000 22.930 125.200 ;
        RECT 18.980 124.400 19.330 125.000 ;
        RECT 23.880 124.450 25.580 126.750 ;
        RECT 26.530 126.600 30.480 126.800 ;
        RECT 30.130 126.000 30.480 126.600 ;
        RECT 26.530 125.800 30.480 126.000 ;
        RECT 30.130 125.200 30.480 125.800 ;
        RECT 26.530 125.000 30.480 125.200 ;
        RECT 18.980 124.200 22.930 124.400 ;
        RECT 18.980 123.600 19.330 124.200 ;
        RECT 18.980 123.400 22.930 123.600 ;
        RECT 18.980 122.800 19.330 123.400 ;
        RECT 18.980 122.600 22.930 122.800 ;
        RECT 18.980 122.000 19.330 122.600 ;
        RECT 6.530 121.400 22.930 122.000 ;
        RECT 9.180 120.800 11.480 120.850 ;
        RECT 17.980 120.800 20.280 120.850 ;
        RECT 23.930 120.800 24.330 124.450 ;
        RECT 5.130 120.400 24.330 120.800 ;
        RECT 25.130 120.800 25.530 124.450 ;
        RECT 30.130 124.400 30.480 125.000 ;
        RECT 26.530 124.200 30.480 124.400 ;
        RECT 30.130 123.600 30.480 124.200 ;
        RECT 26.530 123.400 30.480 123.600 ;
        RECT 30.130 122.800 30.480 123.400 ;
        RECT 26.530 122.600 30.480 122.800 ;
        RECT 30.130 122.000 30.480 122.600 ;
        RECT 31.080 122.000 31.280 129.600 ;
        RECT 31.880 122.000 32.080 129.600 ;
        RECT 32.680 122.000 32.880 129.600 ;
        RECT 33.480 122.000 33.680 129.600 ;
        RECT 34.280 122.000 35.180 138.000 ;
        RECT 35.780 130.400 35.980 138.000 ;
        RECT 36.580 130.400 36.780 138.000 ;
        RECT 37.380 130.400 37.580 138.000 ;
        RECT 38.180 130.400 38.380 138.000 ;
        RECT 38.980 137.400 39.330 138.000 ;
        RECT 38.980 137.200 42.930 137.400 ;
        RECT 38.980 136.600 39.330 137.200 ;
        RECT 38.980 136.400 42.930 136.600 ;
        RECT 38.980 135.800 39.330 136.400 ;
        RECT 38.980 135.600 42.930 135.800 ;
        RECT 38.980 135.000 39.330 135.600 ;
        RECT 43.930 135.550 44.330 139.200 ;
        RECT 45.130 139.200 64.330 139.600 ;
        RECT 45.130 135.550 45.530 139.200 ;
        RECT 49.180 139.150 51.480 139.200 ;
        RECT 57.980 139.150 60.280 139.200 ;
        RECT 46.530 138.000 62.930 138.600 ;
        RECT 50.130 137.400 50.480 138.000 ;
        RECT 46.530 137.200 50.480 137.400 ;
        RECT 50.130 136.600 50.480 137.200 ;
        RECT 46.530 136.400 50.480 136.600 ;
        RECT 50.130 135.800 50.480 136.400 ;
        RECT 46.530 135.600 50.480 135.800 ;
        RECT 38.980 134.800 42.930 135.000 ;
        RECT 38.980 134.200 39.330 134.800 ;
        RECT 38.980 134.000 42.930 134.200 ;
        RECT 38.980 133.400 39.330 134.000 ;
        RECT 38.980 133.200 42.930 133.400 ;
        RECT 43.880 133.250 45.580 135.550 ;
        RECT 50.130 135.000 50.480 135.600 ;
        RECT 46.530 134.800 50.480 135.000 ;
        RECT 50.130 134.200 50.480 134.800 ;
        RECT 46.530 134.000 50.480 134.200 ;
        RECT 50.130 133.400 50.480 134.000 ;
        RECT 38.980 132.600 39.330 133.200 ;
        RECT 38.980 132.400 42.930 132.600 ;
        RECT 38.980 131.800 39.330 132.400 ;
        RECT 38.980 131.600 42.930 131.800 ;
        RECT 38.980 131.000 39.330 131.600 ;
        RECT 38.980 130.800 42.930 131.000 ;
        RECT 38.980 130.400 39.330 130.800 ;
        RECT 35.780 122.000 35.980 129.600 ;
        RECT 36.580 122.000 36.780 129.600 ;
        RECT 37.380 122.000 37.580 129.600 ;
        RECT 38.180 122.000 38.380 129.600 ;
        RECT 38.980 129.200 39.330 129.600 ;
        RECT 38.980 129.000 42.930 129.200 ;
        RECT 38.980 128.400 39.330 129.000 ;
        RECT 38.980 128.200 42.930 128.400 ;
        RECT 38.980 127.600 39.330 128.200 ;
        RECT 38.980 127.400 42.930 127.600 ;
        RECT 38.980 126.800 39.330 127.400 ;
        RECT 38.980 126.600 42.930 126.800 ;
        RECT 43.930 126.750 44.330 133.250 ;
        RECT 45.130 126.750 45.530 133.250 ;
        RECT 46.530 133.200 50.480 133.400 ;
        RECT 50.130 132.600 50.480 133.200 ;
        RECT 46.530 132.400 50.480 132.600 ;
        RECT 50.130 131.800 50.480 132.400 ;
        RECT 46.530 131.600 50.480 131.800 ;
        RECT 50.130 131.000 50.480 131.600 ;
        RECT 46.530 130.800 50.480 131.000 ;
        RECT 50.130 130.400 50.480 130.800 ;
        RECT 51.080 130.400 51.280 138.000 ;
        RECT 51.880 130.400 52.080 138.000 ;
        RECT 52.680 130.400 52.880 138.000 ;
        RECT 53.480 130.400 53.680 138.000 ;
        RECT 50.130 129.200 50.480 129.600 ;
        RECT 46.530 129.000 50.480 129.200 ;
        RECT 50.130 128.400 50.480 129.000 ;
        RECT 46.530 128.200 50.480 128.400 ;
        RECT 50.130 127.600 50.480 128.200 ;
        RECT 46.530 127.400 50.480 127.600 ;
        RECT 50.130 126.800 50.480 127.400 ;
        RECT 38.980 126.000 39.330 126.600 ;
        RECT 38.980 125.800 42.930 126.000 ;
        RECT 38.980 125.200 39.330 125.800 ;
        RECT 38.980 125.000 42.930 125.200 ;
        RECT 38.980 124.400 39.330 125.000 ;
        RECT 43.880 124.450 45.580 126.750 ;
        RECT 46.530 126.600 50.480 126.800 ;
        RECT 50.130 126.000 50.480 126.600 ;
        RECT 46.530 125.800 50.480 126.000 ;
        RECT 50.130 125.200 50.480 125.800 ;
        RECT 46.530 125.000 50.480 125.200 ;
        RECT 38.980 124.200 42.930 124.400 ;
        RECT 38.980 123.600 39.330 124.200 ;
        RECT 38.980 123.400 42.930 123.600 ;
        RECT 38.980 122.800 39.330 123.400 ;
        RECT 38.980 122.600 42.930 122.800 ;
        RECT 38.980 122.000 39.330 122.600 ;
        RECT 26.530 121.400 42.930 122.000 ;
        RECT 29.180 120.800 31.480 120.850 ;
        RECT 37.980 120.800 40.280 120.850 ;
        RECT 43.930 120.800 44.330 124.450 ;
        RECT 25.130 120.400 44.330 120.800 ;
        RECT 45.130 120.800 45.530 124.450 ;
        RECT 50.130 124.400 50.480 125.000 ;
        RECT 46.530 124.200 50.480 124.400 ;
        RECT 50.130 123.600 50.480 124.200 ;
        RECT 46.530 123.400 50.480 123.600 ;
        RECT 50.130 122.800 50.480 123.400 ;
        RECT 46.530 122.600 50.480 122.800 ;
        RECT 50.130 122.000 50.480 122.600 ;
        RECT 51.080 122.000 51.280 129.600 ;
        RECT 51.880 122.000 52.080 129.600 ;
        RECT 52.680 122.000 52.880 129.600 ;
        RECT 53.480 122.000 53.680 129.600 ;
        RECT 54.280 122.000 55.180 138.000 ;
        RECT 55.780 130.400 55.980 138.000 ;
        RECT 56.580 130.400 56.780 138.000 ;
        RECT 57.380 130.400 57.580 138.000 ;
        RECT 58.180 130.400 58.380 138.000 ;
        RECT 58.980 137.400 59.330 138.000 ;
        RECT 58.980 137.200 62.930 137.400 ;
        RECT 58.980 136.600 59.330 137.200 ;
        RECT 58.980 136.400 62.930 136.600 ;
        RECT 58.980 135.800 59.330 136.400 ;
        RECT 58.980 135.600 62.930 135.800 ;
        RECT 58.980 135.000 59.330 135.600 ;
        RECT 63.930 135.550 64.330 139.200 ;
        RECT 65.130 139.200 84.330 139.600 ;
        RECT 65.130 135.550 65.530 139.200 ;
        RECT 69.180 139.150 71.480 139.200 ;
        RECT 77.980 139.150 80.280 139.200 ;
        RECT 66.530 138.000 82.930 138.600 ;
        RECT 70.130 137.400 70.480 138.000 ;
        RECT 66.530 137.200 70.480 137.400 ;
        RECT 70.130 136.600 70.480 137.200 ;
        RECT 66.530 136.400 70.480 136.600 ;
        RECT 70.130 135.800 70.480 136.400 ;
        RECT 66.530 135.600 70.480 135.800 ;
        RECT 58.980 134.800 62.930 135.000 ;
        RECT 58.980 134.200 59.330 134.800 ;
        RECT 58.980 134.000 62.930 134.200 ;
        RECT 58.980 133.400 59.330 134.000 ;
        RECT 58.980 133.200 62.930 133.400 ;
        RECT 63.880 133.250 65.580 135.550 ;
        RECT 70.130 135.000 70.480 135.600 ;
        RECT 66.530 134.800 70.480 135.000 ;
        RECT 70.130 134.200 70.480 134.800 ;
        RECT 66.530 134.000 70.480 134.200 ;
        RECT 70.130 133.400 70.480 134.000 ;
        RECT 58.980 132.600 59.330 133.200 ;
        RECT 58.980 132.400 62.930 132.600 ;
        RECT 58.980 131.800 59.330 132.400 ;
        RECT 58.980 131.600 62.930 131.800 ;
        RECT 58.980 131.000 59.330 131.600 ;
        RECT 58.980 130.800 62.930 131.000 ;
        RECT 58.980 130.400 59.330 130.800 ;
        RECT 55.780 122.000 55.980 129.600 ;
        RECT 56.580 122.000 56.780 129.600 ;
        RECT 57.380 122.000 57.580 129.600 ;
        RECT 58.180 122.000 58.380 129.600 ;
        RECT 58.980 129.200 59.330 129.600 ;
        RECT 58.980 129.000 62.930 129.200 ;
        RECT 58.980 128.400 59.330 129.000 ;
        RECT 58.980 128.200 62.930 128.400 ;
        RECT 58.980 127.600 59.330 128.200 ;
        RECT 58.980 127.400 62.930 127.600 ;
        RECT 58.980 126.800 59.330 127.400 ;
        RECT 58.980 126.600 62.930 126.800 ;
        RECT 63.930 126.750 64.330 133.250 ;
        RECT 65.130 126.750 65.530 133.250 ;
        RECT 66.530 133.200 70.480 133.400 ;
        RECT 70.130 132.600 70.480 133.200 ;
        RECT 66.530 132.400 70.480 132.600 ;
        RECT 70.130 131.800 70.480 132.400 ;
        RECT 66.530 131.600 70.480 131.800 ;
        RECT 70.130 131.000 70.480 131.600 ;
        RECT 66.530 130.800 70.480 131.000 ;
        RECT 70.130 130.400 70.480 130.800 ;
        RECT 71.080 130.400 71.280 138.000 ;
        RECT 71.880 130.400 72.080 138.000 ;
        RECT 72.680 130.400 72.880 138.000 ;
        RECT 73.480 130.400 73.680 138.000 ;
        RECT 70.130 129.200 70.480 129.600 ;
        RECT 66.530 129.000 70.480 129.200 ;
        RECT 70.130 128.400 70.480 129.000 ;
        RECT 66.530 128.200 70.480 128.400 ;
        RECT 70.130 127.600 70.480 128.200 ;
        RECT 66.530 127.400 70.480 127.600 ;
        RECT 70.130 126.800 70.480 127.400 ;
        RECT 58.980 126.000 59.330 126.600 ;
        RECT 58.980 125.800 62.930 126.000 ;
        RECT 58.980 125.200 59.330 125.800 ;
        RECT 58.980 125.000 62.930 125.200 ;
        RECT 58.980 124.400 59.330 125.000 ;
        RECT 63.880 124.450 65.580 126.750 ;
        RECT 66.530 126.600 70.480 126.800 ;
        RECT 70.130 126.000 70.480 126.600 ;
        RECT 66.530 125.800 70.480 126.000 ;
        RECT 70.130 125.200 70.480 125.800 ;
        RECT 66.530 125.000 70.480 125.200 ;
        RECT 58.980 124.200 62.930 124.400 ;
        RECT 58.980 123.600 59.330 124.200 ;
        RECT 58.980 123.400 62.930 123.600 ;
        RECT 58.980 122.800 59.330 123.400 ;
        RECT 58.980 122.600 62.930 122.800 ;
        RECT 58.980 122.000 59.330 122.600 ;
        RECT 46.530 121.400 62.930 122.000 ;
        RECT 49.180 120.800 51.480 120.850 ;
        RECT 57.980 120.800 60.280 120.850 ;
        RECT 63.930 120.800 64.330 124.450 ;
        RECT 45.130 120.400 64.330 120.800 ;
        RECT 65.130 120.800 65.530 124.450 ;
        RECT 70.130 124.400 70.480 125.000 ;
        RECT 66.530 124.200 70.480 124.400 ;
        RECT 70.130 123.600 70.480 124.200 ;
        RECT 66.530 123.400 70.480 123.600 ;
        RECT 70.130 122.800 70.480 123.400 ;
        RECT 66.530 122.600 70.480 122.800 ;
        RECT 70.130 122.000 70.480 122.600 ;
        RECT 71.080 122.000 71.280 129.600 ;
        RECT 71.880 122.000 72.080 129.600 ;
        RECT 72.680 122.000 72.880 129.600 ;
        RECT 73.480 122.000 73.680 129.600 ;
        RECT 74.280 122.000 75.180 138.000 ;
        RECT 75.780 130.400 75.980 138.000 ;
        RECT 76.580 130.400 76.780 138.000 ;
        RECT 77.380 130.400 77.580 138.000 ;
        RECT 78.180 130.400 78.380 138.000 ;
        RECT 78.980 137.400 79.330 138.000 ;
        RECT 78.980 137.200 82.930 137.400 ;
        RECT 78.980 136.600 79.330 137.200 ;
        RECT 78.980 136.400 82.930 136.600 ;
        RECT 78.980 135.800 79.330 136.400 ;
        RECT 78.980 135.600 82.930 135.800 ;
        RECT 78.980 135.000 79.330 135.600 ;
        RECT 83.930 135.550 84.330 139.200 ;
        RECT 85.130 139.200 104.330 139.600 ;
        RECT 85.130 135.550 85.530 139.200 ;
        RECT 89.180 139.150 91.480 139.200 ;
        RECT 97.980 139.150 100.280 139.200 ;
        RECT 86.530 138.000 102.930 138.600 ;
        RECT 90.130 137.400 90.480 138.000 ;
        RECT 86.530 137.200 90.480 137.400 ;
        RECT 90.130 136.600 90.480 137.200 ;
        RECT 86.530 136.400 90.480 136.600 ;
        RECT 90.130 135.800 90.480 136.400 ;
        RECT 86.530 135.600 90.480 135.800 ;
        RECT 78.980 134.800 82.930 135.000 ;
        RECT 78.980 134.200 79.330 134.800 ;
        RECT 78.980 134.000 82.930 134.200 ;
        RECT 78.980 133.400 79.330 134.000 ;
        RECT 78.980 133.200 82.930 133.400 ;
        RECT 83.880 133.250 85.580 135.550 ;
        RECT 90.130 135.000 90.480 135.600 ;
        RECT 86.530 134.800 90.480 135.000 ;
        RECT 90.130 134.200 90.480 134.800 ;
        RECT 86.530 134.000 90.480 134.200 ;
        RECT 90.130 133.400 90.480 134.000 ;
        RECT 78.980 132.600 79.330 133.200 ;
        RECT 78.980 132.400 82.930 132.600 ;
        RECT 78.980 131.800 79.330 132.400 ;
        RECT 78.980 131.600 82.930 131.800 ;
        RECT 78.980 131.000 79.330 131.600 ;
        RECT 78.980 130.800 82.930 131.000 ;
        RECT 78.980 130.400 79.330 130.800 ;
        RECT 75.780 122.000 75.980 129.600 ;
        RECT 76.580 122.000 76.780 129.600 ;
        RECT 77.380 122.000 77.580 129.600 ;
        RECT 78.180 122.000 78.380 129.600 ;
        RECT 78.980 129.200 79.330 129.600 ;
        RECT 78.980 129.000 82.930 129.200 ;
        RECT 78.980 128.400 79.330 129.000 ;
        RECT 78.980 128.200 82.930 128.400 ;
        RECT 78.980 127.600 79.330 128.200 ;
        RECT 78.980 127.400 82.930 127.600 ;
        RECT 78.980 126.800 79.330 127.400 ;
        RECT 78.980 126.600 82.930 126.800 ;
        RECT 83.930 126.750 84.330 133.250 ;
        RECT 85.130 126.750 85.530 133.250 ;
        RECT 86.530 133.200 90.480 133.400 ;
        RECT 90.130 132.600 90.480 133.200 ;
        RECT 86.530 132.400 90.480 132.600 ;
        RECT 90.130 131.800 90.480 132.400 ;
        RECT 86.530 131.600 90.480 131.800 ;
        RECT 90.130 131.000 90.480 131.600 ;
        RECT 86.530 130.800 90.480 131.000 ;
        RECT 90.130 130.400 90.480 130.800 ;
        RECT 91.080 130.400 91.280 138.000 ;
        RECT 91.880 130.400 92.080 138.000 ;
        RECT 92.680 130.400 92.880 138.000 ;
        RECT 93.480 130.400 93.680 138.000 ;
        RECT 90.130 129.200 90.480 129.600 ;
        RECT 86.530 129.000 90.480 129.200 ;
        RECT 90.130 128.400 90.480 129.000 ;
        RECT 86.530 128.200 90.480 128.400 ;
        RECT 90.130 127.600 90.480 128.200 ;
        RECT 86.530 127.400 90.480 127.600 ;
        RECT 90.130 126.800 90.480 127.400 ;
        RECT 78.980 126.000 79.330 126.600 ;
        RECT 78.980 125.800 82.930 126.000 ;
        RECT 78.980 125.200 79.330 125.800 ;
        RECT 78.980 125.000 82.930 125.200 ;
        RECT 78.980 124.400 79.330 125.000 ;
        RECT 83.880 124.450 85.580 126.750 ;
        RECT 86.530 126.600 90.480 126.800 ;
        RECT 90.130 126.000 90.480 126.600 ;
        RECT 86.530 125.800 90.480 126.000 ;
        RECT 90.130 125.200 90.480 125.800 ;
        RECT 86.530 125.000 90.480 125.200 ;
        RECT 78.980 124.200 82.930 124.400 ;
        RECT 78.980 123.600 79.330 124.200 ;
        RECT 78.980 123.400 82.930 123.600 ;
        RECT 78.980 122.800 79.330 123.400 ;
        RECT 78.980 122.600 82.930 122.800 ;
        RECT 78.980 122.000 79.330 122.600 ;
        RECT 66.530 121.400 82.930 122.000 ;
        RECT 69.180 120.800 71.480 120.850 ;
        RECT 77.980 120.800 80.280 120.850 ;
        RECT 83.930 120.800 84.330 124.450 ;
        RECT 65.130 120.400 84.330 120.800 ;
        RECT 85.130 120.800 85.530 124.450 ;
        RECT 90.130 124.400 90.480 125.000 ;
        RECT 86.530 124.200 90.480 124.400 ;
        RECT 90.130 123.600 90.480 124.200 ;
        RECT 86.530 123.400 90.480 123.600 ;
        RECT 90.130 122.800 90.480 123.400 ;
        RECT 86.530 122.600 90.480 122.800 ;
        RECT 90.130 122.000 90.480 122.600 ;
        RECT 91.080 122.000 91.280 129.600 ;
        RECT 91.880 122.000 92.080 129.600 ;
        RECT 92.680 122.000 92.880 129.600 ;
        RECT 93.480 122.000 93.680 129.600 ;
        RECT 94.280 122.000 95.180 138.000 ;
        RECT 95.780 130.400 95.980 138.000 ;
        RECT 96.580 130.400 96.780 138.000 ;
        RECT 97.380 130.400 97.580 138.000 ;
        RECT 98.180 130.400 98.380 138.000 ;
        RECT 98.980 137.400 99.330 138.000 ;
        RECT 98.980 137.200 102.930 137.400 ;
        RECT 98.980 136.600 99.330 137.200 ;
        RECT 98.980 136.400 102.930 136.600 ;
        RECT 98.980 135.800 99.330 136.400 ;
        RECT 98.980 135.600 102.930 135.800 ;
        RECT 98.980 135.000 99.330 135.600 ;
        RECT 103.930 135.550 104.330 139.200 ;
        RECT 105.130 139.200 124.330 139.600 ;
        RECT 105.130 135.550 105.530 139.200 ;
        RECT 109.180 139.150 111.480 139.200 ;
        RECT 117.980 139.150 120.280 139.200 ;
        RECT 106.530 138.000 122.930 138.600 ;
        RECT 110.130 137.400 110.480 138.000 ;
        RECT 106.530 137.200 110.480 137.400 ;
        RECT 110.130 136.600 110.480 137.200 ;
        RECT 106.530 136.400 110.480 136.600 ;
        RECT 110.130 135.800 110.480 136.400 ;
        RECT 106.530 135.600 110.480 135.800 ;
        RECT 98.980 134.800 102.930 135.000 ;
        RECT 98.980 134.200 99.330 134.800 ;
        RECT 98.980 134.000 102.930 134.200 ;
        RECT 98.980 133.400 99.330 134.000 ;
        RECT 98.980 133.200 102.930 133.400 ;
        RECT 103.880 133.250 105.580 135.550 ;
        RECT 110.130 135.000 110.480 135.600 ;
        RECT 106.530 134.800 110.480 135.000 ;
        RECT 110.130 134.200 110.480 134.800 ;
        RECT 106.530 134.000 110.480 134.200 ;
        RECT 110.130 133.400 110.480 134.000 ;
        RECT 98.980 132.600 99.330 133.200 ;
        RECT 98.980 132.400 102.930 132.600 ;
        RECT 98.980 131.800 99.330 132.400 ;
        RECT 98.980 131.600 102.930 131.800 ;
        RECT 98.980 131.000 99.330 131.600 ;
        RECT 98.980 130.800 102.930 131.000 ;
        RECT 98.980 130.400 99.330 130.800 ;
        RECT 95.780 122.000 95.980 129.600 ;
        RECT 96.580 122.000 96.780 129.600 ;
        RECT 97.380 122.000 97.580 129.600 ;
        RECT 98.180 122.000 98.380 129.600 ;
        RECT 98.980 129.200 99.330 129.600 ;
        RECT 98.980 129.000 102.930 129.200 ;
        RECT 98.980 128.400 99.330 129.000 ;
        RECT 98.980 128.200 102.930 128.400 ;
        RECT 98.980 127.600 99.330 128.200 ;
        RECT 98.980 127.400 102.930 127.600 ;
        RECT 98.980 126.800 99.330 127.400 ;
        RECT 98.980 126.600 102.930 126.800 ;
        RECT 103.930 126.750 104.330 133.250 ;
        RECT 105.130 126.750 105.530 133.250 ;
        RECT 106.530 133.200 110.480 133.400 ;
        RECT 110.130 132.600 110.480 133.200 ;
        RECT 106.530 132.400 110.480 132.600 ;
        RECT 110.130 131.800 110.480 132.400 ;
        RECT 106.530 131.600 110.480 131.800 ;
        RECT 110.130 131.000 110.480 131.600 ;
        RECT 106.530 130.800 110.480 131.000 ;
        RECT 110.130 130.400 110.480 130.800 ;
        RECT 111.080 130.400 111.280 138.000 ;
        RECT 111.880 130.400 112.080 138.000 ;
        RECT 112.680 130.400 112.880 138.000 ;
        RECT 113.480 130.400 113.680 138.000 ;
        RECT 110.130 129.200 110.480 129.600 ;
        RECT 106.530 129.000 110.480 129.200 ;
        RECT 110.130 128.400 110.480 129.000 ;
        RECT 106.530 128.200 110.480 128.400 ;
        RECT 110.130 127.600 110.480 128.200 ;
        RECT 106.530 127.400 110.480 127.600 ;
        RECT 110.130 126.800 110.480 127.400 ;
        RECT 98.980 126.000 99.330 126.600 ;
        RECT 98.980 125.800 102.930 126.000 ;
        RECT 98.980 125.200 99.330 125.800 ;
        RECT 98.980 125.000 102.930 125.200 ;
        RECT 98.980 124.400 99.330 125.000 ;
        RECT 103.880 124.450 105.580 126.750 ;
        RECT 106.530 126.600 110.480 126.800 ;
        RECT 110.130 126.000 110.480 126.600 ;
        RECT 106.530 125.800 110.480 126.000 ;
        RECT 110.130 125.200 110.480 125.800 ;
        RECT 106.530 125.000 110.480 125.200 ;
        RECT 98.980 124.200 102.930 124.400 ;
        RECT 98.980 123.600 99.330 124.200 ;
        RECT 98.980 123.400 102.930 123.600 ;
        RECT 98.980 122.800 99.330 123.400 ;
        RECT 98.980 122.600 102.930 122.800 ;
        RECT 98.980 122.000 99.330 122.600 ;
        RECT 86.530 121.400 102.930 122.000 ;
        RECT 89.180 120.800 91.480 120.850 ;
        RECT 97.980 120.800 100.280 120.850 ;
        RECT 103.930 120.800 104.330 124.450 ;
        RECT 85.130 120.400 104.330 120.800 ;
        RECT 105.130 120.800 105.530 124.450 ;
        RECT 110.130 124.400 110.480 125.000 ;
        RECT 106.530 124.200 110.480 124.400 ;
        RECT 110.130 123.600 110.480 124.200 ;
        RECT 106.530 123.400 110.480 123.600 ;
        RECT 110.130 122.800 110.480 123.400 ;
        RECT 106.530 122.600 110.480 122.800 ;
        RECT 110.130 122.000 110.480 122.600 ;
        RECT 111.080 122.000 111.280 129.600 ;
        RECT 111.880 122.000 112.080 129.600 ;
        RECT 112.680 122.000 112.880 129.600 ;
        RECT 113.480 122.000 113.680 129.600 ;
        RECT 114.280 122.000 115.180 138.000 ;
        RECT 115.780 130.400 115.980 138.000 ;
        RECT 116.580 130.400 116.780 138.000 ;
        RECT 117.380 130.400 117.580 138.000 ;
        RECT 118.180 130.400 118.380 138.000 ;
        RECT 118.980 137.400 119.330 138.000 ;
        RECT 118.980 137.200 122.930 137.400 ;
        RECT 118.980 136.600 119.330 137.200 ;
        RECT 118.980 136.400 122.930 136.600 ;
        RECT 118.980 135.800 119.330 136.400 ;
        RECT 118.980 135.600 122.930 135.800 ;
        RECT 118.980 135.000 119.330 135.600 ;
        RECT 123.930 135.550 124.330 139.200 ;
        RECT 125.340 137.220 125.700 137.600 ;
        RECT 125.970 137.220 126.330 137.600 ;
        RECT 126.570 137.220 126.930 137.600 ;
        RECT 125.340 136.630 125.700 137.010 ;
        RECT 125.970 136.630 126.330 137.010 ;
        RECT 126.570 136.630 126.930 137.010 ;
        RECT 118.980 134.800 122.930 135.000 ;
        RECT 118.980 134.200 119.330 134.800 ;
        RECT 118.980 134.000 122.930 134.200 ;
        RECT 118.980 133.400 119.330 134.000 ;
        RECT 118.980 133.200 122.930 133.400 ;
        RECT 123.880 133.250 124.730 135.550 ;
        RECT 118.980 132.600 119.330 133.200 ;
        RECT 118.980 132.400 122.930 132.600 ;
        RECT 118.980 131.800 119.330 132.400 ;
        RECT 118.980 131.600 122.930 131.800 ;
        RECT 118.980 131.000 119.330 131.600 ;
        RECT 118.980 130.800 122.930 131.000 ;
        RECT 118.980 130.400 119.330 130.800 ;
        RECT 115.780 122.000 115.980 129.600 ;
        RECT 116.580 122.000 116.780 129.600 ;
        RECT 117.380 122.000 117.580 129.600 ;
        RECT 118.180 122.000 118.380 129.600 ;
        RECT 118.980 129.200 119.330 129.600 ;
        RECT 118.980 129.000 122.930 129.200 ;
        RECT 118.980 128.400 119.330 129.000 ;
        RECT 118.980 128.200 122.930 128.400 ;
        RECT 118.980 127.600 119.330 128.200 ;
        RECT 118.980 127.400 122.930 127.600 ;
        RECT 118.980 126.800 119.330 127.400 ;
        RECT 118.980 126.600 122.930 126.800 ;
        RECT 123.930 126.750 124.330 133.250 ;
        RECT 118.980 126.000 119.330 126.600 ;
        RECT 118.980 125.800 122.930 126.000 ;
        RECT 118.980 125.200 119.330 125.800 ;
        RECT 118.980 125.000 122.930 125.200 ;
        RECT 118.980 124.400 119.330 125.000 ;
        RECT 123.880 124.450 124.730 126.750 ;
        RECT 118.980 124.200 122.930 124.400 ;
        RECT 118.980 123.600 119.330 124.200 ;
        RECT 118.980 123.400 122.930 123.600 ;
        RECT 118.980 122.800 119.330 123.400 ;
        RECT 118.980 122.600 122.930 122.800 ;
        RECT 118.980 122.000 119.330 122.600 ;
        RECT 106.530 121.400 122.930 122.000 ;
        RECT 109.180 120.800 111.480 120.850 ;
        RECT 117.980 120.800 120.280 120.850 ;
        RECT 123.930 120.800 124.330 124.450 ;
        RECT 125.340 122.415 125.700 122.795 ;
        RECT 125.970 122.415 126.330 122.795 ;
        RECT 126.570 122.415 126.930 122.795 ;
        RECT 125.340 121.825 125.700 122.205 ;
        RECT 125.970 121.825 126.330 122.205 ;
        RECT 126.570 121.825 126.930 122.205 ;
        RECT 105.130 120.400 124.330 120.800 ;
        RECT 9.180 119.600 11.480 120.400 ;
        RECT 17.980 119.600 20.280 120.400 ;
        RECT 29.180 119.600 31.480 120.400 ;
        RECT 37.980 119.600 40.280 120.400 ;
        RECT 49.180 119.600 51.480 120.400 ;
        RECT 57.980 119.600 60.280 120.400 ;
        RECT 69.180 119.600 71.480 120.400 ;
        RECT 77.980 119.600 80.280 120.400 ;
        RECT 89.180 119.600 91.480 120.400 ;
        RECT 97.980 119.600 100.280 120.400 ;
        RECT 109.180 119.600 111.480 120.400 ;
        RECT 117.980 119.600 120.280 120.400 ;
        RECT 5.130 119.200 24.330 119.600 ;
        RECT 2.515 117.640 2.875 118.020 ;
        RECT 3.145 117.640 3.505 118.020 ;
        RECT 3.745 117.640 4.105 118.020 ;
        RECT 2.515 117.050 2.875 117.430 ;
        RECT 3.145 117.050 3.505 117.430 ;
        RECT 3.745 117.050 4.105 117.430 ;
        RECT 5.130 115.550 5.530 119.200 ;
        RECT 9.180 119.150 11.480 119.200 ;
        RECT 17.980 119.150 20.280 119.200 ;
        RECT 6.530 118.000 22.930 118.600 ;
        RECT 10.130 117.400 10.480 118.000 ;
        RECT 6.530 117.200 10.480 117.400 ;
        RECT 10.130 116.600 10.480 117.200 ;
        RECT 6.530 116.400 10.480 116.600 ;
        RECT 10.130 115.800 10.480 116.400 ;
        RECT 6.530 115.600 10.480 115.800 ;
        RECT 4.730 115.545 5.580 115.550 ;
        RECT 2.315 113.250 5.580 115.545 ;
        RECT 10.130 115.000 10.480 115.600 ;
        RECT 6.530 114.800 10.480 115.000 ;
        RECT 10.130 114.200 10.480 114.800 ;
        RECT 6.530 114.000 10.480 114.200 ;
        RECT 10.130 113.400 10.480 114.000 ;
        RECT 5.130 106.750 5.530 113.250 ;
        RECT 6.530 113.200 10.480 113.400 ;
        RECT 10.130 112.600 10.480 113.200 ;
        RECT 6.530 112.400 10.480 112.600 ;
        RECT 10.130 111.800 10.480 112.400 ;
        RECT 6.530 111.600 10.480 111.800 ;
        RECT 10.130 111.000 10.480 111.600 ;
        RECT 6.530 110.800 10.480 111.000 ;
        RECT 10.130 110.400 10.480 110.800 ;
        RECT 11.080 110.400 11.280 118.000 ;
        RECT 11.880 110.400 12.080 118.000 ;
        RECT 12.680 110.400 12.880 118.000 ;
        RECT 13.480 110.400 13.680 118.000 ;
        RECT 10.130 109.200 10.480 109.600 ;
        RECT 6.530 109.000 10.480 109.200 ;
        RECT 10.130 108.400 10.480 109.000 ;
        RECT 6.530 108.200 10.480 108.400 ;
        RECT 10.130 107.600 10.480 108.200 ;
        RECT 6.530 107.400 10.480 107.600 ;
        RECT 10.130 106.800 10.480 107.400 ;
        RECT 4.730 106.745 5.580 106.750 ;
        RECT 2.315 104.450 5.580 106.745 ;
        RECT 6.530 106.600 10.480 106.800 ;
        RECT 10.130 106.000 10.480 106.600 ;
        RECT 6.530 105.800 10.480 106.000 ;
        RECT 10.130 105.200 10.480 105.800 ;
        RECT 6.530 105.000 10.480 105.200 ;
        RECT 2.515 102.750 2.875 103.130 ;
        RECT 3.145 102.750 3.505 103.130 ;
        RECT 3.745 102.750 4.105 103.130 ;
        RECT 2.515 102.160 2.875 102.540 ;
        RECT 3.145 102.160 3.505 102.540 ;
        RECT 3.745 102.160 4.105 102.540 ;
        RECT 5.130 100.800 5.530 104.450 ;
        RECT 10.130 104.400 10.480 105.000 ;
        RECT 6.530 104.200 10.480 104.400 ;
        RECT 10.130 103.600 10.480 104.200 ;
        RECT 6.530 103.400 10.480 103.600 ;
        RECT 10.130 102.800 10.480 103.400 ;
        RECT 6.530 102.600 10.480 102.800 ;
        RECT 10.130 102.000 10.480 102.600 ;
        RECT 11.080 102.000 11.280 109.600 ;
        RECT 11.880 102.000 12.080 109.600 ;
        RECT 12.680 102.000 12.880 109.600 ;
        RECT 13.480 102.000 13.680 109.600 ;
        RECT 14.280 102.000 15.180 118.000 ;
        RECT 15.780 110.400 15.980 118.000 ;
        RECT 16.580 110.400 16.780 118.000 ;
        RECT 17.380 110.400 17.580 118.000 ;
        RECT 18.180 110.400 18.380 118.000 ;
        RECT 18.980 117.400 19.330 118.000 ;
        RECT 18.980 117.200 22.930 117.400 ;
        RECT 18.980 116.600 19.330 117.200 ;
        RECT 18.980 116.400 22.930 116.600 ;
        RECT 18.980 115.800 19.330 116.400 ;
        RECT 18.980 115.600 22.930 115.800 ;
        RECT 18.980 115.000 19.330 115.600 ;
        RECT 23.930 115.550 24.330 119.200 ;
        RECT 25.130 119.200 44.330 119.600 ;
        RECT 25.130 115.550 25.530 119.200 ;
        RECT 29.180 119.150 31.480 119.200 ;
        RECT 37.980 119.150 40.280 119.200 ;
        RECT 26.530 118.000 42.930 118.600 ;
        RECT 30.130 117.400 30.480 118.000 ;
        RECT 26.530 117.200 30.480 117.400 ;
        RECT 30.130 116.600 30.480 117.200 ;
        RECT 26.530 116.400 30.480 116.600 ;
        RECT 30.130 115.800 30.480 116.400 ;
        RECT 26.530 115.600 30.480 115.800 ;
        RECT 18.980 114.800 22.930 115.000 ;
        RECT 18.980 114.200 19.330 114.800 ;
        RECT 18.980 114.000 22.930 114.200 ;
        RECT 18.980 113.400 19.330 114.000 ;
        RECT 18.980 113.200 22.930 113.400 ;
        RECT 23.880 113.250 25.580 115.550 ;
        RECT 30.130 115.000 30.480 115.600 ;
        RECT 26.530 114.800 30.480 115.000 ;
        RECT 30.130 114.200 30.480 114.800 ;
        RECT 26.530 114.000 30.480 114.200 ;
        RECT 30.130 113.400 30.480 114.000 ;
        RECT 18.980 112.600 19.330 113.200 ;
        RECT 18.980 112.400 22.930 112.600 ;
        RECT 18.980 111.800 19.330 112.400 ;
        RECT 18.980 111.600 22.930 111.800 ;
        RECT 18.980 111.000 19.330 111.600 ;
        RECT 18.980 110.800 22.930 111.000 ;
        RECT 18.980 110.400 19.330 110.800 ;
        RECT 15.780 102.000 15.980 109.600 ;
        RECT 16.580 102.000 16.780 109.600 ;
        RECT 17.380 102.000 17.580 109.600 ;
        RECT 18.180 102.000 18.380 109.600 ;
        RECT 18.980 109.200 19.330 109.600 ;
        RECT 18.980 109.000 22.930 109.200 ;
        RECT 18.980 108.400 19.330 109.000 ;
        RECT 18.980 108.200 22.930 108.400 ;
        RECT 18.980 107.600 19.330 108.200 ;
        RECT 18.980 107.400 22.930 107.600 ;
        RECT 18.980 106.800 19.330 107.400 ;
        RECT 18.980 106.600 22.930 106.800 ;
        RECT 23.930 106.750 24.330 113.250 ;
        RECT 25.130 106.750 25.530 113.250 ;
        RECT 26.530 113.200 30.480 113.400 ;
        RECT 30.130 112.600 30.480 113.200 ;
        RECT 26.530 112.400 30.480 112.600 ;
        RECT 30.130 111.800 30.480 112.400 ;
        RECT 26.530 111.600 30.480 111.800 ;
        RECT 30.130 111.000 30.480 111.600 ;
        RECT 26.530 110.800 30.480 111.000 ;
        RECT 30.130 110.400 30.480 110.800 ;
        RECT 31.080 110.400 31.280 118.000 ;
        RECT 31.880 110.400 32.080 118.000 ;
        RECT 32.680 110.400 32.880 118.000 ;
        RECT 33.480 110.400 33.680 118.000 ;
        RECT 30.130 109.200 30.480 109.600 ;
        RECT 26.530 109.000 30.480 109.200 ;
        RECT 30.130 108.400 30.480 109.000 ;
        RECT 26.530 108.200 30.480 108.400 ;
        RECT 30.130 107.600 30.480 108.200 ;
        RECT 26.530 107.400 30.480 107.600 ;
        RECT 30.130 106.800 30.480 107.400 ;
        RECT 18.980 106.000 19.330 106.600 ;
        RECT 18.980 105.800 22.930 106.000 ;
        RECT 18.980 105.200 19.330 105.800 ;
        RECT 18.980 105.000 22.930 105.200 ;
        RECT 18.980 104.400 19.330 105.000 ;
        RECT 23.880 104.450 25.580 106.750 ;
        RECT 26.530 106.600 30.480 106.800 ;
        RECT 30.130 106.000 30.480 106.600 ;
        RECT 26.530 105.800 30.480 106.000 ;
        RECT 30.130 105.200 30.480 105.800 ;
        RECT 26.530 105.000 30.480 105.200 ;
        RECT 18.980 104.200 22.930 104.400 ;
        RECT 18.980 103.600 19.330 104.200 ;
        RECT 18.980 103.400 22.930 103.600 ;
        RECT 18.980 102.800 19.330 103.400 ;
        RECT 18.980 102.600 22.930 102.800 ;
        RECT 18.980 102.000 19.330 102.600 ;
        RECT 6.530 101.400 22.930 102.000 ;
        RECT 9.180 100.800 11.480 100.850 ;
        RECT 17.980 100.800 20.280 100.850 ;
        RECT 23.930 100.800 24.330 104.450 ;
        RECT 5.130 100.400 24.330 100.800 ;
        RECT 25.130 100.800 25.530 104.450 ;
        RECT 30.130 104.400 30.480 105.000 ;
        RECT 26.530 104.200 30.480 104.400 ;
        RECT 30.130 103.600 30.480 104.200 ;
        RECT 26.530 103.400 30.480 103.600 ;
        RECT 30.130 102.800 30.480 103.400 ;
        RECT 26.530 102.600 30.480 102.800 ;
        RECT 30.130 102.000 30.480 102.600 ;
        RECT 31.080 102.000 31.280 109.600 ;
        RECT 31.880 102.000 32.080 109.600 ;
        RECT 32.680 102.000 32.880 109.600 ;
        RECT 33.480 102.000 33.680 109.600 ;
        RECT 34.280 102.000 35.180 118.000 ;
        RECT 35.780 110.400 35.980 118.000 ;
        RECT 36.580 110.400 36.780 118.000 ;
        RECT 37.380 110.400 37.580 118.000 ;
        RECT 38.180 110.400 38.380 118.000 ;
        RECT 38.980 117.400 39.330 118.000 ;
        RECT 38.980 117.200 42.930 117.400 ;
        RECT 38.980 116.600 39.330 117.200 ;
        RECT 38.980 116.400 42.930 116.600 ;
        RECT 38.980 115.800 39.330 116.400 ;
        RECT 38.980 115.600 42.930 115.800 ;
        RECT 38.980 115.000 39.330 115.600 ;
        RECT 43.930 115.550 44.330 119.200 ;
        RECT 45.130 119.200 64.330 119.600 ;
        RECT 45.130 115.550 45.530 119.200 ;
        RECT 49.180 119.150 51.480 119.200 ;
        RECT 57.980 119.150 60.280 119.200 ;
        RECT 46.530 118.000 62.930 118.600 ;
        RECT 50.130 117.400 50.480 118.000 ;
        RECT 46.530 117.200 50.480 117.400 ;
        RECT 50.130 116.600 50.480 117.200 ;
        RECT 46.530 116.400 50.480 116.600 ;
        RECT 50.130 115.800 50.480 116.400 ;
        RECT 46.530 115.600 50.480 115.800 ;
        RECT 38.980 114.800 42.930 115.000 ;
        RECT 38.980 114.200 39.330 114.800 ;
        RECT 38.980 114.000 42.930 114.200 ;
        RECT 38.980 113.400 39.330 114.000 ;
        RECT 38.980 113.200 42.930 113.400 ;
        RECT 43.880 113.250 45.580 115.550 ;
        RECT 50.130 115.000 50.480 115.600 ;
        RECT 46.530 114.800 50.480 115.000 ;
        RECT 50.130 114.200 50.480 114.800 ;
        RECT 46.530 114.000 50.480 114.200 ;
        RECT 50.130 113.400 50.480 114.000 ;
        RECT 38.980 112.600 39.330 113.200 ;
        RECT 38.980 112.400 42.930 112.600 ;
        RECT 38.980 111.800 39.330 112.400 ;
        RECT 38.980 111.600 42.930 111.800 ;
        RECT 38.980 111.000 39.330 111.600 ;
        RECT 38.980 110.800 42.930 111.000 ;
        RECT 38.980 110.400 39.330 110.800 ;
        RECT 35.780 102.000 35.980 109.600 ;
        RECT 36.580 102.000 36.780 109.600 ;
        RECT 37.380 102.000 37.580 109.600 ;
        RECT 38.180 102.000 38.380 109.600 ;
        RECT 38.980 109.200 39.330 109.600 ;
        RECT 38.980 109.000 42.930 109.200 ;
        RECT 38.980 108.400 39.330 109.000 ;
        RECT 38.980 108.200 42.930 108.400 ;
        RECT 38.980 107.600 39.330 108.200 ;
        RECT 38.980 107.400 42.930 107.600 ;
        RECT 38.980 106.800 39.330 107.400 ;
        RECT 38.980 106.600 42.930 106.800 ;
        RECT 43.930 106.750 44.330 113.250 ;
        RECT 45.130 106.750 45.530 113.250 ;
        RECT 46.530 113.200 50.480 113.400 ;
        RECT 50.130 112.600 50.480 113.200 ;
        RECT 46.530 112.400 50.480 112.600 ;
        RECT 50.130 111.800 50.480 112.400 ;
        RECT 46.530 111.600 50.480 111.800 ;
        RECT 50.130 111.000 50.480 111.600 ;
        RECT 46.530 110.800 50.480 111.000 ;
        RECT 50.130 110.400 50.480 110.800 ;
        RECT 51.080 110.400 51.280 118.000 ;
        RECT 51.880 110.400 52.080 118.000 ;
        RECT 52.680 110.400 52.880 118.000 ;
        RECT 53.480 110.400 53.680 118.000 ;
        RECT 50.130 109.200 50.480 109.600 ;
        RECT 46.530 109.000 50.480 109.200 ;
        RECT 50.130 108.400 50.480 109.000 ;
        RECT 46.530 108.200 50.480 108.400 ;
        RECT 50.130 107.600 50.480 108.200 ;
        RECT 46.530 107.400 50.480 107.600 ;
        RECT 50.130 106.800 50.480 107.400 ;
        RECT 38.980 106.000 39.330 106.600 ;
        RECT 38.980 105.800 42.930 106.000 ;
        RECT 38.980 105.200 39.330 105.800 ;
        RECT 38.980 105.000 42.930 105.200 ;
        RECT 38.980 104.400 39.330 105.000 ;
        RECT 43.880 104.450 45.580 106.750 ;
        RECT 46.530 106.600 50.480 106.800 ;
        RECT 50.130 106.000 50.480 106.600 ;
        RECT 46.530 105.800 50.480 106.000 ;
        RECT 50.130 105.200 50.480 105.800 ;
        RECT 46.530 105.000 50.480 105.200 ;
        RECT 38.980 104.200 42.930 104.400 ;
        RECT 38.980 103.600 39.330 104.200 ;
        RECT 38.980 103.400 42.930 103.600 ;
        RECT 38.980 102.800 39.330 103.400 ;
        RECT 38.980 102.600 42.930 102.800 ;
        RECT 38.980 102.000 39.330 102.600 ;
        RECT 26.530 101.400 42.930 102.000 ;
        RECT 29.180 100.800 31.480 100.850 ;
        RECT 37.980 100.800 40.280 100.850 ;
        RECT 43.930 100.800 44.330 104.450 ;
        RECT 25.130 100.400 44.330 100.800 ;
        RECT 45.130 100.800 45.530 104.450 ;
        RECT 50.130 104.400 50.480 105.000 ;
        RECT 46.530 104.200 50.480 104.400 ;
        RECT 50.130 103.600 50.480 104.200 ;
        RECT 46.530 103.400 50.480 103.600 ;
        RECT 50.130 102.800 50.480 103.400 ;
        RECT 46.530 102.600 50.480 102.800 ;
        RECT 50.130 102.000 50.480 102.600 ;
        RECT 51.080 102.000 51.280 109.600 ;
        RECT 51.880 102.000 52.080 109.600 ;
        RECT 52.680 102.000 52.880 109.600 ;
        RECT 53.480 102.000 53.680 109.600 ;
        RECT 54.280 102.000 55.180 118.000 ;
        RECT 55.780 110.400 55.980 118.000 ;
        RECT 56.580 110.400 56.780 118.000 ;
        RECT 57.380 110.400 57.580 118.000 ;
        RECT 58.180 110.400 58.380 118.000 ;
        RECT 58.980 117.400 59.330 118.000 ;
        RECT 58.980 117.200 62.930 117.400 ;
        RECT 58.980 116.600 59.330 117.200 ;
        RECT 58.980 116.400 62.930 116.600 ;
        RECT 58.980 115.800 59.330 116.400 ;
        RECT 58.980 115.600 62.930 115.800 ;
        RECT 58.980 115.000 59.330 115.600 ;
        RECT 63.930 115.550 64.330 119.200 ;
        RECT 65.130 119.200 84.330 119.600 ;
        RECT 65.130 115.550 65.530 119.200 ;
        RECT 69.180 119.150 71.480 119.200 ;
        RECT 77.980 119.150 80.280 119.200 ;
        RECT 66.530 118.000 82.930 118.600 ;
        RECT 70.130 117.400 70.480 118.000 ;
        RECT 66.530 117.200 70.480 117.400 ;
        RECT 70.130 116.600 70.480 117.200 ;
        RECT 66.530 116.400 70.480 116.600 ;
        RECT 70.130 115.800 70.480 116.400 ;
        RECT 66.530 115.600 70.480 115.800 ;
        RECT 58.980 114.800 62.930 115.000 ;
        RECT 58.980 114.200 59.330 114.800 ;
        RECT 58.980 114.000 62.930 114.200 ;
        RECT 58.980 113.400 59.330 114.000 ;
        RECT 58.980 113.200 62.930 113.400 ;
        RECT 63.880 113.250 65.580 115.550 ;
        RECT 70.130 115.000 70.480 115.600 ;
        RECT 66.530 114.800 70.480 115.000 ;
        RECT 70.130 114.200 70.480 114.800 ;
        RECT 66.530 114.000 70.480 114.200 ;
        RECT 70.130 113.400 70.480 114.000 ;
        RECT 58.980 112.600 59.330 113.200 ;
        RECT 58.980 112.400 62.930 112.600 ;
        RECT 58.980 111.800 59.330 112.400 ;
        RECT 58.980 111.600 62.930 111.800 ;
        RECT 58.980 111.000 59.330 111.600 ;
        RECT 58.980 110.800 62.930 111.000 ;
        RECT 58.980 110.400 59.330 110.800 ;
        RECT 55.780 102.000 55.980 109.600 ;
        RECT 56.580 102.000 56.780 109.600 ;
        RECT 57.380 102.000 57.580 109.600 ;
        RECT 58.180 102.000 58.380 109.600 ;
        RECT 58.980 109.200 59.330 109.600 ;
        RECT 58.980 109.000 62.930 109.200 ;
        RECT 58.980 108.400 59.330 109.000 ;
        RECT 58.980 108.200 62.930 108.400 ;
        RECT 58.980 107.600 59.330 108.200 ;
        RECT 58.980 107.400 62.930 107.600 ;
        RECT 58.980 106.800 59.330 107.400 ;
        RECT 58.980 106.600 62.930 106.800 ;
        RECT 63.930 106.750 64.330 113.250 ;
        RECT 65.130 106.750 65.530 113.250 ;
        RECT 66.530 113.200 70.480 113.400 ;
        RECT 70.130 112.600 70.480 113.200 ;
        RECT 66.530 112.400 70.480 112.600 ;
        RECT 70.130 111.800 70.480 112.400 ;
        RECT 66.530 111.600 70.480 111.800 ;
        RECT 70.130 111.000 70.480 111.600 ;
        RECT 66.530 110.800 70.480 111.000 ;
        RECT 70.130 110.400 70.480 110.800 ;
        RECT 71.080 110.400 71.280 118.000 ;
        RECT 71.880 110.400 72.080 118.000 ;
        RECT 72.680 110.400 72.880 118.000 ;
        RECT 73.480 110.400 73.680 118.000 ;
        RECT 70.130 109.200 70.480 109.600 ;
        RECT 66.530 109.000 70.480 109.200 ;
        RECT 70.130 108.400 70.480 109.000 ;
        RECT 66.530 108.200 70.480 108.400 ;
        RECT 70.130 107.600 70.480 108.200 ;
        RECT 66.530 107.400 70.480 107.600 ;
        RECT 70.130 106.800 70.480 107.400 ;
        RECT 58.980 106.000 59.330 106.600 ;
        RECT 58.980 105.800 62.930 106.000 ;
        RECT 58.980 105.200 59.330 105.800 ;
        RECT 58.980 105.000 62.930 105.200 ;
        RECT 58.980 104.400 59.330 105.000 ;
        RECT 63.880 104.450 65.580 106.750 ;
        RECT 66.530 106.600 70.480 106.800 ;
        RECT 70.130 106.000 70.480 106.600 ;
        RECT 66.530 105.800 70.480 106.000 ;
        RECT 70.130 105.200 70.480 105.800 ;
        RECT 66.530 105.000 70.480 105.200 ;
        RECT 58.980 104.200 62.930 104.400 ;
        RECT 58.980 103.600 59.330 104.200 ;
        RECT 58.980 103.400 62.930 103.600 ;
        RECT 58.980 102.800 59.330 103.400 ;
        RECT 58.980 102.600 62.930 102.800 ;
        RECT 58.980 102.000 59.330 102.600 ;
        RECT 46.530 101.400 62.930 102.000 ;
        RECT 49.180 100.800 51.480 100.850 ;
        RECT 57.980 100.800 60.280 100.850 ;
        RECT 63.930 100.800 64.330 104.450 ;
        RECT 45.130 100.400 64.330 100.800 ;
        RECT 65.130 100.800 65.530 104.450 ;
        RECT 70.130 104.400 70.480 105.000 ;
        RECT 66.530 104.200 70.480 104.400 ;
        RECT 70.130 103.600 70.480 104.200 ;
        RECT 66.530 103.400 70.480 103.600 ;
        RECT 70.130 102.800 70.480 103.400 ;
        RECT 66.530 102.600 70.480 102.800 ;
        RECT 70.130 102.000 70.480 102.600 ;
        RECT 71.080 102.000 71.280 109.600 ;
        RECT 71.880 102.000 72.080 109.600 ;
        RECT 72.680 102.000 72.880 109.600 ;
        RECT 73.480 102.000 73.680 109.600 ;
        RECT 74.280 102.000 75.180 118.000 ;
        RECT 75.780 110.400 75.980 118.000 ;
        RECT 76.580 110.400 76.780 118.000 ;
        RECT 77.380 110.400 77.580 118.000 ;
        RECT 78.180 110.400 78.380 118.000 ;
        RECT 78.980 117.400 79.330 118.000 ;
        RECT 78.980 117.200 82.930 117.400 ;
        RECT 78.980 116.600 79.330 117.200 ;
        RECT 78.980 116.400 82.930 116.600 ;
        RECT 78.980 115.800 79.330 116.400 ;
        RECT 78.980 115.600 82.930 115.800 ;
        RECT 78.980 115.000 79.330 115.600 ;
        RECT 83.930 115.550 84.330 119.200 ;
        RECT 85.130 119.200 104.330 119.600 ;
        RECT 85.130 115.550 85.530 119.200 ;
        RECT 89.180 119.150 91.480 119.200 ;
        RECT 97.980 119.150 100.280 119.200 ;
        RECT 86.530 118.000 102.930 118.600 ;
        RECT 90.130 117.400 90.480 118.000 ;
        RECT 86.530 117.200 90.480 117.400 ;
        RECT 90.130 116.600 90.480 117.200 ;
        RECT 86.530 116.400 90.480 116.600 ;
        RECT 90.130 115.800 90.480 116.400 ;
        RECT 86.530 115.600 90.480 115.800 ;
        RECT 78.980 114.800 82.930 115.000 ;
        RECT 78.980 114.200 79.330 114.800 ;
        RECT 78.980 114.000 82.930 114.200 ;
        RECT 78.980 113.400 79.330 114.000 ;
        RECT 78.980 113.200 82.930 113.400 ;
        RECT 83.880 113.250 85.580 115.550 ;
        RECT 90.130 115.000 90.480 115.600 ;
        RECT 86.530 114.800 90.480 115.000 ;
        RECT 90.130 114.200 90.480 114.800 ;
        RECT 86.530 114.000 90.480 114.200 ;
        RECT 90.130 113.400 90.480 114.000 ;
        RECT 78.980 112.600 79.330 113.200 ;
        RECT 78.980 112.400 82.930 112.600 ;
        RECT 78.980 111.800 79.330 112.400 ;
        RECT 78.980 111.600 82.930 111.800 ;
        RECT 78.980 111.000 79.330 111.600 ;
        RECT 78.980 110.800 82.930 111.000 ;
        RECT 78.980 110.400 79.330 110.800 ;
        RECT 75.780 102.000 75.980 109.600 ;
        RECT 76.580 102.000 76.780 109.600 ;
        RECT 77.380 102.000 77.580 109.600 ;
        RECT 78.180 102.000 78.380 109.600 ;
        RECT 78.980 109.200 79.330 109.600 ;
        RECT 78.980 109.000 82.930 109.200 ;
        RECT 78.980 108.400 79.330 109.000 ;
        RECT 78.980 108.200 82.930 108.400 ;
        RECT 78.980 107.600 79.330 108.200 ;
        RECT 78.980 107.400 82.930 107.600 ;
        RECT 78.980 106.800 79.330 107.400 ;
        RECT 78.980 106.600 82.930 106.800 ;
        RECT 83.930 106.750 84.330 113.250 ;
        RECT 85.130 106.750 85.530 113.250 ;
        RECT 86.530 113.200 90.480 113.400 ;
        RECT 90.130 112.600 90.480 113.200 ;
        RECT 86.530 112.400 90.480 112.600 ;
        RECT 90.130 111.800 90.480 112.400 ;
        RECT 86.530 111.600 90.480 111.800 ;
        RECT 90.130 111.000 90.480 111.600 ;
        RECT 86.530 110.800 90.480 111.000 ;
        RECT 90.130 110.400 90.480 110.800 ;
        RECT 91.080 110.400 91.280 118.000 ;
        RECT 91.880 110.400 92.080 118.000 ;
        RECT 92.680 110.400 92.880 118.000 ;
        RECT 93.480 110.400 93.680 118.000 ;
        RECT 90.130 109.200 90.480 109.600 ;
        RECT 86.530 109.000 90.480 109.200 ;
        RECT 90.130 108.400 90.480 109.000 ;
        RECT 86.530 108.200 90.480 108.400 ;
        RECT 90.130 107.600 90.480 108.200 ;
        RECT 86.530 107.400 90.480 107.600 ;
        RECT 90.130 106.800 90.480 107.400 ;
        RECT 78.980 106.000 79.330 106.600 ;
        RECT 78.980 105.800 82.930 106.000 ;
        RECT 78.980 105.200 79.330 105.800 ;
        RECT 78.980 105.000 82.930 105.200 ;
        RECT 78.980 104.400 79.330 105.000 ;
        RECT 83.880 104.450 85.580 106.750 ;
        RECT 86.530 106.600 90.480 106.800 ;
        RECT 90.130 106.000 90.480 106.600 ;
        RECT 86.530 105.800 90.480 106.000 ;
        RECT 90.130 105.200 90.480 105.800 ;
        RECT 86.530 105.000 90.480 105.200 ;
        RECT 78.980 104.200 82.930 104.400 ;
        RECT 78.980 103.600 79.330 104.200 ;
        RECT 78.980 103.400 82.930 103.600 ;
        RECT 78.980 102.800 79.330 103.400 ;
        RECT 78.980 102.600 82.930 102.800 ;
        RECT 78.980 102.000 79.330 102.600 ;
        RECT 66.530 101.400 82.930 102.000 ;
        RECT 69.180 100.800 71.480 100.850 ;
        RECT 77.980 100.800 80.280 100.850 ;
        RECT 83.930 100.800 84.330 104.450 ;
        RECT 65.130 100.400 84.330 100.800 ;
        RECT 85.130 100.800 85.530 104.450 ;
        RECT 90.130 104.400 90.480 105.000 ;
        RECT 86.530 104.200 90.480 104.400 ;
        RECT 90.130 103.600 90.480 104.200 ;
        RECT 86.530 103.400 90.480 103.600 ;
        RECT 90.130 102.800 90.480 103.400 ;
        RECT 86.530 102.600 90.480 102.800 ;
        RECT 90.130 102.000 90.480 102.600 ;
        RECT 91.080 102.000 91.280 109.600 ;
        RECT 91.880 102.000 92.080 109.600 ;
        RECT 92.680 102.000 92.880 109.600 ;
        RECT 93.480 102.000 93.680 109.600 ;
        RECT 94.280 102.000 95.180 118.000 ;
        RECT 95.780 110.400 95.980 118.000 ;
        RECT 96.580 110.400 96.780 118.000 ;
        RECT 97.380 110.400 97.580 118.000 ;
        RECT 98.180 110.400 98.380 118.000 ;
        RECT 98.980 117.400 99.330 118.000 ;
        RECT 98.980 117.200 102.930 117.400 ;
        RECT 98.980 116.600 99.330 117.200 ;
        RECT 98.980 116.400 102.930 116.600 ;
        RECT 98.980 115.800 99.330 116.400 ;
        RECT 98.980 115.600 102.930 115.800 ;
        RECT 98.980 115.000 99.330 115.600 ;
        RECT 103.930 115.550 104.330 119.200 ;
        RECT 105.130 119.200 124.330 119.600 ;
        RECT 105.130 115.550 105.530 119.200 ;
        RECT 109.180 119.150 111.480 119.200 ;
        RECT 117.980 119.150 120.280 119.200 ;
        RECT 106.530 118.000 122.930 118.600 ;
        RECT 110.130 117.400 110.480 118.000 ;
        RECT 106.530 117.200 110.480 117.400 ;
        RECT 110.130 116.600 110.480 117.200 ;
        RECT 106.530 116.400 110.480 116.600 ;
        RECT 110.130 115.800 110.480 116.400 ;
        RECT 106.530 115.600 110.480 115.800 ;
        RECT 98.980 114.800 102.930 115.000 ;
        RECT 98.980 114.200 99.330 114.800 ;
        RECT 98.980 114.000 102.930 114.200 ;
        RECT 98.980 113.400 99.330 114.000 ;
        RECT 98.980 113.200 102.930 113.400 ;
        RECT 103.880 113.250 105.580 115.550 ;
        RECT 110.130 115.000 110.480 115.600 ;
        RECT 106.530 114.800 110.480 115.000 ;
        RECT 110.130 114.200 110.480 114.800 ;
        RECT 106.530 114.000 110.480 114.200 ;
        RECT 110.130 113.400 110.480 114.000 ;
        RECT 98.980 112.600 99.330 113.200 ;
        RECT 98.980 112.400 102.930 112.600 ;
        RECT 98.980 111.800 99.330 112.400 ;
        RECT 98.980 111.600 102.930 111.800 ;
        RECT 98.980 111.000 99.330 111.600 ;
        RECT 98.980 110.800 102.930 111.000 ;
        RECT 98.980 110.400 99.330 110.800 ;
        RECT 95.780 102.000 95.980 109.600 ;
        RECT 96.580 102.000 96.780 109.600 ;
        RECT 97.380 102.000 97.580 109.600 ;
        RECT 98.180 102.000 98.380 109.600 ;
        RECT 98.980 109.200 99.330 109.600 ;
        RECT 98.980 109.000 102.930 109.200 ;
        RECT 98.980 108.400 99.330 109.000 ;
        RECT 98.980 108.200 102.930 108.400 ;
        RECT 98.980 107.600 99.330 108.200 ;
        RECT 98.980 107.400 102.930 107.600 ;
        RECT 98.980 106.800 99.330 107.400 ;
        RECT 98.980 106.600 102.930 106.800 ;
        RECT 103.930 106.750 104.330 113.250 ;
        RECT 105.130 106.750 105.530 113.250 ;
        RECT 106.530 113.200 110.480 113.400 ;
        RECT 110.130 112.600 110.480 113.200 ;
        RECT 106.530 112.400 110.480 112.600 ;
        RECT 110.130 111.800 110.480 112.400 ;
        RECT 106.530 111.600 110.480 111.800 ;
        RECT 110.130 111.000 110.480 111.600 ;
        RECT 106.530 110.800 110.480 111.000 ;
        RECT 110.130 110.400 110.480 110.800 ;
        RECT 111.080 110.400 111.280 118.000 ;
        RECT 111.880 110.400 112.080 118.000 ;
        RECT 112.680 110.400 112.880 118.000 ;
        RECT 113.480 110.400 113.680 118.000 ;
        RECT 110.130 109.200 110.480 109.600 ;
        RECT 106.530 109.000 110.480 109.200 ;
        RECT 110.130 108.400 110.480 109.000 ;
        RECT 106.530 108.200 110.480 108.400 ;
        RECT 110.130 107.600 110.480 108.200 ;
        RECT 106.530 107.400 110.480 107.600 ;
        RECT 110.130 106.800 110.480 107.400 ;
        RECT 98.980 106.000 99.330 106.600 ;
        RECT 98.980 105.800 102.930 106.000 ;
        RECT 98.980 105.200 99.330 105.800 ;
        RECT 98.980 105.000 102.930 105.200 ;
        RECT 98.980 104.400 99.330 105.000 ;
        RECT 103.880 104.450 105.580 106.750 ;
        RECT 106.530 106.600 110.480 106.800 ;
        RECT 110.130 106.000 110.480 106.600 ;
        RECT 106.530 105.800 110.480 106.000 ;
        RECT 110.130 105.200 110.480 105.800 ;
        RECT 106.530 105.000 110.480 105.200 ;
        RECT 98.980 104.200 102.930 104.400 ;
        RECT 98.980 103.600 99.330 104.200 ;
        RECT 98.980 103.400 102.930 103.600 ;
        RECT 98.980 102.800 99.330 103.400 ;
        RECT 98.980 102.600 102.930 102.800 ;
        RECT 98.980 102.000 99.330 102.600 ;
        RECT 86.530 101.400 102.930 102.000 ;
        RECT 89.180 100.800 91.480 100.850 ;
        RECT 97.980 100.800 100.280 100.850 ;
        RECT 103.930 100.800 104.330 104.450 ;
        RECT 85.130 100.400 104.330 100.800 ;
        RECT 105.130 100.800 105.530 104.450 ;
        RECT 110.130 104.400 110.480 105.000 ;
        RECT 106.530 104.200 110.480 104.400 ;
        RECT 110.130 103.600 110.480 104.200 ;
        RECT 106.530 103.400 110.480 103.600 ;
        RECT 110.130 102.800 110.480 103.400 ;
        RECT 106.530 102.600 110.480 102.800 ;
        RECT 110.130 102.000 110.480 102.600 ;
        RECT 111.080 102.000 111.280 109.600 ;
        RECT 111.880 102.000 112.080 109.600 ;
        RECT 112.680 102.000 112.880 109.600 ;
        RECT 113.480 102.000 113.680 109.600 ;
        RECT 114.280 102.000 115.180 118.000 ;
        RECT 115.780 110.400 115.980 118.000 ;
        RECT 116.580 110.400 116.780 118.000 ;
        RECT 117.380 110.400 117.580 118.000 ;
        RECT 118.180 110.400 118.380 118.000 ;
        RECT 118.980 117.400 119.330 118.000 ;
        RECT 118.980 117.200 122.930 117.400 ;
        RECT 118.980 116.600 119.330 117.200 ;
        RECT 118.980 116.400 122.930 116.600 ;
        RECT 118.980 115.800 119.330 116.400 ;
        RECT 118.980 115.600 122.930 115.800 ;
        RECT 118.980 115.000 119.330 115.600 ;
        RECT 123.930 115.550 124.330 119.200 ;
        RECT 125.340 116.830 125.700 117.210 ;
        RECT 125.970 116.830 126.330 117.210 ;
        RECT 126.570 116.830 126.930 117.210 ;
        RECT 125.340 116.240 125.700 116.620 ;
        RECT 125.970 116.240 126.330 116.620 ;
        RECT 126.570 116.240 126.930 116.620 ;
        RECT 118.980 114.800 122.930 115.000 ;
        RECT 118.980 114.200 119.330 114.800 ;
        RECT 118.980 114.000 122.930 114.200 ;
        RECT 118.980 113.400 119.330 114.000 ;
        RECT 118.980 113.200 122.930 113.400 ;
        RECT 123.880 113.250 124.730 115.550 ;
        RECT 118.980 112.600 119.330 113.200 ;
        RECT 118.980 112.400 122.930 112.600 ;
        RECT 118.980 111.800 119.330 112.400 ;
        RECT 118.980 111.600 122.930 111.800 ;
        RECT 118.980 111.000 119.330 111.600 ;
        RECT 118.980 110.800 122.930 111.000 ;
        RECT 118.980 110.400 119.330 110.800 ;
        RECT 115.780 102.000 115.980 109.600 ;
        RECT 116.580 102.000 116.780 109.600 ;
        RECT 117.380 102.000 117.580 109.600 ;
        RECT 118.180 102.000 118.380 109.600 ;
        RECT 118.980 109.200 119.330 109.600 ;
        RECT 118.980 109.000 122.930 109.200 ;
        RECT 118.980 108.400 119.330 109.000 ;
        RECT 118.980 108.200 122.930 108.400 ;
        RECT 118.980 107.600 119.330 108.200 ;
        RECT 118.980 107.400 122.930 107.600 ;
        RECT 118.980 106.800 119.330 107.400 ;
        RECT 118.980 106.600 122.930 106.800 ;
        RECT 123.930 106.750 124.330 113.250 ;
        RECT 118.980 106.000 119.330 106.600 ;
        RECT 118.980 105.800 122.930 106.000 ;
        RECT 118.980 105.200 119.330 105.800 ;
        RECT 118.980 105.000 122.930 105.200 ;
        RECT 118.980 104.400 119.330 105.000 ;
        RECT 123.880 104.450 124.730 106.750 ;
        RECT 118.980 104.200 122.930 104.400 ;
        RECT 118.980 103.600 119.330 104.200 ;
        RECT 118.980 103.400 122.930 103.600 ;
        RECT 118.980 102.800 119.330 103.400 ;
        RECT 118.980 102.600 122.930 102.800 ;
        RECT 118.980 102.000 119.330 102.600 ;
        RECT 106.530 101.400 122.930 102.000 ;
        RECT 109.180 100.800 111.480 100.850 ;
        RECT 117.980 100.800 120.280 100.850 ;
        RECT 123.930 100.800 124.330 104.450 ;
        RECT 125.340 102.615 125.700 102.995 ;
        RECT 125.970 102.615 126.330 102.995 ;
        RECT 126.570 102.615 126.930 102.995 ;
        RECT 125.340 102.025 125.700 102.405 ;
        RECT 125.970 102.025 126.330 102.405 ;
        RECT 126.570 102.025 126.930 102.405 ;
        RECT 105.130 100.400 124.330 100.800 ;
        RECT 9.180 99.600 11.480 100.400 ;
        RECT 17.980 99.600 20.280 100.400 ;
        RECT 29.180 99.600 31.480 100.400 ;
        RECT 37.980 99.600 40.280 100.400 ;
        RECT 49.180 99.600 51.480 100.400 ;
        RECT 57.980 99.600 60.280 100.400 ;
        RECT 69.180 99.600 71.480 100.400 ;
        RECT 77.980 99.600 80.280 100.400 ;
        RECT 89.180 99.600 91.480 100.400 ;
        RECT 97.980 99.600 100.280 100.400 ;
        RECT 109.180 99.600 111.480 100.400 ;
        RECT 117.980 99.600 120.280 100.400 ;
        RECT 5.130 99.200 24.330 99.600 ;
        RECT 2.515 97.340 2.875 97.720 ;
        RECT 3.145 97.340 3.505 97.720 ;
        RECT 3.745 97.340 4.105 97.720 ;
        RECT 2.515 96.750 2.875 97.130 ;
        RECT 3.145 96.750 3.505 97.130 ;
        RECT 3.745 96.750 4.105 97.130 ;
        RECT 5.130 95.550 5.530 99.200 ;
        RECT 9.180 99.150 11.480 99.200 ;
        RECT 17.980 99.150 20.280 99.200 ;
        RECT 6.530 98.000 22.930 98.600 ;
        RECT 10.130 97.400 10.480 98.000 ;
        RECT 6.530 97.200 10.480 97.400 ;
        RECT 10.130 96.600 10.480 97.200 ;
        RECT 6.530 96.400 10.480 96.600 ;
        RECT 10.130 95.800 10.480 96.400 ;
        RECT 6.530 95.600 10.480 95.800 ;
        RECT 4.730 95.545 5.580 95.550 ;
        RECT 2.315 93.250 5.580 95.545 ;
        RECT 10.130 95.000 10.480 95.600 ;
        RECT 6.530 94.800 10.480 95.000 ;
        RECT 10.130 94.200 10.480 94.800 ;
        RECT 6.530 94.000 10.480 94.200 ;
        RECT 10.130 93.400 10.480 94.000 ;
        RECT 5.130 86.750 5.530 93.250 ;
        RECT 6.530 93.200 10.480 93.400 ;
        RECT 10.130 92.600 10.480 93.200 ;
        RECT 6.530 92.400 10.480 92.600 ;
        RECT 10.130 91.800 10.480 92.400 ;
        RECT 6.530 91.600 10.480 91.800 ;
        RECT 10.130 91.000 10.480 91.600 ;
        RECT 6.530 90.800 10.480 91.000 ;
        RECT 10.130 90.400 10.480 90.800 ;
        RECT 11.080 90.400 11.280 98.000 ;
        RECT 11.880 90.400 12.080 98.000 ;
        RECT 12.680 90.400 12.880 98.000 ;
        RECT 13.480 90.400 13.680 98.000 ;
        RECT 10.130 89.200 10.480 89.600 ;
        RECT 6.530 89.000 10.480 89.200 ;
        RECT 10.130 88.400 10.480 89.000 ;
        RECT 6.530 88.200 10.480 88.400 ;
        RECT 10.130 87.600 10.480 88.200 ;
        RECT 6.530 87.400 10.480 87.600 ;
        RECT 10.130 86.800 10.480 87.400 ;
        RECT 2.315 84.455 5.580 86.750 ;
        RECT 6.530 86.600 10.480 86.800 ;
        RECT 10.130 86.000 10.480 86.600 ;
        RECT 6.530 85.800 10.480 86.000 ;
        RECT 10.130 85.200 10.480 85.800 ;
        RECT 6.530 85.000 10.480 85.200 ;
        RECT 4.730 84.450 5.580 84.455 ;
        RECT 2.515 82.965 2.875 83.345 ;
        RECT 3.145 82.965 3.505 83.345 ;
        RECT 3.745 82.965 4.105 83.345 ;
        RECT 2.515 82.375 2.875 82.755 ;
        RECT 3.145 82.375 3.505 82.755 ;
        RECT 3.745 82.375 4.105 82.755 ;
        RECT 5.130 80.800 5.530 84.450 ;
        RECT 10.130 84.400 10.480 85.000 ;
        RECT 6.530 84.200 10.480 84.400 ;
        RECT 10.130 83.600 10.480 84.200 ;
        RECT 6.530 83.400 10.480 83.600 ;
        RECT 10.130 82.800 10.480 83.400 ;
        RECT 6.530 82.600 10.480 82.800 ;
        RECT 10.130 82.000 10.480 82.600 ;
        RECT 11.080 82.000 11.280 89.600 ;
        RECT 11.880 82.000 12.080 89.600 ;
        RECT 12.680 82.000 12.880 89.600 ;
        RECT 13.480 82.000 13.680 89.600 ;
        RECT 14.280 82.000 15.180 98.000 ;
        RECT 15.780 90.400 15.980 98.000 ;
        RECT 16.580 90.400 16.780 98.000 ;
        RECT 17.380 90.400 17.580 98.000 ;
        RECT 18.180 90.400 18.380 98.000 ;
        RECT 18.980 97.400 19.330 98.000 ;
        RECT 18.980 97.200 22.930 97.400 ;
        RECT 18.980 96.600 19.330 97.200 ;
        RECT 18.980 96.400 22.930 96.600 ;
        RECT 18.980 95.800 19.330 96.400 ;
        RECT 18.980 95.600 22.930 95.800 ;
        RECT 18.980 95.000 19.330 95.600 ;
        RECT 23.930 95.550 24.330 99.200 ;
        RECT 25.130 99.200 44.330 99.600 ;
        RECT 25.130 95.550 25.530 99.200 ;
        RECT 29.180 99.150 31.480 99.200 ;
        RECT 37.980 99.150 40.280 99.200 ;
        RECT 26.530 98.000 42.930 98.600 ;
        RECT 30.130 97.400 30.480 98.000 ;
        RECT 26.530 97.200 30.480 97.400 ;
        RECT 30.130 96.600 30.480 97.200 ;
        RECT 26.530 96.400 30.480 96.600 ;
        RECT 30.130 95.800 30.480 96.400 ;
        RECT 26.530 95.600 30.480 95.800 ;
        RECT 18.980 94.800 22.930 95.000 ;
        RECT 18.980 94.200 19.330 94.800 ;
        RECT 18.980 94.000 22.930 94.200 ;
        RECT 18.980 93.400 19.330 94.000 ;
        RECT 18.980 93.200 22.930 93.400 ;
        RECT 23.880 93.250 25.580 95.550 ;
        RECT 30.130 95.000 30.480 95.600 ;
        RECT 26.530 94.800 30.480 95.000 ;
        RECT 30.130 94.200 30.480 94.800 ;
        RECT 26.530 94.000 30.480 94.200 ;
        RECT 30.130 93.400 30.480 94.000 ;
        RECT 18.980 92.600 19.330 93.200 ;
        RECT 18.980 92.400 22.930 92.600 ;
        RECT 18.980 91.800 19.330 92.400 ;
        RECT 18.980 91.600 22.930 91.800 ;
        RECT 18.980 91.000 19.330 91.600 ;
        RECT 18.980 90.800 22.930 91.000 ;
        RECT 18.980 90.400 19.330 90.800 ;
        RECT 15.780 82.000 15.980 89.600 ;
        RECT 16.580 82.000 16.780 89.600 ;
        RECT 17.380 82.000 17.580 89.600 ;
        RECT 18.180 82.000 18.380 89.600 ;
        RECT 18.980 89.200 19.330 89.600 ;
        RECT 18.980 89.000 22.930 89.200 ;
        RECT 18.980 88.400 19.330 89.000 ;
        RECT 18.980 88.200 22.930 88.400 ;
        RECT 18.980 87.600 19.330 88.200 ;
        RECT 18.980 87.400 22.930 87.600 ;
        RECT 18.980 86.800 19.330 87.400 ;
        RECT 18.980 86.600 22.930 86.800 ;
        RECT 23.930 86.750 24.330 93.250 ;
        RECT 25.130 86.750 25.530 93.250 ;
        RECT 26.530 93.200 30.480 93.400 ;
        RECT 30.130 92.600 30.480 93.200 ;
        RECT 26.530 92.400 30.480 92.600 ;
        RECT 30.130 91.800 30.480 92.400 ;
        RECT 26.530 91.600 30.480 91.800 ;
        RECT 30.130 91.000 30.480 91.600 ;
        RECT 26.530 90.800 30.480 91.000 ;
        RECT 30.130 90.400 30.480 90.800 ;
        RECT 31.080 90.400 31.280 98.000 ;
        RECT 31.880 90.400 32.080 98.000 ;
        RECT 32.680 90.400 32.880 98.000 ;
        RECT 33.480 90.400 33.680 98.000 ;
        RECT 30.130 89.200 30.480 89.600 ;
        RECT 26.530 89.000 30.480 89.200 ;
        RECT 30.130 88.400 30.480 89.000 ;
        RECT 26.530 88.200 30.480 88.400 ;
        RECT 30.130 87.600 30.480 88.200 ;
        RECT 26.530 87.400 30.480 87.600 ;
        RECT 30.130 86.800 30.480 87.400 ;
        RECT 18.980 86.000 19.330 86.600 ;
        RECT 18.980 85.800 22.930 86.000 ;
        RECT 18.980 85.200 19.330 85.800 ;
        RECT 18.980 85.000 22.930 85.200 ;
        RECT 18.980 84.400 19.330 85.000 ;
        RECT 23.880 84.450 25.580 86.750 ;
        RECT 26.530 86.600 30.480 86.800 ;
        RECT 30.130 86.000 30.480 86.600 ;
        RECT 26.530 85.800 30.480 86.000 ;
        RECT 30.130 85.200 30.480 85.800 ;
        RECT 26.530 85.000 30.480 85.200 ;
        RECT 18.980 84.200 22.930 84.400 ;
        RECT 18.980 83.600 19.330 84.200 ;
        RECT 18.980 83.400 22.930 83.600 ;
        RECT 18.980 82.800 19.330 83.400 ;
        RECT 18.980 82.600 22.930 82.800 ;
        RECT 18.980 82.000 19.330 82.600 ;
        RECT 6.530 81.400 22.930 82.000 ;
        RECT 9.180 80.800 11.480 80.850 ;
        RECT 17.980 80.800 20.280 80.850 ;
        RECT 23.930 80.800 24.330 84.450 ;
        RECT 5.130 80.400 24.330 80.800 ;
        RECT 25.130 80.800 25.530 84.450 ;
        RECT 30.130 84.400 30.480 85.000 ;
        RECT 26.530 84.200 30.480 84.400 ;
        RECT 30.130 83.600 30.480 84.200 ;
        RECT 26.530 83.400 30.480 83.600 ;
        RECT 30.130 82.800 30.480 83.400 ;
        RECT 26.530 82.600 30.480 82.800 ;
        RECT 30.130 82.000 30.480 82.600 ;
        RECT 31.080 82.000 31.280 89.600 ;
        RECT 31.880 82.000 32.080 89.600 ;
        RECT 32.680 82.000 32.880 89.600 ;
        RECT 33.480 82.000 33.680 89.600 ;
        RECT 34.280 82.000 35.180 98.000 ;
        RECT 35.780 90.400 35.980 98.000 ;
        RECT 36.580 90.400 36.780 98.000 ;
        RECT 37.380 90.400 37.580 98.000 ;
        RECT 38.180 90.400 38.380 98.000 ;
        RECT 38.980 97.400 39.330 98.000 ;
        RECT 38.980 97.200 42.930 97.400 ;
        RECT 38.980 96.600 39.330 97.200 ;
        RECT 38.980 96.400 42.930 96.600 ;
        RECT 38.980 95.800 39.330 96.400 ;
        RECT 38.980 95.600 42.930 95.800 ;
        RECT 38.980 95.000 39.330 95.600 ;
        RECT 43.930 95.550 44.330 99.200 ;
        RECT 45.130 99.200 64.330 99.600 ;
        RECT 45.130 95.550 45.530 99.200 ;
        RECT 49.180 99.150 51.480 99.200 ;
        RECT 57.980 99.150 60.280 99.200 ;
        RECT 46.530 98.000 62.930 98.600 ;
        RECT 50.130 97.400 50.480 98.000 ;
        RECT 46.530 97.200 50.480 97.400 ;
        RECT 50.130 96.600 50.480 97.200 ;
        RECT 46.530 96.400 50.480 96.600 ;
        RECT 50.130 95.800 50.480 96.400 ;
        RECT 46.530 95.600 50.480 95.800 ;
        RECT 38.980 94.800 42.930 95.000 ;
        RECT 38.980 94.200 39.330 94.800 ;
        RECT 38.980 94.000 42.930 94.200 ;
        RECT 38.980 93.400 39.330 94.000 ;
        RECT 38.980 93.200 42.930 93.400 ;
        RECT 43.880 93.250 45.580 95.550 ;
        RECT 50.130 95.000 50.480 95.600 ;
        RECT 46.530 94.800 50.480 95.000 ;
        RECT 50.130 94.200 50.480 94.800 ;
        RECT 46.530 94.000 50.480 94.200 ;
        RECT 50.130 93.400 50.480 94.000 ;
        RECT 38.980 92.600 39.330 93.200 ;
        RECT 38.980 92.400 42.930 92.600 ;
        RECT 38.980 91.800 39.330 92.400 ;
        RECT 38.980 91.600 42.930 91.800 ;
        RECT 38.980 91.000 39.330 91.600 ;
        RECT 38.980 90.800 42.930 91.000 ;
        RECT 38.980 90.400 39.330 90.800 ;
        RECT 35.780 82.000 35.980 89.600 ;
        RECT 36.580 82.000 36.780 89.600 ;
        RECT 37.380 82.000 37.580 89.600 ;
        RECT 38.180 82.000 38.380 89.600 ;
        RECT 38.980 89.200 39.330 89.600 ;
        RECT 38.980 89.000 42.930 89.200 ;
        RECT 38.980 88.400 39.330 89.000 ;
        RECT 38.980 88.200 42.930 88.400 ;
        RECT 38.980 87.600 39.330 88.200 ;
        RECT 38.980 87.400 42.930 87.600 ;
        RECT 38.980 86.800 39.330 87.400 ;
        RECT 38.980 86.600 42.930 86.800 ;
        RECT 43.930 86.750 44.330 93.250 ;
        RECT 45.130 86.750 45.530 93.250 ;
        RECT 46.530 93.200 50.480 93.400 ;
        RECT 50.130 92.600 50.480 93.200 ;
        RECT 46.530 92.400 50.480 92.600 ;
        RECT 50.130 91.800 50.480 92.400 ;
        RECT 46.530 91.600 50.480 91.800 ;
        RECT 50.130 91.000 50.480 91.600 ;
        RECT 46.530 90.800 50.480 91.000 ;
        RECT 50.130 90.400 50.480 90.800 ;
        RECT 51.080 90.400 51.280 98.000 ;
        RECT 51.880 90.400 52.080 98.000 ;
        RECT 52.680 90.400 52.880 98.000 ;
        RECT 53.480 90.400 53.680 98.000 ;
        RECT 50.130 89.200 50.480 89.600 ;
        RECT 46.530 89.000 50.480 89.200 ;
        RECT 50.130 88.400 50.480 89.000 ;
        RECT 46.530 88.200 50.480 88.400 ;
        RECT 50.130 87.600 50.480 88.200 ;
        RECT 46.530 87.400 50.480 87.600 ;
        RECT 50.130 86.800 50.480 87.400 ;
        RECT 38.980 86.000 39.330 86.600 ;
        RECT 38.980 85.800 42.930 86.000 ;
        RECT 38.980 85.200 39.330 85.800 ;
        RECT 38.980 85.000 42.930 85.200 ;
        RECT 38.980 84.400 39.330 85.000 ;
        RECT 43.880 84.450 45.580 86.750 ;
        RECT 46.530 86.600 50.480 86.800 ;
        RECT 50.130 86.000 50.480 86.600 ;
        RECT 46.530 85.800 50.480 86.000 ;
        RECT 50.130 85.200 50.480 85.800 ;
        RECT 46.530 85.000 50.480 85.200 ;
        RECT 38.980 84.200 42.930 84.400 ;
        RECT 38.980 83.600 39.330 84.200 ;
        RECT 38.980 83.400 42.930 83.600 ;
        RECT 38.980 82.800 39.330 83.400 ;
        RECT 38.980 82.600 42.930 82.800 ;
        RECT 38.980 82.000 39.330 82.600 ;
        RECT 26.530 81.400 42.930 82.000 ;
        RECT 29.180 80.800 31.480 80.850 ;
        RECT 37.980 80.800 40.280 80.850 ;
        RECT 43.930 80.800 44.330 84.450 ;
        RECT 25.130 80.400 44.330 80.800 ;
        RECT 45.130 80.800 45.530 84.450 ;
        RECT 50.130 84.400 50.480 85.000 ;
        RECT 46.530 84.200 50.480 84.400 ;
        RECT 50.130 83.600 50.480 84.200 ;
        RECT 46.530 83.400 50.480 83.600 ;
        RECT 50.130 82.800 50.480 83.400 ;
        RECT 46.530 82.600 50.480 82.800 ;
        RECT 50.130 82.000 50.480 82.600 ;
        RECT 51.080 82.000 51.280 89.600 ;
        RECT 51.880 82.000 52.080 89.600 ;
        RECT 52.680 82.000 52.880 89.600 ;
        RECT 53.480 82.000 53.680 89.600 ;
        RECT 54.280 82.000 55.180 98.000 ;
        RECT 55.780 90.400 55.980 98.000 ;
        RECT 56.580 90.400 56.780 98.000 ;
        RECT 57.380 90.400 57.580 98.000 ;
        RECT 58.180 90.400 58.380 98.000 ;
        RECT 58.980 97.400 59.330 98.000 ;
        RECT 58.980 97.200 62.930 97.400 ;
        RECT 58.980 96.600 59.330 97.200 ;
        RECT 58.980 96.400 62.930 96.600 ;
        RECT 58.980 95.800 59.330 96.400 ;
        RECT 58.980 95.600 62.930 95.800 ;
        RECT 58.980 95.000 59.330 95.600 ;
        RECT 63.930 95.550 64.330 99.200 ;
        RECT 65.130 99.200 84.330 99.600 ;
        RECT 65.130 95.550 65.530 99.200 ;
        RECT 69.180 99.150 71.480 99.200 ;
        RECT 77.980 99.150 80.280 99.200 ;
        RECT 66.530 98.000 82.930 98.600 ;
        RECT 70.130 97.400 70.480 98.000 ;
        RECT 66.530 97.200 70.480 97.400 ;
        RECT 70.130 96.600 70.480 97.200 ;
        RECT 66.530 96.400 70.480 96.600 ;
        RECT 70.130 95.800 70.480 96.400 ;
        RECT 66.530 95.600 70.480 95.800 ;
        RECT 58.980 94.800 62.930 95.000 ;
        RECT 58.980 94.200 59.330 94.800 ;
        RECT 58.980 94.000 62.930 94.200 ;
        RECT 58.980 93.400 59.330 94.000 ;
        RECT 58.980 93.200 62.930 93.400 ;
        RECT 63.880 93.250 65.580 95.550 ;
        RECT 70.130 95.000 70.480 95.600 ;
        RECT 66.530 94.800 70.480 95.000 ;
        RECT 70.130 94.200 70.480 94.800 ;
        RECT 66.530 94.000 70.480 94.200 ;
        RECT 70.130 93.400 70.480 94.000 ;
        RECT 58.980 92.600 59.330 93.200 ;
        RECT 58.980 92.400 62.930 92.600 ;
        RECT 58.980 91.800 59.330 92.400 ;
        RECT 58.980 91.600 62.930 91.800 ;
        RECT 58.980 91.000 59.330 91.600 ;
        RECT 58.980 90.800 62.930 91.000 ;
        RECT 58.980 90.400 59.330 90.800 ;
        RECT 55.780 82.000 55.980 89.600 ;
        RECT 56.580 82.000 56.780 89.600 ;
        RECT 57.380 82.000 57.580 89.600 ;
        RECT 58.180 82.000 58.380 89.600 ;
        RECT 58.980 89.200 59.330 89.600 ;
        RECT 58.980 89.000 62.930 89.200 ;
        RECT 58.980 88.400 59.330 89.000 ;
        RECT 58.980 88.200 62.930 88.400 ;
        RECT 58.980 87.600 59.330 88.200 ;
        RECT 58.980 87.400 62.930 87.600 ;
        RECT 58.980 86.800 59.330 87.400 ;
        RECT 58.980 86.600 62.930 86.800 ;
        RECT 63.930 86.750 64.330 93.250 ;
        RECT 65.130 86.750 65.530 93.250 ;
        RECT 66.530 93.200 70.480 93.400 ;
        RECT 70.130 92.600 70.480 93.200 ;
        RECT 66.530 92.400 70.480 92.600 ;
        RECT 70.130 91.800 70.480 92.400 ;
        RECT 66.530 91.600 70.480 91.800 ;
        RECT 70.130 91.000 70.480 91.600 ;
        RECT 66.530 90.800 70.480 91.000 ;
        RECT 70.130 90.400 70.480 90.800 ;
        RECT 71.080 90.400 71.280 98.000 ;
        RECT 71.880 90.400 72.080 98.000 ;
        RECT 72.680 90.400 72.880 98.000 ;
        RECT 73.480 90.400 73.680 98.000 ;
        RECT 70.130 89.200 70.480 89.600 ;
        RECT 66.530 89.000 70.480 89.200 ;
        RECT 70.130 88.400 70.480 89.000 ;
        RECT 66.530 88.200 70.480 88.400 ;
        RECT 70.130 87.600 70.480 88.200 ;
        RECT 66.530 87.400 70.480 87.600 ;
        RECT 70.130 86.800 70.480 87.400 ;
        RECT 58.980 86.000 59.330 86.600 ;
        RECT 58.980 85.800 62.930 86.000 ;
        RECT 58.980 85.200 59.330 85.800 ;
        RECT 58.980 85.000 62.930 85.200 ;
        RECT 58.980 84.400 59.330 85.000 ;
        RECT 63.880 84.450 65.580 86.750 ;
        RECT 66.530 86.600 70.480 86.800 ;
        RECT 70.130 86.000 70.480 86.600 ;
        RECT 66.530 85.800 70.480 86.000 ;
        RECT 70.130 85.200 70.480 85.800 ;
        RECT 66.530 85.000 70.480 85.200 ;
        RECT 58.980 84.200 62.930 84.400 ;
        RECT 58.980 83.600 59.330 84.200 ;
        RECT 58.980 83.400 62.930 83.600 ;
        RECT 58.980 82.800 59.330 83.400 ;
        RECT 58.980 82.600 62.930 82.800 ;
        RECT 58.980 82.000 59.330 82.600 ;
        RECT 46.530 81.400 62.930 82.000 ;
        RECT 49.180 80.800 51.480 80.850 ;
        RECT 57.980 80.800 60.280 80.850 ;
        RECT 63.930 80.800 64.330 84.450 ;
        RECT 45.130 80.400 64.330 80.800 ;
        RECT 65.130 80.800 65.530 84.450 ;
        RECT 70.130 84.400 70.480 85.000 ;
        RECT 66.530 84.200 70.480 84.400 ;
        RECT 70.130 83.600 70.480 84.200 ;
        RECT 66.530 83.400 70.480 83.600 ;
        RECT 70.130 82.800 70.480 83.400 ;
        RECT 66.530 82.600 70.480 82.800 ;
        RECT 70.130 82.000 70.480 82.600 ;
        RECT 71.080 82.000 71.280 89.600 ;
        RECT 71.880 82.000 72.080 89.600 ;
        RECT 72.680 82.000 72.880 89.600 ;
        RECT 73.480 82.000 73.680 89.600 ;
        RECT 74.280 82.000 75.180 98.000 ;
        RECT 75.780 90.400 75.980 98.000 ;
        RECT 76.580 90.400 76.780 98.000 ;
        RECT 77.380 90.400 77.580 98.000 ;
        RECT 78.180 90.400 78.380 98.000 ;
        RECT 78.980 97.400 79.330 98.000 ;
        RECT 78.980 97.200 82.930 97.400 ;
        RECT 78.980 96.600 79.330 97.200 ;
        RECT 78.980 96.400 82.930 96.600 ;
        RECT 78.980 95.800 79.330 96.400 ;
        RECT 78.980 95.600 82.930 95.800 ;
        RECT 78.980 95.000 79.330 95.600 ;
        RECT 83.930 95.550 84.330 99.200 ;
        RECT 85.130 99.200 104.330 99.600 ;
        RECT 85.130 95.550 85.530 99.200 ;
        RECT 89.180 99.150 91.480 99.200 ;
        RECT 97.980 99.150 100.280 99.200 ;
        RECT 86.530 98.000 102.930 98.600 ;
        RECT 90.130 97.400 90.480 98.000 ;
        RECT 86.530 97.200 90.480 97.400 ;
        RECT 90.130 96.600 90.480 97.200 ;
        RECT 86.530 96.400 90.480 96.600 ;
        RECT 90.130 95.800 90.480 96.400 ;
        RECT 86.530 95.600 90.480 95.800 ;
        RECT 78.980 94.800 82.930 95.000 ;
        RECT 78.980 94.200 79.330 94.800 ;
        RECT 78.980 94.000 82.930 94.200 ;
        RECT 78.980 93.400 79.330 94.000 ;
        RECT 78.980 93.200 82.930 93.400 ;
        RECT 83.880 93.250 85.580 95.550 ;
        RECT 90.130 95.000 90.480 95.600 ;
        RECT 86.530 94.800 90.480 95.000 ;
        RECT 90.130 94.200 90.480 94.800 ;
        RECT 86.530 94.000 90.480 94.200 ;
        RECT 90.130 93.400 90.480 94.000 ;
        RECT 78.980 92.600 79.330 93.200 ;
        RECT 78.980 92.400 82.930 92.600 ;
        RECT 78.980 91.800 79.330 92.400 ;
        RECT 78.980 91.600 82.930 91.800 ;
        RECT 78.980 91.000 79.330 91.600 ;
        RECT 78.980 90.800 82.930 91.000 ;
        RECT 78.980 90.400 79.330 90.800 ;
        RECT 75.780 82.000 75.980 89.600 ;
        RECT 76.580 82.000 76.780 89.600 ;
        RECT 77.380 82.000 77.580 89.600 ;
        RECT 78.180 82.000 78.380 89.600 ;
        RECT 78.980 89.200 79.330 89.600 ;
        RECT 78.980 89.000 82.930 89.200 ;
        RECT 78.980 88.400 79.330 89.000 ;
        RECT 78.980 88.200 82.930 88.400 ;
        RECT 78.980 87.600 79.330 88.200 ;
        RECT 78.980 87.400 82.930 87.600 ;
        RECT 78.980 86.800 79.330 87.400 ;
        RECT 78.980 86.600 82.930 86.800 ;
        RECT 83.930 86.750 84.330 93.250 ;
        RECT 85.130 86.750 85.530 93.250 ;
        RECT 86.530 93.200 90.480 93.400 ;
        RECT 90.130 92.600 90.480 93.200 ;
        RECT 86.530 92.400 90.480 92.600 ;
        RECT 90.130 91.800 90.480 92.400 ;
        RECT 86.530 91.600 90.480 91.800 ;
        RECT 90.130 91.000 90.480 91.600 ;
        RECT 86.530 90.800 90.480 91.000 ;
        RECT 90.130 90.400 90.480 90.800 ;
        RECT 91.080 90.400 91.280 98.000 ;
        RECT 91.880 90.400 92.080 98.000 ;
        RECT 92.680 90.400 92.880 98.000 ;
        RECT 93.480 90.400 93.680 98.000 ;
        RECT 90.130 89.200 90.480 89.600 ;
        RECT 86.530 89.000 90.480 89.200 ;
        RECT 90.130 88.400 90.480 89.000 ;
        RECT 86.530 88.200 90.480 88.400 ;
        RECT 90.130 87.600 90.480 88.200 ;
        RECT 86.530 87.400 90.480 87.600 ;
        RECT 90.130 86.800 90.480 87.400 ;
        RECT 78.980 86.000 79.330 86.600 ;
        RECT 78.980 85.800 82.930 86.000 ;
        RECT 78.980 85.200 79.330 85.800 ;
        RECT 78.980 85.000 82.930 85.200 ;
        RECT 78.980 84.400 79.330 85.000 ;
        RECT 83.880 84.450 85.580 86.750 ;
        RECT 86.530 86.600 90.480 86.800 ;
        RECT 90.130 86.000 90.480 86.600 ;
        RECT 86.530 85.800 90.480 86.000 ;
        RECT 90.130 85.200 90.480 85.800 ;
        RECT 86.530 85.000 90.480 85.200 ;
        RECT 78.980 84.200 82.930 84.400 ;
        RECT 78.980 83.600 79.330 84.200 ;
        RECT 78.980 83.400 82.930 83.600 ;
        RECT 78.980 82.800 79.330 83.400 ;
        RECT 78.980 82.600 82.930 82.800 ;
        RECT 78.980 82.000 79.330 82.600 ;
        RECT 66.530 81.400 82.930 82.000 ;
        RECT 69.180 80.800 71.480 80.850 ;
        RECT 77.980 80.800 80.280 80.850 ;
        RECT 83.930 80.800 84.330 84.450 ;
        RECT 65.130 80.400 84.330 80.800 ;
        RECT 85.130 80.800 85.530 84.450 ;
        RECT 90.130 84.400 90.480 85.000 ;
        RECT 86.530 84.200 90.480 84.400 ;
        RECT 90.130 83.600 90.480 84.200 ;
        RECT 86.530 83.400 90.480 83.600 ;
        RECT 90.130 82.800 90.480 83.400 ;
        RECT 86.530 82.600 90.480 82.800 ;
        RECT 90.130 82.000 90.480 82.600 ;
        RECT 91.080 82.000 91.280 89.600 ;
        RECT 91.880 82.000 92.080 89.600 ;
        RECT 92.680 82.000 92.880 89.600 ;
        RECT 93.480 82.000 93.680 89.600 ;
        RECT 94.280 82.000 95.180 98.000 ;
        RECT 95.780 90.400 95.980 98.000 ;
        RECT 96.580 90.400 96.780 98.000 ;
        RECT 97.380 90.400 97.580 98.000 ;
        RECT 98.180 90.400 98.380 98.000 ;
        RECT 98.980 97.400 99.330 98.000 ;
        RECT 98.980 97.200 102.930 97.400 ;
        RECT 98.980 96.600 99.330 97.200 ;
        RECT 98.980 96.400 102.930 96.600 ;
        RECT 98.980 95.800 99.330 96.400 ;
        RECT 98.980 95.600 102.930 95.800 ;
        RECT 98.980 95.000 99.330 95.600 ;
        RECT 103.930 95.550 104.330 99.200 ;
        RECT 105.130 99.200 124.330 99.600 ;
        RECT 105.130 95.550 105.530 99.200 ;
        RECT 109.180 99.150 111.480 99.200 ;
        RECT 117.980 99.150 120.280 99.200 ;
        RECT 106.530 98.000 122.930 98.600 ;
        RECT 110.130 97.400 110.480 98.000 ;
        RECT 106.530 97.200 110.480 97.400 ;
        RECT 110.130 96.600 110.480 97.200 ;
        RECT 106.530 96.400 110.480 96.600 ;
        RECT 110.130 95.800 110.480 96.400 ;
        RECT 106.530 95.600 110.480 95.800 ;
        RECT 98.980 94.800 102.930 95.000 ;
        RECT 98.980 94.200 99.330 94.800 ;
        RECT 98.980 94.000 102.930 94.200 ;
        RECT 98.980 93.400 99.330 94.000 ;
        RECT 98.980 93.200 102.930 93.400 ;
        RECT 103.880 93.250 105.580 95.550 ;
        RECT 110.130 95.000 110.480 95.600 ;
        RECT 106.530 94.800 110.480 95.000 ;
        RECT 110.130 94.200 110.480 94.800 ;
        RECT 106.530 94.000 110.480 94.200 ;
        RECT 110.130 93.400 110.480 94.000 ;
        RECT 98.980 92.600 99.330 93.200 ;
        RECT 98.980 92.400 102.930 92.600 ;
        RECT 98.980 91.800 99.330 92.400 ;
        RECT 98.980 91.600 102.930 91.800 ;
        RECT 98.980 91.000 99.330 91.600 ;
        RECT 98.980 90.800 102.930 91.000 ;
        RECT 98.980 90.400 99.330 90.800 ;
        RECT 95.780 82.000 95.980 89.600 ;
        RECT 96.580 82.000 96.780 89.600 ;
        RECT 97.380 82.000 97.580 89.600 ;
        RECT 98.180 82.000 98.380 89.600 ;
        RECT 98.980 89.200 99.330 89.600 ;
        RECT 98.980 89.000 102.930 89.200 ;
        RECT 98.980 88.400 99.330 89.000 ;
        RECT 98.980 88.200 102.930 88.400 ;
        RECT 98.980 87.600 99.330 88.200 ;
        RECT 98.980 87.400 102.930 87.600 ;
        RECT 98.980 86.800 99.330 87.400 ;
        RECT 98.980 86.600 102.930 86.800 ;
        RECT 103.930 86.750 104.330 93.250 ;
        RECT 105.130 86.750 105.530 93.250 ;
        RECT 106.530 93.200 110.480 93.400 ;
        RECT 110.130 92.600 110.480 93.200 ;
        RECT 106.530 92.400 110.480 92.600 ;
        RECT 110.130 91.800 110.480 92.400 ;
        RECT 106.530 91.600 110.480 91.800 ;
        RECT 110.130 91.000 110.480 91.600 ;
        RECT 106.530 90.800 110.480 91.000 ;
        RECT 110.130 90.400 110.480 90.800 ;
        RECT 111.080 90.400 111.280 98.000 ;
        RECT 111.880 90.400 112.080 98.000 ;
        RECT 112.680 90.400 112.880 98.000 ;
        RECT 113.480 90.400 113.680 98.000 ;
        RECT 110.130 89.200 110.480 89.600 ;
        RECT 106.530 89.000 110.480 89.200 ;
        RECT 110.130 88.400 110.480 89.000 ;
        RECT 106.530 88.200 110.480 88.400 ;
        RECT 110.130 87.600 110.480 88.200 ;
        RECT 106.530 87.400 110.480 87.600 ;
        RECT 110.130 86.800 110.480 87.400 ;
        RECT 98.980 86.000 99.330 86.600 ;
        RECT 98.980 85.800 102.930 86.000 ;
        RECT 98.980 85.200 99.330 85.800 ;
        RECT 98.980 85.000 102.930 85.200 ;
        RECT 98.980 84.400 99.330 85.000 ;
        RECT 103.880 84.450 105.580 86.750 ;
        RECT 106.530 86.600 110.480 86.800 ;
        RECT 110.130 86.000 110.480 86.600 ;
        RECT 106.530 85.800 110.480 86.000 ;
        RECT 110.130 85.200 110.480 85.800 ;
        RECT 106.530 85.000 110.480 85.200 ;
        RECT 98.980 84.200 102.930 84.400 ;
        RECT 98.980 83.600 99.330 84.200 ;
        RECT 98.980 83.400 102.930 83.600 ;
        RECT 98.980 82.800 99.330 83.400 ;
        RECT 98.980 82.600 102.930 82.800 ;
        RECT 98.980 82.000 99.330 82.600 ;
        RECT 86.530 81.400 102.930 82.000 ;
        RECT 89.180 80.800 91.480 80.850 ;
        RECT 97.980 80.800 100.280 80.850 ;
        RECT 103.930 80.800 104.330 84.450 ;
        RECT 85.130 80.400 104.330 80.800 ;
        RECT 105.130 80.800 105.530 84.450 ;
        RECT 110.130 84.400 110.480 85.000 ;
        RECT 106.530 84.200 110.480 84.400 ;
        RECT 110.130 83.600 110.480 84.200 ;
        RECT 106.530 83.400 110.480 83.600 ;
        RECT 110.130 82.800 110.480 83.400 ;
        RECT 106.530 82.600 110.480 82.800 ;
        RECT 110.130 82.000 110.480 82.600 ;
        RECT 111.080 82.000 111.280 89.600 ;
        RECT 111.880 82.000 112.080 89.600 ;
        RECT 112.680 82.000 112.880 89.600 ;
        RECT 113.480 82.000 113.680 89.600 ;
        RECT 114.280 82.000 115.180 98.000 ;
        RECT 115.780 90.400 115.980 98.000 ;
        RECT 116.580 90.400 116.780 98.000 ;
        RECT 117.380 90.400 117.580 98.000 ;
        RECT 118.180 90.400 118.380 98.000 ;
        RECT 118.980 97.400 119.330 98.000 ;
        RECT 118.980 97.200 122.930 97.400 ;
        RECT 118.980 96.600 119.330 97.200 ;
        RECT 118.980 96.400 122.930 96.600 ;
        RECT 118.980 95.800 119.330 96.400 ;
        RECT 118.980 95.600 122.930 95.800 ;
        RECT 118.980 95.000 119.330 95.600 ;
        RECT 123.930 95.550 124.330 99.200 ;
        RECT 125.340 96.740 125.700 97.120 ;
        RECT 125.970 96.740 126.330 97.120 ;
        RECT 126.570 96.740 126.930 97.120 ;
        RECT 125.340 96.150 125.700 96.530 ;
        RECT 125.970 96.150 126.330 96.530 ;
        RECT 126.570 96.150 126.930 96.530 ;
        RECT 118.980 94.800 122.930 95.000 ;
        RECT 118.980 94.200 119.330 94.800 ;
        RECT 118.980 94.000 122.930 94.200 ;
        RECT 118.980 93.400 119.330 94.000 ;
        RECT 118.980 93.200 122.930 93.400 ;
        RECT 123.880 93.250 124.730 95.550 ;
        RECT 118.980 92.600 119.330 93.200 ;
        RECT 118.980 92.400 122.930 92.600 ;
        RECT 118.980 91.800 119.330 92.400 ;
        RECT 118.980 91.600 122.930 91.800 ;
        RECT 118.980 91.000 119.330 91.600 ;
        RECT 118.980 90.800 122.930 91.000 ;
        RECT 118.980 90.400 119.330 90.800 ;
        RECT 115.780 82.000 115.980 89.600 ;
        RECT 116.580 82.000 116.780 89.600 ;
        RECT 117.380 82.000 117.580 89.600 ;
        RECT 118.180 82.000 118.380 89.600 ;
        RECT 118.980 89.200 119.330 89.600 ;
        RECT 118.980 89.000 122.930 89.200 ;
        RECT 118.980 88.400 119.330 89.000 ;
        RECT 118.980 88.200 122.930 88.400 ;
        RECT 118.980 87.600 119.330 88.200 ;
        RECT 118.980 87.400 122.930 87.600 ;
        RECT 118.980 86.800 119.330 87.400 ;
        RECT 118.980 86.600 122.930 86.800 ;
        RECT 123.930 86.750 124.330 93.250 ;
        RECT 118.980 86.000 119.330 86.600 ;
        RECT 118.980 85.800 122.930 86.000 ;
        RECT 118.980 85.200 119.330 85.800 ;
        RECT 118.980 85.000 122.930 85.200 ;
        RECT 118.980 84.400 119.330 85.000 ;
        RECT 123.880 84.450 124.730 86.750 ;
        RECT 118.980 84.200 122.930 84.400 ;
        RECT 118.980 83.600 119.330 84.200 ;
        RECT 118.980 83.400 122.930 83.600 ;
        RECT 118.980 82.800 119.330 83.400 ;
        RECT 118.980 82.600 122.930 82.800 ;
        RECT 118.980 82.000 119.330 82.600 ;
        RECT 106.530 81.400 122.930 82.000 ;
        RECT 109.180 80.800 111.480 80.850 ;
        RECT 117.980 80.800 120.280 80.850 ;
        RECT 123.930 80.800 124.330 84.450 ;
        RECT 125.340 82.535 125.700 82.915 ;
        RECT 125.970 82.535 126.330 82.915 ;
        RECT 126.570 82.535 126.930 82.915 ;
        RECT 125.340 81.945 125.700 82.325 ;
        RECT 125.970 81.945 126.330 82.325 ;
        RECT 126.570 81.945 126.930 82.325 ;
        RECT 105.130 80.400 124.330 80.800 ;
        RECT 9.180 79.600 11.480 80.400 ;
        RECT 17.980 79.600 20.280 80.400 ;
        RECT 29.180 79.600 31.480 80.400 ;
        RECT 37.980 79.600 40.280 80.400 ;
        RECT 49.180 79.600 51.480 80.400 ;
        RECT 57.980 79.600 60.280 80.400 ;
        RECT 69.180 79.600 71.480 80.400 ;
        RECT 77.980 79.600 80.280 80.400 ;
        RECT 89.180 79.600 91.480 80.400 ;
        RECT 97.980 79.600 100.280 80.400 ;
        RECT 109.180 79.600 111.480 80.400 ;
        RECT 117.980 79.600 120.280 80.400 ;
        RECT 5.130 79.200 24.330 79.600 ;
        RECT 2.515 77.460 2.875 77.840 ;
        RECT 3.145 77.460 3.505 77.840 ;
        RECT 3.745 77.460 4.105 77.840 ;
        RECT 2.515 76.870 2.875 77.250 ;
        RECT 3.145 76.870 3.505 77.250 ;
        RECT 3.745 76.870 4.105 77.250 ;
        RECT 5.130 75.550 5.530 79.200 ;
        RECT 9.180 79.150 11.480 79.200 ;
        RECT 17.980 79.150 20.280 79.200 ;
        RECT 6.530 78.000 22.930 78.600 ;
        RECT 10.130 77.400 10.480 78.000 ;
        RECT 6.530 77.200 10.480 77.400 ;
        RECT 10.130 76.600 10.480 77.200 ;
        RECT 6.530 76.400 10.480 76.600 ;
        RECT 10.130 75.800 10.480 76.400 ;
        RECT 6.530 75.600 10.480 75.800 ;
        RECT 4.730 75.545 5.580 75.550 ;
        RECT 2.315 73.250 5.580 75.545 ;
        RECT 10.130 75.000 10.480 75.600 ;
        RECT 6.530 74.800 10.480 75.000 ;
        RECT 10.130 74.200 10.480 74.800 ;
        RECT 6.530 74.000 10.480 74.200 ;
        RECT 10.130 73.400 10.480 74.000 ;
        RECT 5.130 66.750 5.530 73.250 ;
        RECT 6.530 73.200 10.480 73.400 ;
        RECT 10.130 72.600 10.480 73.200 ;
        RECT 6.530 72.400 10.480 72.600 ;
        RECT 10.130 71.800 10.480 72.400 ;
        RECT 6.530 71.600 10.480 71.800 ;
        RECT 10.130 71.000 10.480 71.600 ;
        RECT 6.530 70.800 10.480 71.000 ;
        RECT 10.130 70.400 10.480 70.800 ;
        RECT 11.080 70.400 11.280 78.000 ;
        RECT 11.880 70.400 12.080 78.000 ;
        RECT 12.680 70.400 12.880 78.000 ;
        RECT 13.480 70.400 13.680 78.000 ;
        RECT 10.130 69.200 10.480 69.600 ;
        RECT 6.530 69.000 10.480 69.200 ;
        RECT 10.130 68.400 10.480 69.000 ;
        RECT 6.530 68.200 10.480 68.400 ;
        RECT 10.130 67.600 10.480 68.200 ;
        RECT 6.530 67.400 10.480 67.600 ;
        RECT 10.130 66.800 10.480 67.400 ;
        RECT 4.730 66.745 5.580 66.750 ;
        RECT 2.315 64.450 5.580 66.745 ;
        RECT 6.530 66.600 10.480 66.800 ;
        RECT 10.130 66.000 10.480 66.600 ;
        RECT 6.530 65.800 10.480 66.000 ;
        RECT 10.130 65.200 10.480 65.800 ;
        RECT 6.530 65.000 10.480 65.200 ;
        RECT 2.515 63.130 2.875 63.510 ;
        RECT 3.145 63.130 3.505 63.510 ;
        RECT 3.745 63.130 4.105 63.510 ;
        RECT 2.515 62.540 2.875 62.920 ;
        RECT 3.145 62.540 3.505 62.920 ;
        RECT 3.745 62.540 4.105 62.920 ;
        RECT 5.130 60.800 5.530 64.450 ;
        RECT 10.130 64.400 10.480 65.000 ;
        RECT 6.530 64.200 10.480 64.400 ;
        RECT 10.130 63.600 10.480 64.200 ;
        RECT 6.530 63.400 10.480 63.600 ;
        RECT 10.130 62.800 10.480 63.400 ;
        RECT 6.530 62.600 10.480 62.800 ;
        RECT 10.130 62.000 10.480 62.600 ;
        RECT 11.080 62.000 11.280 69.600 ;
        RECT 11.880 62.000 12.080 69.600 ;
        RECT 12.680 62.000 12.880 69.600 ;
        RECT 13.480 62.000 13.680 69.600 ;
        RECT 14.280 62.000 15.180 78.000 ;
        RECT 15.780 70.400 15.980 78.000 ;
        RECT 16.580 70.400 16.780 78.000 ;
        RECT 17.380 70.400 17.580 78.000 ;
        RECT 18.180 70.400 18.380 78.000 ;
        RECT 18.980 77.400 19.330 78.000 ;
        RECT 18.980 77.200 22.930 77.400 ;
        RECT 18.980 76.600 19.330 77.200 ;
        RECT 18.980 76.400 22.930 76.600 ;
        RECT 18.980 75.800 19.330 76.400 ;
        RECT 18.980 75.600 22.930 75.800 ;
        RECT 18.980 75.000 19.330 75.600 ;
        RECT 23.930 75.550 24.330 79.200 ;
        RECT 25.130 79.200 44.330 79.600 ;
        RECT 25.130 75.550 25.530 79.200 ;
        RECT 29.180 79.150 31.480 79.200 ;
        RECT 37.980 79.150 40.280 79.200 ;
        RECT 26.530 78.000 42.930 78.600 ;
        RECT 30.130 77.400 30.480 78.000 ;
        RECT 26.530 77.200 30.480 77.400 ;
        RECT 30.130 76.600 30.480 77.200 ;
        RECT 26.530 76.400 30.480 76.600 ;
        RECT 30.130 75.800 30.480 76.400 ;
        RECT 26.530 75.600 30.480 75.800 ;
        RECT 18.980 74.800 22.930 75.000 ;
        RECT 18.980 74.200 19.330 74.800 ;
        RECT 18.980 74.000 22.930 74.200 ;
        RECT 18.980 73.400 19.330 74.000 ;
        RECT 18.980 73.200 22.930 73.400 ;
        RECT 23.880 73.250 25.580 75.550 ;
        RECT 30.130 75.000 30.480 75.600 ;
        RECT 26.530 74.800 30.480 75.000 ;
        RECT 30.130 74.200 30.480 74.800 ;
        RECT 26.530 74.000 30.480 74.200 ;
        RECT 30.130 73.400 30.480 74.000 ;
        RECT 18.980 72.600 19.330 73.200 ;
        RECT 18.980 72.400 22.930 72.600 ;
        RECT 18.980 71.800 19.330 72.400 ;
        RECT 18.980 71.600 22.930 71.800 ;
        RECT 18.980 71.000 19.330 71.600 ;
        RECT 18.980 70.800 22.930 71.000 ;
        RECT 18.980 70.400 19.330 70.800 ;
        RECT 15.780 62.000 15.980 69.600 ;
        RECT 16.580 62.000 16.780 69.600 ;
        RECT 17.380 62.000 17.580 69.600 ;
        RECT 18.180 62.000 18.380 69.600 ;
        RECT 18.980 69.200 19.330 69.600 ;
        RECT 18.980 69.000 22.930 69.200 ;
        RECT 18.980 68.400 19.330 69.000 ;
        RECT 18.980 68.200 22.930 68.400 ;
        RECT 18.980 67.600 19.330 68.200 ;
        RECT 18.980 67.400 22.930 67.600 ;
        RECT 18.980 66.800 19.330 67.400 ;
        RECT 18.980 66.600 22.930 66.800 ;
        RECT 23.930 66.750 24.330 73.250 ;
        RECT 25.130 66.750 25.530 73.250 ;
        RECT 26.530 73.200 30.480 73.400 ;
        RECT 30.130 72.600 30.480 73.200 ;
        RECT 26.530 72.400 30.480 72.600 ;
        RECT 30.130 71.800 30.480 72.400 ;
        RECT 26.530 71.600 30.480 71.800 ;
        RECT 30.130 71.000 30.480 71.600 ;
        RECT 26.530 70.800 30.480 71.000 ;
        RECT 30.130 70.400 30.480 70.800 ;
        RECT 31.080 70.400 31.280 78.000 ;
        RECT 31.880 70.400 32.080 78.000 ;
        RECT 32.680 70.400 32.880 78.000 ;
        RECT 33.480 70.400 33.680 78.000 ;
        RECT 30.130 69.200 30.480 69.600 ;
        RECT 26.530 69.000 30.480 69.200 ;
        RECT 30.130 68.400 30.480 69.000 ;
        RECT 26.530 68.200 30.480 68.400 ;
        RECT 30.130 67.600 30.480 68.200 ;
        RECT 26.530 67.400 30.480 67.600 ;
        RECT 30.130 66.800 30.480 67.400 ;
        RECT 18.980 66.000 19.330 66.600 ;
        RECT 18.980 65.800 22.930 66.000 ;
        RECT 18.980 65.200 19.330 65.800 ;
        RECT 18.980 65.000 22.930 65.200 ;
        RECT 18.980 64.400 19.330 65.000 ;
        RECT 23.880 64.450 25.580 66.750 ;
        RECT 26.530 66.600 30.480 66.800 ;
        RECT 30.130 66.000 30.480 66.600 ;
        RECT 26.530 65.800 30.480 66.000 ;
        RECT 30.130 65.200 30.480 65.800 ;
        RECT 26.530 65.000 30.480 65.200 ;
        RECT 18.980 64.200 22.930 64.400 ;
        RECT 18.980 63.600 19.330 64.200 ;
        RECT 18.980 63.400 22.930 63.600 ;
        RECT 18.980 62.800 19.330 63.400 ;
        RECT 18.980 62.600 22.930 62.800 ;
        RECT 18.980 62.000 19.330 62.600 ;
        RECT 6.530 61.400 22.930 62.000 ;
        RECT 9.180 60.800 11.480 60.850 ;
        RECT 17.980 60.800 20.280 60.850 ;
        RECT 23.930 60.800 24.330 64.450 ;
        RECT 5.130 60.400 24.330 60.800 ;
        RECT 25.130 60.800 25.530 64.450 ;
        RECT 30.130 64.400 30.480 65.000 ;
        RECT 26.530 64.200 30.480 64.400 ;
        RECT 30.130 63.600 30.480 64.200 ;
        RECT 26.530 63.400 30.480 63.600 ;
        RECT 30.130 62.800 30.480 63.400 ;
        RECT 26.530 62.600 30.480 62.800 ;
        RECT 30.130 62.000 30.480 62.600 ;
        RECT 31.080 62.000 31.280 69.600 ;
        RECT 31.880 62.000 32.080 69.600 ;
        RECT 32.680 62.000 32.880 69.600 ;
        RECT 33.480 62.000 33.680 69.600 ;
        RECT 34.280 62.000 35.180 78.000 ;
        RECT 35.780 70.400 35.980 78.000 ;
        RECT 36.580 70.400 36.780 78.000 ;
        RECT 37.380 70.400 37.580 78.000 ;
        RECT 38.180 70.400 38.380 78.000 ;
        RECT 38.980 77.400 39.330 78.000 ;
        RECT 38.980 77.200 42.930 77.400 ;
        RECT 38.980 76.600 39.330 77.200 ;
        RECT 38.980 76.400 42.930 76.600 ;
        RECT 38.980 75.800 39.330 76.400 ;
        RECT 38.980 75.600 42.930 75.800 ;
        RECT 38.980 75.000 39.330 75.600 ;
        RECT 43.930 75.550 44.330 79.200 ;
        RECT 45.130 79.200 64.330 79.600 ;
        RECT 45.130 75.550 45.530 79.200 ;
        RECT 49.180 79.150 51.480 79.200 ;
        RECT 57.980 79.150 60.280 79.200 ;
        RECT 46.530 78.000 62.930 78.600 ;
        RECT 50.130 77.400 50.480 78.000 ;
        RECT 46.530 77.200 50.480 77.400 ;
        RECT 50.130 76.600 50.480 77.200 ;
        RECT 46.530 76.400 50.480 76.600 ;
        RECT 50.130 75.800 50.480 76.400 ;
        RECT 46.530 75.600 50.480 75.800 ;
        RECT 38.980 74.800 42.930 75.000 ;
        RECT 38.980 74.200 39.330 74.800 ;
        RECT 38.980 74.000 42.930 74.200 ;
        RECT 38.980 73.400 39.330 74.000 ;
        RECT 38.980 73.200 42.930 73.400 ;
        RECT 43.880 73.250 45.580 75.550 ;
        RECT 50.130 75.000 50.480 75.600 ;
        RECT 46.530 74.800 50.480 75.000 ;
        RECT 50.130 74.200 50.480 74.800 ;
        RECT 46.530 74.000 50.480 74.200 ;
        RECT 50.130 73.400 50.480 74.000 ;
        RECT 38.980 72.600 39.330 73.200 ;
        RECT 38.980 72.400 42.930 72.600 ;
        RECT 38.980 71.800 39.330 72.400 ;
        RECT 38.980 71.600 42.930 71.800 ;
        RECT 38.980 71.000 39.330 71.600 ;
        RECT 38.980 70.800 42.930 71.000 ;
        RECT 38.980 70.400 39.330 70.800 ;
        RECT 35.780 62.000 35.980 69.600 ;
        RECT 36.580 62.000 36.780 69.600 ;
        RECT 37.380 62.000 37.580 69.600 ;
        RECT 38.180 62.000 38.380 69.600 ;
        RECT 38.980 69.200 39.330 69.600 ;
        RECT 38.980 69.000 42.930 69.200 ;
        RECT 38.980 68.400 39.330 69.000 ;
        RECT 38.980 68.200 42.930 68.400 ;
        RECT 38.980 67.600 39.330 68.200 ;
        RECT 38.980 67.400 42.930 67.600 ;
        RECT 38.980 66.800 39.330 67.400 ;
        RECT 38.980 66.600 42.930 66.800 ;
        RECT 43.930 66.750 44.330 73.250 ;
        RECT 45.130 66.750 45.530 73.250 ;
        RECT 46.530 73.200 50.480 73.400 ;
        RECT 50.130 72.600 50.480 73.200 ;
        RECT 46.530 72.400 50.480 72.600 ;
        RECT 50.130 71.800 50.480 72.400 ;
        RECT 46.530 71.600 50.480 71.800 ;
        RECT 50.130 71.000 50.480 71.600 ;
        RECT 46.530 70.800 50.480 71.000 ;
        RECT 50.130 70.400 50.480 70.800 ;
        RECT 51.080 70.400 51.280 78.000 ;
        RECT 51.880 70.400 52.080 78.000 ;
        RECT 52.680 70.400 52.880 78.000 ;
        RECT 53.480 70.400 53.680 78.000 ;
        RECT 50.130 69.200 50.480 69.600 ;
        RECT 46.530 69.000 50.480 69.200 ;
        RECT 50.130 68.400 50.480 69.000 ;
        RECT 46.530 68.200 50.480 68.400 ;
        RECT 50.130 67.600 50.480 68.200 ;
        RECT 46.530 67.400 50.480 67.600 ;
        RECT 50.130 66.800 50.480 67.400 ;
        RECT 38.980 66.000 39.330 66.600 ;
        RECT 38.980 65.800 42.930 66.000 ;
        RECT 38.980 65.200 39.330 65.800 ;
        RECT 38.980 65.000 42.930 65.200 ;
        RECT 38.980 64.400 39.330 65.000 ;
        RECT 43.880 64.450 45.580 66.750 ;
        RECT 46.530 66.600 50.480 66.800 ;
        RECT 50.130 66.000 50.480 66.600 ;
        RECT 46.530 65.800 50.480 66.000 ;
        RECT 50.130 65.200 50.480 65.800 ;
        RECT 46.530 65.000 50.480 65.200 ;
        RECT 38.980 64.200 42.930 64.400 ;
        RECT 38.980 63.600 39.330 64.200 ;
        RECT 38.980 63.400 42.930 63.600 ;
        RECT 38.980 62.800 39.330 63.400 ;
        RECT 38.980 62.600 42.930 62.800 ;
        RECT 38.980 62.000 39.330 62.600 ;
        RECT 26.530 61.400 42.930 62.000 ;
        RECT 29.180 60.800 31.480 60.850 ;
        RECT 37.980 60.800 40.280 60.850 ;
        RECT 43.930 60.800 44.330 64.450 ;
        RECT 25.130 60.400 44.330 60.800 ;
        RECT 45.130 60.800 45.530 64.450 ;
        RECT 50.130 64.400 50.480 65.000 ;
        RECT 46.530 64.200 50.480 64.400 ;
        RECT 50.130 63.600 50.480 64.200 ;
        RECT 46.530 63.400 50.480 63.600 ;
        RECT 50.130 62.800 50.480 63.400 ;
        RECT 46.530 62.600 50.480 62.800 ;
        RECT 50.130 62.000 50.480 62.600 ;
        RECT 51.080 62.000 51.280 69.600 ;
        RECT 51.880 62.000 52.080 69.600 ;
        RECT 52.680 62.000 52.880 69.600 ;
        RECT 53.480 62.000 53.680 69.600 ;
        RECT 54.280 62.000 55.180 78.000 ;
        RECT 55.780 70.400 55.980 78.000 ;
        RECT 56.580 70.400 56.780 78.000 ;
        RECT 57.380 70.400 57.580 78.000 ;
        RECT 58.180 70.400 58.380 78.000 ;
        RECT 58.980 77.400 59.330 78.000 ;
        RECT 58.980 77.200 62.930 77.400 ;
        RECT 58.980 76.600 59.330 77.200 ;
        RECT 58.980 76.400 62.930 76.600 ;
        RECT 58.980 75.800 59.330 76.400 ;
        RECT 58.980 75.600 62.930 75.800 ;
        RECT 58.980 75.000 59.330 75.600 ;
        RECT 63.930 75.550 64.330 79.200 ;
        RECT 65.130 79.200 84.330 79.600 ;
        RECT 65.130 75.550 65.530 79.200 ;
        RECT 69.180 79.150 71.480 79.200 ;
        RECT 77.980 79.150 80.280 79.200 ;
        RECT 66.530 78.000 82.930 78.600 ;
        RECT 70.130 77.400 70.480 78.000 ;
        RECT 66.530 77.200 70.480 77.400 ;
        RECT 70.130 76.600 70.480 77.200 ;
        RECT 66.530 76.400 70.480 76.600 ;
        RECT 70.130 75.800 70.480 76.400 ;
        RECT 66.530 75.600 70.480 75.800 ;
        RECT 58.980 74.800 62.930 75.000 ;
        RECT 58.980 74.200 59.330 74.800 ;
        RECT 58.980 74.000 62.930 74.200 ;
        RECT 58.980 73.400 59.330 74.000 ;
        RECT 58.980 73.200 62.930 73.400 ;
        RECT 63.880 73.250 65.580 75.550 ;
        RECT 70.130 75.000 70.480 75.600 ;
        RECT 66.530 74.800 70.480 75.000 ;
        RECT 70.130 74.200 70.480 74.800 ;
        RECT 66.530 74.000 70.480 74.200 ;
        RECT 70.130 73.400 70.480 74.000 ;
        RECT 58.980 72.600 59.330 73.200 ;
        RECT 58.980 72.400 62.930 72.600 ;
        RECT 58.980 71.800 59.330 72.400 ;
        RECT 58.980 71.600 62.930 71.800 ;
        RECT 58.980 71.000 59.330 71.600 ;
        RECT 58.980 70.800 62.930 71.000 ;
        RECT 58.980 70.400 59.330 70.800 ;
        RECT 55.780 62.000 55.980 69.600 ;
        RECT 56.580 62.000 56.780 69.600 ;
        RECT 57.380 62.000 57.580 69.600 ;
        RECT 58.180 62.000 58.380 69.600 ;
        RECT 58.980 69.200 59.330 69.600 ;
        RECT 58.980 69.000 62.930 69.200 ;
        RECT 58.980 68.400 59.330 69.000 ;
        RECT 58.980 68.200 62.930 68.400 ;
        RECT 58.980 67.600 59.330 68.200 ;
        RECT 58.980 67.400 62.930 67.600 ;
        RECT 58.980 66.800 59.330 67.400 ;
        RECT 58.980 66.600 62.930 66.800 ;
        RECT 63.930 66.750 64.330 73.250 ;
        RECT 65.130 66.750 65.530 73.250 ;
        RECT 66.530 73.200 70.480 73.400 ;
        RECT 70.130 72.600 70.480 73.200 ;
        RECT 66.530 72.400 70.480 72.600 ;
        RECT 70.130 71.800 70.480 72.400 ;
        RECT 66.530 71.600 70.480 71.800 ;
        RECT 70.130 71.000 70.480 71.600 ;
        RECT 66.530 70.800 70.480 71.000 ;
        RECT 70.130 70.400 70.480 70.800 ;
        RECT 71.080 70.400 71.280 78.000 ;
        RECT 71.880 70.400 72.080 78.000 ;
        RECT 72.680 70.400 72.880 78.000 ;
        RECT 73.480 70.400 73.680 78.000 ;
        RECT 70.130 69.200 70.480 69.600 ;
        RECT 66.530 69.000 70.480 69.200 ;
        RECT 70.130 68.400 70.480 69.000 ;
        RECT 66.530 68.200 70.480 68.400 ;
        RECT 70.130 67.600 70.480 68.200 ;
        RECT 66.530 67.400 70.480 67.600 ;
        RECT 70.130 66.800 70.480 67.400 ;
        RECT 58.980 66.000 59.330 66.600 ;
        RECT 58.980 65.800 62.930 66.000 ;
        RECT 58.980 65.200 59.330 65.800 ;
        RECT 58.980 65.000 62.930 65.200 ;
        RECT 58.980 64.400 59.330 65.000 ;
        RECT 63.880 64.450 65.580 66.750 ;
        RECT 66.530 66.600 70.480 66.800 ;
        RECT 70.130 66.000 70.480 66.600 ;
        RECT 66.530 65.800 70.480 66.000 ;
        RECT 70.130 65.200 70.480 65.800 ;
        RECT 66.530 65.000 70.480 65.200 ;
        RECT 58.980 64.200 62.930 64.400 ;
        RECT 58.980 63.600 59.330 64.200 ;
        RECT 58.980 63.400 62.930 63.600 ;
        RECT 58.980 62.800 59.330 63.400 ;
        RECT 58.980 62.600 62.930 62.800 ;
        RECT 58.980 62.000 59.330 62.600 ;
        RECT 46.530 61.400 62.930 62.000 ;
        RECT 49.180 60.800 51.480 60.850 ;
        RECT 57.980 60.800 60.280 60.850 ;
        RECT 63.930 60.800 64.330 64.450 ;
        RECT 45.130 60.400 64.330 60.800 ;
        RECT 65.130 60.800 65.530 64.450 ;
        RECT 70.130 64.400 70.480 65.000 ;
        RECT 66.530 64.200 70.480 64.400 ;
        RECT 70.130 63.600 70.480 64.200 ;
        RECT 66.530 63.400 70.480 63.600 ;
        RECT 70.130 62.800 70.480 63.400 ;
        RECT 66.530 62.600 70.480 62.800 ;
        RECT 70.130 62.000 70.480 62.600 ;
        RECT 71.080 62.000 71.280 69.600 ;
        RECT 71.880 62.000 72.080 69.600 ;
        RECT 72.680 62.000 72.880 69.600 ;
        RECT 73.480 62.000 73.680 69.600 ;
        RECT 74.280 62.000 75.180 78.000 ;
        RECT 75.780 70.400 75.980 78.000 ;
        RECT 76.580 70.400 76.780 78.000 ;
        RECT 77.380 70.400 77.580 78.000 ;
        RECT 78.180 70.400 78.380 78.000 ;
        RECT 78.980 77.400 79.330 78.000 ;
        RECT 78.980 77.200 82.930 77.400 ;
        RECT 78.980 76.600 79.330 77.200 ;
        RECT 78.980 76.400 82.930 76.600 ;
        RECT 78.980 75.800 79.330 76.400 ;
        RECT 78.980 75.600 82.930 75.800 ;
        RECT 78.980 75.000 79.330 75.600 ;
        RECT 83.930 75.550 84.330 79.200 ;
        RECT 85.130 79.200 104.330 79.600 ;
        RECT 85.130 75.550 85.530 79.200 ;
        RECT 89.180 79.150 91.480 79.200 ;
        RECT 97.980 79.150 100.280 79.200 ;
        RECT 86.530 78.000 102.930 78.600 ;
        RECT 90.130 77.400 90.480 78.000 ;
        RECT 86.530 77.200 90.480 77.400 ;
        RECT 90.130 76.600 90.480 77.200 ;
        RECT 86.530 76.400 90.480 76.600 ;
        RECT 90.130 75.800 90.480 76.400 ;
        RECT 86.530 75.600 90.480 75.800 ;
        RECT 78.980 74.800 82.930 75.000 ;
        RECT 78.980 74.200 79.330 74.800 ;
        RECT 78.980 74.000 82.930 74.200 ;
        RECT 78.980 73.400 79.330 74.000 ;
        RECT 78.980 73.200 82.930 73.400 ;
        RECT 83.880 73.250 85.580 75.550 ;
        RECT 90.130 75.000 90.480 75.600 ;
        RECT 86.530 74.800 90.480 75.000 ;
        RECT 90.130 74.200 90.480 74.800 ;
        RECT 86.530 74.000 90.480 74.200 ;
        RECT 90.130 73.400 90.480 74.000 ;
        RECT 78.980 72.600 79.330 73.200 ;
        RECT 78.980 72.400 82.930 72.600 ;
        RECT 78.980 71.800 79.330 72.400 ;
        RECT 78.980 71.600 82.930 71.800 ;
        RECT 78.980 71.000 79.330 71.600 ;
        RECT 78.980 70.800 82.930 71.000 ;
        RECT 78.980 70.400 79.330 70.800 ;
        RECT 75.780 62.000 75.980 69.600 ;
        RECT 76.580 62.000 76.780 69.600 ;
        RECT 77.380 62.000 77.580 69.600 ;
        RECT 78.180 62.000 78.380 69.600 ;
        RECT 78.980 69.200 79.330 69.600 ;
        RECT 78.980 69.000 82.930 69.200 ;
        RECT 78.980 68.400 79.330 69.000 ;
        RECT 78.980 68.200 82.930 68.400 ;
        RECT 78.980 67.600 79.330 68.200 ;
        RECT 78.980 67.400 82.930 67.600 ;
        RECT 78.980 66.800 79.330 67.400 ;
        RECT 78.980 66.600 82.930 66.800 ;
        RECT 83.930 66.750 84.330 73.250 ;
        RECT 85.130 66.750 85.530 73.250 ;
        RECT 86.530 73.200 90.480 73.400 ;
        RECT 90.130 72.600 90.480 73.200 ;
        RECT 86.530 72.400 90.480 72.600 ;
        RECT 90.130 71.800 90.480 72.400 ;
        RECT 86.530 71.600 90.480 71.800 ;
        RECT 90.130 71.000 90.480 71.600 ;
        RECT 86.530 70.800 90.480 71.000 ;
        RECT 90.130 70.400 90.480 70.800 ;
        RECT 91.080 70.400 91.280 78.000 ;
        RECT 91.880 70.400 92.080 78.000 ;
        RECT 92.680 70.400 92.880 78.000 ;
        RECT 93.480 70.400 93.680 78.000 ;
        RECT 90.130 69.200 90.480 69.600 ;
        RECT 86.530 69.000 90.480 69.200 ;
        RECT 90.130 68.400 90.480 69.000 ;
        RECT 86.530 68.200 90.480 68.400 ;
        RECT 90.130 67.600 90.480 68.200 ;
        RECT 86.530 67.400 90.480 67.600 ;
        RECT 90.130 66.800 90.480 67.400 ;
        RECT 78.980 66.000 79.330 66.600 ;
        RECT 78.980 65.800 82.930 66.000 ;
        RECT 78.980 65.200 79.330 65.800 ;
        RECT 78.980 65.000 82.930 65.200 ;
        RECT 78.980 64.400 79.330 65.000 ;
        RECT 83.880 64.450 85.580 66.750 ;
        RECT 86.530 66.600 90.480 66.800 ;
        RECT 90.130 66.000 90.480 66.600 ;
        RECT 86.530 65.800 90.480 66.000 ;
        RECT 90.130 65.200 90.480 65.800 ;
        RECT 86.530 65.000 90.480 65.200 ;
        RECT 78.980 64.200 82.930 64.400 ;
        RECT 78.980 63.600 79.330 64.200 ;
        RECT 78.980 63.400 82.930 63.600 ;
        RECT 78.980 62.800 79.330 63.400 ;
        RECT 78.980 62.600 82.930 62.800 ;
        RECT 78.980 62.000 79.330 62.600 ;
        RECT 66.530 61.400 82.930 62.000 ;
        RECT 69.180 60.800 71.480 60.850 ;
        RECT 77.980 60.800 80.280 60.850 ;
        RECT 83.930 60.800 84.330 64.450 ;
        RECT 65.130 60.400 84.330 60.800 ;
        RECT 85.130 60.800 85.530 64.450 ;
        RECT 90.130 64.400 90.480 65.000 ;
        RECT 86.530 64.200 90.480 64.400 ;
        RECT 90.130 63.600 90.480 64.200 ;
        RECT 86.530 63.400 90.480 63.600 ;
        RECT 90.130 62.800 90.480 63.400 ;
        RECT 86.530 62.600 90.480 62.800 ;
        RECT 90.130 62.000 90.480 62.600 ;
        RECT 91.080 62.000 91.280 69.600 ;
        RECT 91.880 62.000 92.080 69.600 ;
        RECT 92.680 62.000 92.880 69.600 ;
        RECT 93.480 62.000 93.680 69.600 ;
        RECT 94.280 62.000 95.180 78.000 ;
        RECT 95.780 70.400 95.980 78.000 ;
        RECT 96.580 70.400 96.780 78.000 ;
        RECT 97.380 70.400 97.580 78.000 ;
        RECT 98.180 70.400 98.380 78.000 ;
        RECT 98.980 77.400 99.330 78.000 ;
        RECT 98.980 77.200 102.930 77.400 ;
        RECT 98.980 76.600 99.330 77.200 ;
        RECT 98.980 76.400 102.930 76.600 ;
        RECT 98.980 75.800 99.330 76.400 ;
        RECT 98.980 75.600 102.930 75.800 ;
        RECT 98.980 75.000 99.330 75.600 ;
        RECT 103.930 75.550 104.330 79.200 ;
        RECT 105.130 79.200 124.330 79.600 ;
        RECT 105.130 75.550 105.530 79.200 ;
        RECT 109.180 79.150 111.480 79.200 ;
        RECT 117.980 79.150 120.280 79.200 ;
        RECT 106.530 78.000 122.930 78.600 ;
        RECT 110.130 77.400 110.480 78.000 ;
        RECT 106.530 77.200 110.480 77.400 ;
        RECT 110.130 76.600 110.480 77.200 ;
        RECT 106.530 76.400 110.480 76.600 ;
        RECT 110.130 75.800 110.480 76.400 ;
        RECT 106.530 75.600 110.480 75.800 ;
        RECT 98.980 74.800 102.930 75.000 ;
        RECT 98.980 74.200 99.330 74.800 ;
        RECT 98.980 74.000 102.930 74.200 ;
        RECT 98.980 73.400 99.330 74.000 ;
        RECT 98.980 73.200 102.930 73.400 ;
        RECT 103.880 73.250 105.580 75.550 ;
        RECT 110.130 75.000 110.480 75.600 ;
        RECT 106.530 74.800 110.480 75.000 ;
        RECT 110.130 74.200 110.480 74.800 ;
        RECT 106.530 74.000 110.480 74.200 ;
        RECT 110.130 73.400 110.480 74.000 ;
        RECT 98.980 72.600 99.330 73.200 ;
        RECT 98.980 72.400 102.930 72.600 ;
        RECT 98.980 71.800 99.330 72.400 ;
        RECT 98.980 71.600 102.930 71.800 ;
        RECT 98.980 71.000 99.330 71.600 ;
        RECT 98.980 70.800 102.930 71.000 ;
        RECT 98.980 70.400 99.330 70.800 ;
        RECT 95.780 62.000 95.980 69.600 ;
        RECT 96.580 62.000 96.780 69.600 ;
        RECT 97.380 62.000 97.580 69.600 ;
        RECT 98.180 62.000 98.380 69.600 ;
        RECT 98.980 69.200 99.330 69.600 ;
        RECT 98.980 69.000 102.930 69.200 ;
        RECT 98.980 68.400 99.330 69.000 ;
        RECT 98.980 68.200 102.930 68.400 ;
        RECT 98.980 67.600 99.330 68.200 ;
        RECT 98.980 67.400 102.930 67.600 ;
        RECT 98.980 66.800 99.330 67.400 ;
        RECT 98.980 66.600 102.930 66.800 ;
        RECT 103.930 66.750 104.330 73.250 ;
        RECT 105.130 66.750 105.530 73.250 ;
        RECT 106.530 73.200 110.480 73.400 ;
        RECT 110.130 72.600 110.480 73.200 ;
        RECT 106.530 72.400 110.480 72.600 ;
        RECT 110.130 71.800 110.480 72.400 ;
        RECT 106.530 71.600 110.480 71.800 ;
        RECT 110.130 71.000 110.480 71.600 ;
        RECT 106.530 70.800 110.480 71.000 ;
        RECT 110.130 70.400 110.480 70.800 ;
        RECT 111.080 70.400 111.280 78.000 ;
        RECT 111.880 70.400 112.080 78.000 ;
        RECT 112.680 70.400 112.880 78.000 ;
        RECT 113.480 70.400 113.680 78.000 ;
        RECT 110.130 69.200 110.480 69.600 ;
        RECT 106.530 69.000 110.480 69.200 ;
        RECT 110.130 68.400 110.480 69.000 ;
        RECT 106.530 68.200 110.480 68.400 ;
        RECT 110.130 67.600 110.480 68.200 ;
        RECT 106.530 67.400 110.480 67.600 ;
        RECT 110.130 66.800 110.480 67.400 ;
        RECT 98.980 66.000 99.330 66.600 ;
        RECT 98.980 65.800 102.930 66.000 ;
        RECT 98.980 65.200 99.330 65.800 ;
        RECT 98.980 65.000 102.930 65.200 ;
        RECT 98.980 64.400 99.330 65.000 ;
        RECT 103.880 64.450 105.580 66.750 ;
        RECT 106.530 66.600 110.480 66.800 ;
        RECT 110.130 66.000 110.480 66.600 ;
        RECT 106.530 65.800 110.480 66.000 ;
        RECT 110.130 65.200 110.480 65.800 ;
        RECT 106.530 65.000 110.480 65.200 ;
        RECT 98.980 64.200 102.930 64.400 ;
        RECT 98.980 63.600 99.330 64.200 ;
        RECT 98.980 63.400 102.930 63.600 ;
        RECT 98.980 62.800 99.330 63.400 ;
        RECT 98.980 62.600 102.930 62.800 ;
        RECT 98.980 62.000 99.330 62.600 ;
        RECT 86.530 61.400 102.930 62.000 ;
        RECT 89.180 60.800 91.480 60.850 ;
        RECT 97.980 60.800 100.280 60.850 ;
        RECT 103.930 60.800 104.330 64.450 ;
        RECT 85.130 60.400 104.330 60.800 ;
        RECT 105.130 60.800 105.530 64.450 ;
        RECT 110.130 64.400 110.480 65.000 ;
        RECT 106.530 64.200 110.480 64.400 ;
        RECT 110.130 63.600 110.480 64.200 ;
        RECT 106.530 63.400 110.480 63.600 ;
        RECT 110.130 62.800 110.480 63.400 ;
        RECT 106.530 62.600 110.480 62.800 ;
        RECT 110.130 62.000 110.480 62.600 ;
        RECT 111.080 62.000 111.280 69.600 ;
        RECT 111.880 62.000 112.080 69.600 ;
        RECT 112.680 62.000 112.880 69.600 ;
        RECT 113.480 62.000 113.680 69.600 ;
        RECT 114.280 62.000 115.180 78.000 ;
        RECT 115.780 70.400 115.980 78.000 ;
        RECT 116.580 70.400 116.780 78.000 ;
        RECT 117.380 70.400 117.580 78.000 ;
        RECT 118.180 70.400 118.380 78.000 ;
        RECT 118.980 77.400 119.330 78.000 ;
        RECT 118.980 77.200 122.930 77.400 ;
        RECT 118.980 76.600 119.330 77.200 ;
        RECT 118.980 76.400 122.930 76.600 ;
        RECT 118.980 75.800 119.330 76.400 ;
        RECT 118.980 75.600 122.930 75.800 ;
        RECT 118.980 75.000 119.330 75.600 ;
        RECT 123.930 75.550 124.330 79.200 ;
        RECT 125.340 76.680 125.700 77.060 ;
        RECT 125.970 76.680 126.330 77.060 ;
        RECT 126.570 76.680 126.930 77.060 ;
        RECT 125.340 76.090 125.700 76.470 ;
        RECT 125.970 76.090 126.330 76.470 ;
        RECT 126.570 76.090 126.930 76.470 ;
        RECT 118.980 74.800 122.930 75.000 ;
        RECT 118.980 74.200 119.330 74.800 ;
        RECT 118.980 74.000 122.930 74.200 ;
        RECT 118.980 73.400 119.330 74.000 ;
        RECT 118.980 73.200 122.930 73.400 ;
        RECT 123.880 73.250 124.730 75.550 ;
        RECT 118.980 72.600 119.330 73.200 ;
        RECT 118.980 72.400 122.930 72.600 ;
        RECT 118.980 71.800 119.330 72.400 ;
        RECT 118.980 71.600 122.930 71.800 ;
        RECT 118.980 71.000 119.330 71.600 ;
        RECT 118.980 70.800 122.930 71.000 ;
        RECT 118.980 70.400 119.330 70.800 ;
        RECT 115.780 62.000 115.980 69.600 ;
        RECT 116.580 62.000 116.780 69.600 ;
        RECT 117.380 62.000 117.580 69.600 ;
        RECT 118.180 62.000 118.380 69.600 ;
        RECT 118.980 69.200 119.330 69.600 ;
        RECT 118.980 69.000 122.930 69.200 ;
        RECT 118.980 68.400 119.330 69.000 ;
        RECT 118.980 68.200 122.930 68.400 ;
        RECT 118.980 67.600 119.330 68.200 ;
        RECT 118.980 67.400 122.930 67.600 ;
        RECT 118.980 66.800 119.330 67.400 ;
        RECT 118.980 66.600 122.930 66.800 ;
        RECT 123.930 66.750 124.330 73.250 ;
        RECT 118.980 66.000 119.330 66.600 ;
        RECT 118.980 65.800 122.930 66.000 ;
        RECT 118.980 65.200 119.330 65.800 ;
        RECT 118.980 65.000 122.930 65.200 ;
        RECT 118.980 64.400 119.330 65.000 ;
        RECT 123.880 64.450 124.730 66.750 ;
        RECT 118.980 64.200 122.930 64.400 ;
        RECT 118.980 63.600 119.330 64.200 ;
        RECT 118.980 63.400 122.930 63.600 ;
        RECT 118.980 62.800 119.330 63.400 ;
        RECT 118.980 62.600 122.930 62.800 ;
        RECT 118.980 62.000 119.330 62.600 ;
        RECT 106.530 61.400 122.930 62.000 ;
        RECT 109.180 60.800 111.480 60.850 ;
        RECT 117.980 60.800 120.280 60.850 ;
        RECT 123.930 60.800 124.330 64.450 ;
        RECT 125.340 62.875 125.700 63.255 ;
        RECT 125.970 62.875 126.330 63.255 ;
        RECT 126.570 62.875 126.930 63.255 ;
        RECT 125.340 62.285 125.700 62.665 ;
        RECT 125.970 62.285 126.330 62.665 ;
        RECT 126.570 62.285 126.930 62.665 ;
        RECT 105.130 60.400 124.330 60.800 ;
        RECT 9.180 59.600 11.480 60.400 ;
        RECT 17.980 59.600 20.280 60.400 ;
        RECT 29.180 59.600 31.480 60.400 ;
        RECT 37.980 59.600 40.280 60.400 ;
        RECT 49.180 59.600 51.480 60.400 ;
        RECT 57.980 59.600 60.280 60.400 ;
        RECT 69.180 59.600 71.480 60.400 ;
        RECT 77.980 59.600 80.280 60.400 ;
        RECT 89.180 59.600 91.480 60.400 ;
        RECT 97.980 59.600 100.280 60.400 ;
        RECT 109.180 59.600 111.480 60.400 ;
        RECT 117.980 59.600 120.280 60.400 ;
        RECT 5.130 59.200 24.330 59.600 ;
        RECT 2.515 57.050 2.875 57.430 ;
        RECT 3.145 57.050 3.505 57.430 ;
        RECT 3.745 57.050 4.105 57.430 ;
        RECT 2.515 56.460 2.875 56.840 ;
        RECT 3.145 56.460 3.505 56.840 ;
        RECT 3.745 56.460 4.105 56.840 ;
        RECT 5.130 55.550 5.530 59.200 ;
        RECT 9.180 59.150 11.480 59.200 ;
        RECT 17.980 59.150 20.280 59.200 ;
        RECT 6.530 58.000 22.930 58.600 ;
        RECT 10.130 57.400 10.480 58.000 ;
        RECT 6.530 57.200 10.480 57.400 ;
        RECT 10.130 56.600 10.480 57.200 ;
        RECT 6.530 56.400 10.480 56.600 ;
        RECT 10.130 55.800 10.480 56.400 ;
        RECT 6.530 55.600 10.480 55.800 ;
        RECT 4.730 55.545 5.580 55.550 ;
        RECT 2.315 53.250 5.580 55.545 ;
        RECT 10.130 55.000 10.480 55.600 ;
        RECT 6.530 54.800 10.480 55.000 ;
        RECT 10.130 54.200 10.480 54.800 ;
        RECT 6.530 54.000 10.480 54.200 ;
        RECT 10.130 53.400 10.480 54.000 ;
        RECT 5.130 46.750 5.530 53.250 ;
        RECT 6.530 53.200 10.480 53.400 ;
        RECT 10.130 52.600 10.480 53.200 ;
        RECT 6.530 52.400 10.480 52.600 ;
        RECT 10.130 51.800 10.480 52.400 ;
        RECT 6.530 51.600 10.480 51.800 ;
        RECT 10.130 51.000 10.480 51.600 ;
        RECT 6.530 50.800 10.480 51.000 ;
        RECT 10.130 50.400 10.480 50.800 ;
        RECT 11.080 50.400 11.280 58.000 ;
        RECT 11.880 50.400 12.080 58.000 ;
        RECT 12.680 50.400 12.880 58.000 ;
        RECT 13.480 50.400 13.680 58.000 ;
        RECT 10.130 49.200 10.480 49.600 ;
        RECT 6.530 49.000 10.480 49.200 ;
        RECT 10.130 48.400 10.480 49.000 ;
        RECT 6.530 48.200 10.480 48.400 ;
        RECT 10.130 47.600 10.480 48.200 ;
        RECT 6.530 47.400 10.480 47.600 ;
        RECT 10.130 46.800 10.480 47.400 ;
        RECT 4.730 46.745 5.580 46.750 ;
        RECT 2.315 44.450 5.580 46.745 ;
        RECT 6.530 46.600 10.480 46.800 ;
        RECT 10.130 46.000 10.480 46.600 ;
        RECT 6.530 45.800 10.480 46.000 ;
        RECT 10.130 45.200 10.480 45.800 ;
        RECT 6.530 45.000 10.480 45.200 ;
        RECT 2.515 42.725 2.875 43.105 ;
        RECT 3.145 42.725 3.505 43.105 ;
        RECT 3.745 42.725 4.105 43.105 ;
        RECT 2.515 42.135 2.875 42.515 ;
        RECT 3.145 42.135 3.505 42.515 ;
        RECT 3.745 42.135 4.105 42.515 ;
        RECT 5.130 40.800 5.530 44.450 ;
        RECT 10.130 44.400 10.480 45.000 ;
        RECT 6.530 44.200 10.480 44.400 ;
        RECT 10.130 43.600 10.480 44.200 ;
        RECT 6.530 43.400 10.480 43.600 ;
        RECT 10.130 42.800 10.480 43.400 ;
        RECT 6.530 42.600 10.480 42.800 ;
        RECT 10.130 42.000 10.480 42.600 ;
        RECT 11.080 42.000 11.280 49.600 ;
        RECT 11.880 42.000 12.080 49.600 ;
        RECT 12.680 42.000 12.880 49.600 ;
        RECT 13.480 42.000 13.680 49.600 ;
        RECT 14.280 42.000 15.180 58.000 ;
        RECT 15.780 50.400 15.980 58.000 ;
        RECT 16.580 50.400 16.780 58.000 ;
        RECT 17.380 50.400 17.580 58.000 ;
        RECT 18.180 50.400 18.380 58.000 ;
        RECT 18.980 57.400 19.330 58.000 ;
        RECT 18.980 57.200 22.930 57.400 ;
        RECT 18.980 56.600 19.330 57.200 ;
        RECT 18.980 56.400 22.930 56.600 ;
        RECT 18.980 55.800 19.330 56.400 ;
        RECT 18.980 55.600 22.930 55.800 ;
        RECT 18.980 55.000 19.330 55.600 ;
        RECT 23.930 55.550 24.330 59.200 ;
        RECT 25.130 59.200 44.330 59.600 ;
        RECT 25.130 55.550 25.530 59.200 ;
        RECT 29.180 59.150 31.480 59.200 ;
        RECT 37.980 59.150 40.280 59.200 ;
        RECT 26.530 58.000 42.930 58.600 ;
        RECT 30.130 57.400 30.480 58.000 ;
        RECT 26.530 57.200 30.480 57.400 ;
        RECT 30.130 56.600 30.480 57.200 ;
        RECT 26.530 56.400 30.480 56.600 ;
        RECT 30.130 55.800 30.480 56.400 ;
        RECT 26.530 55.600 30.480 55.800 ;
        RECT 18.980 54.800 22.930 55.000 ;
        RECT 18.980 54.200 19.330 54.800 ;
        RECT 18.980 54.000 22.930 54.200 ;
        RECT 18.980 53.400 19.330 54.000 ;
        RECT 18.980 53.200 22.930 53.400 ;
        RECT 23.880 53.250 25.580 55.550 ;
        RECT 30.130 55.000 30.480 55.600 ;
        RECT 26.530 54.800 30.480 55.000 ;
        RECT 30.130 54.200 30.480 54.800 ;
        RECT 26.530 54.000 30.480 54.200 ;
        RECT 30.130 53.400 30.480 54.000 ;
        RECT 18.980 52.600 19.330 53.200 ;
        RECT 18.980 52.400 22.930 52.600 ;
        RECT 18.980 51.800 19.330 52.400 ;
        RECT 18.980 51.600 22.930 51.800 ;
        RECT 18.980 51.000 19.330 51.600 ;
        RECT 18.980 50.800 22.930 51.000 ;
        RECT 18.980 50.400 19.330 50.800 ;
        RECT 15.780 42.000 15.980 49.600 ;
        RECT 16.580 42.000 16.780 49.600 ;
        RECT 17.380 42.000 17.580 49.600 ;
        RECT 18.180 42.000 18.380 49.600 ;
        RECT 18.980 49.200 19.330 49.600 ;
        RECT 18.980 49.000 22.930 49.200 ;
        RECT 18.980 48.400 19.330 49.000 ;
        RECT 18.980 48.200 22.930 48.400 ;
        RECT 18.980 47.600 19.330 48.200 ;
        RECT 18.980 47.400 22.930 47.600 ;
        RECT 18.980 46.800 19.330 47.400 ;
        RECT 18.980 46.600 22.930 46.800 ;
        RECT 23.930 46.750 24.330 53.250 ;
        RECT 25.130 46.750 25.530 53.250 ;
        RECT 26.530 53.200 30.480 53.400 ;
        RECT 30.130 52.600 30.480 53.200 ;
        RECT 26.530 52.400 30.480 52.600 ;
        RECT 30.130 51.800 30.480 52.400 ;
        RECT 26.530 51.600 30.480 51.800 ;
        RECT 30.130 51.000 30.480 51.600 ;
        RECT 26.530 50.800 30.480 51.000 ;
        RECT 30.130 50.400 30.480 50.800 ;
        RECT 31.080 50.400 31.280 58.000 ;
        RECT 31.880 50.400 32.080 58.000 ;
        RECT 32.680 50.400 32.880 58.000 ;
        RECT 33.480 50.400 33.680 58.000 ;
        RECT 30.130 49.200 30.480 49.600 ;
        RECT 26.530 49.000 30.480 49.200 ;
        RECT 30.130 48.400 30.480 49.000 ;
        RECT 26.530 48.200 30.480 48.400 ;
        RECT 30.130 47.600 30.480 48.200 ;
        RECT 26.530 47.400 30.480 47.600 ;
        RECT 30.130 46.800 30.480 47.400 ;
        RECT 18.980 46.000 19.330 46.600 ;
        RECT 18.980 45.800 22.930 46.000 ;
        RECT 18.980 45.200 19.330 45.800 ;
        RECT 18.980 45.000 22.930 45.200 ;
        RECT 18.980 44.400 19.330 45.000 ;
        RECT 23.880 44.450 25.580 46.750 ;
        RECT 26.530 46.600 30.480 46.800 ;
        RECT 30.130 46.000 30.480 46.600 ;
        RECT 26.530 45.800 30.480 46.000 ;
        RECT 30.130 45.200 30.480 45.800 ;
        RECT 26.530 45.000 30.480 45.200 ;
        RECT 18.980 44.200 22.930 44.400 ;
        RECT 18.980 43.600 19.330 44.200 ;
        RECT 18.980 43.400 22.930 43.600 ;
        RECT 18.980 42.800 19.330 43.400 ;
        RECT 18.980 42.600 22.930 42.800 ;
        RECT 18.980 42.000 19.330 42.600 ;
        RECT 6.530 41.400 22.930 42.000 ;
        RECT 9.180 40.800 11.480 40.850 ;
        RECT 17.980 40.800 20.280 40.850 ;
        RECT 23.930 40.800 24.330 44.450 ;
        RECT 5.130 40.400 24.330 40.800 ;
        RECT 25.130 40.800 25.530 44.450 ;
        RECT 30.130 44.400 30.480 45.000 ;
        RECT 26.530 44.200 30.480 44.400 ;
        RECT 30.130 43.600 30.480 44.200 ;
        RECT 26.530 43.400 30.480 43.600 ;
        RECT 30.130 42.800 30.480 43.400 ;
        RECT 26.530 42.600 30.480 42.800 ;
        RECT 30.130 42.000 30.480 42.600 ;
        RECT 31.080 42.000 31.280 49.600 ;
        RECT 31.880 42.000 32.080 49.600 ;
        RECT 32.680 42.000 32.880 49.600 ;
        RECT 33.480 42.000 33.680 49.600 ;
        RECT 34.280 42.000 35.180 58.000 ;
        RECT 35.780 50.400 35.980 58.000 ;
        RECT 36.580 50.400 36.780 58.000 ;
        RECT 37.380 50.400 37.580 58.000 ;
        RECT 38.180 50.400 38.380 58.000 ;
        RECT 38.980 57.400 39.330 58.000 ;
        RECT 38.980 57.200 42.930 57.400 ;
        RECT 38.980 56.600 39.330 57.200 ;
        RECT 38.980 56.400 42.930 56.600 ;
        RECT 38.980 55.800 39.330 56.400 ;
        RECT 38.980 55.600 42.930 55.800 ;
        RECT 38.980 55.000 39.330 55.600 ;
        RECT 43.930 55.550 44.330 59.200 ;
        RECT 45.130 59.200 64.330 59.600 ;
        RECT 45.130 55.550 45.530 59.200 ;
        RECT 49.180 59.150 51.480 59.200 ;
        RECT 57.980 59.150 60.280 59.200 ;
        RECT 46.530 58.000 62.930 58.600 ;
        RECT 50.130 57.400 50.480 58.000 ;
        RECT 46.530 57.200 50.480 57.400 ;
        RECT 50.130 56.600 50.480 57.200 ;
        RECT 46.530 56.400 50.480 56.600 ;
        RECT 50.130 55.800 50.480 56.400 ;
        RECT 46.530 55.600 50.480 55.800 ;
        RECT 38.980 54.800 42.930 55.000 ;
        RECT 38.980 54.200 39.330 54.800 ;
        RECT 38.980 54.000 42.930 54.200 ;
        RECT 38.980 53.400 39.330 54.000 ;
        RECT 38.980 53.200 42.930 53.400 ;
        RECT 43.880 53.250 45.580 55.550 ;
        RECT 50.130 55.000 50.480 55.600 ;
        RECT 46.530 54.800 50.480 55.000 ;
        RECT 50.130 54.200 50.480 54.800 ;
        RECT 46.530 54.000 50.480 54.200 ;
        RECT 50.130 53.400 50.480 54.000 ;
        RECT 38.980 52.600 39.330 53.200 ;
        RECT 38.980 52.400 42.930 52.600 ;
        RECT 38.980 51.800 39.330 52.400 ;
        RECT 38.980 51.600 42.930 51.800 ;
        RECT 38.980 51.000 39.330 51.600 ;
        RECT 38.980 50.800 42.930 51.000 ;
        RECT 38.980 50.400 39.330 50.800 ;
        RECT 35.780 42.000 35.980 49.600 ;
        RECT 36.580 42.000 36.780 49.600 ;
        RECT 37.380 42.000 37.580 49.600 ;
        RECT 38.180 42.000 38.380 49.600 ;
        RECT 38.980 49.200 39.330 49.600 ;
        RECT 38.980 49.000 42.930 49.200 ;
        RECT 38.980 48.400 39.330 49.000 ;
        RECT 38.980 48.200 42.930 48.400 ;
        RECT 38.980 47.600 39.330 48.200 ;
        RECT 38.980 47.400 42.930 47.600 ;
        RECT 38.980 46.800 39.330 47.400 ;
        RECT 38.980 46.600 42.930 46.800 ;
        RECT 43.930 46.750 44.330 53.250 ;
        RECT 45.130 46.750 45.530 53.250 ;
        RECT 46.530 53.200 50.480 53.400 ;
        RECT 50.130 52.600 50.480 53.200 ;
        RECT 46.530 52.400 50.480 52.600 ;
        RECT 50.130 51.800 50.480 52.400 ;
        RECT 46.530 51.600 50.480 51.800 ;
        RECT 50.130 51.000 50.480 51.600 ;
        RECT 46.530 50.800 50.480 51.000 ;
        RECT 50.130 50.400 50.480 50.800 ;
        RECT 51.080 50.400 51.280 58.000 ;
        RECT 51.880 50.400 52.080 58.000 ;
        RECT 52.680 50.400 52.880 58.000 ;
        RECT 53.480 50.400 53.680 58.000 ;
        RECT 50.130 49.200 50.480 49.600 ;
        RECT 46.530 49.000 50.480 49.200 ;
        RECT 50.130 48.400 50.480 49.000 ;
        RECT 46.530 48.200 50.480 48.400 ;
        RECT 50.130 47.600 50.480 48.200 ;
        RECT 46.530 47.400 50.480 47.600 ;
        RECT 50.130 46.800 50.480 47.400 ;
        RECT 38.980 46.000 39.330 46.600 ;
        RECT 38.980 45.800 42.930 46.000 ;
        RECT 38.980 45.200 39.330 45.800 ;
        RECT 38.980 45.000 42.930 45.200 ;
        RECT 38.980 44.400 39.330 45.000 ;
        RECT 43.880 44.450 45.580 46.750 ;
        RECT 46.530 46.600 50.480 46.800 ;
        RECT 50.130 46.000 50.480 46.600 ;
        RECT 46.530 45.800 50.480 46.000 ;
        RECT 50.130 45.200 50.480 45.800 ;
        RECT 46.530 45.000 50.480 45.200 ;
        RECT 38.980 44.200 42.930 44.400 ;
        RECT 38.980 43.600 39.330 44.200 ;
        RECT 38.980 43.400 42.930 43.600 ;
        RECT 38.980 42.800 39.330 43.400 ;
        RECT 38.980 42.600 42.930 42.800 ;
        RECT 38.980 42.000 39.330 42.600 ;
        RECT 26.530 41.400 42.930 42.000 ;
        RECT 29.180 40.800 31.480 40.850 ;
        RECT 37.980 40.800 40.280 40.850 ;
        RECT 43.930 40.800 44.330 44.450 ;
        RECT 25.130 40.400 44.330 40.800 ;
        RECT 45.130 40.800 45.530 44.450 ;
        RECT 50.130 44.400 50.480 45.000 ;
        RECT 46.530 44.200 50.480 44.400 ;
        RECT 50.130 43.600 50.480 44.200 ;
        RECT 46.530 43.400 50.480 43.600 ;
        RECT 50.130 42.800 50.480 43.400 ;
        RECT 46.530 42.600 50.480 42.800 ;
        RECT 50.130 42.000 50.480 42.600 ;
        RECT 51.080 42.000 51.280 49.600 ;
        RECT 51.880 42.000 52.080 49.600 ;
        RECT 52.680 42.000 52.880 49.600 ;
        RECT 53.480 42.000 53.680 49.600 ;
        RECT 54.280 42.000 55.180 58.000 ;
        RECT 55.780 50.400 55.980 58.000 ;
        RECT 56.580 50.400 56.780 58.000 ;
        RECT 57.380 50.400 57.580 58.000 ;
        RECT 58.180 50.400 58.380 58.000 ;
        RECT 58.980 57.400 59.330 58.000 ;
        RECT 58.980 57.200 62.930 57.400 ;
        RECT 58.980 56.600 59.330 57.200 ;
        RECT 58.980 56.400 62.930 56.600 ;
        RECT 58.980 55.800 59.330 56.400 ;
        RECT 58.980 55.600 62.930 55.800 ;
        RECT 58.980 55.000 59.330 55.600 ;
        RECT 63.930 55.550 64.330 59.200 ;
        RECT 65.130 59.200 84.330 59.600 ;
        RECT 65.130 55.550 65.530 59.200 ;
        RECT 69.180 59.150 71.480 59.200 ;
        RECT 77.980 59.150 80.280 59.200 ;
        RECT 66.530 58.000 82.930 58.600 ;
        RECT 70.130 57.400 70.480 58.000 ;
        RECT 66.530 57.200 70.480 57.400 ;
        RECT 70.130 56.600 70.480 57.200 ;
        RECT 66.530 56.400 70.480 56.600 ;
        RECT 70.130 55.800 70.480 56.400 ;
        RECT 66.530 55.600 70.480 55.800 ;
        RECT 58.980 54.800 62.930 55.000 ;
        RECT 58.980 54.200 59.330 54.800 ;
        RECT 58.980 54.000 62.930 54.200 ;
        RECT 58.980 53.400 59.330 54.000 ;
        RECT 58.980 53.200 62.930 53.400 ;
        RECT 63.880 53.250 65.580 55.550 ;
        RECT 70.130 55.000 70.480 55.600 ;
        RECT 66.530 54.800 70.480 55.000 ;
        RECT 70.130 54.200 70.480 54.800 ;
        RECT 66.530 54.000 70.480 54.200 ;
        RECT 70.130 53.400 70.480 54.000 ;
        RECT 58.980 52.600 59.330 53.200 ;
        RECT 58.980 52.400 62.930 52.600 ;
        RECT 58.980 51.800 59.330 52.400 ;
        RECT 58.980 51.600 62.930 51.800 ;
        RECT 58.980 51.000 59.330 51.600 ;
        RECT 58.980 50.800 62.930 51.000 ;
        RECT 58.980 50.400 59.330 50.800 ;
        RECT 55.780 42.000 55.980 49.600 ;
        RECT 56.580 42.000 56.780 49.600 ;
        RECT 57.380 42.000 57.580 49.600 ;
        RECT 58.180 42.000 58.380 49.600 ;
        RECT 58.980 49.200 59.330 49.600 ;
        RECT 58.980 49.000 62.930 49.200 ;
        RECT 58.980 48.400 59.330 49.000 ;
        RECT 58.980 48.200 62.930 48.400 ;
        RECT 58.980 47.600 59.330 48.200 ;
        RECT 58.980 47.400 62.930 47.600 ;
        RECT 58.980 46.800 59.330 47.400 ;
        RECT 58.980 46.600 62.930 46.800 ;
        RECT 63.930 46.750 64.330 53.250 ;
        RECT 65.130 46.750 65.530 53.250 ;
        RECT 66.530 53.200 70.480 53.400 ;
        RECT 70.130 52.600 70.480 53.200 ;
        RECT 66.530 52.400 70.480 52.600 ;
        RECT 70.130 51.800 70.480 52.400 ;
        RECT 66.530 51.600 70.480 51.800 ;
        RECT 70.130 51.000 70.480 51.600 ;
        RECT 66.530 50.800 70.480 51.000 ;
        RECT 70.130 50.400 70.480 50.800 ;
        RECT 71.080 50.400 71.280 58.000 ;
        RECT 71.880 50.400 72.080 58.000 ;
        RECT 72.680 50.400 72.880 58.000 ;
        RECT 73.480 50.400 73.680 58.000 ;
        RECT 70.130 49.200 70.480 49.600 ;
        RECT 66.530 49.000 70.480 49.200 ;
        RECT 70.130 48.400 70.480 49.000 ;
        RECT 66.530 48.200 70.480 48.400 ;
        RECT 70.130 47.600 70.480 48.200 ;
        RECT 66.530 47.400 70.480 47.600 ;
        RECT 70.130 46.800 70.480 47.400 ;
        RECT 58.980 46.000 59.330 46.600 ;
        RECT 58.980 45.800 62.930 46.000 ;
        RECT 58.980 45.200 59.330 45.800 ;
        RECT 58.980 45.000 62.930 45.200 ;
        RECT 58.980 44.400 59.330 45.000 ;
        RECT 63.880 44.450 65.580 46.750 ;
        RECT 66.530 46.600 70.480 46.800 ;
        RECT 70.130 46.000 70.480 46.600 ;
        RECT 66.530 45.800 70.480 46.000 ;
        RECT 70.130 45.200 70.480 45.800 ;
        RECT 66.530 45.000 70.480 45.200 ;
        RECT 58.980 44.200 62.930 44.400 ;
        RECT 58.980 43.600 59.330 44.200 ;
        RECT 58.980 43.400 62.930 43.600 ;
        RECT 58.980 42.800 59.330 43.400 ;
        RECT 58.980 42.600 62.930 42.800 ;
        RECT 58.980 42.000 59.330 42.600 ;
        RECT 46.530 41.400 62.930 42.000 ;
        RECT 49.180 40.800 51.480 40.850 ;
        RECT 57.980 40.800 60.280 40.850 ;
        RECT 63.930 40.800 64.330 44.450 ;
        RECT 45.130 40.400 64.330 40.800 ;
        RECT 65.130 40.800 65.530 44.450 ;
        RECT 70.130 44.400 70.480 45.000 ;
        RECT 66.530 44.200 70.480 44.400 ;
        RECT 70.130 43.600 70.480 44.200 ;
        RECT 66.530 43.400 70.480 43.600 ;
        RECT 70.130 42.800 70.480 43.400 ;
        RECT 66.530 42.600 70.480 42.800 ;
        RECT 70.130 42.000 70.480 42.600 ;
        RECT 71.080 42.000 71.280 49.600 ;
        RECT 71.880 42.000 72.080 49.600 ;
        RECT 72.680 42.000 72.880 49.600 ;
        RECT 73.480 42.000 73.680 49.600 ;
        RECT 74.280 42.000 75.180 58.000 ;
        RECT 75.780 50.400 75.980 58.000 ;
        RECT 76.580 50.400 76.780 58.000 ;
        RECT 77.380 50.400 77.580 58.000 ;
        RECT 78.180 50.400 78.380 58.000 ;
        RECT 78.980 57.400 79.330 58.000 ;
        RECT 78.980 57.200 82.930 57.400 ;
        RECT 78.980 56.600 79.330 57.200 ;
        RECT 78.980 56.400 82.930 56.600 ;
        RECT 78.980 55.800 79.330 56.400 ;
        RECT 78.980 55.600 82.930 55.800 ;
        RECT 78.980 55.000 79.330 55.600 ;
        RECT 83.930 55.550 84.330 59.200 ;
        RECT 85.130 59.200 104.330 59.600 ;
        RECT 85.130 55.550 85.530 59.200 ;
        RECT 89.180 59.150 91.480 59.200 ;
        RECT 97.980 59.150 100.280 59.200 ;
        RECT 86.530 58.000 102.930 58.600 ;
        RECT 90.130 57.400 90.480 58.000 ;
        RECT 86.530 57.200 90.480 57.400 ;
        RECT 90.130 56.600 90.480 57.200 ;
        RECT 86.530 56.400 90.480 56.600 ;
        RECT 90.130 55.800 90.480 56.400 ;
        RECT 86.530 55.600 90.480 55.800 ;
        RECT 78.980 54.800 82.930 55.000 ;
        RECT 78.980 54.200 79.330 54.800 ;
        RECT 78.980 54.000 82.930 54.200 ;
        RECT 78.980 53.400 79.330 54.000 ;
        RECT 78.980 53.200 82.930 53.400 ;
        RECT 83.880 53.250 85.580 55.550 ;
        RECT 90.130 55.000 90.480 55.600 ;
        RECT 86.530 54.800 90.480 55.000 ;
        RECT 90.130 54.200 90.480 54.800 ;
        RECT 86.530 54.000 90.480 54.200 ;
        RECT 90.130 53.400 90.480 54.000 ;
        RECT 78.980 52.600 79.330 53.200 ;
        RECT 78.980 52.400 82.930 52.600 ;
        RECT 78.980 51.800 79.330 52.400 ;
        RECT 78.980 51.600 82.930 51.800 ;
        RECT 78.980 51.000 79.330 51.600 ;
        RECT 78.980 50.800 82.930 51.000 ;
        RECT 78.980 50.400 79.330 50.800 ;
        RECT 75.780 42.000 75.980 49.600 ;
        RECT 76.580 42.000 76.780 49.600 ;
        RECT 77.380 42.000 77.580 49.600 ;
        RECT 78.180 42.000 78.380 49.600 ;
        RECT 78.980 49.200 79.330 49.600 ;
        RECT 78.980 49.000 82.930 49.200 ;
        RECT 78.980 48.400 79.330 49.000 ;
        RECT 78.980 48.200 82.930 48.400 ;
        RECT 78.980 47.600 79.330 48.200 ;
        RECT 78.980 47.400 82.930 47.600 ;
        RECT 78.980 46.800 79.330 47.400 ;
        RECT 78.980 46.600 82.930 46.800 ;
        RECT 83.930 46.750 84.330 53.250 ;
        RECT 85.130 46.750 85.530 53.250 ;
        RECT 86.530 53.200 90.480 53.400 ;
        RECT 90.130 52.600 90.480 53.200 ;
        RECT 86.530 52.400 90.480 52.600 ;
        RECT 90.130 51.800 90.480 52.400 ;
        RECT 86.530 51.600 90.480 51.800 ;
        RECT 90.130 51.000 90.480 51.600 ;
        RECT 86.530 50.800 90.480 51.000 ;
        RECT 90.130 50.400 90.480 50.800 ;
        RECT 91.080 50.400 91.280 58.000 ;
        RECT 91.880 50.400 92.080 58.000 ;
        RECT 92.680 50.400 92.880 58.000 ;
        RECT 93.480 50.400 93.680 58.000 ;
        RECT 90.130 49.200 90.480 49.600 ;
        RECT 86.530 49.000 90.480 49.200 ;
        RECT 90.130 48.400 90.480 49.000 ;
        RECT 86.530 48.200 90.480 48.400 ;
        RECT 90.130 47.600 90.480 48.200 ;
        RECT 86.530 47.400 90.480 47.600 ;
        RECT 90.130 46.800 90.480 47.400 ;
        RECT 78.980 46.000 79.330 46.600 ;
        RECT 78.980 45.800 82.930 46.000 ;
        RECT 78.980 45.200 79.330 45.800 ;
        RECT 78.980 45.000 82.930 45.200 ;
        RECT 78.980 44.400 79.330 45.000 ;
        RECT 83.880 44.450 85.580 46.750 ;
        RECT 86.530 46.600 90.480 46.800 ;
        RECT 90.130 46.000 90.480 46.600 ;
        RECT 86.530 45.800 90.480 46.000 ;
        RECT 90.130 45.200 90.480 45.800 ;
        RECT 86.530 45.000 90.480 45.200 ;
        RECT 78.980 44.200 82.930 44.400 ;
        RECT 78.980 43.600 79.330 44.200 ;
        RECT 78.980 43.400 82.930 43.600 ;
        RECT 78.980 42.800 79.330 43.400 ;
        RECT 78.980 42.600 82.930 42.800 ;
        RECT 78.980 42.000 79.330 42.600 ;
        RECT 66.530 41.400 82.930 42.000 ;
        RECT 69.180 40.800 71.480 40.850 ;
        RECT 77.980 40.800 80.280 40.850 ;
        RECT 83.930 40.800 84.330 44.450 ;
        RECT 65.130 40.400 84.330 40.800 ;
        RECT 85.130 40.800 85.530 44.450 ;
        RECT 90.130 44.400 90.480 45.000 ;
        RECT 86.530 44.200 90.480 44.400 ;
        RECT 90.130 43.600 90.480 44.200 ;
        RECT 86.530 43.400 90.480 43.600 ;
        RECT 90.130 42.800 90.480 43.400 ;
        RECT 86.530 42.600 90.480 42.800 ;
        RECT 90.130 42.000 90.480 42.600 ;
        RECT 91.080 42.000 91.280 49.600 ;
        RECT 91.880 42.000 92.080 49.600 ;
        RECT 92.680 42.000 92.880 49.600 ;
        RECT 93.480 42.000 93.680 49.600 ;
        RECT 94.280 42.000 95.180 58.000 ;
        RECT 95.780 50.400 95.980 58.000 ;
        RECT 96.580 50.400 96.780 58.000 ;
        RECT 97.380 50.400 97.580 58.000 ;
        RECT 98.180 50.400 98.380 58.000 ;
        RECT 98.980 57.400 99.330 58.000 ;
        RECT 98.980 57.200 102.930 57.400 ;
        RECT 98.980 56.600 99.330 57.200 ;
        RECT 98.980 56.400 102.930 56.600 ;
        RECT 98.980 55.800 99.330 56.400 ;
        RECT 98.980 55.600 102.930 55.800 ;
        RECT 98.980 55.000 99.330 55.600 ;
        RECT 103.930 55.550 104.330 59.200 ;
        RECT 105.130 59.200 124.330 59.600 ;
        RECT 105.130 55.550 105.530 59.200 ;
        RECT 109.180 59.150 111.480 59.200 ;
        RECT 117.980 59.150 120.280 59.200 ;
        RECT 106.530 58.000 122.930 58.600 ;
        RECT 110.130 57.400 110.480 58.000 ;
        RECT 106.530 57.200 110.480 57.400 ;
        RECT 110.130 56.600 110.480 57.200 ;
        RECT 106.530 56.400 110.480 56.600 ;
        RECT 110.130 55.800 110.480 56.400 ;
        RECT 106.530 55.600 110.480 55.800 ;
        RECT 98.980 54.800 102.930 55.000 ;
        RECT 98.980 54.200 99.330 54.800 ;
        RECT 98.980 54.000 102.930 54.200 ;
        RECT 98.980 53.400 99.330 54.000 ;
        RECT 98.980 53.200 102.930 53.400 ;
        RECT 103.880 53.250 105.580 55.550 ;
        RECT 110.130 55.000 110.480 55.600 ;
        RECT 106.530 54.800 110.480 55.000 ;
        RECT 110.130 54.200 110.480 54.800 ;
        RECT 106.530 54.000 110.480 54.200 ;
        RECT 110.130 53.400 110.480 54.000 ;
        RECT 98.980 52.600 99.330 53.200 ;
        RECT 98.980 52.400 102.930 52.600 ;
        RECT 98.980 51.800 99.330 52.400 ;
        RECT 98.980 51.600 102.930 51.800 ;
        RECT 98.980 51.000 99.330 51.600 ;
        RECT 98.980 50.800 102.930 51.000 ;
        RECT 98.980 50.400 99.330 50.800 ;
        RECT 95.780 42.000 95.980 49.600 ;
        RECT 96.580 42.000 96.780 49.600 ;
        RECT 97.380 42.000 97.580 49.600 ;
        RECT 98.180 42.000 98.380 49.600 ;
        RECT 98.980 49.200 99.330 49.600 ;
        RECT 98.980 49.000 102.930 49.200 ;
        RECT 98.980 48.400 99.330 49.000 ;
        RECT 98.980 48.200 102.930 48.400 ;
        RECT 98.980 47.600 99.330 48.200 ;
        RECT 98.980 47.400 102.930 47.600 ;
        RECT 98.980 46.800 99.330 47.400 ;
        RECT 98.980 46.600 102.930 46.800 ;
        RECT 103.930 46.750 104.330 53.250 ;
        RECT 105.130 46.750 105.530 53.250 ;
        RECT 106.530 53.200 110.480 53.400 ;
        RECT 110.130 52.600 110.480 53.200 ;
        RECT 106.530 52.400 110.480 52.600 ;
        RECT 110.130 51.800 110.480 52.400 ;
        RECT 106.530 51.600 110.480 51.800 ;
        RECT 110.130 51.000 110.480 51.600 ;
        RECT 106.530 50.800 110.480 51.000 ;
        RECT 110.130 50.400 110.480 50.800 ;
        RECT 111.080 50.400 111.280 58.000 ;
        RECT 111.880 50.400 112.080 58.000 ;
        RECT 112.680 50.400 112.880 58.000 ;
        RECT 113.480 50.400 113.680 58.000 ;
        RECT 110.130 49.200 110.480 49.600 ;
        RECT 106.530 49.000 110.480 49.200 ;
        RECT 110.130 48.400 110.480 49.000 ;
        RECT 106.530 48.200 110.480 48.400 ;
        RECT 110.130 47.600 110.480 48.200 ;
        RECT 106.530 47.400 110.480 47.600 ;
        RECT 110.130 46.800 110.480 47.400 ;
        RECT 98.980 46.000 99.330 46.600 ;
        RECT 98.980 45.800 102.930 46.000 ;
        RECT 98.980 45.200 99.330 45.800 ;
        RECT 98.980 45.000 102.930 45.200 ;
        RECT 98.980 44.400 99.330 45.000 ;
        RECT 103.880 44.450 105.580 46.750 ;
        RECT 106.530 46.600 110.480 46.800 ;
        RECT 110.130 46.000 110.480 46.600 ;
        RECT 106.530 45.800 110.480 46.000 ;
        RECT 110.130 45.200 110.480 45.800 ;
        RECT 106.530 45.000 110.480 45.200 ;
        RECT 98.980 44.200 102.930 44.400 ;
        RECT 98.980 43.600 99.330 44.200 ;
        RECT 98.980 43.400 102.930 43.600 ;
        RECT 98.980 42.800 99.330 43.400 ;
        RECT 98.980 42.600 102.930 42.800 ;
        RECT 98.980 42.000 99.330 42.600 ;
        RECT 86.530 41.400 102.930 42.000 ;
        RECT 89.180 40.800 91.480 40.850 ;
        RECT 97.980 40.800 100.280 40.850 ;
        RECT 103.930 40.800 104.330 44.450 ;
        RECT 85.130 40.400 104.330 40.800 ;
        RECT 105.130 40.800 105.530 44.450 ;
        RECT 110.130 44.400 110.480 45.000 ;
        RECT 106.530 44.200 110.480 44.400 ;
        RECT 110.130 43.600 110.480 44.200 ;
        RECT 106.530 43.400 110.480 43.600 ;
        RECT 110.130 42.800 110.480 43.400 ;
        RECT 106.530 42.600 110.480 42.800 ;
        RECT 110.130 42.000 110.480 42.600 ;
        RECT 111.080 42.000 111.280 49.600 ;
        RECT 111.880 42.000 112.080 49.600 ;
        RECT 112.680 42.000 112.880 49.600 ;
        RECT 113.480 42.000 113.680 49.600 ;
        RECT 114.280 42.000 115.180 58.000 ;
        RECT 115.780 50.400 115.980 58.000 ;
        RECT 116.580 50.400 116.780 58.000 ;
        RECT 117.380 50.400 117.580 58.000 ;
        RECT 118.180 50.400 118.380 58.000 ;
        RECT 118.980 57.400 119.330 58.000 ;
        RECT 118.980 57.200 122.930 57.400 ;
        RECT 118.980 56.600 119.330 57.200 ;
        RECT 118.980 56.400 122.930 56.600 ;
        RECT 118.980 55.800 119.330 56.400 ;
        RECT 118.980 55.600 122.930 55.800 ;
        RECT 118.980 55.000 119.330 55.600 ;
        RECT 123.930 55.550 124.330 59.200 ;
        RECT 125.340 56.805 125.700 57.185 ;
        RECT 125.970 56.805 126.330 57.185 ;
        RECT 126.570 56.805 126.930 57.185 ;
        RECT 125.340 56.215 125.700 56.595 ;
        RECT 125.970 56.215 126.330 56.595 ;
        RECT 126.570 56.215 126.930 56.595 ;
        RECT 118.980 54.800 122.930 55.000 ;
        RECT 118.980 54.200 119.330 54.800 ;
        RECT 118.980 54.000 122.930 54.200 ;
        RECT 118.980 53.400 119.330 54.000 ;
        RECT 118.980 53.200 122.930 53.400 ;
        RECT 123.880 53.250 124.730 55.550 ;
        RECT 118.980 52.600 119.330 53.200 ;
        RECT 118.980 52.400 122.930 52.600 ;
        RECT 118.980 51.800 119.330 52.400 ;
        RECT 118.980 51.600 122.930 51.800 ;
        RECT 118.980 51.000 119.330 51.600 ;
        RECT 118.980 50.800 122.930 51.000 ;
        RECT 118.980 50.400 119.330 50.800 ;
        RECT 115.780 42.000 115.980 49.600 ;
        RECT 116.580 42.000 116.780 49.600 ;
        RECT 117.380 42.000 117.580 49.600 ;
        RECT 118.180 42.000 118.380 49.600 ;
        RECT 118.980 49.200 119.330 49.600 ;
        RECT 118.980 49.000 122.930 49.200 ;
        RECT 118.980 48.400 119.330 49.000 ;
        RECT 118.980 48.200 122.930 48.400 ;
        RECT 118.980 47.600 119.330 48.200 ;
        RECT 118.980 47.400 122.930 47.600 ;
        RECT 118.980 46.800 119.330 47.400 ;
        RECT 118.980 46.600 122.930 46.800 ;
        RECT 123.930 46.750 124.330 53.250 ;
        RECT 118.980 46.000 119.330 46.600 ;
        RECT 118.980 45.800 122.930 46.000 ;
        RECT 118.980 45.200 119.330 45.800 ;
        RECT 118.980 45.000 122.930 45.200 ;
        RECT 118.980 44.400 119.330 45.000 ;
        RECT 123.880 44.450 124.730 46.750 ;
        RECT 118.980 44.200 122.930 44.400 ;
        RECT 118.980 43.600 119.330 44.200 ;
        RECT 118.980 43.400 122.930 43.600 ;
        RECT 118.980 42.800 119.330 43.400 ;
        RECT 118.980 42.600 122.930 42.800 ;
        RECT 118.980 42.000 119.330 42.600 ;
        RECT 106.530 41.400 122.930 42.000 ;
        RECT 109.180 40.800 111.480 40.850 ;
        RECT 117.980 40.800 120.280 40.850 ;
        RECT 123.930 40.800 124.330 44.450 ;
        RECT 125.340 42.590 125.700 42.970 ;
        RECT 125.970 42.590 126.330 42.970 ;
        RECT 126.570 42.590 126.930 42.970 ;
        RECT 125.340 42.000 125.700 42.380 ;
        RECT 125.970 42.000 126.330 42.380 ;
        RECT 126.570 42.000 126.930 42.380 ;
        RECT 105.130 40.400 124.330 40.800 ;
        RECT 9.180 39.600 11.480 40.400 ;
        RECT 17.980 39.600 20.280 40.400 ;
        RECT 29.180 39.600 31.480 40.400 ;
        RECT 37.980 39.600 40.280 40.400 ;
        RECT 49.180 39.600 51.480 40.400 ;
        RECT 57.980 39.600 60.280 40.400 ;
        RECT 69.180 39.600 71.480 40.400 ;
        RECT 77.980 39.600 80.280 40.400 ;
        RECT 89.180 39.600 91.480 40.400 ;
        RECT 97.980 39.600 100.280 40.400 ;
        RECT 109.180 39.600 111.480 40.400 ;
        RECT 117.980 39.600 120.280 40.400 ;
        RECT 5.130 39.200 24.330 39.600 ;
        RECT 2.515 37.115 2.875 37.495 ;
        RECT 3.145 37.115 3.505 37.495 ;
        RECT 3.745 37.115 4.105 37.495 ;
        RECT 2.515 36.525 2.875 36.905 ;
        RECT 3.145 36.525 3.505 36.905 ;
        RECT 3.745 36.525 4.105 36.905 ;
        RECT 5.130 35.550 5.530 39.200 ;
        RECT 9.180 39.150 11.480 39.200 ;
        RECT 17.980 39.150 20.280 39.200 ;
        RECT 6.530 38.000 22.930 38.600 ;
        RECT 10.130 37.400 10.480 38.000 ;
        RECT 6.530 37.200 10.480 37.400 ;
        RECT 10.130 36.600 10.480 37.200 ;
        RECT 6.530 36.400 10.480 36.600 ;
        RECT 10.130 35.800 10.480 36.400 ;
        RECT 6.530 35.600 10.480 35.800 ;
        RECT 2.315 33.255 5.580 35.550 ;
        RECT 10.130 35.000 10.480 35.600 ;
        RECT 6.530 34.800 10.480 35.000 ;
        RECT 10.130 34.200 10.480 34.800 ;
        RECT 6.530 34.000 10.480 34.200 ;
        RECT 10.130 33.400 10.480 34.000 ;
        RECT 4.730 33.250 5.580 33.255 ;
        RECT 5.130 26.750 5.530 33.250 ;
        RECT 6.530 33.200 10.480 33.400 ;
        RECT 10.130 32.600 10.480 33.200 ;
        RECT 6.530 32.400 10.480 32.600 ;
        RECT 10.130 31.800 10.480 32.400 ;
        RECT 6.530 31.600 10.480 31.800 ;
        RECT 10.130 31.000 10.480 31.600 ;
        RECT 6.530 30.800 10.480 31.000 ;
        RECT 10.130 30.400 10.480 30.800 ;
        RECT 11.080 30.400 11.280 38.000 ;
        RECT 11.880 30.400 12.080 38.000 ;
        RECT 12.680 30.400 12.880 38.000 ;
        RECT 13.480 30.400 13.680 38.000 ;
        RECT 10.130 29.200 10.480 29.600 ;
        RECT 6.530 29.000 10.480 29.200 ;
        RECT 10.130 28.400 10.480 29.000 ;
        RECT 6.530 28.200 10.480 28.400 ;
        RECT 10.130 27.600 10.480 28.200 ;
        RECT 6.530 27.400 10.480 27.600 ;
        RECT 10.130 26.800 10.480 27.400 ;
        RECT 4.730 26.740 5.580 26.750 ;
        RECT 2.315 24.450 5.580 26.740 ;
        RECT 6.530 26.600 10.480 26.800 ;
        RECT 10.130 26.000 10.480 26.600 ;
        RECT 6.530 25.800 10.480 26.000 ;
        RECT 10.130 25.200 10.480 25.800 ;
        RECT 6.530 25.000 10.480 25.200 ;
        RECT 2.315 24.445 4.730 24.450 ;
        RECT 2.515 22.815 2.875 23.195 ;
        RECT 3.145 22.815 3.505 23.195 ;
        RECT 3.745 22.815 4.105 23.195 ;
        RECT 2.515 22.225 2.875 22.605 ;
        RECT 3.145 22.225 3.505 22.605 ;
        RECT 3.745 22.225 4.105 22.605 ;
        RECT 5.130 20.800 5.530 24.450 ;
        RECT 10.130 24.400 10.480 25.000 ;
        RECT 6.530 24.200 10.480 24.400 ;
        RECT 10.130 23.600 10.480 24.200 ;
        RECT 6.530 23.400 10.480 23.600 ;
        RECT 10.130 22.800 10.480 23.400 ;
        RECT 6.530 22.600 10.480 22.800 ;
        RECT 10.130 22.000 10.480 22.600 ;
        RECT 11.080 22.000 11.280 29.600 ;
        RECT 11.880 22.000 12.080 29.600 ;
        RECT 12.680 22.000 12.880 29.600 ;
        RECT 13.480 22.000 13.680 29.600 ;
        RECT 14.280 22.000 15.180 38.000 ;
        RECT 15.780 30.400 15.980 38.000 ;
        RECT 16.580 30.400 16.780 38.000 ;
        RECT 17.380 30.400 17.580 38.000 ;
        RECT 18.180 30.400 18.380 38.000 ;
        RECT 18.980 37.400 19.330 38.000 ;
        RECT 18.980 37.200 22.930 37.400 ;
        RECT 18.980 36.600 19.330 37.200 ;
        RECT 18.980 36.400 22.930 36.600 ;
        RECT 18.980 35.800 19.330 36.400 ;
        RECT 18.980 35.600 22.930 35.800 ;
        RECT 18.980 35.000 19.330 35.600 ;
        RECT 23.930 35.550 24.330 39.200 ;
        RECT 25.130 39.200 44.330 39.600 ;
        RECT 25.130 35.550 25.530 39.200 ;
        RECT 29.180 39.150 31.480 39.200 ;
        RECT 37.980 39.150 40.280 39.200 ;
        RECT 26.530 38.000 42.930 38.600 ;
        RECT 30.130 37.400 30.480 38.000 ;
        RECT 26.530 37.200 30.480 37.400 ;
        RECT 30.130 36.600 30.480 37.200 ;
        RECT 26.530 36.400 30.480 36.600 ;
        RECT 30.130 35.800 30.480 36.400 ;
        RECT 26.530 35.600 30.480 35.800 ;
        RECT 18.980 34.800 22.930 35.000 ;
        RECT 18.980 34.200 19.330 34.800 ;
        RECT 18.980 34.000 22.930 34.200 ;
        RECT 18.980 33.400 19.330 34.000 ;
        RECT 18.980 33.200 22.930 33.400 ;
        RECT 23.880 33.250 25.580 35.550 ;
        RECT 30.130 35.000 30.480 35.600 ;
        RECT 26.530 34.800 30.480 35.000 ;
        RECT 30.130 34.200 30.480 34.800 ;
        RECT 26.530 34.000 30.480 34.200 ;
        RECT 30.130 33.400 30.480 34.000 ;
        RECT 18.980 32.600 19.330 33.200 ;
        RECT 18.980 32.400 22.930 32.600 ;
        RECT 18.980 31.800 19.330 32.400 ;
        RECT 18.980 31.600 22.930 31.800 ;
        RECT 18.980 31.000 19.330 31.600 ;
        RECT 18.980 30.800 22.930 31.000 ;
        RECT 18.980 30.400 19.330 30.800 ;
        RECT 15.780 22.000 15.980 29.600 ;
        RECT 16.580 22.000 16.780 29.600 ;
        RECT 17.380 22.000 17.580 29.600 ;
        RECT 18.180 22.000 18.380 29.600 ;
        RECT 18.980 29.200 19.330 29.600 ;
        RECT 18.980 29.000 22.930 29.200 ;
        RECT 18.980 28.400 19.330 29.000 ;
        RECT 18.980 28.200 22.930 28.400 ;
        RECT 18.980 27.600 19.330 28.200 ;
        RECT 18.980 27.400 22.930 27.600 ;
        RECT 18.980 26.800 19.330 27.400 ;
        RECT 18.980 26.600 22.930 26.800 ;
        RECT 23.930 26.750 24.330 33.250 ;
        RECT 25.130 26.750 25.530 33.250 ;
        RECT 26.530 33.200 30.480 33.400 ;
        RECT 30.130 32.600 30.480 33.200 ;
        RECT 26.530 32.400 30.480 32.600 ;
        RECT 30.130 31.800 30.480 32.400 ;
        RECT 26.530 31.600 30.480 31.800 ;
        RECT 30.130 31.000 30.480 31.600 ;
        RECT 26.530 30.800 30.480 31.000 ;
        RECT 30.130 30.400 30.480 30.800 ;
        RECT 31.080 30.400 31.280 38.000 ;
        RECT 31.880 30.400 32.080 38.000 ;
        RECT 32.680 30.400 32.880 38.000 ;
        RECT 33.480 30.400 33.680 38.000 ;
        RECT 30.130 29.200 30.480 29.600 ;
        RECT 26.530 29.000 30.480 29.200 ;
        RECT 30.130 28.400 30.480 29.000 ;
        RECT 26.530 28.200 30.480 28.400 ;
        RECT 30.130 27.600 30.480 28.200 ;
        RECT 26.530 27.400 30.480 27.600 ;
        RECT 30.130 26.800 30.480 27.400 ;
        RECT 18.980 26.000 19.330 26.600 ;
        RECT 18.980 25.800 22.930 26.000 ;
        RECT 18.980 25.200 19.330 25.800 ;
        RECT 18.980 25.000 22.930 25.200 ;
        RECT 18.980 24.400 19.330 25.000 ;
        RECT 23.880 24.450 25.580 26.750 ;
        RECT 26.530 26.600 30.480 26.800 ;
        RECT 30.130 26.000 30.480 26.600 ;
        RECT 26.530 25.800 30.480 26.000 ;
        RECT 30.130 25.200 30.480 25.800 ;
        RECT 26.530 25.000 30.480 25.200 ;
        RECT 18.980 24.200 22.930 24.400 ;
        RECT 18.980 23.600 19.330 24.200 ;
        RECT 18.980 23.400 22.930 23.600 ;
        RECT 18.980 22.800 19.330 23.400 ;
        RECT 18.980 22.600 22.930 22.800 ;
        RECT 18.980 22.000 19.330 22.600 ;
        RECT 6.530 21.400 22.930 22.000 ;
        RECT 9.180 20.800 11.480 20.850 ;
        RECT 17.980 20.800 20.280 20.850 ;
        RECT 23.930 20.800 24.330 24.450 ;
        RECT 5.130 20.400 24.330 20.800 ;
        RECT 25.130 20.800 25.530 24.450 ;
        RECT 30.130 24.400 30.480 25.000 ;
        RECT 26.530 24.200 30.480 24.400 ;
        RECT 30.130 23.600 30.480 24.200 ;
        RECT 26.530 23.400 30.480 23.600 ;
        RECT 30.130 22.800 30.480 23.400 ;
        RECT 26.530 22.600 30.480 22.800 ;
        RECT 30.130 22.000 30.480 22.600 ;
        RECT 31.080 22.000 31.280 29.600 ;
        RECT 31.880 22.000 32.080 29.600 ;
        RECT 32.680 22.000 32.880 29.600 ;
        RECT 33.480 22.000 33.680 29.600 ;
        RECT 34.280 22.000 35.180 38.000 ;
        RECT 35.780 30.400 35.980 38.000 ;
        RECT 36.580 30.400 36.780 38.000 ;
        RECT 37.380 30.400 37.580 38.000 ;
        RECT 38.180 30.400 38.380 38.000 ;
        RECT 38.980 37.400 39.330 38.000 ;
        RECT 38.980 37.200 42.930 37.400 ;
        RECT 38.980 36.600 39.330 37.200 ;
        RECT 38.980 36.400 42.930 36.600 ;
        RECT 38.980 35.800 39.330 36.400 ;
        RECT 38.980 35.600 42.930 35.800 ;
        RECT 38.980 35.000 39.330 35.600 ;
        RECT 43.930 35.550 44.330 39.200 ;
        RECT 45.130 39.200 64.330 39.600 ;
        RECT 45.130 35.550 45.530 39.200 ;
        RECT 49.180 39.150 51.480 39.200 ;
        RECT 57.980 39.150 60.280 39.200 ;
        RECT 46.530 38.000 62.930 38.600 ;
        RECT 50.130 37.400 50.480 38.000 ;
        RECT 46.530 37.200 50.480 37.400 ;
        RECT 50.130 36.600 50.480 37.200 ;
        RECT 46.530 36.400 50.480 36.600 ;
        RECT 50.130 35.800 50.480 36.400 ;
        RECT 46.530 35.600 50.480 35.800 ;
        RECT 38.980 34.800 42.930 35.000 ;
        RECT 38.980 34.200 39.330 34.800 ;
        RECT 38.980 34.000 42.930 34.200 ;
        RECT 38.980 33.400 39.330 34.000 ;
        RECT 38.980 33.200 42.930 33.400 ;
        RECT 43.880 33.250 45.580 35.550 ;
        RECT 50.130 35.000 50.480 35.600 ;
        RECT 46.530 34.800 50.480 35.000 ;
        RECT 50.130 34.200 50.480 34.800 ;
        RECT 46.530 34.000 50.480 34.200 ;
        RECT 50.130 33.400 50.480 34.000 ;
        RECT 38.980 32.600 39.330 33.200 ;
        RECT 38.980 32.400 42.930 32.600 ;
        RECT 38.980 31.800 39.330 32.400 ;
        RECT 38.980 31.600 42.930 31.800 ;
        RECT 38.980 31.000 39.330 31.600 ;
        RECT 38.980 30.800 42.930 31.000 ;
        RECT 38.980 30.400 39.330 30.800 ;
        RECT 35.780 22.000 35.980 29.600 ;
        RECT 36.580 22.000 36.780 29.600 ;
        RECT 37.380 22.000 37.580 29.600 ;
        RECT 38.180 22.000 38.380 29.600 ;
        RECT 38.980 29.200 39.330 29.600 ;
        RECT 38.980 29.000 42.930 29.200 ;
        RECT 38.980 28.400 39.330 29.000 ;
        RECT 38.980 28.200 42.930 28.400 ;
        RECT 38.980 27.600 39.330 28.200 ;
        RECT 38.980 27.400 42.930 27.600 ;
        RECT 38.980 26.800 39.330 27.400 ;
        RECT 38.980 26.600 42.930 26.800 ;
        RECT 43.930 26.750 44.330 33.250 ;
        RECT 45.130 26.750 45.530 33.250 ;
        RECT 46.530 33.200 50.480 33.400 ;
        RECT 50.130 32.600 50.480 33.200 ;
        RECT 46.530 32.400 50.480 32.600 ;
        RECT 50.130 31.800 50.480 32.400 ;
        RECT 46.530 31.600 50.480 31.800 ;
        RECT 50.130 31.000 50.480 31.600 ;
        RECT 46.530 30.800 50.480 31.000 ;
        RECT 50.130 30.400 50.480 30.800 ;
        RECT 51.080 30.400 51.280 38.000 ;
        RECT 51.880 30.400 52.080 38.000 ;
        RECT 52.680 30.400 52.880 38.000 ;
        RECT 53.480 30.400 53.680 38.000 ;
        RECT 50.130 29.200 50.480 29.600 ;
        RECT 46.530 29.000 50.480 29.200 ;
        RECT 50.130 28.400 50.480 29.000 ;
        RECT 46.530 28.200 50.480 28.400 ;
        RECT 50.130 27.600 50.480 28.200 ;
        RECT 46.530 27.400 50.480 27.600 ;
        RECT 50.130 26.800 50.480 27.400 ;
        RECT 38.980 26.000 39.330 26.600 ;
        RECT 38.980 25.800 42.930 26.000 ;
        RECT 38.980 25.200 39.330 25.800 ;
        RECT 38.980 25.000 42.930 25.200 ;
        RECT 38.980 24.400 39.330 25.000 ;
        RECT 43.880 24.450 45.580 26.750 ;
        RECT 46.530 26.600 50.480 26.800 ;
        RECT 50.130 26.000 50.480 26.600 ;
        RECT 46.530 25.800 50.480 26.000 ;
        RECT 50.130 25.200 50.480 25.800 ;
        RECT 46.530 25.000 50.480 25.200 ;
        RECT 38.980 24.200 42.930 24.400 ;
        RECT 38.980 23.600 39.330 24.200 ;
        RECT 38.980 23.400 42.930 23.600 ;
        RECT 38.980 22.800 39.330 23.400 ;
        RECT 38.980 22.600 42.930 22.800 ;
        RECT 38.980 22.000 39.330 22.600 ;
        RECT 26.530 21.400 42.930 22.000 ;
        RECT 29.180 20.800 31.480 20.850 ;
        RECT 37.980 20.800 40.280 20.850 ;
        RECT 43.930 20.800 44.330 24.450 ;
        RECT 25.130 20.400 44.330 20.800 ;
        RECT 45.130 20.800 45.530 24.450 ;
        RECT 50.130 24.400 50.480 25.000 ;
        RECT 46.530 24.200 50.480 24.400 ;
        RECT 50.130 23.600 50.480 24.200 ;
        RECT 46.530 23.400 50.480 23.600 ;
        RECT 50.130 22.800 50.480 23.400 ;
        RECT 46.530 22.600 50.480 22.800 ;
        RECT 50.130 22.000 50.480 22.600 ;
        RECT 51.080 22.000 51.280 29.600 ;
        RECT 51.880 22.000 52.080 29.600 ;
        RECT 52.680 22.000 52.880 29.600 ;
        RECT 53.480 22.000 53.680 29.600 ;
        RECT 54.280 22.000 55.180 38.000 ;
        RECT 55.780 30.400 55.980 38.000 ;
        RECT 56.580 30.400 56.780 38.000 ;
        RECT 57.380 30.400 57.580 38.000 ;
        RECT 58.180 30.400 58.380 38.000 ;
        RECT 58.980 37.400 59.330 38.000 ;
        RECT 58.980 37.200 62.930 37.400 ;
        RECT 58.980 36.600 59.330 37.200 ;
        RECT 58.980 36.400 62.930 36.600 ;
        RECT 58.980 35.800 59.330 36.400 ;
        RECT 58.980 35.600 62.930 35.800 ;
        RECT 58.980 35.000 59.330 35.600 ;
        RECT 63.930 35.550 64.330 39.200 ;
        RECT 65.130 39.200 84.330 39.600 ;
        RECT 65.130 35.550 65.530 39.200 ;
        RECT 69.180 39.150 71.480 39.200 ;
        RECT 77.980 39.150 80.280 39.200 ;
        RECT 66.530 38.000 82.930 38.600 ;
        RECT 70.130 37.400 70.480 38.000 ;
        RECT 66.530 37.200 70.480 37.400 ;
        RECT 70.130 36.600 70.480 37.200 ;
        RECT 66.530 36.400 70.480 36.600 ;
        RECT 70.130 35.800 70.480 36.400 ;
        RECT 66.530 35.600 70.480 35.800 ;
        RECT 58.980 34.800 62.930 35.000 ;
        RECT 58.980 34.200 59.330 34.800 ;
        RECT 58.980 34.000 62.930 34.200 ;
        RECT 58.980 33.400 59.330 34.000 ;
        RECT 58.980 33.200 62.930 33.400 ;
        RECT 63.880 33.250 65.580 35.550 ;
        RECT 70.130 35.000 70.480 35.600 ;
        RECT 66.530 34.800 70.480 35.000 ;
        RECT 70.130 34.200 70.480 34.800 ;
        RECT 66.530 34.000 70.480 34.200 ;
        RECT 70.130 33.400 70.480 34.000 ;
        RECT 58.980 32.600 59.330 33.200 ;
        RECT 58.980 32.400 62.930 32.600 ;
        RECT 58.980 31.800 59.330 32.400 ;
        RECT 58.980 31.600 62.930 31.800 ;
        RECT 58.980 31.000 59.330 31.600 ;
        RECT 58.980 30.800 62.930 31.000 ;
        RECT 58.980 30.400 59.330 30.800 ;
        RECT 55.780 22.000 55.980 29.600 ;
        RECT 56.580 22.000 56.780 29.600 ;
        RECT 57.380 22.000 57.580 29.600 ;
        RECT 58.180 22.000 58.380 29.600 ;
        RECT 58.980 29.200 59.330 29.600 ;
        RECT 58.980 29.000 62.930 29.200 ;
        RECT 58.980 28.400 59.330 29.000 ;
        RECT 58.980 28.200 62.930 28.400 ;
        RECT 58.980 27.600 59.330 28.200 ;
        RECT 58.980 27.400 62.930 27.600 ;
        RECT 58.980 26.800 59.330 27.400 ;
        RECT 58.980 26.600 62.930 26.800 ;
        RECT 63.930 26.750 64.330 33.250 ;
        RECT 65.130 26.750 65.530 33.250 ;
        RECT 66.530 33.200 70.480 33.400 ;
        RECT 70.130 32.600 70.480 33.200 ;
        RECT 66.530 32.400 70.480 32.600 ;
        RECT 70.130 31.800 70.480 32.400 ;
        RECT 66.530 31.600 70.480 31.800 ;
        RECT 70.130 31.000 70.480 31.600 ;
        RECT 66.530 30.800 70.480 31.000 ;
        RECT 70.130 30.400 70.480 30.800 ;
        RECT 71.080 30.400 71.280 38.000 ;
        RECT 71.880 30.400 72.080 38.000 ;
        RECT 72.680 30.400 72.880 38.000 ;
        RECT 73.480 30.400 73.680 38.000 ;
        RECT 70.130 29.200 70.480 29.600 ;
        RECT 66.530 29.000 70.480 29.200 ;
        RECT 70.130 28.400 70.480 29.000 ;
        RECT 66.530 28.200 70.480 28.400 ;
        RECT 70.130 27.600 70.480 28.200 ;
        RECT 66.530 27.400 70.480 27.600 ;
        RECT 70.130 26.800 70.480 27.400 ;
        RECT 58.980 26.000 59.330 26.600 ;
        RECT 58.980 25.800 62.930 26.000 ;
        RECT 58.980 25.200 59.330 25.800 ;
        RECT 58.980 25.000 62.930 25.200 ;
        RECT 58.980 24.400 59.330 25.000 ;
        RECT 63.880 24.450 65.580 26.750 ;
        RECT 66.530 26.600 70.480 26.800 ;
        RECT 70.130 26.000 70.480 26.600 ;
        RECT 66.530 25.800 70.480 26.000 ;
        RECT 70.130 25.200 70.480 25.800 ;
        RECT 66.530 25.000 70.480 25.200 ;
        RECT 58.980 24.200 62.930 24.400 ;
        RECT 58.980 23.600 59.330 24.200 ;
        RECT 58.980 23.400 62.930 23.600 ;
        RECT 58.980 22.800 59.330 23.400 ;
        RECT 58.980 22.600 62.930 22.800 ;
        RECT 58.980 22.000 59.330 22.600 ;
        RECT 46.530 21.400 62.930 22.000 ;
        RECT 49.180 20.800 51.480 20.850 ;
        RECT 57.980 20.800 60.280 20.850 ;
        RECT 63.930 20.800 64.330 24.450 ;
        RECT 45.130 20.400 64.330 20.800 ;
        RECT 65.130 20.800 65.530 24.450 ;
        RECT 70.130 24.400 70.480 25.000 ;
        RECT 66.530 24.200 70.480 24.400 ;
        RECT 70.130 23.600 70.480 24.200 ;
        RECT 66.530 23.400 70.480 23.600 ;
        RECT 70.130 22.800 70.480 23.400 ;
        RECT 66.530 22.600 70.480 22.800 ;
        RECT 70.130 22.000 70.480 22.600 ;
        RECT 71.080 22.000 71.280 29.600 ;
        RECT 71.880 22.000 72.080 29.600 ;
        RECT 72.680 22.000 72.880 29.600 ;
        RECT 73.480 22.000 73.680 29.600 ;
        RECT 74.280 22.000 75.180 38.000 ;
        RECT 75.780 30.400 75.980 38.000 ;
        RECT 76.580 30.400 76.780 38.000 ;
        RECT 77.380 30.400 77.580 38.000 ;
        RECT 78.180 30.400 78.380 38.000 ;
        RECT 78.980 37.400 79.330 38.000 ;
        RECT 78.980 37.200 82.930 37.400 ;
        RECT 78.980 36.600 79.330 37.200 ;
        RECT 78.980 36.400 82.930 36.600 ;
        RECT 78.980 35.800 79.330 36.400 ;
        RECT 78.980 35.600 82.930 35.800 ;
        RECT 78.980 35.000 79.330 35.600 ;
        RECT 83.930 35.550 84.330 39.200 ;
        RECT 85.130 39.200 104.330 39.600 ;
        RECT 85.130 35.550 85.530 39.200 ;
        RECT 89.180 39.150 91.480 39.200 ;
        RECT 97.980 39.150 100.280 39.200 ;
        RECT 86.530 38.000 102.930 38.600 ;
        RECT 90.130 37.400 90.480 38.000 ;
        RECT 86.530 37.200 90.480 37.400 ;
        RECT 90.130 36.600 90.480 37.200 ;
        RECT 86.530 36.400 90.480 36.600 ;
        RECT 90.130 35.800 90.480 36.400 ;
        RECT 86.530 35.600 90.480 35.800 ;
        RECT 78.980 34.800 82.930 35.000 ;
        RECT 78.980 34.200 79.330 34.800 ;
        RECT 78.980 34.000 82.930 34.200 ;
        RECT 78.980 33.400 79.330 34.000 ;
        RECT 78.980 33.200 82.930 33.400 ;
        RECT 83.880 33.250 85.580 35.550 ;
        RECT 90.130 35.000 90.480 35.600 ;
        RECT 86.530 34.800 90.480 35.000 ;
        RECT 90.130 34.200 90.480 34.800 ;
        RECT 86.530 34.000 90.480 34.200 ;
        RECT 90.130 33.400 90.480 34.000 ;
        RECT 78.980 32.600 79.330 33.200 ;
        RECT 78.980 32.400 82.930 32.600 ;
        RECT 78.980 31.800 79.330 32.400 ;
        RECT 78.980 31.600 82.930 31.800 ;
        RECT 78.980 31.000 79.330 31.600 ;
        RECT 78.980 30.800 82.930 31.000 ;
        RECT 78.980 30.400 79.330 30.800 ;
        RECT 75.780 22.000 75.980 29.600 ;
        RECT 76.580 22.000 76.780 29.600 ;
        RECT 77.380 22.000 77.580 29.600 ;
        RECT 78.180 22.000 78.380 29.600 ;
        RECT 78.980 29.200 79.330 29.600 ;
        RECT 78.980 29.000 82.930 29.200 ;
        RECT 78.980 28.400 79.330 29.000 ;
        RECT 78.980 28.200 82.930 28.400 ;
        RECT 78.980 27.600 79.330 28.200 ;
        RECT 78.980 27.400 82.930 27.600 ;
        RECT 78.980 26.800 79.330 27.400 ;
        RECT 78.980 26.600 82.930 26.800 ;
        RECT 83.930 26.750 84.330 33.250 ;
        RECT 85.130 26.750 85.530 33.250 ;
        RECT 86.530 33.200 90.480 33.400 ;
        RECT 90.130 32.600 90.480 33.200 ;
        RECT 86.530 32.400 90.480 32.600 ;
        RECT 90.130 31.800 90.480 32.400 ;
        RECT 86.530 31.600 90.480 31.800 ;
        RECT 90.130 31.000 90.480 31.600 ;
        RECT 86.530 30.800 90.480 31.000 ;
        RECT 90.130 30.400 90.480 30.800 ;
        RECT 91.080 30.400 91.280 38.000 ;
        RECT 91.880 30.400 92.080 38.000 ;
        RECT 92.680 30.400 92.880 38.000 ;
        RECT 93.480 30.400 93.680 38.000 ;
        RECT 90.130 29.200 90.480 29.600 ;
        RECT 86.530 29.000 90.480 29.200 ;
        RECT 90.130 28.400 90.480 29.000 ;
        RECT 86.530 28.200 90.480 28.400 ;
        RECT 90.130 27.600 90.480 28.200 ;
        RECT 86.530 27.400 90.480 27.600 ;
        RECT 90.130 26.800 90.480 27.400 ;
        RECT 78.980 26.000 79.330 26.600 ;
        RECT 78.980 25.800 82.930 26.000 ;
        RECT 78.980 25.200 79.330 25.800 ;
        RECT 78.980 25.000 82.930 25.200 ;
        RECT 78.980 24.400 79.330 25.000 ;
        RECT 83.880 24.450 85.580 26.750 ;
        RECT 86.530 26.600 90.480 26.800 ;
        RECT 90.130 26.000 90.480 26.600 ;
        RECT 86.530 25.800 90.480 26.000 ;
        RECT 90.130 25.200 90.480 25.800 ;
        RECT 86.530 25.000 90.480 25.200 ;
        RECT 78.980 24.200 82.930 24.400 ;
        RECT 78.980 23.600 79.330 24.200 ;
        RECT 78.980 23.400 82.930 23.600 ;
        RECT 78.980 22.800 79.330 23.400 ;
        RECT 78.980 22.600 82.930 22.800 ;
        RECT 78.980 22.000 79.330 22.600 ;
        RECT 66.530 21.400 82.930 22.000 ;
        RECT 69.180 20.800 71.480 20.850 ;
        RECT 77.980 20.800 80.280 20.850 ;
        RECT 83.930 20.800 84.330 24.450 ;
        RECT 65.130 20.400 84.330 20.800 ;
        RECT 85.130 20.800 85.530 24.450 ;
        RECT 90.130 24.400 90.480 25.000 ;
        RECT 86.530 24.200 90.480 24.400 ;
        RECT 90.130 23.600 90.480 24.200 ;
        RECT 86.530 23.400 90.480 23.600 ;
        RECT 90.130 22.800 90.480 23.400 ;
        RECT 86.530 22.600 90.480 22.800 ;
        RECT 90.130 22.000 90.480 22.600 ;
        RECT 91.080 22.000 91.280 29.600 ;
        RECT 91.880 22.000 92.080 29.600 ;
        RECT 92.680 22.000 92.880 29.600 ;
        RECT 93.480 22.000 93.680 29.600 ;
        RECT 94.280 22.000 95.180 38.000 ;
        RECT 95.780 30.400 95.980 38.000 ;
        RECT 96.580 30.400 96.780 38.000 ;
        RECT 97.380 30.400 97.580 38.000 ;
        RECT 98.180 30.400 98.380 38.000 ;
        RECT 98.980 37.400 99.330 38.000 ;
        RECT 98.980 37.200 102.930 37.400 ;
        RECT 98.980 36.600 99.330 37.200 ;
        RECT 98.980 36.400 102.930 36.600 ;
        RECT 98.980 35.800 99.330 36.400 ;
        RECT 98.980 35.600 102.930 35.800 ;
        RECT 98.980 35.000 99.330 35.600 ;
        RECT 103.930 35.550 104.330 39.200 ;
        RECT 105.130 39.200 124.330 39.600 ;
        RECT 105.130 35.550 105.530 39.200 ;
        RECT 109.180 39.150 111.480 39.200 ;
        RECT 117.980 39.150 120.280 39.200 ;
        RECT 106.530 38.000 122.930 38.600 ;
        RECT 110.130 37.400 110.480 38.000 ;
        RECT 106.530 37.200 110.480 37.400 ;
        RECT 110.130 36.600 110.480 37.200 ;
        RECT 106.530 36.400 110.480 36.600 ;
        RECT 110.130 35.800 110.480 36.400 ;
        RECT 106.530 35.600 110.480 35.800 ;
        RECT 98.980 34.800 102.930 35.000 ;
        RECT 98.980 34.200 99.330 34.800 ;
        RECT 98.980 34.000 102.930 34.200 ;
        RECT 98.980 33.400 99.330 34.000 ;
        RECT 98.980 33.200 102.930 33.400 ;
        RECT 103.880 33.250 105.580 35.550 ;
        RECT 110.130 35.000 110.480 35.600 ;
        RECT 106.530 34.800 110.480 35.000 ;
        RECT 110.130 34.200 110.480 34.800 ;
        RECT 106.530 34.000 110.480 34.200 ;
        RECT 110.130 33.400 110.480 34.000 ;
        RECT 98.980 32.600 99.330 33.200 ;
        RECT 98.980 32.400 102.930 32.600 ;
        RECT 98.980 31.800 99.330 32.400 ;
        RECT 98.980 31.600 102.930 31.800 ;
        RECT 98.980 31.000 99.330 31.600 ;
        RECT 98.980 30.800 102.930 31.000 ;
        RECT 98.980 30.400 99.330 30.800 ;
        RECT 95.780 22.000 95.980 29.600 ;
        RECT 96.580 22.000 96.780 29.600 ;
        RECT 97.380 22.000 97.580 29.600 ;
        RECT 98.180 22.000 98.380 29.600 ;
        RECT 98.980 29.200 99.330 29.600 ;
        RECT 98.980 29.000 102.930 29.200 ;
        RECT 98.980 28.400 99.330 29.000 ;
        RECT 98.980 28.200 102.930 28.400 ;
        RECT 98.980 27.600 99.330 28.200 ;
        RECT 98.980 27.400 102.930 27.600 ;
        RECT 98.980 26.800 99.330 27.400 ;
        RECT 98.980 26.600 102.930 26.800 ;
        RECT 103.930 26.750 104.330 33.250 ;
        RECT 105.130 26.750 105.530 33.250 ;
        RECT 106.530 33.200 110.480 33.400 ;
        RECT 110.130 32.600 110.480 33.200 ;
        RECT 106.530 32.400 110.480 32.600 ;
        RECT 110.130 31.800 110.480 32.400 ;
        RECT 106.530 31.600 110.480 31.800 ;
        RECT 110.130 31.000 110.480 31.600 ;
        RECT 106.530 30.800 110.480 31.000 ;
        RECT 110.130 30.400 110.480 30.800 ;
        RECT 111.080 30.400 111.280 38.000 ;
        RECT 111.880 30.400 112.080 38.000 ;
        RECT 112.680 30.400 112.880 38.000 ;
        RECT 113.480 30.400 113.680 38.000 ;
        RECT 110.130 29.200 110.480 29.600 ;
        RECT 106.530 29.000 110.480 29.200 ;
        RECT 110.130 28.400 110.480 29.000 ;
        RECT 106.530 28.200 110.480 28.400 ;
        RECT 110.130 27.600 110.480 28.200 ;
        RECT 106.530 27.400 110.480 27.600 ;
        RECT 110.130 26.800 110.480 27.400 ;
        RECT 98.980 26.000 99.330 26.600 ;
        RECT 98.980 25.800 102.930 26.000 ;
        RECT 98.980 25.200 99.330 25.800 ;
        RECT 98.980 25.000 102.930 25.200 ;
        RECT 98.980 24.400 99.330 25.000 ;
        RECT 103.880 24.450 105.580 26.750 ;
        RECT 106.530 26.600 110.480 26.800 ;
        RECT 110.130 26.000 110.480 26.600 ;
        RECT 106.530 25.800 110.480 26.000 ;
        RECT 110.130 25.200 110.480 25.800 ;
        RECT 106.530 25.000 110.480 25.200 ;
        RECT 98.980 24.200 102.930 24.400 ;
        RECT 98.980 23.600 99.330 24.200 ;
        RECT 98.980 23.400 102.930 23.600 ;
        RECT 98.980 22.800 99.330 23.400 ;
        RECT 98.980 22.600 102.930 22.800 ;
        RECT 98.980 22.000 99.330 22.600 ;
        RECT 86.530 21.400 102.930 22.000 ;
        RECT 89.180 20.800 91.480 20.850 ;
        RECT 97.980 20.800 100.280 20.850 ;
        RECT 103.930 20.800 104.330 24.450 ;
        RECT 85.130 20.400 104.330 20.800 ;
        RECT 105.130 20.800 105.530 24.450 ;
        RECT 110.130 24.400 110.480 25.000 ;
        RECT 106.530 24.200 110.480 24.400 ;
        RECT 110.130 23.600 110.480 24.200 ;
        RECT 106.530 23.400 110.480 23.600 ;
        RECT 110.130 22.800 110.480 23.400 ;
        RECT 106.530 22.600 110.480 22.800 ;
        RECT 110.130 22.000 110.480 22.600 ;
        RECT 111.080 22.000 111.280 29.600 ;
        RECT 111.880 22.000 112.080 29.600 ;
        RECT 112.680 22.000 112.880 29.600 ;
        RECT 113.480 22.000 113.680 29.600 ;
        RECT 114.280 22.000 115.180 38.000 ;
        RECT 115.780 30.400 115.980 38.000 ;
        RECT 116.580 30.400 116.780 38.000 ;
        RECT 117.380 30.400 117.580 38.000 ;
        RECT 118.180 30.400 118.380 38.000 ;
        RECT 118.980 37.400 119.330 38.000 ;
        RECT 118.980 37.200 122.930 37.400 ;
        RECT 118.980 36.600 119.330 37.200 ;
        RECT 118.980 36.400 122.930 36.600 ;
        RECT 118.980 35.800 119.330 36.400 ;
        RECT 118.980 35.600 122.930 35.800 ;
        RECT 118.980 35.000 119.330 35.600 ;
        RECT 123.930 35.550 124.330 39.200 ;
        RECT 125.340 36.805 125.700 37.185 ;
        RECT 125.970 36.805 126.330 37.185 ;
        RECT 126.570 36.805 126.930 37.185 ;
        RECT 125.340 36.215 125.700 36.595 ;
        RECT 125.970 36.215 126.330 36.595 ;
        RECT 126.570 36.215 126.930 36.595 ;
        RECT 118.980 34.800 122.930 35.000 ;
        RECT 118.980 34.200 119.330 34.800 ;
        RECT 118.980 34.000 122.930 34.200 ;
        RECT 118.980 33.400 119.330 34.000 ;
        RECT 118.980 33.200 122.930 33.400 ;
        RECT 123.880 33.250 124.730 35.550 ;
        RECT 118.980 32.600 119.330 33.200 ;
        RECT 118.980 32.400 122.930 32.600 ;
        RECT 118.980 31.800 119.330 32.400 ;
        RECT 118.980 31.600 122.930 31.800 ;
        RECT 118.980 31.000 119.330 31.600 ;
        RECT 118.980 30.800 122.930 31.000 ;
        RECT 118.980 30.400 119.330 30.800 ;
        RECT 115.780 22.000 115.980 29.600 ;
        RECT 116.580 22.000 116.780 29.600 ;
        RECT 117.380 22.000 117.580 29.600 ;
        RECT 118.180 22.000 118.380 29.600 ;
        RECT 118.980 29.200 119.330 29.600 ;
        RECT 118.980 29.000 122.930 29.200 ;
        RECT 118.980 28.400 119.330 29.000 ;
        RECT 118.980 28.200 122.930 28.400 ;
        RECT 118.980 27.600 119.330 28.200 ;
        RECT 118.980 27.400 122.930 27.600 ;
        RECT 118.980 26.800 119.330 27.400 ;
        RECT 118.980 26.600 122.930 26.800 ;
        RECT 123.930 26.750 124.330 33.250 ;
        RECT 118.980 26.000 119.330 26.600 ;
        RECT 118.980 25.800 122.930 26.000 ;
        RECT 118.980 25.200 119.330 25.800 ;
        RECT 118.980 25.000 122.930 25.200 ;
        RECT 118.980 24.400 119.330 25.000 ;
        RECT 123.880 24.450 124.730 26.750 ;
        RECT 118.980 24.200 122.930 24.400 ;
        RECT 118.980 23.600 119.330 24.200 ;
        RECT 118.980 23.400 122.930 23.600 ;
        RECT 118.980 22.800 119.330 23.400 ;
        RECT 118.980 22.600 122.930 22.800 ;
        RECT 118.980 22.000 119.330 22.600 ;
        RECT 106.530 21.400 122.930 22.000 ;
        RECT 109.180 20.800 111.480 20.850 ;
        RECT 117.980 20.800 120.280 20.850 ;
        RECT 123.930 20.800 124.330 24.450 ;
        RECT 125.340 22.590 125.700 22.970 ;
        RECT 125.970 22.590 126.330 22.970 ;
        RECT 126.570 22.590 126.930 22.970 ;
        RECT 125.340 22.000 125.700 22.380 ;
        RECT 125.970 22.000 126.330 22.380 ;
        RECT 126.570 22.000 126.930 22.380 ;
        RECT 105.130 20.400 124.330 20.800 ;
        RECT 9.180 19.600 11.480 20.400 ;
        RECT 17.980 19.600 20.280 20.400 ;
        RECT 29.180 19.600 31.480 20.400 ;
        RECT 37.980 19.600 40.280 20.400 ;
        RECT 49.180 19.600 51.480 20.400 ;
        RECT 57.980 19.600 60.280 20.400 ;
        RECT 69.180 19.600 71.480 20.400 ;
        RECT 77.980 19.600 80.280 20.400 ;
        RECT 89.180 19.600 91.480 20.400 ;
        RECT 97.980 19.600 100.280 20.400 ;
        RECT 109.180 19.600 111.480 20.400 ;
        RECT 117.980 19.600 120.280 20.400 ;
        RECT 5.130 19.200 24.330 19.600 ;
        RECT 2.515 17.260 2.875 17.640 ;
        RECT 3.145 17.260 3.505 17.640 ;
        RECT 3.745 17.260 4.105 17.640 ;
        RECT 2.515 16.670 2.875 17.050 ;
        RECT 3.145 16.670 3.505 17.050 ;
        RECT 3.745 16.670 4.105 17.050 ;
        RECT 5.130 15.550 5.530 19.200 ;
        RECT 9.180 19.150 11.480 19.200 ;
        RECT 17.980 19.150 20.280 19.200 ;
        RECT 6.530 18.000 22.930 18.600 ;
        RECT 10.130 17.400 10.480 18.000 ;
        RECT 6.530 17.200 10.480 17.400 ;
        RECT 10.130 16.600 10.480 17.200 ;
        RECT 6.530 16.400 10.480 16.600 ;
        RECT 10.130 15.800 10.480 16.400 ;
        RECT 6.530 15.600 10.480 15.800 ;
        RECT 2.315 13.255 5.580 15.550 ;
        RECT 10.130 15.000 10.480 15.600 ;
        RECT 6.530 14.800 10.480 15.000 ;
        RECT 10.130 14.200 10.480 14.800 ;
        RECT 6.530 14.000 10.480 14.200 ;
        RECT 10.130 13.400 10.480 14.000 ;
        RECT 4.730 13.250 5.580 13.255 ;
        RECT 5.130 6.750 5.530 13.250 ;
        RECT 6.530 13.200 10.480 13.400 ;
        RECT 10.130 12.600 10.480 13.200 ;
        RECT 6.530 12.400 10.480 12.600 ;
        RECT 10.130 11.800 10.480 12.400 ;
        RECT 6.530 11.600 10.480 11.800 ;
        RECT 10.130 11.000 10.480 11.600 ;
        RECT 6.530 10.800 10.480 11.000 ;
        RECT 10.130 10.400 10.480 10.800 ;
        RECT 11.080 10.400 11.280 18.000 ;
        RECT 11.880 10.400 12.080 18.000 ;
        RECT 12.680 10.400 12.880 18.000 ;
        RECT 13.480 10.400 13.680 18.000 ;
        RECT 10.130 9.200 10.480 9.600 ;
        RECT 6.530 9.000 10.480 9.200 ;
        RECT 10.130 8.400 10.480 9.000 ;
        RECT 6.530 8.200 10.480 8.400 ;
        RECT 10.130 7.600 10.480 8.200 ;
        RECT 6.530 7.400 10.480 7.600 ;
        RECT 10.130 6.800 10.480 7.400 ;
        RECT 4.730 6.745 5.580 6.750 ;
        RECT 2.315 4.450 5.580 6.745 ;
        RECT 6.530 6.600 10.480 6.800 ;
        RECT 10.130 6.000 10.480 6.600 ;
        RECT 6.530 5.800 10.480 6.000 ;
        RECT 10.130 5.200 10.480 5.800 ;
        RECT 6.530 5.000 10.480 5.200 ;
        RECT 2.515 3.145 2.875 3.525 ;
        RECT 3.145 3.145 3.505 3.525 ;
        RECT 3.745 3.145 4.105 3.525 ;
        RECT 2.515 2.555 2.875 2.935 ;
        RECT 3.145 2.555 3.505 2.935 ;
        RECT 3.745 2.555 4.105 2.935 ;
        RECT 5.130 0.800 5.530 4.450 ;
        RECT 10.130 4.400 10.480 5.000 ;
        RECT 6.530 4.200 10.480 4.400 ;
        RECT 10.130 3.600 10.480 4.200 ;
        RECT 6.530 3.400 10.480 3.600 ;
        RECT 10.130 2.800 10.480 3.400 ;
        RECT 6.530 2.600 10.480 2.800 ;
        RECT 10.130 2.000 10.480 2.600 ;
        RECT 11.080 2.000 11.280 9.600 ;
        RECT 11.880 2.000 12.080 9.600 ;
        RECT 12.680 2.000 12.880 9.600 ;
        RECT 13.480 2.000 13.680 9.600 ;
        RECT 14.280 2.000 15.180 18.000 ;
        RECT 15.780 10.400 15.980 18.000 ;
        RECT 16.580 10.400 16.780 18.000 ;
        RECT 17.380 10.400 17.580 18.000 ;
        RECT 18.180 10.400 18.380 18.000 ;
        RECT 18.980 17.400 19.330 18.000 ;
        RECT 18.980 17.200 22.930 17.400 ;
        RECT 18.980 16.600 19.330 17.200 ;
        RECT 18.980 16.400 22.930 16.600 ;
        RECT 18.980 15.800 19.330 16.400 ;
        RECT 18.980 15.600 22.930 15.800 ;
        RECT 18.980 15.000 19.330 15.600 ;
        RECT 23.930 15.550 24.330 19.200 ;
        RECT 25.130 19.200 44.330 19.600 ;
        RECT 25.130 15.550 25.530 19.200 ;
        RECT 29.180 19.150 31.480 19.200 ;
        RECT 37.980 19.150 40.280 19.200 ;
        RECT 26.530 18.000 42.930 18.600 ;
        RECT 30.130 17.400 30.480 18.000 ;
        RECT 26.530 17.200 30.480 17.400 ;
        RECT 30.130 16.600 30.480 17.200 ;
        RECT 26.530 16.400 30.480 16.600 ;
        RECT 30.130 15.800 30.480 16.400 ;
        RECT 26.530 15.600 30.480 15.800 ;
        RECT 18.980 14.800 22.930 15.000 ;
        RECT 18.980 14.200 19.330 14.800 ;
        RECT 18.980 14.000 22.930 14.200 ;
        RECT 18.980 13.400 19.330 14.000 ;
        RECT 18.980 13.200 22.930 13.400 ;
        RECT 23.880 13.250 25.580 15.550 ;
        RECT 30.130 15.000 30.480 15.600 ;
        RECT 26.530 14.800 30.480 15.000 ;
        RECT 30.130 14.200 30.480 14.800 ;
        RECT 26.530 14.000 30.480 14.200 ;
        RECT 30.130 13.400 30.480 14.000 ;
        RECT 18.980 12.600 19.330 13.200 ;
        RECT 18.980 12.400 22.930 12.600 ;
        RECT 18.980 11.800 19.330 12.400 ;
        RECT 18.980 11.600 22.930 11.800 ;
        RECT 18.980 11.000 19.330 11.600 ;
        RECT 18.980 10.800 22.930 11.000 ;
        RECT 18.980 10.400 19.330 10.800 ;
        RECT 15.780 2.000 15.980 9.600 ;
        RECT 16.580 2.000 16.780 9.600 ;
        RECT 17.380 2.000 17.580 9.600 ;
        RECT 18.180 2.000 18.380 9.600 ;
        RECT 18.980 9.200 19.330 9.600 ;
        RECT 18.980 9.000 22.930 9.200 ;
        RECT 18.980 8.400 19.330 9.000 ;
        RECT 18.980 8.200 22.930 8.400 ;
        RECT 18.980 7.600 19.330 8.200 ;
        RECT 18.980 7.400 22.930 7.600 ;
        RECT 18.980 6.800 19.330 7.400 ;
        RECT 18.980 6.600 22.930 6.800 ;
        RECT 23.930 6.750 24.330 13.250 ;
        RECT 25.130 6.750 25.530 13.250 ;
        RECT 26.530 13.200 30.480 13.400 ;
        RECT 30.130 12.600 30.480 13.200 ;
        RECT 26.530 12.400 30.480 12.600 ;
        RECT 30.130 11.800 30.480 12.400 ;
        RECT 26.530 11.600 30.480 11.800 ;
        RECT 30.130 11.000 30.480 11.600 ;
        RECT 26.530 10.800 30.480 11.000 ;
        RECT 30.130 10.400 30.480 10.800 ;
        RECT 31.080 10.400 31.280 18.000 ;
        RECT 31.880 10.400 32.080 18.000 ;
        RECT 32.680 10.400 32.880 18.000 ;
        RECT 33.480 10.400 33.680 18.000 ;
        RECT 30.130 9.200 30.480 9.600 ;
        RECT 26.530 9.000 30.480 9.200 ;
        RECT 30.130 8.400 30.480 9.000 ;
        RECT 26.530 8.200 30.480 8.400 ;
        RECT 30.130 7.600 30.480 8.200 ;
        RECT 26.530 7.400 30.480 7.600 ;
        RECT 30.130 6.800 30.480 7.400 ;
        RECT 18.980 6.000 19.330 6.600 ;
        RECT 18.980 5.800 22.930 6.000 ;
        RECT 18.980 5.200 19.330 5.800 ;
        RECT 18.980 5.000 22.930 5.200 ;
        RECT 18.980 4.400 19.330 5.000 ;
        RECT 23.880 4.450 25.580 6.750 ;
        RECT 26.530 6.600 30.480 6.800 ;
        RECT 30.130 6.000 30.480 6.600 ;
        RECT 26.530 5.800 30.480 6.000 ;
        RECT 30.130 5.200 30.480 5.800 ;
        RECT 26.530 5.000 30.480 5.200 ;
        RECT 18.980 4.200 22.930 4.400 ;
        RECT 18.980 3.600 19.330 4.200 ;
        RECT 18.980 3.400 22.930 3.600 ;
        RECT 18.980 2.800 19.330 3.400 ;
        RECT 18.980 2.600 22.930 2.800 ;
        RECT 18.980 2.000 19.330 2.600 ;
        RECT 6.530 1.400 22.930 2.000 ;
        RECT 9.180 0.800 11.480 0.850 ;
        RECT 17.980 0.800 20.280 0.850 ;
        RECT 23.930 0.800 24.330 4.450 ;
        RECT 5.130 0.400 24.330 0.800 ;
        RECT 25.130 0.800 25.530 4.450 ;
        RECT 30.130 4.400 30.480 5.000 ;
        RECT 26.530 4.200 30.480 4.400 ;
        RECT 30.130 3.600 30.480 4.200 ;
        RECT 26.530 3.400 30.480 3.600 ;
        RECT 30.130 2.800 30.480 3.400 ;
        RECT 26.530 2.600 30.480 2.800 ;
        RECT 30.130 2.000 30.480 2.600 ;
        RECT 31.080 2.000 31.280 9.600 ;
        RECT 31.880 2.000 32.080 9.600 ;
        RECT 32.680 2.000 32.880 9.600 ;
        RECT 33.480 2.000 33.680 9.600 ;
        RECT 34.280 2.000 35.180 18.000 ;
        RECT 35.780 10.400 35.980 18.000 ;
        RECT 36.580 10.400 36.780 18.000 ;
        RECT 37.380 10.400 37.580 18.000 ;
        RECT 38.180 10.400 38.380 18.000 ;
        RECT 38.980 17.400 39.330 18.000 ;
        RECT 38.980 17.200 42.930 17.400 ;
        RECT 38.980 16.600 39.330 17.200 ;
        RECT 38.980 16.400 42.930 16.600 ;
        RECT 38.980 15.800 39.330 16.400 ;
        RECT 38.980 15.600 42.930 15.800 ;
        RECT 38.980 15.000 39.330 15.600 ;
        RECT 43.930 15.550 44.330 19.200 ;
        RECT 45.130 19.200 64.330 19.600 ;
        RECT 45.130 15.550 45.530 19.200 ;
        RECT 49.180 19.150 51.480 19.200 ;
        RECT 57.980 19.150 60.280 19.200 ;
        RECT 46.530 18.000 62.930 18.600 ;
        RECT 50.130 17.400 50.480 18.000 ;
        RECT 46.530 17.200 50.480 17.400 ;
        RECT 50.130 16.600 50.480 17.200 ;
        RECT 46.530 16.400 50.480 16.600 ;
        RECT 50.130 15.800 50.480 16.400 ;
        RECT 46.530 15.600 50.480 15.800 ;
        RECT 38.980 14.800 42.930 15.000 ;
        RECT 38.980 14.200 39.330 14.800 ;
        RECT 38.980 14.000 42.930 14.200 ;
        RECT 38.980 13.400 39.330 14.000 ;
        RECT 38.980 13.200 42.930 13.400 ;
        RECT 43.880 13.250 45.580 15.550 ;
        RECT 50.130 15.000 50.480 15.600 ;
        RECT 46.530 14.800 50.480 15.000 ;
        RECT 50.130 14.200 50.480 14.800 ;
        RECT 46.530 14.000 50.480 14.200 ;
        RECT 50.130 13.400 50.480 14.000 ;
        RECT 38.980 12.600 39.330 13.200 ;
        RECT 38.980 12.400 42.930 12.600 ;
        RECT 38.980 11.800 39.330 12.400 ;
        RECT 38.980 11.600 42.930 11.800 ;
        RECT 38.980 11.000 39.330 11.600 ;
        RECT 38.980 10.800 42.930 11.000 ;
        RECT 38.980 10.400 39.330 10.800 ;
        RECT 35.780 2.000 35.980 9.600 ;
        RECT 36.580 2.000 36.780 9.600 ;
        RECT 37.380 2.000 37.580 9.600 ;
        RECT 38.180 2.000 38.380 9.600 ;
        RECT 38.980 9.200 39.330 9.600 ;
        RECT 38.980 9.000 42.930 9.200 ;
        RECT 38.980 8.400 39.330 9.000 ;
        RECT 38.980 8.200 42.930 8.400 ;
        RECT 38.980 7.600 39.330 8.200 ;
        RECT 38.980 7.400 42.930 7.600 ;
        RECT 38.980 6.800 39.330 7.400 ;
        RECT 38.980 6.600 42.930 6.800 ;
        RECT 43.930 6.750 44.330 13.250 ;
        RECT 45.130 6.750 45.530 13.250 ;
        RECT 46.530 13.200 50.480 13.400 ;
        RECT 50.130 12.600 50.480 13.200 ;
        RECT 46.530 12.400 50.480 12.600 ;
        RECT 50.130 11.800 50.480 12.400 ;
        RECT 46.530 11.600 50.480 11.800 ;
        RECT 50.130 11.000 50.480 11.600 ;
        RECT 46.530 10.800 50.480 11.000 ;
        RECT 50.130 10.400 50.480 10.800 ;
        RECT 51.080 10.400 51.280 18.000 ;
        RECT 51.880 10.400 52.080 18.000 ;
        RECT 52.680 10.400 52.880 18.000 ;
        RECT 53.480 10.400 53.680 18.000 ;
        RECT 50.130 9.200 50.480 9.600 ;
        RECT 46.530 9.000 50.480 9.200 ;
        RECT 50.130 8.400 50.480 9.000 ;
        RECT 46.530 8.200 50.480 8.400 ;
        RECT 50.130 7.600 50.480 8.200 ;
        RECT 46.530 7.400 50.480 7.600 ;
        RECT 50.130 6.800 50.480 7.400 ;
        RECT 38.980 6.000 39.330 6.600 ;
        RECT 38.980 5.800 42.930 6.000 ;
        RECT 38.980 5.200 39.330 5.800 ;
        RECT 38.980 5.000 42.930 5.200 ;
        RECT 38.980 4.400 39.330 5.000 ;
        RECT 43.880 4.450 45.580 6.750 ;
        RECT 46.530 6.600 50.480 6.800 ;
        RECT 50.130 6.000 50.480 6.600 ;
        RECT 46.530 5.800 50.480 6.000 ;
        RECT 50.130 5.200 50.480 5.800 ;
        RECT 46.530 5.000 50.480 5.200 ;
        RECT 38.980 4.200 42.930 4.400 ;
        RECT 38.980 3.600 39.330 4.200 ;
        RECT 38.980 3.400 42.930 3.600 ;
        RECT 38.980 2.800 39.330 3.400 ;
        RECT 38.980 2.600 42.930 2.800 ;
        RECT 38.980 2.000 39.330 2.600 ;
        RECT 26.530 1.400 42.930 2.000 ;
        RECT 29.180 0.800 31.480 0.850 ;
        RECT 37.980 0.800 40.280 0.850 ;
        RECT 43.930 0.800 44.330 4.450 ;
        RECT 25.130 0.400 44.330 0.800 ;
        RECT 45.130 0.800 45.530 4.450 ;
        RECT 50.130 4.400 50.480 5.000 ;
        RECT 46.530 4.200 50.480 4.400 ;
        RECT 50.130 3.600 50.480 4.200 ;
        RECT 46.530 3.400 50.480 3.600 ;
        RECT 50.130 2.800 50.480 3.400 ;
        RECT 46.530 2.600 50.480 2.800 ;
        RECT 50.130 2.000 50.480 2.600 ;
        RECT 51.080 2.000 51.280 9.600 ;
        RECT 51.880 2.000 52.080 9.600 ;
        RECT 52.680 2.000 52.880 9.600 ;
        RECT 53.480 2.000 53.680 9.600 ;
        RECT 54.280 2.000 55.180 18.000 ;
        RECT 55.780 10.400 55.980 18.000 ;
        RECT 56.580 10.400 56.780 18.000 ;
        RECT 57.380 10.400 57.580 18.000 ;
        RECT 58.180 10.400 58.380 18.000 ;
        RECT 58.980 17.400 59.330 18.000 ;
        RECT 58.980 17.200 62.930 17.400 ;
        RECT 58.980 16.600 59.330 17.200 ;
        RECT 58.980 16.400 62.930 16.600 ;
        RECT 58.980 15.800 59.330 16.400 ;
        RECT 58.980 15.600 62.930 15.800 ;
        RECT 58.980 15.000 59.330 15.600 ;
        RECT 63.930 15.550 64.330 19.200 ;
        RECT 65.130 19.200 84.330 19.600 ;
        RECT 65.130 15.550 65.530 19.200 ;
        RECT 69.180 19.150 71.480 19.200 ;
        RECT 77.980 19.150 80.280 19.200 ;
        RECT 66.530 18.000 82.930 18.600 ;
        RECT 70.130 17.400 70.480 18.000 ;
        RECT 66.530 17.200 70.480 17.400 ;
        RECT 70.130 16.600 70.480 17.200 ;
        RECT 66.530 16.400 70.480 16.600 ;
        RECT 70.130 15.800 70.480 16.400 ;
        RECT 66.530 15.600 70.480 15.800 ;
        RECT 58.980 14.800 62.930 15.000 ;
        RECT 58.980 14.200 59.330 14.800 ;
        RECT 58.980 14.000 62.930 14.200 ;
        RECT 58.980 13.400 59.330 14.000 ;
        RECT 58.980 13.200 62.930 13.400 ;
        RECT 63.880 13.250 65.580 15.550 ;
        RECT 70.130 15.000 70.480 15.600 ;
        RECT 66.530 14.800 70.480 15.000 ;
        RECT 70.130 14.200 70.480 14.800 ;
        RECT 66.530 14.000 70.480 14.200 ;
        RECT 70.130 13.400 70.480 14.000 ;
        RECT 58.980 12.600 59.330 13.200 ;
        RECT 58.980 12.400 62.930 12.600 ;
        RECT 58.980 11.800 59.330 12.400 ;
        RECT 58.980 11.600 62.930 11.800 ;
        RECT 58.980 11.000 59.330 11.600 ;
        RECT 58.980 10.800 62.930 11.000 ;
        RECT 58.980 10.400 59.330 10.800 ;
        RECT 55.780 2.000 55.980 9.600 ;
        RECT 56.580 2.000 56.780 9.600 ;
        RECT 57.380 2.000 57.580 9.600 ;
        RECT 58.180 2.000 58.380 9.600 ;
        RECT 58.980 9.200 59.330 9.600 ;
        RECT 58.980 9.000 62.930 9.200 ;
        RECT 58.980 8.400 59.330 9.000 ;
        RECT 58.980 8.200 62.930 8.400 ;
        RECT 58.980 7.600 59.330 8.200 ;
        RECT 58.980 7.400 62.930 7.600 ;
        RECT 58.980 6.800 59.330 7.400 ;
        RECT 58.980 6.600 62.930 6.800 ;
        RECT 63.930 6.750 64.330 13.250 ;
        RECT 65.130 6.750 65.530 13.250 ;
        RECT 66.530 13.200 70.480 13.400 ;
        RECT 70.130 12.600 70.480 13.200 ;
        RECT 66.530 12.400 70.480 12.600 ;
        RECT 70.130 11.800 70.480 12.400 ;
        RECT 66.530 11.600 70.480 11.800 ;
        RECT 70.130 11.000 70.480 11.600 ;
        RECT 66.530 10.800 70.480 11.000 ;
        RECT 70.130 10.400 70.480 10.800 ;
        RECT 71.080 10.400 71.280 18.000 ;
        RECT 71.880 10.400 72.080 18.000 ;
        RECT 72.680 10.400 72.880 18.000 ;
        RECT 73.480 10.400 73.680 18.000 ;
        RECT 70.130 9.200 70.480 9.600 ;
        RECT 66.530 9.000 70.480 9.200 ;
        RECT 70.130 8.400 70.480 9.000 ;
        RECT 66.530 8.200 70.480 8.400 ;
        RECT 70.130 7.600 70.480 8.200 ;
        RECT 66.530 7.400 70.480 7.600 ;
        RECT 70.130 6.800 70.480 7.400 ;
        RECT 58.980 6.000 59.330 6.600 ;
        RECT 58.980 5.800 62.930 6.000 ;
        RECT 58.980 5.200 59.330 5.800 ;
        RECT 58.980 5.000 62.930 5.200 ;
        RECT 58.980 4.400 59.330 5.000 ;
        RECT 63.880 4.450 65.580 6.750 ;
        RECT 66.530 6.600 70.480 6.800 ;
        RECT 70.130 6.000 70.480 6.600 ;
        RECT 66.530 5.800 70.480 6.000 ;
        RECT 70.130 5.200 70.480 5.800 ;
        RECT 66.530 5.000 70.480 5.200 ;
        RECT 58.980 4.200 62.930 4.400 ;
        RECT 58.980 3.600 59.330 4.200 ;
        RECT 58.980 3.400 62.930 3.600 ;
        RECT 58.980 2.800 59.330 3.400 ;
        RECT 58.980 2.600 62.930 2.800 ;
        RECT 58.980 2.000 59.330 2.600 ;
        RECT 46.530 1.400 62.930 2.000 ;
        RECT 49.180 0.800 51.480 0.850 ;
        RECT 57.980 0.800 60.280 0.850 ;
        RECT 63.930 0.800 64.330 4.450 ;
        RECT 45.130 0.400 64.330 0.800 ;
        RECT 65.130 0.800 65.530 4.450 ;
        RECT 70.130 4.400 70.480 5.000 ;
        RECT 66.530 4.200 70.480 4.400 ;
        RECT 70.130 3.600 70.480 4.200 ;
        RECT 66.530 3.400 70.480 3.600 ;
        RECT 70.130 2.800 70.480 3.400 ;
        RECT 66.530 2.600 70.480 2.800 ;
        RECT 70.130 2.000 70.480 2.600 ;
        RECT 71.080 2.000 71.280 9.600 ;
        RECT 71.880 2.000 72.080 9.600 ;
        RECT 72.680 2.000 72.880 9.600 ;
        RECT 73.480 2.000 73.680 9.600 ;
        RECT 74.280 2.000 75.180 18.000 ;
        RECT 75.780 10.400 75.980 18.000 ;
        RECT 76.580 10.400 76.780 18.000 ;
        RECT 77.380 10.400 77.580 18.000 ;
        RECT 78.180 10.400 78.380 18.000 ;
        RECT 78.980 17.400 79.330 18.000 ;
        RECT 78.980 17.200 82.930 17.400 ;
        RECT 78.980 16.600 79.330 17.200 ;
        RECT 78.980 16.400 82.930 16.600 ;
        RECT 78.980 15.800 79.330 16.400 ;
        RECT 78.980 15.600 82.930 15.800 ;
        RECT 78.980 15.000 79.330 15.600 ;
        RECT 83.930 15.550 84.330 19.200 ;
        RECT 85.130 19.200 104.330 19.600 ;
        RECT 85.130 15.550 85.530 19.200 ;
        RECT 89.180 19.150 91.480 19.200 ;
        RECT 97.980 19.150 100.280 19.200 ;
        RECT 86.530 18.000 102.930 18.600 ;
        RECT 90.130 17.400 90.480 18.000 ;
        RECT 86.530 17.200 90.480 17.400 ;
        RECT 90.130 16.600 90.480 17.200 ;
        RECT 86.530 16.400 90.480 16.600 ;
        RECT 90.130 15.800 90.480 16.400 ;
        RECT 86.530 15.600 90.480 15.800 ;
        RECT 78.980 14.800 82.930 15.000 ;
        RECT 78.980 14.200 79.330 14.800 ;
        RECT 78.980 14.000 82.930 14.200 ;
        RECT 78.980 13.400 79.330 14.000 ;
        RECT 78.980 13.200 82.930 13.400 ;
        RECT 83.880 13.250 85.580 15.550 ;
        RECT 90.130 15.000 90.480 15.600 ;
        RECT 86.530 14.800 90.480 15.000 ;
        RECT 90.130 14.200 90.480 14.800 ;
        RECT 86.530 14.000 90.480 14.200 ;
        RECT 90.130 13.400 90.480 14.000 ;
        RECT 78.980 12.600 79.330 13.200 ;
        RECT 78.980 12.400 82.930 12.600 ;
        RECT 78.980 11.800 79.330 12.400 ;
        RECT 78.980 11.600 82.930 11.800 ;
        RECT 78.980 11.000 79.330 11.600 ;
        RECT 78.980 10.800 82.930 11.000 ;
        RECT 78.980 10.400 79.330 10.800 ;
        RECT 75.780 2.000 75.980 9.600 ;
        RECT 76.580 2.000 76.780 9.600 ;
        RECT 77.380 2.000 77.580 9.600 ;
        RECT 78.180 2.000 78.380 9.600 ;
        RECT 78.980 9.200 79.330 9.600 ;
        RECT 78.980 9.000 82.930 9.200 ;
        RECT 78.980 8.400 79.330 9.000 ;
        RECT 78.980 8.200 82.930 8.400 ;
        RECT 78.980 7.600 79.330 8.200 ;
        RECT 78.980 7.400 82.930 7.600 ;
        RECT 78.980 6.800 79.330 7.400 ;
        RECT 78.980 6.600 82.930 6.800 ;
        RECT 83.930 6.750 84.330 13.250 ;
        RECT 85.130 6.750 85.530 13.250 ;
        RECT 86.530 13.200 90.480 13.400 ;
        RECT 90.130 12.600 90.480 13.200 ;
        RECT 86.530 12.400 90.480 12.600 ;
        RECT 90.130 11.800 90.480 12.400 ;
        RECT 86.530 11.600 90.480 11.800 ;
        RECT 90.130 11.000 90.480 11.600 ;
        RECT 86.530 10.800 90.480 11.000 ;
        RECT 90.130 10.400 90.480 10.800 ;
        RECT 91.080 10.400 91.280 18.000 ;
        RECT 91.880 10.400 92.080 18.000 ;
        RECT 92.680 10.400 92.880 18.000 ;
        RECT 93.480 10.400 93.680 18.000 ;
        RECT 90.130 9.200 90.480 9.600 ;
        RECT 86.530 9.000 90.480 9.200 ;
        RECT 90.130 8.400 90.480 9.000 ;
        RECT 86.530 8.200 90.480 8.400 ;
        RECT 90.130 7.600 90.480 8.200 ;
        RECT 86.530 7.400 90.480 7.600 ;
        RECT 90.130 6.800 90.480 7.400 ;
        RECT 78.980 6.000 79.330 6.600 ;
        RECT 78.980 5.800 82.930 6.000 ;
        RECT 78.980 5.200 79.330 5.800 ;
        RECT 78.980 5.000 82.930 5.200 ;
        RECT 78.980 4.400 79.330 5.000 ;
        RECT 83.880 4.450 85.580 6.750 ;
        RECT 86.530 6.600 90.480 6.800 ;
        RECT 90.130 6.000 90.480 6.600 ;
        RECT 86.530 5.800 90.480 6.000 ;
        RECT 90.130 5.200 90.480 5.800 ;
        RECT 86.530 5.000 90.480 5.200 ;
        RECT 78.980 4.200 82.930 4.400 ;
        RECT 78.980 3.600 79.330 4.200 ;
        RECT 78.980 3.400 82.930 3.600 ;
        RECT 78.980 2.800 79.330 3.400 ;
        RECT 78.980 2.600 82.930 2.800 ;
        RECT 78.980 2.000 79.330 2.600 ;
        RECT 66.530 1.400 82.930 2.000 ;
        RECT 69.180 0.800 71.480 0.850 ;
        RECT 77.980 0.800 80.280 0.850 ;
        RECT 83.930 0.800 84.330 4.450 ;
        RECT 65.130 0.400 84.330 0.800 ;
        RECT 85.130 0.800 85.530 4.450 ;
        RECT 90.130 4.400 90.480 5.000 ;
        RECT 86.530 4.200 90.480 4.400 ;
        RECT 90.130 3.600 90.480 4.200 ;
        RECT 86.530 3.400 90.480 3.600 ;
        RECT 90.130 2.800 90.480 3.400 ;
        RECT 86.530 2.600 90.480 2.800 ;
        RECT 90.130 2.000 90.480 2.600 ;
        RECT 91.080 2.000 91.280 9.600 ;
        RECT 91.880 2.000 92.080 9.600 ;
        RECT 92.680 2.000 92.880 9.600 ;
        RECT 93.480 2.000 93.680 9.600 ;
        RECT 94.280 2.000 95.180 18.000 ;
        RECT 95.780 10.400 95.980 18.000 ;
        RECT 96.580 10.400 96.780 18.000 ;
        RECT 97.380 10.400 97.580 18.000 ;
        RECT 98.180 10.400 98.380 18.000 ;
        RECT 98.980 17.400 99.330 18.000 ;
        RECT 98.980 17.200 102.930 17.400 ;
        RECT 98.980 16.600 99.330 17.200 ;
        RECT 98.980 16.400 102.930 16.600 ;
        RECT 98.980 15.800 99.330 16.400 ;
        RECT 98.980 15.600 102.930 15.800 ;
        RECT 98.980 15.000 99.330 15.600 ;
        RECT 103.930 15.550 104.330 19.200 ;
        RECT 105.130 19.200 124.330 19.600 ;
        RECT 105.130 15.550 105.530 19.200 ;
        RECT 109.180 19.150 111.480 19.200 ;
        RECT 117.980 19.150 120.280 19.200 ;
        RECT 106.530 18.000 122.930 18.600 ;
        RECT 110.130 17.400 110.480 18.000 ;
        RECT 106.530 17.200 110.480 17.400 ;
        RECT 110.130 16.600 110.480 17.200 ;
        RECT 106.530 16.400 110.480 16.600 ;
        RECT 110.130 15.800 110.480 16.400 ;
        RECT 106.530 15.600 110.480 15.800 ;
        RECT 98.980 14.800 102.930 15.000 ;
        RECT 98.980 14.200 99.330 14.800 ;
        RECT 98.980 14.000 102.930 14.200 ;
        RECT 98.980 13.400 99.330 14.000 ;
        RECT 98.980 13.200 102.930 13.400 ;
        RECT 103.880 13.250 105.580 15.550 ;
        RECT 110.130 15.000 110.480 15.600 ;
        RECT 106.530 14.800 110.480 15.000 ;
        RECT 110.130 14.200 110.480 14.800 ;
        RECT 106.530 14.000 110.480 14.200 ;
        RECT 110.130 13.400 110.480 14.000 ;
        RECT 98.980 12.600 99.330 13.200 ;
        RECT 98.980 12.400 102.930 12.600 ;
        RECT 98.980 11.800 99.330 12.400 ;
        RECT 98.980 11.600 102.930 11.800 ;
        RECT 98.980 11.000 99.330 11.600 ;
        RECT 98.980 10.800 102.930 11.000 ;
        RECT 98.980 10.400 99.330 10.800 ;
        RECT 95.780 2.000 95.980 9.600 ;
        RECT 96.580 2.000 96.780 9.600 ;
        RECT 97.380 2.000 97.580 9.600 ;
        RECT 98.180 2.000 98.380 9.600 ;
        RECT 98.980 9.200 99.330 9.600 ;
        RECT 98.980 9.000 102.930 9.200 ;
        RECT 98.980 8.400 99.330 9.000 ;
        RECT 98.980 8.200 102.930 8.400 ;
        RECT 98.980 7.600 99.330 8.200 ;
        RECT 98.980 7.400 102.930 7.600 ;
        RECT 98.980 6.800 99.330 7.400 ;
        RECT 98.980 6.600 102.930 6.800 ;
        RECT 103.930 6.750 104.330 13.250 ;
        RECT 105.130 6.750 105.530 13.250 ;
        RECT 106.530 13.200 110.480 13.400 ;
        RECT 110.130 12.600 110.480 13.200 ;
        RECT 106.530 12.400 110.480 12.600 ;
        RECT 110.130 11.800 110.480 12.400 ;
        RECT 106.530 11.600 110.480 11.800 ;
        RECT 110.130 11.000 110.480 11.600 ;
        RECT 106.530 10.800 110.480 11.000 ;
        RECT 110.130 10.400 110.480 10.800 ;
        RECT 111.080 10.400 111.280 18.000 ;
        RECT 111.880 10.400 112.080 18.000 ;
        RECT 112.680 10.400 112.880 18.000 ;
        RECT 113.480 10.400 113.680 18.000 ;
        RECT 110.130 9.200 110.480 9.600 ;
        RECT 106.530 9.000 110.480 9.200 ;
        RECT 110.130 8.400 110.480 9.000 ;
        RECT 106.530 8.200 110.480 8.400 ;
        RECT 110.130 7.600 110.480 8.200 ;
        RECT 106.530 7.400 110.480 7.600 ;
        RECT 110.130 6.800 110.480 7.400 ;
        RECT 98.980 6.000 99.330 6.600 ;
        RECT 98.980 5.800 102.930 6.000 ;
        RECT 98.980 5.200 99.330 5.800 ;
        RECT 98.980 5.000 102.930 5.200 ;
        RECT 98.980 4.400 99.330 5.000 ;
        RECT 103.880 4.450 105.580 6.750 ;
        RECT 106.530 6.600 110.480 6.800 ;
        RECT 110.130 6.000 110.480 6.600 ;
        RECT 106.530 5.800 110.480 6.000 ;
        RECT 110.130 5.200 110.480 5.800 ;
        RECT 106.530 5.000 110.480 5.200 ;
        RECT 98.980 4.200 102.930 4.400 ;
        RECT 98.980 3.600 99.330 4.200 ;
        RECT 98.980 3.400 102.930 3.600 ;
        RECT 98.980 2.800 99.330 3.400 ;
        RECT 98.980 2.600 102.930 2.800 ;
        RECT 98.980 2.000 99.330 2.600 ;
        RECT 86.530 1.400 102.930 2.000 ;
        RECT 89.180 0.800 91.480 0.850 ;
        RECT 97.980 0.800 100.280 0.850 ;
        RECT 103.930 0.800 104.330 4.450 ;
        RECT 85.130 0.400 104.330 0.800 ;
        RECT 105.130 0.800 105.530 4.450 ;
        RECT 110.130 4.400 110.480 5.000 ;
        RECT 106.530 4.200 110.480 4.400 ;
        RECT 110.130 3.600 110.480 4.200 ;
        RECT 106.530 3.400 110.480 3.600 ;
        RECT 110.130 2.800 110.480 3.400 ;
        RECT 106.530 2.600 110.480 2.800 ;
        RECT 110.130 2.000 110.480 2.600 ;
        RECT 111.080 2.000 111.280 9.600 ;
        RECT 111.880 2.000 112.080 9.600 ;
        RECT 112.680 2.000 112.880 9.600 ;
        RECT 113.480 2.000 113.680 9.600 ;
        RECT 114.280 2.000 115.180 18.000 ;
        RECT 115.780 10.400 115.980 18.000 ;
        RECT 116.580 10.400 116.780 18.000 ;
        RECT 117.380 10.400 117.580 18.000 ;
        RECT 118.180 10.400 118.380 18.000 ;
        RECT 118.980 17.400 119.330 18.000 ;
        RECT 118.980 17.200 122.930 17.400 ;
        RECT 118.980 16.600 119.330 17.200 ;
        RECT 118.980 16.400 122.930 16.600 ;
        RECT 118.980 15.800 119.330 16.400 ;
        RECT 118.980 15.600 122.930 15.800 ;
        RECT 118.980 15.000 119.330 15.600 ;
        RECT 123.930 15.550 124.330 19.200 ;
        RECT 125.340 16.805 125.700 17.185 ;
        RECT 125.970 16.805 126.330 17.185 ;
        RECT 126.570 16.805 126.930 17.185 ;
        RECT 125.340 16.215 125.700 16.595 ;
        RECT 125.970 16.215 126.330 16.595 ;
        RECT 126.570 16.215 126.930 16.595 ;
        RECT 118.980 14.800 122.930 15.000 ;
        RECT 118.980 14.200 119.330 14.800 ;
        RECT 118.980 14.000 122.930 14.200 ;
        RECT 118.980 13.400 119.330 14.000 ;
        RECT 118.980 13.200 122.930 13.400 ;
        RECT 123.880 13.250 124.730 15.550 ;
        RECT 118.980 12.600 119.330 13.200 ;
        RECT 118.980 12.400 122.930 12.600 ;
        RECT 118.980 11.800 119.330 12.400 ;
        RECT 118.980 11.600 122.930 11.800 ;
        RECT 118.980 11.000 119.330 11.600 ;
        RECT 118.980 10.800 122.930 11.000 ;
        RECT 118.980 10.400 119.330 10.800 ;
        RECT 115.780 2.000 115.980 9.600 ;
        RECT 116.580 2.000 116.780 9.600 ;
        RECT 117.380 2.000 117.580 9.600 ;
        RECT 118.180 2.000 118.380 9.600 ;
        RECT 118.980 9.200 119.330 9.600 ;
        RECT 118.980 9.000 122.930 9.200 ;
        RECT 118.980 8.400 119.330 9.000 ;
        RECT 118.980 8.200 122.930 8.400 ;
        RECT 118.980 7.600 119.330 8.200 ;
        RECT 118.980 7.400 122.930 7.600 ;
        RECT 118.980 6.800 119.330 7.400 ;
        RECT 118.980 6.600 122.930 6.800 ;
        RECT 123.930 6.750 124.330 13.250 ;
        RECT 118.980 6.000 119.330 6.600 ;
        RECT 118.980 5.800 122.930 6.000 ;
        RECT 118.980 5.200 119.330 5.800 ;
        RECT 118.980 5.000 122.930 5.200 ;
        RECT 118.980 4.400 119.330 5.000 ;
        RECT 123.880 4.450 124.730 6.750 ;
        RECT 118.980 4.200 122.930 4.400 ;
        RECT 118.980 3.600 119.330 4.200 ;
        RECT 118.980 3.400 122.930 3.600 ;
        RECT 118.980 2.800 119.330 3.400 ;
        RECT 118.980 2.600 122.930 2.800 ;
        RECT 118.980 2.000 119.330 2.600 ;
        RECT 106.530 1.400 122.930 2.000 ;
        RECT 109.180 0.800 111.480 0.850 ;
        RECT 117.980 0.800 120.280 0.850 ;
        RECT 123.930 0.800 124.330 4.450 ;
        RECT 125.340 2.590 125.700 2.970 ;
        RECT 125.970 2.590 126.330 2.970 ;
        RECT 126.570 2.590 126.930 2.970 ;
        RECT 125.340 2.000 125.700 2.380 ;
        RECT 125.970 2.000 126.330 2.380 ;
        RECT 126.570 2.000 126.930 2.380 ;
        RECT 105.130 0.400 124.330 0.800 ;
        RECT 9.180 0.000 11.480 0.400 ;
        RECT 17.980 0.000 20.280 0.400 ;
        RECT 29.180 0.000 31.480 0.400 ;
        RECT 37.980 0.000 40.280 0.400 ;
        RECT 49.180 0.000 51.480 0.400 ;
        RECT 57.980 0.000 60.280 0.400 ;
        RECT 69.180 0.000 71.480 0.400 ;
        RECT 77.980 0.000 80.280 0.400 ;
        RECT 89.180 0.000 91.480 0.400 ;
        RECT 97.980 0.000 100.280 0.400 ;
        RECT 109.180 0.000 111.480 0.400 ;
        RECT 117.980 0.000 120.280 0.400 ;
      LAYER mcon ;
        RECT 6.830 338.100 7.430 338.600 ;
        RECT 7.630 338.100 8.230 338.600 ;
        RECT 8.430 338.100 9.030 338.600 ;
        RECT 9.230 338.100 9.830 338.600 ;
        RECT 10.030 338.100 10.630 338.600 ;
        RECT 18.830 338.100 19.430 338.600 ;
        RECT 19.630 338.100 20.230 338.600 ;
        RECT 20.430 338.100 21.030 338.600 ;
        RECT 21.230 338.100 21.830 338.600 ;
        RECT 22.030 338.100 22.580 338.600 ;
        RECT 2.520 334.920 2.880 335.300 ;
        RECT 3.130 334.920 3.490 335.300 ;
        RECT 3.760 334.920 4.120 335.300 ;
        RECT 2.520 334.185 2.880 334.565 ;
        RECT 3.130 334.185 3.490 334.565 ;
        RECT 3.760 334.185 4.120 334.565 ;
        RECT 2.520 333.500 2.880 333.880 ;
        RECT 3.130 333.500 3.490 333.880 ;
        RECT 3.760 333.500 4.120 333.880 ;
        RECT 2.520 326.120 2.880 326.500 ;
        RECT 3.130 326.120 3.490 326.500 ;
        RECT 3.760 326.120 4.120 326.500 ;
        RECT 2.520 325.385 2.880 325.765 ;
        RECT 3.130 325.385 3.490 325.765 ;
        RECT 3.760 325.385 4.120 325.765 ;
        RECT 2.520 324.700 2.880 325.080 ;
        RECT 3.130 324.700 3.490 325.080 ;
        RECT 3.760 324.700 4.120 325.080 ;
        RECT 26.830 338.100 27.430 338.600 ;
        RECT 27.630 338.100 28.230 338.600 ;
        RECT 28.430 338.100 29.030 338.600 ;
        RECT 29.230 338.100 29.830 338.600 ;
        RECT 30.030 338.100 30.630 338.600 ;
        RECT 38.830 338.100 39.430 338.600 ;
        RECT 39.630 338.100 40.230 338.600 ;
        RECT 40.430 338.100 41.030 338.600 ;
        RECT 41.230 338.100 41.830 338.600 ;
        RECT 42.030 338.100 42.580 338.600 ;
        RECT 6.830 321.400 7.430 321.900 ;
        RECT 7.630 321.400 8.230 321.900 ;
        RECT 8.430 321.400 9.030 321.900 ;
        RECT 9.230 321.400 9.830 321.900 ;
        RECT 10.030 321.400 10.630 321.900 ;
        RECT 18.830 321.400 19.430 321.900 ;
        RECT 19.630 321.400 20.230 321.900 ;
        RECT 20.430 321.400 21.030 321.900 ;
        RECT 21.230 321.400 21.830 321.900 ;
        RECT 22.030 321.400 22.580 321.900 ;
        RECT 46.830 338.100 47.430 338.600 ;
        RECT 47.630 338.100 48.230 338.600 ;
        RECT 48.430 338.100 49.030 338.600 ;
        RECT 49.230 338.100 49.830 338.600 ;
        RECT 50.030 338.100 50.630 338.600 ;
        RECT 58.830 338.100 59.430 338.600 ;
        RECT 59.630 338.100 60.230 338.600 ;
        RECT 60.430 338.100 61.030 338.600 ;
        RECT 61.230 338.100 61.830 338.600 ;
        RECT 62.030 338.100 62.580 338.600 ;
        RECT 26.830 321.400 27.430 321.900 ;
        RECT 27.630 321.400 28.230 321.900 ;
        RECT 28.430 321.400 29.030 321.900 ;
        RECT 29.230 321.400 29.830 321.900 ;
        RECT 30.030 321.400 30.630 321.900 ;
        RECT 38.830 321.400 39.430 321.900 ;
        RECT 39.630 321.400 40.230 321.900 ;
        RECT 40.430 321.400 41.030 321.900 ;
        RECT 41.230 321.400 41.830 321.900 ;
        RECT 42.030 321.400 42.580 321.900 ;
        RECT 66.830 338.100 67.430 338.600 ;
        RECT 67.630 338.100 68.230 338.600 ;
        RECT 68.430 338.100 69.030 338.600 ;
        RECT 69.230 338.100 69.830 338.600 ;
        RECT 70.030 338.100 70.630 338.600 ;
        RECT 78.830 338.100 79.430 338.600 ;
        RECT 79.630 338.100 80.230 338.600 ;
        RECT 80.430 338.100 81.030 338.600 ;
        RECT 81.230 338.100 81.830 338.600 ;
        RECT 82.030 338.100 82.580 338.600 ;
        RECT 46.830 321.400 47.430 321.900 ;
        RECT 47.630 321.400 48.230 321.900 ;
        RECT 48.430 321.400 49.030 321.900 ;
        RECT 49.230 321.400 49.830 321.900 ;
        RECT 50.030 321.400 50.630 321.900 ;
        RECT 58.830 321.400 59.430 321.900 ;
        RECT 59.630 321.400 60.230 321.900 ;
        RECT 60.430 321.400 61.030 321.900 ;
        RECT 61.230 321.400 61.830 321.900 ;
        RECT 62.030 321.400 62.580 321.900 ;
        RECT 86.830 338.100 87.430 338.600 ;
        RECT 87.630 338.100 88.230 338.600 ;
        RECT 88.430 338.100 89.030 338.600 ;
        RECT 89.230 338.100 89.830 338.600 ;
        RECT 90.030 338.100 90.630 338.600 ;
        RECT 98.830 338.100 99.430 338.600 ;
        RECT 99.630 338.100 100.230 338.600 ;
        RECT 100.430 338.100 101.030 338.600 ;
        RECT 101.230 338.100 101.830 338.600 ;
        RECT 102.030 338.100 102.580 338.600 ;
        RECT 66.830 321.400 67.430 321.900 ;
        RECT 67.630 321.400 68.230 321.900 ;
        RECT 68.430 321.400 69.030 321.900 ;
        RECT 69.230 321.400 69.830 321.900 ;
        RECT 70.030 321.400 70.630 321.900 ;
        RECT 78.830 321.400 79.430 321.900 ;
        RECT 79.630 321.400 80.230 321.900 ;
        RECT 80.430 321.400 81.030 321.900 ;
        RECT 81.230 321.400 81.830 321.900 ;
        RECT 82.030 321.400 82.580 321.900 ;
        RECT 106.830 338.100 107.430 338.600 ;
        RECT 107.630 338.100 108.230 338.600 ;
        RECT 108.430 338.100 109.030 338.600 ;
        RECT 109.230 338.100 109.830 338.600 ;
        RECT 110.030 338.100 110.630 338.600 ;
        RECT 118.830 338.100 119.430 338.600 ;
        RECT 119.630 338.100 120.230 338.600 ;
        RECT 120.430 338.100 121.030 338.600 ;
        RECT 121.230 338.100 121.830 338.600 ;
        RECT 122.030 338.100 122.580 338.600 ;
        RECT 86.830 321.400 87.430 321.900 ;
        RECT 87.630 321.400 88.230 321.900 ;
        RECT 88.430 321.400 89.030 321.900 ;
        RECT 89.230 321.400 89.830 321.900 ;
        RECT 90.030 321.400 90.630 321.900 ;
        RECT 98.830 321.400 99.430 321.900 ;
        RECT 99.630 321.400 100.230 321.900 ;
        RECT 100.430 321.400 101.030 321.900 ;
        RECT 101.230 321.400 101.830 321.900 ;
        RECT 102.030 321.400 102.580 321.900 ;
        RECT 106.830 321.400 107.430 321.900 ;
        RECT 107.630 321.400 108.230 321.900 ;
        RECT 108.430 321.400 109.030 321.900 ;
        RECT 109.230 321.400 109.830 321.900 ;
        RECT 110.030 321.400 110.630 321.900 ;
        RECT 118.830 321.400 119.430 321.900 ;
        RECT 119.630 321.400 120.230 321.900 ;
        RECT 120.430 321.400 121.030 321.900 ;
        RECT 121.230 321.400 121.830 321.900 ;
        RECT 122.030 321.400 122.580 321.900 ;
        RECT 6.830 318.100 7.430 318.600 ;
        RECT 7.630 318.100 8.230 318.600 ;
        RECT 8.430 318.100 9.030 318.600 ;
        RECT 9.230 318.100 9.830 318.600 ;
        RECT 10.030 318.100 10.630 318.600 ;
        RECT 18.830 318.100 19.430 318.600 ;
        RECT 19.630 318.100 20.230 318.600 ;
        RECT 20.430 318.100 21.030 318.600 ;
        RECT 21.230 318.100 21.830 318.600 ;
        RECT 22.030 318.100 22.580 318.600 ;
        RECT 2.520 314.920 2.880 315.300 ;
        RECT 3.130 314.920 3.490 315.300 ;
        RECT 3.760 314.920 4.120 315.300 ;
        RECT 2.520 314.185 2.880 314.565 ;
        RECT 3.130 314.185 3.490 314.565 ;
        RECT 3.760 314.185 4.120 314.565 ;
        RECT 2.520 313.500 2.880 313.880 ;
        RECT 3.130 313.500 3.490 313.880 ;
        RECT 3.760 313.500 4.120 313.880 ;
        RECT 2.520 306.125 2.880 306.505 ;
        RECT 3.130 306.125 3.490 306.505 ;
        RECT 3.760 306.125 4.120 306.505 ;
        RECT 2.520 305.390 2.880 305.770 ;
        RECT 3.130 305.390 3.490 305.770 ;
        RECT 3.760 305.390 4.120 305.770 ;
        RECT 2.520 304.705 2.880 305.085 ;
        RECT 3.130 304.705 3.490 305.085 ;
        RECT 3.760 304.705 4.120 305.085 ;
        RECT 26.830 318.100 27.430 318.600 ;
        RECT 27.630 318.100 28.230 318.600 ;
        RECT 28.430 318.100 29.030 318.600 ;
        RECT 29.230 318.100 29.830 318.600 ;
        RECT 30.030 318.100 30.630 318.600 ;
        RECT 38.830 318.100 39.430 318.600 ;
        RECT 39.630 318.100 40.230 318.600 ;
        RECT 40.430 318.100 41.030 318.600 ;
        RECT 41.230 318.100 41.830 318.600 ;
        RECT 42.030 318.100 42.580 318.600 ;
        RECT 6.830 301.400 7.430 301.900 ;
        RECT 7.630 301.400 8.230 301.900 ;
        RECT 8.430 301.400 9.030 301.900 ;
        RECT 9.230 301.400 9.830 301.900 ;
        RECT 10.030 301.400 10.630 301.900 ;
        RECT 18.830 301.400 19.430 301.900 ;
        RECT 19.630 301.400 20.230 301.900 ;
        RECT 20.430 301.400 21.030 301.900 ;
        RECT 21.230 301.400 21.830 301.900 ;
        RECT 22.030 301.400 22.580 301.900 ;
        RECT 46.830 318.100 47.430 318.600 ;
        RECT 47.630 318.100 48.230 318.600 ;
        RECT 48.430 318.100 49.030 318.600 ;
        RECT 49.230 318.100 49.830 318.600 ;
        RECT 50.030 318.100 50.630 318.600 ;
        RECT 58.830 318.100 59.430 318.600 ;
        RECT 59.630 318.100 60.230 318.600 ;
        RECT 60.430 318.100 61.030 318.600 ;
        RECT 61.230 318.100 61.830 318.600 ;
        RECT 62.030 318.100 62.580 318.600 ;
        RECT 26.830 301.400 27.430 301.900 ;
        RECT 27.630 301.400 28.230 301.900 ;
        RECT 28.430 301.400 29.030 301.900 ;
        RECT 29.230 301.400 29.830 301.900 ;
        RECT 30.030 301.400 30.630 301.900 ;
        RECT 38.830 301.400 39.430 301.900 ;
        RECT 39.630 301.400 40.230 301.900 ;
        RECT 40.430 301.400 41.030 301.900 ;
        RECT 41.230 301.400 41.830 301.900 ;
        RECT 42.030 301.400 42.580 301.900 ;
        RECT 66.830 318.100 67.430 318.600 ;
        RECT 67.630 318.100 68.230 318.600 ;
        RECT 68.430 318.100 69.030 318.600 ;
        RECT 69.230 318.100 69.830 318.600 ;
        RECT 70.030 318.100 70.630 318.600 ;
        RECT 78.830 318.100 79.430 318.600 ;
        RECT 79.630 318.100 80.230 318.600 ;
        RECT 80.430 318.100 81.030 318.600 ;
        RECT 81.230 318.100 81.830 318.600 ;
        RECT 82.030 318.100 82.580 318.600 ;
        RECT 46.830 301.400 47.430 301.900 ;
        RECT 47.630 301.400 48.230 301.900 ;
        RECT 48.430 301.400 49.030 301.900 ;
        RECT 49.230 301.400 49.830 301.900 ;
        RECT 50.030 301.400 50.630 301.900 ;
        RECT 58.830 301.400 59.430 301.900 ;
        RECT 59.630 301.400 60.230 301.900 ;
        RECT 60.430 301.400 61.030 301.900 ;
        RECT 61.230 301.400 61.830 301.900 ;
        RECT 62.030 301.400 62.580 301.900 ;
        RECT 86.830 318.100 87.430 318.600 ;
        RECT 87.630 318.100 88.230 318.600 ;
        RECT 88.430 318.100 89.030 318.600 ;
        RECT 89.230 318.100 89.830 318.600 ;
        RECT 90.030 318.100 90.630 318.600 ;
        RECT 98.830 318.100 99.430 318.600 ;
        RECT 99.630 318.100 100.230 318.600 ;
        RECT 100.430 318.100 101.030 318.600 ;
        RECT 101.230 318.100 101.830 318.600 ;
        RECT 102.030 318.100 102.580 318.600 ;
        RECT 66.830 301.400 67.430 301.900 ;
        RECT 67.630 301.400 68.230 301.900 ;
        RECT 68.430 301.400 69.030 301.900 ;
        RECT 69.230 301.400 69.830 301.900 ;
        RECT 70.030 301.400 70.630 301.900 ;
        RECT 78.830 301.400 79.430 301.900 ;
        RECT 79.630 301.400 80.230 301.900 ;
        RECT 80.430 301.400 81.030 301.900 ;
        RECT 81.230 301.400 81.830 301.900 ;
        RECT 82.030 301.400 82.580 301.900 ;
        RECT 106.830 318.100 107.430 318.600 ;
        RECT 107.630 318.100 108.230 318.600 ;
        RECT 108.430 318.100 109.030 318.600 ;
        RECT 109.230 318.100 109.830 318.600 ;
        RECT 110.030 318.100 110.630 318.600 ;
        RECT 118.830 318.100 119.430 318.600 ;
        RECT 119.630 318.100 120.230 318.600 ;
        RECT 120.430 318.100 121.030 318.600 ;
        RECT 121.230 318.100 121.830 318.600 ;
        RECT 122.030 318.100 122.580 318.600 ;
        RECT 86.830 301.400 87.430 301.900 ;
        RECT 87.630 301.400 88.230 301.900 ;
        RECT 88.430 301.400 89.030 301.900 ;
        RECT 89.230 301.400 89.830 301.900 ;
        RECT 90.030 301.400 90.630 301.900 ;
        RECT 98.830 301.400 99.430 301.900 ;
        RECT 99.630 301.400 100.230 301.900 ;
        RECT 100.430 301.400 101.030 301.900 ;
        RECT 101.230 301.400 101.830 301.900 ;
        RECT 102.030 301.400 102.580 301.900 ;
        RECT 106.830 301.400 107.430 301.900 ;
        RECT 107.630 301.400 108.230 301.900 ;
        RECT 108.430 301.400 109.030 301.900 ;
        RECT 109.230 301.400 109.830 301.900 ;
        RECT 110.030 301.400 110.630 301.900 ;
        RECT 118.830 301.400 119.430 301.900 ;
        RECT 119.630 301.400 120.230 301.900 ;
        RECT 120.430 301.400 121.030 301.900 ;
        RECT 121.230 301.400 121.830 301.900 ;
        RECT 122.030 301.400 122.580 301.900 ;
        RECT 6.830 298.100 7.430 298.600 ;
        RECT 7.630 298.100 8.230 298.600 ;
        RECT 8.430 298.100 9.030 298.600 ;
        RECT 9.230 298.100 9.830 298.600 ;
        RECT 10.030 298.100 10.630 298.600 ;
        RECT 18.830 298.100 19.430 298.600 ;
        RECT 19.630 298.100 20.230 298.600 ;
        RECT 20.430 298.100 21.030 298.600 ;
        RECT 21.230 298.100 21.830 298.600 ;
        RECT 22.030 298.100 22.580 298.600 ;
        RECT 2.520 294.920 2.880 295.300 ;
        RECT 3.130 294.920 3.490 295.300 ;
        RECT 3.760 294.920 4.120 295.300 ;
        RECT 2.520 294.185 2.880 294.565 ;
        RECT 3.130 294.185 3.490 294.565 ;
        RECT 3.760 294.185 4.120 294.565 ;
        RECT 2.520 293.500 2.880 293.880 ;
        RECT 3.130 293.500 3.490 293.880 ;
        RECT 3.760 293.500 4.120 293.880 ;
        RECT 2.520 286.125 2.880 286.505 ;
        RECT 3.130 286.125 3.490 286.505 ;
        RECT 3.760 286.125 4.120 286.505 ;
        RECT 2.520 285.390 2.880 285.770 ;
        RECT 3.130 285.390 3.490 285.770 ;
        RECT 3.760 285.390 4.120 285.770 ;
        RECT 2.520 284.705 2.880 285.085 ;
        RECT 3.130 284.705 3.490 285.085 ;
        RECT 3.760 284.705 4.120 285.085 ;
        RECT 26.830 298.100 27.430 298.600 ;
        RECT 27.630 298.100 28.230 298.600 ;
        RECT 28.430 298.100 29.030 298.600 ;
        RECT 29.230 298.100 29.830 298.600 ;
        RECT 30.030 298.100 30.630 298.600 ;
        RECT 38.830 298.100 39.430 298.600 ;
        RECT 39.630 298.100 40.230 298.600 ;
        RECT 40.430 298.100 41.030 298.600 ;
        RECT 41.230 298.100 41.830 298.600 ;
        RECT 42.030 298.100 42.580 298.600 ;
        RECT 6.830 281.400 7.430 281.900 ;
        RECT 7.630 281.400 8.230 281.900 ;
        RECT 8.430 281.400 9.030 281.900 ;
        RECT 9.230 281.400 9.830 281.900 ;
        RECT 10.030 281.400 10.630 281.900 ;
        RECT 18.830 281.400 19.430 281.900 ;
        RECT 19.630 281.400 20.230 281.900 ;
        RECT 20.430 281.400 21.030 281.900 ;
        RECT 21.230 281.400 21.830 281.900 ;
        RECT 22.030 281.400 22.580 281.900 ;
        RECT 46.830 298.100 47.430 298.600 ;
        RECT 47.630 298.100 48.230 298.600 ;
        RECT 48.430 298.100 49.030 298.600 ;
        RECT 49.230 298.100 49.830 298.600 ;
        RECT 50.030 298.100 50.630 298.600 ;
        RECT 58.830 298.100 59.430 298.600 ;
        RECT 59.630 298.100 60.230 298.600 ;
        RECT 60.430 298.100 61.030 298.600 ;
        RECT 61.230 298.100 61.830 298.600 ;
        RECT 62.030 298.100 62.580 298.600 ;
        RECT 26.830 281.400 27.430 281.900 ;
        RECT 27.630 281.400 28.230 281.900 ;
        RECT 28.430 281.400 29.030 281.900 ;
        RECT 29.230 281.400 29.830 281.900 ;
        RECT 30.030 281.400 30.630 281.900 ;
        RECT 38.830 281.400 39.430 281.900 ;
        RECT 39.630 281.400 40.230 281.900 ;
        RECT 40.430 281.400 41.030 281.900 ;
        RECT 41.230 281.400 41.830 281.900 ;
        RECT 42.030 281.400 42.580 281.900 ;
        RECT 66.830 298.100 67.430 298.600 ;
        RECT 67.630 298.100 68.230 298.600 ;
        RECT 68.430 298.100 69.030 298.600 ;
        RECT 69.230 298.100 69.830 298.600 ;
        RECT 70.030 298.100 70.630 298.600 ;
        RECT 78.830 298.100 79.430 298.600 ;
        RECT 79.630 298.100 80.230 298.600 ;
        RECT 80.430 298.100 81.030 298.600 ;
        RECT 81.230 298.100 81.830 298.600 ;
        RECT 82.030 298.100 82.580 298.600 ;
        RECT 46.830 281.400 47.430 281.900 ;
        RECT 47.630 281.400 48.230 281.900 ;
        RECT 48.430 281.400 49.030 281.900 ;
        RECT 49.230 281.400 49.830 281.900 ;
        RECT 50.030 281.400 50.630 281.900 ;
        RECT 58.830 281.400 59.430 281.900 ;
        RECT 59.630 281.400 60.230 281.900 ;
        RECT 60.430 281.400 61.030 281.900 ;
        RECT 61.230 281.400 61.830 281.900 ;
        RECT 62.030 281.400 62.580 281.900 ;
        RECT 86.830 298.100 87.430 298.600 ;
        RECT 87.630 298.100 88.230 298.600 ;
        RECT 88.430 298.100 89.030 298.600 ;
        RECT 89.230 298.100 89.830 298.600 ;
        RECT 90.030 298.100 90.630 298.600 ;
        RECT 98.830 298.100 99.430 298.600 ;
        RECT 99.630 298.100 100.230 298.600 ;
        RECT 100.430 298.100 101.030 298.600 ;
        RECT 101.230 298.100 101.830 298.600 ;
        RECT 102.030 298.100 102.580 298.600 ;
        RECT 66.830 281.400 67.430 281.900 ;
        RECT 67.630 281.400 68.230 281.900 ;
        RECT 68.430 281.400 69.030 281.900 ;
        RECT 69.230 281.400 69.830 281.900 ;
        RECT 70.030 281.400 70.630 281.900 ;
        RECT 78.830 281.400 79.430 281.900 ;
        RECT 79.630 281.400 80.230 281.900 ;
        RECT 80.430 281.400 81.030 281.900 ;
        RECT 81.230 281.400 81.830 281.900 ;
        RECT 82.030 281.400 82.580 281.900 ;
        RECT 106.830 298.100 107.430 298.600 ;
        RECT 107.630 298.100 108.230 298.600 ;
        RECT 108.430 298.100 109.030 298.600 ;
        RECT 109.230 298.100 109.830 298.600 ;
        RECT 110.030 298.100 110.630 298.600 ;
        RECT 118.830 298.100 119.430 298.600 ;
        RECT 119.630 298.100 120.230 298.600 ;
        RECT 120.430 298.100 121.030 298.600 ;
        RECT 121.230 298.100 121.830 298.600 ;
        RECT 122.030 298.100 122.580 298.600 ;
        RECT 86.830 281.400 87.430 281.900 ;
        RECT 87.630 281.400 88.230 281.900 ;
        RECT 88.430 281.400 89.030 281.900 ;
        RECT 89.230 281.400 89.830 281.900 ;
        RECT 90.030 281.400 90.630 281.900 ;
        RECT 98.830 281.400 99.430 281.900 ;
        RECT 99.630 281.400 100.230 281.900 ;
        RECT 100.430 281.400 101.030 281.900 ;
        RECT 101.230 281.400 101.830 281.900 ;
        RECT 102.030 281.400 102.580 281.900 ;
        RECT 106.830 281.400 107.430 281.900 ;
        RECT 107.630 281.400 108.230 281.900 ;
        RECT 108.430 281.400 109.030 281.900 ;
        RECT 109.230 281.400 109.830 281.900 ;
        RECT 110.030 281.400 110.630 281.900 ;
        RECT 118.830 281.400 119.430 281.900 ;
        RECT 119.630 281.400 120.230 281.900 ;
        RECT 120.430 281.400 121.030 281.900 ;
        RECT 121.230 281.400 121.830 281.900 ;
        RECT 122.030 281.400 122.580 281.900 ;
        RECT 6.830 278.100 7.430 278.600 ;
        RECT 7.630 278.100 8.230 278.600 ;
        RECT 8.430 278.100 9.030 278.600 ;
        RECT 9.230 278.100 9.830 278.600 ;
        RECT 10.030 278.100 10.630 278.600 ;
        RECT 18.830 278.100 19.430 278.600 ;
        RECT 19.630 278.100 20.230 278.600 ;
        RECT 20.430 278.100 21.030 278.600 ;
        RECT 21.230 278.100 21.830 278.600 ;
        RECT 22.030 278.100 22.580 278.600 ;
        RECT 2.520 274.920 2.880 275.300 ;
        RECT 3.130 274.920 3.490 275.300 ;
        RECT 3.760 274.920 4.120 275.300 ;
        RECT 2.520 274.185 2.880 274.565 ;
        RECT 3.130 274.185 3.490 274.565 ;
        RECT 3.760 274.185 4.120 274.565 ;
        RECT 2.520 273.500 2.880 273.880 ;
        RECT 3.130 273.500 3.490 273.880 ;
        RECT 3.760 273.500 4.120 273.880 ;
        RECT 2.520 266.115 2.880 266.495 ;
        RECT 3.130 266.115 3.490 266.495 ;
        RECT 3.760 266.115 4.120 266.495 ;
        RECT 2.520 265.380 2.880 265.760 ;
        RECT 3.130 265.380 3.490 265.760 ;
        RECT 3.760 265.380 4.120 265.760 ;
        RECT 2.520 264.695 2.880 265.075 ;
        RECT 3.130 264.695 3.490 265.075 ;
        RECT 3.760 264.695 4.120 265.075 ;
        RECT 26.830 278.100 27.430 278.600 ;
        RECT 27.630 278.100 28.230 278.600 ;
        RECT 28.430 278.100 29.030 278.600 ;
        RECT 29.230 278.100 29.830 278.600 ;
        RECT 30.030 278.100 30.630 278.600 ;
        RECT 38.830 278.100 39.430 278.600 ;
        RECT 39.630 278.100 40.230 278.600 ;
        RECT 40.430 278.100 41.030 278.600 ;
        RECT 41.230 278.100 41.830 278.600 ;
        RECT 42.030 278.100 42.580 278.600 ;
        RECT 6.830 261.400 7.430 261.900 ;
        RECT 7.630 261.400 8.230 261.900 ;
        RECT 8.430 261.400 9.030 261.900 ;
        RECT 9.230 261.400 9.830 261.900 ;
        RECT 10.030 261.400 10.630 261.900 ;
        RECT 18.830 261.400 19.430 261.900 ;
        RECT 19.630 261.400 20.230 261.900 ;
        RECT 20.430 261.400 21.030 261.900 ;
        RECT 21.230 261.400 21.830 261.900 ;
        RECT 22.030 261.400 22.580 261.900 ;
        RECT 46.830 278.100 47.430 278.600 ;
        RECT 47.630 278.100 48.230 278.600 ;
        RECT 48.430 278.100 49.030 278.600 ;
        RECT 49.230 278.100 49.830 278.600 ;
        RECT 50.030 278.100 50.630 278.600 ;
        RECT 58.830 278.100 59.430 278.600 ;
        RECT 59.630 278.100 60.230 278.600 ;
        RECT 60.430 278.100 61.030 278.600 ;
        RECT 61.230 278.100 61.830 278.600 ;
        RECT 62.030 278.100 62.580 278.600 ;
        RECT 26.830 261.400 27.430 261.900 ;
        RECT 27.630 261.400 28.230 261.900 ;
        RECT 28.430 261.400 29.030 261.900 ;
        RECT 29.230 261.400 29.830 261.900 ;
        RECT 30.030 261.400 30.630 261.900 ;
        RECT 38.830 261.400 39.430 261.900 ;
        RECT 39.630 261.400 40.230 261.900 ;
        RECT 40.430 261.400 41.030 261.900 ;
        RECT 41.230 261.400 41.830 261.900 ;
        RECT 42.030 261.400 42.580 261.900 ;
        RECT 66.830 278.100 67.430 278.600 ;
        RECT 67.630 278.100 68.230 278.600 ;
        RECT 68.430 278.100 69.030 278.600 ;
        RECT 69.230 278.100 69.830 278.600 ;
        RECT 70.030 278.100 70.630 278.600 ;
        RECT 78.830 278.100 79.430 278.600 ;
        RECT 79.630 278.100 80.230 278.600 ;
        RECT 80.430 278.100 81.030 278.600 ;
        RECT 81.230 278.100 81.830 278.600 ;
        RECT 82.030 278.100 82.580 278.600 ;
        RECT 46.830 261.400 47.430 261.900 ;
        RECT 47.630 261.400 48.230 261.900 ;
        RECT 48.430 261.400 49.030 261.900 ;
        RECT 49.230 261.400 49.830 261.900 ;
        RECT 50.030 261.400 50.630 261.900 ;
        RECT 58.830 261.400 59.430 261.900 ;
        RECT 59.630 261.400 60.230 261.900 ;
        RECT 60.430 261.400 61.030 261.900 ;
        RECT 61.230 261.400 61.830 261.900 ;
        RECT 62.030 261.400 62.580 261.900 ;
        RECT 86.830 278.100 87.430 278.600 ;
        RECT 87.630 278.100 88.230 278.600 ;
        RECT 88.430 278.100 89.030 278.600 ;
        RECT 89.230 278.100 89.830 278.600 ;
        RECT 90.030 278.100 90.630 278.600 ;
        RECT 98.830 278.100 99.430 278.600 ;
        RECT 99.630 278.100 100.230 278.600 ;
        RECT 100.430 278.100 101.030 278.600 ;
        RECT 101.230 278.100 101.830 278.600 ;
        RECT 102.030 278.100 102.580 278.600 ;
        RECT 66.830 261.400 67.430 261.900 ;
        RECT 67.630 261.400 68.230 261.900 ;
        RECT 68.430 261.400 69.030 261.900 ;
        RECT 69.230 261.400 69.830 261.900 ;
        RECT 70.030 261.400 70.630 261.900 ;
        RECT 78.830 261.400 79.430 261.900 ;
        RECT 79.630 261.400 80.230 261.900 ;
        RECT 80.430 261.400 81.030 261.900 ;
        RECT 81.230 261.400 81.830 261.900 ;
        RECT 82.030 261.400 82.580 261.900 ;
        RECT 106.830 278.100 107.430 278.600 ;
        RECT 107.630 278.100 108.230 278.600 ;
        RECT 108.430 278.100 109.030 278.600 ;
        RECT 109.230 278.100 109.830 278.600 ;
        RECT 110.030 278.100 110.630 278.600 ;
        RECT 118.830 278.100 119.430 278.600 ;
        RECT 119.630 278.100 120.230 278.600 ;
        RECT 120.430 278.100 121.030 278.600 ;
        RECT 121.230 278.100 121.830 278.600 ;
        RECT 122.030 278.100 122.580 278.600 ;
        RECT 86.830 261.400 87.430 261.900 ;
        RECT 87.630 261.400 88.230 261.900 ;
        RECT 88.430 261.400 89.030 261.900 ;
        RECT 89.230 261.400 89.830 261.900 ;
        RECT 90.030 261.400 90.630 261.900 ;
        RECT 98.830 261.400 99.430 261.900 ;
        RECT 99.630 261.400 100.230 261.900 ;
        RECT 100.430 261.400 101.030 261.900 ;
        RECT 101.230 261.400 101.830 261.900 ;
        RECT 102.030 261.400 102.580 261.900 ;
        RECT 106.830 261.400 107.430 261.900 ;
        RECT 107.630 261.400 108.230 261.900 ;
        RECT 108.430 261.400 109.030 261.900 ;
        RECT 109.230 261.400 109.830 261.900 ;
        RECT 110.030 261.400 110.630 261.900 ;
        RECT 118.830 261.400 119.430 261.900 ;
        RECT 119.630 261.400 120.230 261.900 ;
        RECT 120.430 261.400 121.030 261.900 ;
        RECT 121.230 261.400 121.830 261.900 ;
        RECT 122.030 261.400 122.580 261.900 ;
        RECT 6.830 258.100 7.430 258.600 ;
        RECT 7.630 258.100 8.230 258.600 ;
        RECT 8.430 258.100 9.030 258.600 ;
        RECT 9.230 258.100 9.830 258.600 ;
        RECT 10.030 258.100 10.630 258.600 ;
        RECT 18.830 258.100 19.430 258.600 ;
        RECT 19.630 258.100 20.230 258.600 ;
        RECT 20.430 258.100 21.030 258.600 ;
        RECT 21.230 258.100 21.830 258.600 ;
        RECT 22.030 258.100 22.580 258.600 ;
        RECT 2.520 254.920 2.880 255.300 ;
        RECT 3.130 254.920 3.490 255.300 ;
        RECT 3.760 254.920 4.120 255.300 ;
        RECT 2.520 254.185 2.880 254.565 ;
        RECT 3.130 254.185 3.490 254.565 ;
        RECT 3.760 254.185 4.120 254.565 ;
        RECT 2.520 253.500 2.880 253.880 ;
        RECT 3.130 253.500 3.490 253.880 ;
        RECT 3.760 253.500 4.120 253.880 ;
        RECT 2.520 246.125 2.880 246.505 ;
        RECT 3.130 246.125 3.490 246.505 ;
        RECT 3.760 246.125 4.120 246.505 ;
        RECT 2.520 245.390 2.880 245.770 ;
        RECT 3.130 245.390 3.490 245.770 ;
        RECT 3.760 245.390 4.120 245.770 ;
        RECT 2.520 244.705 2.880 245.085 ;
        RECT 3.130 244.705 3.490 245.085 ;
        RECT 3.760 244.705 4.120 245.085 ;
        RECT 26.830 258.100 27.430 258.600 ;
        RECT 27.630 258.100 28.230 258.600 ;
        RECT 28.430 258.100 29.030 258.600 ;
        RECT 29.230 258.100 29.830 258.600 ;
        RECT 30.030 258.100 30.630 258.600 ;
        RECT 38.830 258.100 39.430 258.600 ;
        RECT 39.630 258.100 40.230 258.600 ;
        RECT 40.430 258.100 41.030 258.600 ;
        RECT 41.230 258.100 41.830 258.600 ;
        RECT 42.030 258.100 42.580 258.600 ;
        RECT 6.830 241.400 7.430 241.900 ;
        RECT 7.630 241.400 8.230 241.900 ;
        RECT 8.430 241.400 9.030 241.900 ;
        RECT 9.230 241.400 9.830 241.900 ;
        RECT 10.030 241.400 10.630 241.900 ;
        RECT 18.830 241.400 19.430 241.900 ;
        RECT 19.630 241.400 20.230 241.900 ;
        RECT 20.430 241.400 21.030 241.900 ;
        RECT 21.230 241.400 21.830 241.900 ;
        RECT 22.030 241.400 22.580 241.900 ;
        RECT 46.830 258.100 47.430 258.600 ;
        RECT 47.630 258.100 48.230 258.600 ;
        RECT 48.430 258.100 49.030 258.600 ;
        RECT 49.230 258.100 49.830 258.600 ;
        RECT 50.030 258.100 50.630 258.600 ;
        RECT 58.830 258.100 59.430 258.600 ;
        RECT 59.630 258.100 60.230 258.600 ;
        RECT 60.430 258.100 61.030 258.600 ;
        RECT 61.230 258.100 61.830 258.600 ;
        RECT 62.030 258.100 62.580 258.600 ;
        RECT 26.830 241.400 27.430 241.900 ;
        RECT 27.630 241.400 28.230 241.900 ;
        RECT 28.430 241.400 29.030 241.900 ;
        RECT 29.230 241.400 29.830 241.900 ;
        RECT 30.030 241.400 30.630 241.900 ;
        RECT 38.830 241.400 39.430 241.900 ;
        RECT 39.630 241.400 40.230 241.900 ;
        RECT 40.430 241.400 41.030 241.900 ;
        RECT 41.230 241.400 41.830 241.900 ;
        RECT 42.030 241.400 42.580 241.900 ;
        RECT 66.830 258.100 67.430 258.600 ;
        RECT 67.630 258.100 68.230 258.600 ;
        RECT 68.430 258.100 69.030 258.600 ;
        RECT 69.230 258.100 69.830 258.600 ;
        RECT 70.030 258.100 70.630 258.600 ;
        RECT 78.830 258.100 79.430 258.600 ;
        RECT 79.630 258.100 80.230 258.600 ;
        RECT 80.430 258.100 81.030 258.600 ;
        RECT 81.230 258.100 81.830 258.600 ;
        RECT 82.030 258.100 82.580 258.600 ;
        RECT 46.830 241.400 47.430 241.900 ;
        RECT 47.630 241.400 48.230 241.900 ;
        RECT 48.430 241.400 49.030 241.900 ;
        RECT 49.230 241.400 49.830 241.900 ;
        RECT 50.030 241.400 50.630 241.900 ;
        RECT 58.830 241.400 59.430 241.900 ;
        RECT 59.630 241.400 60.230 241.900 ;
        RECT 60.430 241.400 61.030 241.900 ;
        RECT 61.230 241.400 61.830 241.900 ;
        RECT 62.030 241.400 62.580 241.900 ;
        RECT 86.830 258.100 87.430 258.600 ;
        RECT 87.630 258.100 88.230 258.600 ;
        RECT 88.430 258.100 89.030 258.600 ;
        RECT 89.230 258.100 89.830 258.600 ;
        RECT 90.030 258.100 90.630 258.600 ;
        RECT 98.830 258.100 99.430 258.600 ;
        RECT 99.630 258.100 100.230 258.600 ;
        RECT 100.430 258.100 101.030 258.600 ;
        RECT 101.230 258.100 101.830 258.600 ;
        RECT 102.030 258.100 102.580 258.600 ;
        RECT 66.830 241.400 67.430 241.900 ;
        RECT 67.630 241.400 68.230 241.900 ;
        RECT 68.430 241.400 69.030 241.900 ;
        RECT 69.230 241.400 69.830 241.900 ;
        RECT 70.030 241.400 70.630 241.900 ;
        RECT 78.830 241.400 79.430 241.900 ;
        RECT 79.630 241.400 80.230 241.900 ;
        RECT 80.430 241.400 81.030 241.900 ;
        RECT 81.230 241.400 81.830 241.900 ;
        RECT 82.030 241.400 82.580 241.900 ;
        RECT 106.830 258.100 107.430 258.600 ;
        RECT 107.630 258.100 108.230 258.600 ;
        RECT 108.430 258.100 109.030 258.600 ;
        RECT 109.230 258.100 109.830 258.600 ;
        RECT 110.030 258.100 110.630 258.600 ;
        RECT 118.830 258.100 119.430 258.600 ;
        RECT 119.630 258.100 120.230 258.600 ;
        RECT 120.430 258.100 121.030 258.600 ;
        RECT 121.230 258.100 121.830 258.600 ;
        RECT 122.030 258.100 122.580 258.600 ;
        RECT 86.830 241.400 87.430 241.900 ;
        RECT 87.630 241.400 88.230 241.900 ;
        RECT 88.430 241.400 89.030 241.900 ;
        RECT 89.230 241.400 89.830 241.900 ;
        RECT 90.030 241.400 90.630 241.900 ;
        RECT 98.830 241.400 99.430 241.900 ;
        RECT 99.630 241.400 100.230 241.900 ;
        RECT 100.430 241.400 101.030 241.900 ;
        RECT 101.230 241.400 101.830 241.900 ;
        RECT 102.030 241.400 102.580 241.900 ;
        RECT 106.830 241.400 107.430 241.900 ;
        RECT 107.630 241.400 108.230 241.900 ;
        RECT 108.430 241.400 109.030 241.900 ;
        RECT 109.230 241.400 109.830 241.900 ;
        RECT 110.030 241.400 110.630 241.900 ;
        RECT 118.830 241.400 119.430 241.900 ;
        RECT 119.630 241.400 120.230 241.900 ;
        RECT 120.430 241.400 121.030 241.900 ;
        RECT 121.230 241.400 121.830 241.900 ;
        RECT 122.030 241.400 122.580 241.900 ;
        RECT 6.830 238.100 7.430 238.600 ;
        RECT 7.630 238.100 8.230 238.600 ;
        RECT 8.430 238.100 9.030 238.600 ;
        RECT 9.230 238.100 9.830 238.600 ;
        RECT 10.030 238.100 10.630 238.600 ;
        RECT 18.830 238.100 19.430 238.600 ;
        RECT 19.630 238.100 20.230 238.600 ;
        RECT 20.430 238.100 21.030 238.600 ;
        RECT 21.230 238.100 21.830 238.600 ;
        RECT 22.030 238.100 22.580 238.600 ;
        RECT 2.520 234.920 2.880 235.300 ;
        RECT 3.130 234.920 3.490 235.300 ;
        RECT 3.760 234.920 4.120 235.300 ;
        RECT 2.520 234.185 2.880 234.565 ;
        RECT 3.130 234.185 3.490 234.565 ;
        RECT 3.760 234.185 4.120 234.565 ;
        RECT 2.520 233.500 2.880 233.880 ;
        RECT 3.130 233.500 3.490 233.880 ;
        RECT 3.760 233.500 4.120 233.880 ;
        RECT 2.520 226.125 2.880 226.505 ;
        RECT 3.130 226.125 3.490 226.505 ;
        RECT 3.760 226.125 4.120 226.505 ;
        RECT 2.520 225.390 2.880 225.770 ;
        RECT 3.130 225.390 3.490 225.770 ;
        RECT 3.760 225.390 4.120 225.770 ;
        RECT 2.520 224.705 2.880 225.085 ;
        RECT 3.130 224.705 3.490 225.085 ;
        RECT 3.760 224.705 4.120 225.085 ;
        RECT 26.830 238.100 27.430 238.600 ;
        RECT 27.630 238.100 28.230 238.600 ;
        RECT 28.430 238.100 29.030 238.600 ;
        RECT 29.230 238.100 29.830 238.600 ;
        RECT 30.030 238.100 30.630 238.600 ;
        RECT 38.830 238.100 39.430 238.600 ;
        RECT 39.630 238.100 40.230 238.600 ;
        RECT 40.430 238.100 41.030 238.600 ;
        RECT 41.230 238.100 41.830 238.600 ;
        RECT 42.030 238.100 42.580 238.600 ;
        RECT 6.830 221.400 7.430 221.900 ;
        RECT 7.630 221.400 8.230 221.900 ;
        RECT 8.430 221.400 9.030 221.900 ;
        RECT 9.230 221.400 9.830 221.900 ;
        RECT 10.030 221.400 10.630 221.900 ;
        RECT 18.830 221.400 19.430 221.900 ;
        RECT 19.630 221.400 20.230 221.900 ;
        RECT 20.430 221.400 21.030 221.900 ;
        RECT 21.230 221.400 21.830 221.900 ;
        RECT 22.030 221.400 22.580 221.900 ;
        RECT 46.830 238.100 47.430 238.600 ;
        RECT 47.630 238.100 48.230 238.600 ;
        RECT 48.430 238.100 49.030 238.600 ;
        RECT 49.230 238.100 49.830 238.600 ;
        RECT 50.030 238.100 50.630 238.600 ;
        RECT 58.830 238.100 59.430 238.600 ;
        RECT 59.630 238.100 60.230 238.600 ;
        RECT 60.430 238.100 61.030 238.600 ;
        RECT 61.230 238.100 61.830 238.600 ;
        RECT 62.030 238.100 62.580 238.600 ;
        RECT 26.830 221.400 27.430 221.900 ;
        RECT 27.630 221.400 28.230 221.900 ;
        RECT 28.430 221.400 29.030 221.900 ;
        RECT 29.230 221.400 29.830 221.900 ;
        RECT 30.030 221.400 30.630 221.900 ;
        RECT 38.830 221.400 39.430 221.900 ;
        RECT 39.630 221.400 40.230 221.900 ;
        RECT 40.430 221.400 41.030 221.900 ;
        RECT 41.230 221.400 41.830 221.900 ;
        RECT 42.030 221.400 42.580 221.900 ;
        RECT 66.830 238.100 67.430 238.600 ;
        RECT 67.630 238.100 68.230 238.600 ;
        RECT 68.430 238.100 69.030 238.600 ;
        RECT 69.230 238.100 69.830 238.600 ;
        RECT 70.030 238.100 70.630 238.600 ;
        RECT 78.830 238.100 79.430 238.600 ;
        RECT 79.630 238.100 80.230 238.600 ;
        RECT 80.430 238.100 81.030 238.600 ;
        RECT 81.230 238.100 81.830 238.600 ;
        RECT 82.030 238.100 82.580 238.600 ;
        RECT 46.830 221.400 47.430 221.900 ;
        RECT 47.630 221.400 48.230 221.900 ;
        RECT 48.430 221.400 49.030 221.900 ;
        RECT 49.230 221.400 49.830 221.900 ;
        RECT 50.030 221.400 50.630 221.900 ;
        RECT 58.830 221.400 59.430 221.900 ;
        RECT 59.630 221.400 60.230 221.900 ;
        RECT 60.430 221.400 61.030 221.900 ;
        RECT 61.230 221.400 61.830 221.900 ;
        RECT 62.030 221.400 62.580 221.900 ;
        RECT 86.830 238.100 87.430 238.600 ;
        RECT 87.630 238.100 88.230 238.600 ;
        RECT 88.430 238.100 89.030 238.600 ;
        RECT 89.230 238.100 89.830 238.600 ;
        RECT 90.030 238.100 90.630 238.600 ;
        RECT 98.830 238.100 99.430 238.600 ;
        RECT 99.630 238.100 100.230 238.600 ;
        RECT 100.430 238.100 101.030 238.600 ;
        RECT 101.230 238.100 101.830 238.600 ;
        RECT 102.030 238.100 102.580 238.600 ;
        RECT 66.830 221.400 67.430 221.900 ;
        RECT 67.630 221.400 68.230 221.900 ;
        RECT 68.430 221.400 69.030 221.900 ;
        RECT 69.230 221.400 69.830 221.900 ;
        RECT 70.030 221.400 70.630 221.900 ;
        RECT 78.830 221.400 79.430 221.900 ;
        RECT 79.630 221.400 80.230 221.900 ;
        RECT 80.430 221.400 81.030 221.900 ;
        RECT 81.230 221.400 81.830 221.900 ;
        RECT 82.030 221.400 82.580 221.900 ;
        RECT 106.830 238.100 107.430 238.600 ;
        RECT 107.630 238.100 108.230 238.600 ;
        RECT 108.430 238.100 109.030 238.600 ;
        RECT 109.230 238.100 109.830 238.600 ;
        RECT 110.030 238.100 110.630 238.600 ;
        RECT 118.830 238.100 119.430 238.600 ;
        RECT 119.630 238.100 120.230 238.600 ;
        RECT 120.430 238.100 121.030 238.600 ;
        RECT 121.230 238.100 121.830 238.600 ;
        RECT 122.030 238.100 122.580 238.600 ;
        RECT 86.830 221.400 87.430 221.900 ;
        RECT 87.630 221.400 88.230 221.900 ;
        RECT 88.430 221.400 89.030 221.900 ;
        RECT 89.230 221.400 89.830 221.900 ;
        RECT 90.030 221.400 90.630 221.900 ;
        RECT 98.830 221.400 99.430 221.900 ;
        RECT 99.630 221.400 100.230 221.900 ;
        RECT 100.430 221.400 101.030 221.900 ;
        RECT 101.230 221.400 101.830 221.900 ;
        RECT 102.030 221.400 102.580 221.900 ;
        RECT 106.830 221.400 107.430 221.900 ;
        RECT 107.630 221.400 108.230 221.900 ;
        RECT 108.430 221.400 109.030 221.900 ;
        RECT 109.230 221.400 109.830 221.900 ;
        RECT 110.030 221.400 110.630 221.900 ;
        RECT 118.830 221.400 119.430 221.900 ;
        RECT 119.630 221.400 120.230 221.900 ;
        RECT 120.430 221.400 121.030 221.900 ;
        RECT 121.230 221.400 121.830 221.900 ;
        RECT 122.030 221.400 122.580 221.900 ;
        RECT 6.830 218.100 7.430 218.600 ;
        RECT 7.630 218.100 8.230 218.600 ;
        RECT 8.430 218.100 9.030 218.600 ;
        RECT 9.230 218.100 9.830 218.600 ;
        RECT 10.030 218.100 10.630 218.600 ;
        RECT 18.830 218.100 19.430 218.600 ;
        RECT 19.630 218.100 20.230 218.600 ;
        RECT 20.430 218.100 21.030 218.600 ;
        RECT 21.230 218.100 21.830 218.600 ;
        RECT 22.030 218.100 22.580 218.600 ;
        RECT 2.520 214.920 2.880 215.300 ;
        RECT 3.130 214.920 3.490 215.300 ;
        RECT 3.760 214.920 4.120 215.300 ;
        RECT 2.520 214.185 2.880 214.565 ;
        RECT 3.130 214.185 3.490 214.565 ;
        RECT 3.760 214.185 4.120 214.565 ;
        RECT 2.520 213.500 2.880 213.880 ;
        RECT 3.130 213.500 3.490 213.880 ;
        RECT 3.760 213.500 4.120 213.880 ;
        RECT 2.520 206.120 2.880 206.500 ;
        RECT 3.130 206.120 3.490 206.500 ;
        RECT 3.760 206.120 4.120 206.500 ;
        RECT 2.520 205.385 2.880 205.765 ;
        RECT 3.130 205.385 3.490 205.765 ;
        RECT 3.760 205.385 4.120 205.765 ;
        RECT 2.520 204.700 2.880 205.080 ;
        RECT 3.130 204.700 3.490 205.080 ;
        RECT 3.760 204.700 4.120 205.080 ;
        RECT 26.830 218.100 27.430 218.600 ;
        RECT 27.630 218.100 28.230 218.600 ;
        RECT 28.430 218.100 29.030 218.600 ;
        RECT 29.230 218.100 29.830 218.600 ;
        RECT 30.030 218.100 30.630 218.600 ;
        RECT 38.830 218.100 39.430 218.600 ;
        RECT 39.630 218.100 40.230 218.600 ;
        RECT 40.430 218.100 41.030 218.600 ;
        RECT 41.230 218.100 41.830 218.600 ;
        RECT 42.030 218.100 42.580 218.600 ;
        RECT 6.830 201.400 7.430 201.900 ;
        RECT 7.630 201.400 8.230 201.900 ;
        RECT 8.430 201.400 9.030 201.900 ;
        RECT 9.230 201.400 9.830 201.900 ;
        RECT 10.030 201.400 10.630 201.900 ;
        RECT 18.830 201.400 19.430 201.900 ;
        RECT 19.630 201.400 20.230 201.900 ;
        RECT 20.430 201.400 21.030 201.900 ;
        RECT 21.230 201.400 21.830 201.900 ;
        RECT 22.030 201.400 22.580 201.900 ;
        RECT 46.830 218.100 47.430 218.600 ;
        RECT 47.630 218.100 48.230 218.600 ;
        RECT 48.430 218.100 49.030 218.600 ;
        RECT 49.230 218.100 49.830 218.600 ;
        RECT 50.030 218.100 50.630 218.600 ;
        RECT 58.830 218.100 59.430 218.600 ;
        RECT 59.630 218.100 60.230 218.600 ;
        RECT 60.430 218.100 61.030 218.600 ;
        RECT 61.230 218.100 61.830 218.600 ;
        RECT 62.030 218.100 62.580 218.600 ;
        RECT 26.830 201.400 27.430 201.900 ;
        RECT 27.630 201.400 28.230 201.900 ;
        RECT 28.430 201.400 29.030 201.900 ;
        RECT 29.230 201.400 29.830 201.900 ;
        RECT 30.030 201.400 30.630 201.900 ;
        RECT 38.830 201.400 39.430 201.900 ;
        RECT 39.630 201.400 40.230 201.900 ;
        RECT 40.430 201.400 41.030 201.900 ;
        RECT 41.230 201.400 41.830 201.900 ;
        RECT 42.030 201.400 42.580 201.900 ;
        RECT 66.830 218.100 67.430 218.600 ;
        RECT 67.630 218.100 68.230 218.600 ;
        RECT 68.430 218.100 69.030 218.600 ;
        RECT 69.230 218.100 69.830 218.600 ;
        RECT 70.030 218.100 70.630 218.600 ;
        RECT 78.830 218.100 79.430 218.600 ;
        RECT 79.630 218.100 80.230 218.600 ;
        RECT 80.430 218.100 81.030 218.600 ;
        RECT 81.230 218.100 81.830 218.600 ;
        RECT 82.030 218.100 82.580 218.600 ;
        RECT 46.830 201.400 47.430 201.900 ;
        RECT 47.630 201.400 48.230 201.900 ;
        RECT 48.430 201.400 49.030 201.900 ;
        RECT 49.230 201.400 49.830 201.900 ;
        RECT 50.030 201.400 50.630 201.900 ;
        RECT 58.830 201.400 59.430 201.900 ;
        RECT 59.630 201.400 60.230 201.900 ;
        RECT 60.430 201.400 61.030 201.900 ;
        RECT 61.230 201.400 61.830 201.900 ;
        RECT 62.030 201.400 62.580 201.900 ;
        RECT 86.830 218.100 87.430 218.600 ;
        RECT 87.630 218.100 88.230 218.600 ;
        RECT 88.430 218.100 89.030 218.600 ;
        RECT 89.230 218.100 89.830 218.600 ;
        RECT 90.030 218.100 90.630 218.600 ;
        RECT 98.830 218.100 99.430 218.600 ;
        RECT 99.630 218.100 100.230 218.600 ;
        RECT 100.430 218.100 101.030 218.600 ;
        RECT 101.230 218.100 101.830 218.600 ;
        RECT 102.030 218.100 102.580 218.600 ;
        RECT 66.830 201.400 67.430 201.900 ;
        RECT 67.630 201.400 68.230 201.900 ;
        RECT 68.430 201.400 69.030 201.900 ;
        RECT 69.230 201.400 69.830 201.900 ;
        RECT 70.030 201.400 70.630 201.900 ;
        RECT 78.830 201.400 79.430 201.900 ;
        RECT 79.630 201.400 80.230 201.900 ;
        RECT 80.430 201.400 81.030 201.900 ;
        RECT 81.230 201.400 81.830 201.900 ;
        RECT 82.030 201.400 82.580 201.900 ;
        RECT 106.830 218.100 107.430 218.600 ;
        RECT 107.630 218.100 108.230 218.600 ;
        RECT 108.430 218.100 109.030 218.600 ;
        RECT 109.230 218.100 109.830 218.600 ;
        RECT 110.030 218.100 110.630 218.600 ;
        RECT 118.830 218.100 119.430 218.600 ;
        RECT 119.630 218.100 120.230 218.600 ;
        RECT 120.430 218.100 121.030 218.600 ;
        RECT 121.230 218.100 121.830 218.600 ;
        RECT 122.030 218.100 122.580 218.600 ;
        RECT 86.830 201.400 87.430 201.900 ;
        RECT 87.630 201.400 88.230 201.900 ;
        RECT 88.430 201.400 89.030 201.900 ;
        RECT 89.230 201.400 89.830 201.900 ;
        RECT 90.030 201.400 90.630 201.900 ;
        RECT 98.830 201.400 99.430 201.900 ;
        RECT 99.630 201.400 100.230 201.900 ;
        RECT 100.430 201.400 101.030 201.900 ;
        RECT 101.230 201.400 101.830 201.900 ;
        RECT 102.030 201.400 102.580 201.900 ;
        RECT 106.830 201.400 107.430 201.900 ;
        RECT 107.630 201.400 108.230 201.900 ;
        RECT 108.430 201.400 109.030 201.900 ;
        RECT 109.230 201.400 109.830 201.900 ;
        RECT 110.030 201.400 110.630 201.900 ;
        RECT 118.830 201.400 119.430 201.900 ;
        RECT 119.630 201.400 120.230 201.900 ;
        RECT 120.430 201.400 121.030 201.900 ;
        RECT 121.230 201.400 121.830 201.900 ;
        RECT 122.030 201.400 122.580 201.900 ;
        RECT 4.845 175.310 5.205 175.685 ;
        RECT 5.630 175.315 5.830 175.690 ;
        RECT 7.245 175.375 7.415 175.545 ;
        RECT 4.860 174.730 5.220 175.105 ;
        RECT 5.630 174.745 5.990 175.120 ;
        RECT 8.020 175.295 8.190 175.625 ;
        RECT 9.600 175.345 9.770 175.620 ;
        RECT 15.010 175.370 15.180 175.540 ;
        RECT 15.470 175.370 15.640 175.540 ;
        RECT 15.930 175.370 16.100 175.540 ;
        RECT 16.390 175.370 16.560 175.540 ;
        RECT 16.850 175.370 17.020 175.540 ;
        RECT 17.310 175.370 17.480 175.540 ;
        RECT 17.770 175.370 17.940 175.540 ;
        RECT 18.230 175.370 18.400 175.540 ;
        RECT 18.690 175.370 18.860 175.540 ;
        RECT 19.150 175.370 19.320 175.540 ;
        RECT 19.610 175.370 19.780 175.540 ;
        RECT 20.070 175.370 20.240 175.540 ;
        RECT 20.530 175.370 20.700 175.540 ;
        RECT 20.990 175.370 21.160 175.540 ;
        RECT 21.450 175.370 21.620 175.540 ;
        RECT 21.910 175.370 22.080 175.540 ;
        RECT 22.370 175.370 22.540 175.540 ;
        RECT 22.830 175.370 23.000 175.540 ;
        RECT 23.290 175.370 23.460 175.540 ;
        RECT 8.020 174.445 8.190 174.720 ;
        RECT 9.600 174.445 9.770 174.720 ;
        RECT 44.735 174.760 45.335 175.260 ;
        RECT 45.535 174.760 46.135 175.260 ;
        RECT 46.335 174.760 46.935 175.260 ;
        RECT 47.135 174.760 47.735 175.260 ;
        RECT 47.935 174.760 48.535 175.260 ;
        RECT 56.735 174.760 57.335 175.260 ;
        RECT 57.535 174.760 58.135 175.260 ;
        RECT 58.335 174.760 58.935 175.260 ;
        RECT 59.135 174.760 59.735 175.260 ;
        RECT 59.935 174.760 60.485 175.260 ;
        RECT 6.730 169.930 6.900 170.100 ;
        RECT 7.190 169.930 7.360 170.100 ;
        RECT 7.650 169.930 7.820 170.100 ;
        RECT 8.110 169.930 8.280 170.100 ;
        RECT 8.570 169.930 8.740 170.100 ;
        RECT 9.030 169.930 9.200 170.100 ;
        RECT 9.490 169.930 9.660 170.100 ;
        RECT 9.950 169.930 10.120 170.100 ;
        RECT 10.410 169.930 10.580 170.100 ;
        RECT 10.870 169.930 11.040 170.100 ;
        RECT 11.330 169.930 11.500 170.100 ;
        RECT 11.790 169.930 11.960 170.100 ;
        RECT 12.250 169.930 12.420 170.100 ;
        RECT 12.710 169.930 12.880 170.100 ;
        RECT 13.170 169.930 13.340 170.100 ;
        RECT 13.630 169.930 13.800 170.100 ;
        RECT 14.090 169.930 14.260 170.100 ;
        RECT 14.550 169.930 14.720 170.100 ;
        RECT 15.010 169.930 15.180 170.100 ;
        RECT 15.470 169.930 15.640 170.100 ;
        RECT 15.930 169.930 16.100 170.100 ;
        RECT 16.390 169.930 16.560 170.100 ;
        RECT 16.850 169.930 17.020 170.100 ;
        RECT 17.310 169.930 17.480 170.100 ;
        RECT 17.770 169.930 17.940 170.100 ;
        RECT 18.230 169.930 18.400 170.100 ;
        RECT 18.690 169.930 18.860 170.100 ;
        RECT 19.150 169.930 19.320 170.100 ;
        RECT 19.610 169.930 19.780 170.100 ;
        RECT 20.070 169.930 20.240 170.100 ;
        RECT 20.530 169.930 20.700 170.100 ;
        RECT 20.990 169.930 21.160 170.100 ;
        RECT 21.450 169.930 21.620 170.100 ;
        RECT 21.910 169.930 22.080 170.100 ;
        RECT 22.370 169.930 22.540 170.100 ;
        RECT 22.830 169.930 23.000 170.100 ;
        RECT 23.290 169.930 23.460 170.100 ;
        RECT 23.750 169.930 23.920 170.100 ;
        RECT 4.875 164.955 5.350 165.395 ;
        RECT 5.540 164.955 6.015 165.395 ;
        RECT 4.875 164.305 5.350 164.745 ;
        RECT 5.545 164.305 6.020 164.745 ;
        RECT 7.650 164.490 7.820 164.660 ;
        RECT 15.010 164.490 15.180 164.660 ;
        RECT 15.470 164.490 15.640 164.660 ;
        RECT 15.930 164.490 16.100 164.660 ;
        RECT 16.390 164.490 16.560 164.660 ;
        RECT 16.850 164.490 17.020 164.660 ;
        RECT 17.310 164.490 17.480 164.660 ;
        RECT 17.770 164.490 17.940 164.660 ;
        RECT 18.230 164.490 18.400 164.660 ;
        RECT 18.690 164.490 18.860 164.660 ;
        RECT 19.150 164.490 19.320 164.660 ;
        RECT 19.610 164.490 19.780 164.660 ;
        RECT 20.070 164.490 20.240 164.660 ;
        RECT 20.530 164.490 20.700 164.660 ;
        RECT 20.990 164.490 21.160 164.660 ;
        RECT 21.450 164.490 21.620 164.660 ;
        RECT 21.910 164.490 22.080 164.660 ;
        RECT 22.370 164.490 22.540 164.660 ;
        RECT 22.830 164.490 23.000 164.660 ;
        RECT 23.290 164.490 23.460 164.660 ;
        RECT 64.735 174.760 65.335 175.260 ;
        RECT 65.535 174.760 66.135 175.260 ;
        RECT 66.335 174.760 66.935 175.260 ;
        RECT 67.135 174.760 67.735 175.260 ;
        RECT 67.935 174.760 68.535 175.260 ;
        RECT 76.735 174.760 77.335 175.260 ;
        RECT 77.535 174.760 78.135 175.260 ;
        RECT 78.335 174.760 78.935 175.260 ;
        RECT 79.135 174.760 79.735 175.260 ;
        RECT 79.935 174.760 80.485 175.260 ;
        RECT 44.735 158.060 45.335 158.560 ;
        RECT 45.535 158.060 46.135 158.560 ;
        RECT 46.335 158.060 46.935 158.560 ;
        RECT 47.135 158.060 47.735 158.560 ;
        RECT 47.935 158.060 48.535 158.560 ;
        RECT 56.735 158.060 57.335 158.560 ;
        RECT 57.535 158.060 58.135 158.560 ;
        RECT 58.335 158.060 58.935 158.560 ;
        RECT 59.135 158.060 59.735 158.560 ;
        RECT 59.935 158.060 60.485 158.560 ;
        RECT 84.735 174.760 85.335 175.260 ;
        RECT 85.535 174.760 86.135 175.260 ;
        RECT 86.335 174.760 86.935 175.260 ;
        RECT 87.135 174.760 87.735 175.260 ;
        RECT 87.935 174.760 88.535 175.260 ;
        RECT 96.735 174.760 97.335 175.260 ;
        RECT 97.535 174.760 98.135 175.260 ;
        RECT 98.335 174.760 98.935 175.260 ;
        RECT 99.135 174.760 99.735 175.260 ;
        RECT 99.935 174.760 100.485 175.260 ;
        RECT 64.735 158.060 65.335 158.560 ;
        RECT 65.535 158.060 66.135 158.560 ;
        RECT 66.335 158.060 66.935 158.560 ;
        RECT 67.135 158.060 67.735 158.560 ;
        RECT 67.935 158.060 68.535 158.560 ;
        RECT 76.735 158.060 77.335 158.560 ;
        RECT 77.535 158.060 78.135 158.560 ;
        RECT 78.335 158.060 78.935 158.560 ;
        RECT 79.135 158.060 79.735 158.560 ;
        RECT 79.935 158.060 80.485 158.560 ;
        RECT 104.735 174.760 105.335 175.260 ;
        RECT 105.535 174.760 106.135 175.260 ;
        RECT 106.335 174.760 106.935 175.260 ;
        RECT 107.135 174.760 107.735 175.260 ;
        RECT 107.935 174.760 108.535 175.260 ;
        RECT 116.735 174.760 117.335 175.260 ;
        RECT 117.535 174.760 118.135 175.260 ;
        RECT 118.335 174.760 118.935 175.260 ;
        RECT 119.135 174.760 119.735 175.260 ;
        RECT 119.935 174.760 120.485 175.260 ;
        RECT 84.735 158.060 85.335 158.560 ;
        RECT 85.535 158.060 86.135 158.560 ;
        RECT 86.335 158.060 86.935 158.560 ;
        RECT 87.135 158.060 87.735 158.560 ;
        RECT 87.935 158.060 88.535 158.560 ;
        RECT 96.735 158.060 97.335 158.560 ;
        RECT 97.535 158.060 98.135 158.560 ;
        RECT 98.335 158.060 98.935 158.560 ;
        RECT 99.135 158.060 99.735 158.560 ;
        RECT 99.935 158.060 100.485 158.560 ;
        RECT 125.345 171.580 125.705 171.960 ;
        RECT 125.955 171.580 126.315 171.960 ;
        RECT 126.585 171.580 126.945 171.960 ;
        RECT 125.345 170.845 125.705 171.225 ;
        RECT 125.955 170.845 126.315 171.225 ;
        RECT 126.585 170.845 126.945 171.225 ;
        RECT 125.345 170.160 125.705 170.540 ;
        RECT 125.955 170.160 126.315 170.540 ;
        RECT 126.585 170.160 126.945 170.540 ;
        RECT 125.345 162.780 125.705 163.160 ;
        RECT 125.955 162.780 126.315 163.160 ;
        RECT 126.585 162.780 126.945 163.160 ;
        RECT 125.345 162.045 125.705 162.425 ;
        RECT 125.955 162.045 126.315 162.425 ;
        RECT 126.585 162.045 126.945 162.425 ;
        RECT 125.345 161.360 125.705 161.740 ;
        RECT 125.955 161.360 126.315 161.740 ;
        RECT 126.585 161.360 126.945 161.740 ;
        RECT 104.735 158.060 105.335 158.560 ;
        RECT 105.535 158.060 106.135 158.560 ;
        RECT 106.335 158.060 106.935 158.560 ;
        RECT 107.135 158.060 107.735 158.560 ;
        RECT 107.935 158.060 108.535 158.560 ;
        RECT 116.735 158.060 117.335 158.560 ;
        RECT 117.535 158.060 118.135 158.560 ;
        RECT 118.335 158.060 118.935 158.560 ;
        RECT 119.135 158.060 119.735 158.560 ;
        RECT 119.935 158.060 120.485 158.560 ;
        RECT 6.830 138.100 7.430 138.600 ;
        RECT 7.630 138.100 8.230 138.600 ;
        RECT 8.430 138.100 9.030 138.600 ;
        RECT 9.230 138.100 9.830 138.600 ;
        RECT 10.030 138.100 10.630 138.600 ;
        RECT 18.830 138.100 19.430 138.600 ;
        RECT 19.630 138.100 20.230 138.600 ;
        RECT 20.430 138.100 21.030 138.600 ;
        RECT 21.230 138.100 21.830 138.600 ;
        RECT 22.030 138.100 22.580 138.600 ;
        RECT 2.520 134.925 2.880 135.305 ;
        RECT 3.130 134.925 3.490 135.305 ;
        RECT 3.760 134.925 4.120 135.305 ;
        RECT 2.520 134.190 2.880 134.570 ;
        RECT 3.130 134.190 3.490 134.570 ;
        RECT 3.760 134.190 4.120 134.570 ;
        RECT 2.520 133.505 2.880 133.885 ;
        RECT 3.130 133.505 3.490 133.885 ;
        RECT 3.760 133.505 4.120 133.885 ;
        RECT 2.520 126.090 2.880 126.470 ;
        RECT 3.130 126.090 3.490 126.470 ;
        RECT 3.760 126.090 4.120 126.470 ;
        RECT 2.520 125.355 2.880 125.735 ;
        RECT 3.130 125.355 3.490 125.735 ;
        RECT 3.760 125.355 4.120 125.735 ;
        RECT 2.520 124.670 2.880 125.050 ;
        RECT 3.130 124.670 3.490 125.050 ;
        RECT 3.760 124.670 4.120 125.050 ;
        RECT 26.830 138.100 27.430 138.600 ;
        RECT 27.630 138.100 28.230 138.600 ;
        RECT 28.430 138.100 29.030 138.600 ;
        RECT 29.230 138.100 29.830 138.600 ;
        RECT 30.030 138.100 30.630 138.600 ;
        RECT 38.830 138.100 39.430 138.600 ;
        RECT 39.630 138.100 40.230 138.600 ;
        RECT 40.430 138.100 41.030 138.600 ;
        RECT 41.230 138.100 41.830 138.600 ;
        RECT 42.030 138.100 42.580 138.600 ;
        RECT 6.830 121.400 7.430 121.900 ;
        RECT 7.630 121.400 8.230 121.900 ;
        RECT 8.430 121.400 9.030 121.900 ;
        RECT 9.230 121.400 9.830 121.900 ;
        RECT 10.030 121.400 10.630 121.900 ;
        RECT 18.830 121.400 19.430 121.900 ;
        RECT 19.630 121.400 20.230 121.900 ;
        RECT 20.430 121.400 21.030 121.900 ;
        RECT 21.230 121.400 21.830 121.900 ;
        RECT 22.030 121.400 22.580 121.900 ;
        RECT 46.830 138.100 47.430 138.600 ;
        RECT 47.630 138.100 48.230 138.600 ;
        RECT 48.430 138.100 49.030 138.600 ;
        RECT 49.230 138.100 49.830 138.600 ;
        RECT 50.030 138.100 50.630 138.600 ;
        RECT 58.830 138.100 59.430 138.600 ;
        RECT 59.630 138.100 60.230 138.600 ;
        RECT 60.430 138.100 61.030 138.600 ;
        RECT 61.230 138.100 61.830 138.600 ;
        RECT 62.030 138.100 62.580 138.600 ;
        RECT 26.830 121.400 27.430 121.900 ;
        RECT 27.630 121.400 28.230 121.900 ;
        RECT 28.430 121.400 29.030 121.900 ;
        RECT 29.230 121.400 29.830 121.900 ;
        RECT 30.030 121.400 30.630 121.900 ;
        RECT 38.830 121.400 39.430 121.900 ;
        RECT 39.630 121.400 40.230 121.900 ;
        RECT 40.430 121.400 41.030 121.900 ;
        RECT 41.230 121.400 41.830 121.900 ;
        RECT 42.030 121.400 42.580 121.900 ;
        RECT 66.830 138.100 67.430 138.600 ;
        RECT 67.630 138.100 68.230 138.600 ;
        RECT 68.430 138.100 69.030 138.600 ;
        RECT 69.230 138.100 69.830 138.600 ;
        RECT 70.030 138.100 70.630 138.600 ;
        RECT 78.830 138.100 79.430 138.600 ;
        RECT 79.630 138.100 80.230 138.600 ;
        RECT 80.430 138.100 81.030 138.600 ;
        RECT 81.230 138.100 81.830 138.600 ;
        RECT 82.030 138.100 82.580 138.600 ;
        RECT 46.830 121.400 47.430 121.900 ;
        RECT 47.630 121.400 48.230 121.900 ;
        RECT 48.430 121.400 49.030 121.900 ;
        RECT 49.230 121.400 49.830 121.900 ;
        RECT 50.030 121.400 50.630 121.900 ;
        RECT 58.830 121.400 59.430 121.900 ;
        RECT 59.630 121.400 60.230 121.900 ;
        RECT 60.430 121.400 61.030 121.900 ;
        RECT 61.230 121.400 61.830 121.900 ;
        RECT 62.030 121.400 62.580 121.900 ;
        RECT 86.830 138.100 87.430 138.600 ;
        RECT 87.630 138.100 88.230 138.600 ;
        RECT 88.430 138.100 89.030 138.600 ;
        RECT 89.230 138.100 89.830 138.600 ;
        RECT 90.030 138.100 90.630 138.600 ;
        RECT 98.830 138.100 99.430 138.600 ;
        RECT 99.630 138.100 100.230 138.600 ;
        RECT 100.430 138.100 101.030 138.600 ;
        RECT 101.230 138.100 101.830 138.600 ;
        RECT 102.030 138.100 102.580 138.600 ;
        RECT 66.830 121.400 67.430 121.900 ;
        RECT 67.630 121.400 68.230 121.900 ;
        RECT 68.430 121.400 69.030 121.900 ;
        RECT 69.230 121.400 69.830 121.900 ;
        RECT 70.030 121.400 70.630 121.900 ;
        RECT 78.830 121.400 79.430 121.900 ;
        RECT 79.630 121.400 80.230 121.900 ;
        RECT 80.430 121.400 81.030 121.900 ;
        RECT 81.230 121.400 81.830 121.900 ;
        RECT 82.030 121.400 82.580 121.900 ;
        RECT 106.830 138.100 107.430 138.600 ;
        RECT 107.630 138.100 108.230 138.600 ;
        RECT 108.430 138.100 109.030 138.600 ;
        RECT 109.230 138.100 109.830 138.600 ;
        RECT 110.030 138.100 110.630 138.600 ;
        RECT 118.830 138.100 119.430 138.600 ;
        RECT 119.630 138.100 120.230 138.600 ;
        RECT 120.430 138.100 121.030 138.600 ;
        RECT 121.230 138.100 121.830 138.600 ;
        RECT 122.030 138.100 122.580 138.600 ;
        RECT 86.830 121.400 87.430 121.900 ;
        RECT 87.630 121.400 88.230 121.900 ;
        RECT 88.430 121.400 89.030 121.900 ;
        RECT 89.230 121.400 89.830 121.900 ;
        RECT 90.030 121.400 90.630 121.900 ;
        RECT 98.830 121.400 99.430 121.900 ;
        RECT 99.630 121.400 100.230 121.900 ;
        RECT 100.430 121.400 101.030 121.900 ;
        RECT 101.230 121.400 101.830 121.900 ;
        RECT 102.030 121.400 102.580 121.900 ;
        RECT 106.830 121.400 107.430 121.900 ;
        RECT 107.630 121.400 108.230 121.900 ;
        RECT 108.430 121.400 109.030 121.900 ;
        RECT 109.230 121.400 109.830 121.900 ;
        RECT 110.030 121.400 110.630 121.900 ;
        RECT 118.830 121.400 119.430 121.900 ;
        RECT 119.630 121.400 120.230 121.900 ;
        RECT 120.430 121.400 121.030 121.900 ;
        RECT 121.230 121.400 121.830 121.900 ;
        RECT 122.030 121.400 122.580 121.900 ;
        RECT 6.830 118.100 7.430 118.600 ;
        RECT 7.630 118.100 8.230 118.600 ;
        RECT 8.430 118.100 9.030 118.600 ;
        RECT 9.230 118.100 9.830 118.600 ;
        RECT 10.030 118.100 10.630 118.600 ;
        RECT 18.830 118.100 19.430 118.600 ;
        RECT 19.630 118.100 20.230 118.600 ;
        RECT 20.430 118.100 21.030 118.600 ;
        RECT 21.230 118.100 21.830 118.600 ;
        RECT 22.030 118.100 22.580 118.600 ;
        RECT 2.520 114.920 2.880 115.300 ;
        RECT 3.130 114.920 3.490 115.300 ;
        RECT 3.760 114.920 4.120 115.300 ;
        RECT 2.520 114.185 2.880 114.565 ;
        RECT 3.130 114.185 3.490 114.565 ;
        RECT 3.760 114.185 4.120 114.565 ;
        RECT 2.520 113.500 2.880 113.880 ;
        RECT 3.130 113.500 3.490 113.880 ;
        RECT 3.760 113.500 4.120 113.880 ;
        RECT 2.520 106.120 2.880 106.500 ;
        RECT 3.130 106.120 3.490 106.500 ;
        RECT 3.760 106.120 4.120 106.500 ;
        RECT 2.520 105.385 2.880 105.765 ;
        RECT 3.130 105.385 3.490 105.765 ;
        RECT 3.760 105.385 4.120 105.765 ;
        RECT 2.520 104.700 2.880 105.080 ;
        RECT 3.130 104.700 3.490 105.080 ;
        RECT 3.760 104.700 4.120 105.080 ;
        RECT 26.830 118.100 27.430 118.600 ;
        RECT 27.630 118.100 28.230 118.600 ;
        RECT 28.430 118.100 29.030 118.600 ;
        RECT 29.230 118.100 29.830 118.600 ;
        RECT 30.030 118.100 30.630 118.600 ;
        RECT 38.830 118.100 39.430 118.600 ;
        RECT 39.630 118.100 40.230 118.600 ;
        RECT 40.430 118.100 41.030 118.600 ;
        RECT 41.230 118.100 41.830 118.600 ;
        RECT 42.030 118.100 42.580 118.600 ;
        RECT 6.830 101.400 7.430 101.900 ;
        RECT 7.630 101.400 8.230 101.900 ;
        RECT 8.430 101.400 9.030 101.900 ;
        RECT 9.230 101.400 9.830 101.900 ;
        RECT 10.030 101.400 10.630 101.900 ;
        RECT 18.830 101.400 19.430 101.900 ;
        RECT 19.630 101.400 20.230 101.900 ;
        RECT 20.430 101.400 21.030 101.900 ;
        RECT 21.230 101.400 21.830 101.900 ;
        RECT 22.030 101.400 22.580 101.900 ;
        RECT 46.830 118.100 47.430 118.600 ;
        RECT 47.630 118.100 48.230 118.600 ;
        RECT 48.430 118.100 49.030 118.600 ;
        RECT 49.230 118.100 49.830 118.600 ;
        RECT 50.030 118.100 50.630 118.600 ;
        RECT 58.830 118.100 59.430 118.600 ;
        RECT 59.630 118.100 60.230 118.600 ;
        RECT 60.430 118.100 61.030 118.600 ;
        RECT 61.230 118.100 61.830 118.600 ;
        RECT 62.030 118.100 62.580 118.600 ;
        RECT 26.830 101.400 27.430 101.900 ;
        RECT 27.630 101.400 28.230 101.900 ;
        RECT 28.430 101.400 29.030 101.900 ;
        RECT 29.230 101.400 29.830 101.900 ;
        RECT 30.030 101.400 30.630 101.900 ;
        RECT 38.830 101.400 39.430 101.900 ;
        RECT 39.630 101.400 40.230 101.900 ;
        RECT 40.430 101.400 41.030 101.900 ;
        RECT 41.230 101.400 41.830 101.900 ;
        RECT 42.030 101.400 42.580 101.900 ;
        RECT 66.830 118.100 67.430 118.600 ;
        RECT 67.630 118.100 68.230 118.600 ;
        RECT 68.430 118.100 69.030 118.600 ;
        RECT 69.230 118.100 69.830 118.600 ;
        RECT 70.030 118.100 70.630 118.600 ;
        RECT 78.830 118.100 79.430 118.600 ;
        RECT 79.630 118.100 80.230 118.600 ;
        RECT 80.430 118.100 81.030 118.600 ;
        RECT 81.230 118.100 81.830 118.600 ;
        RECT 82.030 118.100 82.580 118.600 ;
        RECT 46.830 101.400 47.430 101.900 ;
        RECT 47.630 101.400 48.230 101.900 ;
        RECT 48.430 101.400 49.030 101.900 ;
        RECT 49.230 101.400 49.830 101.900 ;
        RECT 50.030 101.400 50.630 101.900 ;
        RECT 58.830 101.400 59.430 101.900 ;
        RECT 59.630 101.400 60.230 101.900 ;
        RECT 60.430 101.400 61.030 101.900 ;
        RECT 61.230 101.400 61.830 101.900 ;
        RECT 62.030 101.400 62.580 101.900 ;
        RECT 86.830 118.100 87.430 118.600 ;
        RECT 87.630 118.100 88.230 118.600 ;
        RECT 88.430 118.100 89.030 118.600 ;
        RECT 89.230 118.100 89.830 118.600 ;
        RECT 90.030 118.100 90.630 118.600 ;
        RECT 98.830 118.100 99.430 118.600 ;
        RECT 99.630 118.100 100.230 118.600 ;
        RECT 100.430 118.100 101.030 118.600 ;
        RECT 101.230 118.100 101.830 118.600 ;
        RECT 102.030 118.100 102.580 118.600 ;
        RECT 66.830 101.400 67.430 101.900 ;
        RECT 67.630 101.400 68.230 101.900 ;
        RECT 68.430 101.400 69.030 101.900 ;
        RECT 69.230 101.400 69.830 101.900 ;
        RECT 70.030 101.400 70.630 101.900 ;
        RECT 78.830 101.400 79.430 101.900 ;
        RECT 79.630 101.400 80.230 101.900 ;
        RECT 80.430 101.400 81.030 101.900 ;
        RECT 81.230 101.400 81.830 101.900 ;
        RECT 82.030 101.400 82.580 101.900 ;
        RECT 106.830 118.100 107.430 118.600 ;
        RECT 107.630 118.100 108.230 118.600 ;
        RECT 108.430 118.100 109.030 118.600 ;
        RECT 109.230 118.100 109.830 118.600 ;
        RECT 110.030 118.100 110.630 118.600 ;
        RECT 118.830 118.100 119.430 118.600 ;
        RECT 119.630 118.100 120.230 118.600 ;
        RECT 120.430 118.100 121.030 118.600 ;
        RECT 121.230 118.100 121.830 118.600 ;
        RECT 122.030 118.100 122.580 118.600 ;
        RECT 86.830 101.400 87.430 101.900 ;
        RECT 87.630 101.400 88.230 101.900 ;
        RECT 88.430 101.400 89.030 101.900 ;
        RECT 89.230 101.400 89.830 101.900 ;
        RECT 90.030 101.400 90.630 101.900 ;
        RECT 98.830 101.400 99.430 101.900 ;
        RECT 99.630 101.400 100.230 101.900 ;
        RECT 100.430 101.400 101.030 101.900 ;
        RECT 101.230 101.400 101.830 101.900 ;
        RECT 102.030 101.400 102.580 101.900 ;
        RECT 106.830 101.400 107.430 101.900 ;
        RECT 107.630 101.400 108.230 101.900 ;
        RECT 108.430 101.400 109.030 101.900 ;
        RECT 109.230 101.400 109.830 101.900 ;
        RECT 110.030 101.400 110.630 101.900 ;
        RECT 118.830 101.400 119.430 101.900 ;
        RECT 119.630 101.400 120.230 101.900 ;
        RECT 120.430 101.400 121.030 101.900 ;
        RECT 121.230 101.400 121.830 101.900 ;
        RECT 122.030 101.400 122.580 101.900 ;
        RECT 6.830 98.100 7.430 98.600 ;
        RECT 7.630 98.100 8.230 98.600 ;
        RECT 8.430 98.100 9.030 98.600 ;
        RECT 9.230 98.100 9.830 98.600 ;
        RECT 10.030 98.100 10.630 98.600 ;
        RECT 18.830 98.100 19.430 98.600 ;
        RECT 19.630 98.100 20.230 98.600 ;
        RECT 20.430 98.100 21.030 98.600 ;
        RECT 21.230 98.100 21.830 98.600 ;
        RECT 22.030 98.100 22.580 98.600 ;
        RECT 2.520 94.920 2.880 95.300 ;
        RECT 3.130 94.920 3.490 95.300 ;
        RECT 3.760 94.920 4.120 95.300 ;
        RECT 2.520 94.185 2.880 94.565 ;
        RECT 3.130 94.185 3.490 94.565 ;
        RECT 3.760 94.185 4.120 94.565 ;
        RECT 2.520 93.500 2.880 93.880 ;
        RECT 3.130 93.500 3.490 93.880 ;
        RECT 3.760 93.500 4.120 93.880 ;
        RECT 2.520 86.125 2.880 86.505 ;
        RECT 3.130 86.125 3.490 86.505 ;
        RECT 3.760 86.125 4.120 86.505 ;
        RECT 2.520 85.390 2.880 85.770 ;
        RECT 3.130 85.390 3.490 85.770 ;
        RECT 3.760 85.390 4.120 85.770 ;
        RECT 2.520 84.705 2.880 85.085 ;
        RECT 3.130 84.705 3.490 85.085 ;
        RECT 3.760 84.705 4.120 85.085 ;
        RECT 26.830 98.100 27.430 98.600 ;
        RECT 27.630 98.100 28.230 98.600 ;
        RECT 28.430 98.100 29.030 98.600 ;
        RECT 29.230 98.100 29.830 98.600 ;
        RECT 30.030 98.100 30.630 98.600 ;
        RECT 38.830 98.100 39.430 98.600 ;
        RECT 39.630 98.100 40.230 98.600 ;
        RECT 40.430 98.100 41.030 98.600 ;
        RECT 41.230 98.100 41.830 98.600 ;
        RECT 42.030 98.100 42.580 98.600 ;
        RECT 6.830 81.400 7.430 81.900 ;
        RECT 7.630 81.400 8.230 81.900 ;
        RECT 8.430 81.400 9.030 81.900 ;
        RECT 9.230 81.400 9.830 81.900 ;
        RECT 10.030 81.400 10.630 81.900 ;
        RECT 18.830 81.400 19.430 81.900 ;
        RECT 19.630 81.400 20.230 81.900 ;
        RECT 20.430 81.400 21.030 81.900 ;
        RECT 21.230 81.400 21.830 81.900 ;
        RECT 22.030 81.400 22.580 81.900 ;
        RECT 46.830 98.100 47.430 98.600 ;
        RECT 47.630 98.100 48.230 98.600 ;
        RECT 48.430 98.100 49.030 98.600 ;
        RECT 49.230 98.100 49.830 98.600 ;
        RECT 50.030 98.100 50.630 98.600 ;
        RECT 58.830 98.100 59.430 98.600 ;
        RECT 59.630 98.100 60.230 98.600 ;
        RECT 60.430 98.100 61.030 98.600 ;
        RECT 61.230 98.100 61.830 98.600 ;
        RECT 62.030 98.100 62.580 98.600 ;
        RECT 26.830 81.400 27.430 81.900 ;
        RECT 27.630 81.400 28.230 81.900 ;
        RECT 28.430 81.400 29.030 81.900 ;
        RECT 29.230 81.400 29.830 81.900 ;
        RECT 30.030 81.400 30.630 81.900 ;
        RECT 38.830 81.400 39.430 81.900 ;
        RECT 39.630 81.400 40.230 81.900 ;
        RECT 40.430 81.400 41.030 81.900 ;
        RECT 41.230 81.400 41.830 81.900 ;
        RECT 42.030 81.400 42.580 81.900 ;
        RECT 66.830 98.100 67.430 98.600 ;
        RECT 67.630 98.100 68.230 98.600 ;
        RECT 68.430 98.100 69.030 98.600 ;
        RECT 69.230 98.100 69.830 98.600 ;
        RECT 70.030 98.100 70.630 98.600 ;
        RECT 78.830 98.100 79.430 98.600 ;
        RECT 79.630 98.100 80.230 98.600 ;
        RECT 80.430 98.100 81.030 98.600 ;
        RECT 81.230 98.100 81.830 98.600 ;
        RECT 82.030 98.100 82.580 98.600 ;
        RECT 46.830 81.400 47.430 81.900 ;
        RECT 47.630 81.400 48.230 81.900 ;
        RECT 48.430 81.400 49.030 81.900 ;
        RECT 49.230 81.400 49.830 81.900 ;
        RECT 50.030 81.400 50.630 81.900 ;
        RECT 58.830 81.400 59.430 81.900 ;
        RECT 59.630 81.400 60.230 81.900 ;
        RECT 60.430 81.400 61.030 81.900 ;
        RECT 61.230 81.400 61.830 81.900 ;
        RECT 62.030 81.400 62.580 81.900 ;
        RECT 86.830 98.100 87.430 98.600 ;
        RECT 87.630 98.100 88.230 98.600 ;
        RECT 88.430 98.100 89.030 98.600 ;
        RECT 89.230 98.100 89.830 98.600 ;
        RECT 90.030 98.100 90.630 98.600 ;
        RECT 98.830 98.100 99.430 98.600 ;
        RECT 99.630 98.100 100.230 98.600 ;
        RECT 100.430 98.100 101.030 98.600 ;
        RECT 101.230 98.100 101.830 98.600 ;
        RECT 102.030 98.100 102.580 98.600 ;
        RECT 66.830 81.400 67.430 81.900 ;
        RECT 67.630 81.400 68.230 81.900 ;
        RECT 68.430 81.400 69.030 81.900 ;
        RECT 69.230 81.400 69.830 81.900 ;
        RECT 70.030 81.400 70.630 81.900 ;
        RECT 78.830 81.400 79.430 81.900 ;
        RECT 79.630 81.400 80.230 81.900 ;
        RECT 80.430 81.400 81.030 81.900 ;
        RECT 81.230 81.400 81.830 81.900 ;
        RECT 82.030 81.400 82.580 81.900 ;
        RECT 106.830 98.100 107.430 98.600 ;
        RECT 107.630 98.100 108.230 98.600 ;
        RECT 108.430 98.100 109.030 98.600 ;
        RECT 109.230 98.100 109.830 98.600 ;
        RECT 110.030 98.100 110.630 98.600 ;
        RECT 118.830 98.100 119.430 98.600 ;
        RECT 119.630 98.100 120.230 98.600 ;
        RECT 120.430 98.100 121.030 98.600 ;
        RECT 121.230 98.100 121.830 98.600 ;
        RECT 122.030 98.100 122.580 98.600 ;
        RECT 86.830 81.400 87.430 81.900 ;
        RECT 87.630 81.400 88.230 81.900 ;
        RECT 88.430 81.400 89.030 81.900 ;
        RECT 89.230 81.400 89.830 81.900 ;
        RECT 90.030 81.400 90.630 81.900 ;
        RECT 98.830 81.400 99.430 81.900 ;
        RECT 99.630 81.400 100.230 81.900 ;
        RECT 100.430 81.400 101.030 81.900 ;
        RECT 101.230 81.400 101.830 81.900 ;
        RECT 102.030 81.400 102.580 81.900 ;
        RECT 106.830 81.400 107.430 81.900 ;
        RECT 107.630 81.400 108.230 81.900 ;
        RECT 108.430 81.400 109.030 81.900 ;
        RECT 109.230 81.400 109.830 81.900 ;
        RECT 110.030 81.400 110.630 81.900 ;
        RECT 118.830 81.400 119.430 81.900 ;
        RECT 119.630 81.400 120.230 81.900 ;
        RECT 120.430 81.400 121.030 81.900 ;
        RECT 121.230 81.400 121.830 81.900 ;
        RECT 122.030 81.400 122.580 81.900 ;
        RECT 6.830 78.100 7.430 78.600 ;
        RECT 7.630 78.100 8.230 78.600 ;
        RECT 8.430 78.100 9.030 78.600 ;
        RECT 9.230 78.100 9.830 78.600 ;
        RECT 10.030 78.100 10.630 78.600 ;
        RECT 18.830 78.100 19.430 78.600 ;
        RECT 19.630 78.100 20.230 78.600 ;
        RECT 20.430 78.100 21.030 78.600 ;
        RECT 21.230 78.100 21.830 78.600 ;
        RECT 22.030 78.100 22.580 78.600 ;
        RECT 2.520 74.920 2.880 75.300 ;
        RECT 3.130 74.920 3.490 75.300 ;
        RECT 3.760 74.920 4.120 75.300 ;
        RECT 2.520 74.185 2.880 74.565 ;
        RECT 3.130 74.185 3.490 74.565 ;
        RECT 3.760 74.185 4.120 74.565 ;
        RECT 2.520 73.500 2.880 73.880 ;
        RECT 3.130 73.500 3.490 73.880 ;
        RECT 3.760 73.500 4.120 73.880 ;
        RECT 2.520 66.120 2.880 66.500 ;
        RECT 3.130 66.120 3.490 66.500 ;
        RECT 3.760 66.120 4.120 66.500 ;
        RECT 2.520 65.385 2.880 65.765 ;
        RECT 3.130 65.385 3.490 65.765 ;
        RECT 3.760 65.385 4.120 65.765 ;
        RECT 2.520 64.700 2.880 65.080 ;
        RECT 3.130 64.700 3.490 65.080 ;
        RECT 3.760 64.700 4.120 65.080 ;
        RECT 26.830 78.100 27.430 78.600 ;
        RECT 27.630 78.100 28.230 78.600 ;
        RECT 28.430 78.100 29.030 78.600 ;
        RECT 29.230 78.100 29.830 78.600 ;
        RECT 30.030 78.100 30.630 78.600 ;
        RECT 38.830 78.100 39.430 78.600 ;
        RECT 39.630 78.100 40.230 78.600 ;
        RECT 40.430 78.100 41.030 78.600 ;
        RECT 41.230 78.100 41.830 78.600 ;
        RECT 42.030 78.100 42.580 78.600 ;
        RECT 6.830 61.400 7.430 61.900 ;
        RECT 7.630 61.400 8.230 61.900 ;
        RECT 8.430 61.400 9.030 61.900 ;
        RECT 9.230 61.400 9.830 61.900 ;
        RECT 10.030 61.400 10.630 61.900 ;
        RECT 18.830 61.400 19.430 61.900 ;
        RECT 19.630 61.400 20.230 61.900 ;
        RECT 20.430 61.400 21.030 61.900 ;
        RECT 21.230 61.400 21.830 61.900 ;
        RECT 22.030 61.400 22.580 61.900 ;
        RECT 46.830 78.100 47.430 78.600 ;
        RECT 47.630 78.100 48.230 78.600 ;
        RECT 48.430 78.100 49.030 78.600 ;
        RECT 49.230 78.100 49.830 78.600 ;
        RECT 50.030 78.100 50.630 78.600 ;
        RECT 58.830 78.100 59.430 78.600 ;
        RECT 59.630 78.100 60.230 78.600 ;
        RECT 60.430 78.100 61.030 78.600 ;
        RECT 61.230 78.100 61.830 78.600 ;
        RECT 62.030 78.100 62.580 78.600 ;
        RECT 26.830 61.400 27.430 61.900 ;
        RECT 27.630 61.400 28.230 61.900 ;
        RECT 28.430 61.400 29.030 61.900 ;
        RECT 29.230 61.400 29.830 61.900 ;
        RECT 30.030 61.400 30.630 61.900 ;
        RECT 38.830 61.400 39.430 61.900 ;
        RECT 39.630 61.400 40.230 61.900 ;
        RECT 40.430 61.400 41.030 61.900 ;
        RECT 41.230 61.400 41.830 61.900 ;
        RECT 42.030 61.400 42.580 61.900 ;
        RECT 66.830 78.100 67.430 78.600 ;
        RECT 67.630 78.100 68.230 78.600 ;
        RECT 68.430 78.100 69.030 78.600 ;
        RECT 69.230 78.100 69.830 78.600 ;
        RECT 70.030 78.100 70.630 78.600 ;
        RECT 78.830 78.100 79.430 78.600 ;
        RECT 79.630 78.100 80.230 78.600 ;
        RECT 80.430 78.100 81.030 78.600 ;
        RECT 81.230 78.100 81.830 78.600 ;
        RECT 82.030 78.100 82.580 78.600 ;
        RECT 46.830 61.400 47.430 61.900 ;
        RECT 47.630 61.400 48.230 61.900 ;
        RECT 48.430 61.400 49.030 61.900 ;
        RECT 49.230 61.400 49.830 61.900 ;
        RECT 50.030 61.400 50.630 61.900 ;
        RECT 58.830 61.400 59.430 61.900 ;
        RECT 59.630 61.400 60.230 61.900 ;
        RECT 60.430 61.400 61.030 61.900 ;
        RECT 61.230 61.400 61.830 61.900 ;
        RECT 62.030 61.400 62.580 61.900 ;
        RECT 86.830 78.100 87.430 78.600 ;
        RECT 87.630 78.100 88.230 78.600 ;
        RECT 88.430 78.100 89.030 78.600 ;
        RECT 89.230 78.100 89.830 78.600 ;
        RECT 90.030 78.100 90.630 78.600 ;
        RECT 98.830 78.100 99.430 78.600 ;
        RECT 99.630 78.100 100.230 78.600 ;
        RECT 100.430 78.100 101.030 78.600 ;
        RECT 101.230 78.100 101.830 78.600 ;
        RECT 102.030 78.100 102.580 78.600 ;
        RECT 66.830 61.400 67.430 61.900 ;
        RECT 67.630 61.400 68.230 61.900 ;
        RECT 68.430 61.400 69.030 61.900 ;
        RECT 69.230 61.400 69.830 61.900 ;
        RECT 70.030 61.400 70.630 61.900 ;
        RECT 78.830 61.400 79.430 61.900 ;
        RECT 79.630 61.400 80.230 61.900 ;
        RECT 80.430 61.400 81.030 61.900 ;
        RECT 81.230 61.400 81.830 61.900 ;
        RECT 82.030 61.400 82.580 61.900 ;
        RECT 106.830 78.100 107.430 78.600 ;
        RECT 107.630 78.100 108.230 78.600 ;
        RECT 108.430 78.100 109.030 78.600 ;
        RECT 109.230 78.100 109.830 78.600 ;
        RECT 110.030 78.100 110.630 78.600 ;
        RECT 118.830 78.100 119.430 78.600 ;
        RECT 119.630 78.100 120.230 78.600 ;
        RECT 120.430 78.100 121.030 78.600 ;
        RECT 121.230 78.100 121.830 78.600 ;
        RECT 122.030 78.100 122.580 78.600 ;
        RECT 86.830 61.400 87.430 61.900 ;
        RECT 87.630 61.400 88.230 61.900 ;
        RECT 88.430 61.400 89.030 61.900 ;
        RECT 89.230 61.400 89.830 61.900 ;
        RECT 90.030 61.400 90.630 61.900 ;
        RECT 98.830 61.400 99.430 61.900 ;
        RECT 99.630 61.400 100.230 61.900 ;
        RECT 100.430 61.400 101.030 61.900 ;
        RECT 101.230 61.400 101.830 61.900 ;
        RECT 102.030 61.400 102.580 61.900 ;
        RECT 106.830 61.400 107.430 61.900 ;
        RECT 107.630 61.400 108.230 61.900 ;
        RECT 108.430 61.400 109.030 61.900 ;
        RECT 109.230 61.400 109.830 61.900 ;
        RECT 110.030 61.400 110.630 61.900 ;
        RECT 118.830 61.400 119.430 61.900 ;
        RECT 119.630 61.400 120.230 61.900 ;
        RECT 120.430 61.400 121.030 61.900 ;
        RECT 121.230 61.400 121.830 61.900 ;
        RECT 122.030 61.400 122.580 61.900 ;
        RECT 6.830 58.100 7.430 58.600 ;
        RECT 7.630 58.100 8.230 58.600 ;
        RECT 8.430 58.100 9.030 58.600 ;
        RECT 9.230 58.100 9.830 58.600 ;
        RECT 10.030 58.100 10.630 58.600 ;
        RECT 18.830 58.100 19.430 58.600 ;
        RECT 19.630 58.100 20.230 58.600 ;
        RECT 20.430 58.100 21.030 58.600 ;
        RECT 21.230 58.100 21.830 58.600 ;
        RECT 22.030 58.100 22.580 58.600 ;
        RECT 2.520 54.920 2.880 55.300 ;
        RECT 3.130 54.920 3.490 55.300 ;
        RECT 3.760 54.920 4.120 55.300 ;
        RECT 2.520 54.185 2.880 54.565 ;
        RECT 3.130 54.185 3.490 54.565 ;
        RECT 3.760 54.185 4.120 54.565 ;
        RECT 2.520 53.500 2.880 53.880 ;
        RECT 3.130 53.500 3.490 53.880 ;
        RECT 3.760 53.500 4.120 53.880 ;
        RECT 2.520 46.120 2.880 46.500 ;
        RECT 3.130 46.120 3.490 46.500 ;
        RECT 3.760 46.120 4.120 46.500 ;
        RECT 2.520 45.385 2.880 45.765 ;
        RECT 3.130 45.385 3.490 45.765 ;
        RECT 3.760 45.385 4.120 45.765 ;
        RECT 2.520 44.700 2.880 45.080 ;
        RECT 3.130 44.700 3.490 45.080 ;
        RECT 3.760 44.700 4.120 45.080 ;
        RECT 26.830 58.100 27.430 58.600 ;
        RECT 27.630 58.100 28.230 58.600 ;
        RECT 28.430 58.100 29.030 58.600 ;
        RECT 29.230 58.100 29.830 58.600 ;
        RECT 30.030 58.100 30.630 58.600 ;
        RECT 38.830 58.100 39.430 58.600 ;
        RECT 39.630 58.100 40.230 58.600 ;
        RECT 40.430 58.100 41.030 58.600 ;
        RECT 41.230 58.100 41.830 58.600 ;
        RECT 42.030 58.100 42.580 58.600 ;
        RECT 6.830 41.400 7.430 41.900 ;
        RECT 7.630 41.400 8.230 41.900 ;
        RECT 8.430 41.400 9.030 41.900 ;
        RECT 9.230 41.400 9.830 41.900 ;
        RECT 10.030 41.400 10.630 41.900 ;
        RECT 18.830 41.400 19.430 41.900 ;
        RECT 19.630 41.400 20.230 41.900 ;
        RECT 20.430 41.400 21.030 41.900 ;
        RECT 21.230 41.400 21.830 41.900 ;
        RECT 22.030 41.400 22.580 41.900 ;
        RECT 46.830 58.100 47.430 58.600 ;
        RECT 47.630 58.100 48.230 58.600 ;
        RECT 48.430 58.100 49.030 58.600 ;
        RECT 49.230 58.100 49.830 58.600 ;
        RECT 50.030 58.100 50.630 58.600 ;
        RECT 58.830 58.100 59.430 58.600 ;
        RECT 59.630 58.100 60.230 58.600 ;
        RECT 60.430 58.100 61.030 58.600 ;
        RECT 61.230 58.100 61.830 58.600 ;
        RECT 62.030 58.100 62.580 58.600 ;
        RECT 26.830 41.400 27.430 41.900 ;
        RECT 27.630 41.400 28.230 41.900 ;
        RECT 28.430 41.400 29.030 41.900 ;
        RECT 29.230 41.400 29.830 41.900 ;
        RECT 30.030 41.400 30.630 41.900 ;
        RECT 38.830 41.400 39.430 41.900 ;
        RECT 39.630 41.400 40.230 41.900 ;
        RECT 40.430 41.400 41.030 41.900 ;
        RECT 41.230 41.400 41.830 41.900 ;
        RECT 42.030 41.400 42.580 41.900 ;
        RECT 66.830 58.100 67.430 58.600 ;
        RECT 67.630 58.100 68.230 58.600 ;
        RECT 68.430 58.100 69.030 58.600 ;
        RECT 69.230 58.100 69.830 58.600 ;
        RECT 70.030 58.100 70.630 58.600 ;
        RECT 78.830 58.100 79.430 58.600 ;
        RECT 79.630 58.100 80.230 58.600 ;
        RECT 80.430 58.100 81.030 58.600 ;
        RECT 81.230 58.100 81.830 58.600 ;
        RECT 82.030 58.100 82.580 58.600 ;
        RECT 46.830 41.400 47.430 41.900 ;
        RECT 47.630 41.400 48.230 41.900 ;
        RECT 48.430 41.400 49.030 41.900 ;
        RECT 49.230 41.400 49.830 41.900 ;
        RECT 50.030 41.400 50.630 41.900 ;
        RECT 58.830 41.400 59.430 41.900 ;
        RECT 59.630 41.400 60.230 41.900 ;
        RECT 60.430 41.400 61.030 41.900 ;
        RECT 61.230 41.400 61.830 41.900 ;
        RECT 62.030 41.400 62.580 41.900 ;
        RECT 86.830 58.100 87.430 58.600 ;
        RECT 87.630 58.100 88.230 58.600 ;
        RECT 88.430 58.100 89.030 58.600 ;
        RECT 89.230 58.100 89.830 58.600 ;
        RECT 90.030 58.100 90.630 58.600 ;
        RECT 98.830 58.100 99.430 58.600 ;
        RECT 99.630 58.100 100.230 58.600 ;
        RECT 100.430 58.100 101.030 58.600 ;
        RECT 101.230 58.100 101.830 58.600 ;
        RECT 102.030 58.100 102.580 58.600 ;
        RECT 66.830 41.400 67.430 41.900 ;
        RECT 67.630 41.400 68.230 41.900 ;
        RECT 68.430 41.400 69.030 41.900 ;
        RECT 69.230 41.400 69.830 41.900 ;
        RECT 70.030 41.400 70.630 41.900 ;
        RECT 78.830 41.400 79.430 41.900 ;
        RECT 79.630 41.400 80.230 41.900 ;
        RECT 80.430 41.400 81.030 41.900 ;
        RECT 81.230 41.400 81.830 41.900 ;
        RECT 82.030 41.400 82.580 41.900 ;
        RECT 106.830 58.100 107.430 58.600 ;
        RECT 107.630 58.100 108.230 58.600 ;
        RECT 108.430 58.100 109.030 58.600 ;
        RECT 109.230 58.100 109.830 58.600 ;
        RECT 110.030 58.100 110.630 58.600 ;
        RECT 118.830 58.100 119.430 58.600 ;
        RECT 119.630 58.100 120.230 58.600 ;
        RECT 120.430 58.100 121.030 58.600 ;
        RECT 121.230 58.100 121.830 58.600 ;
        RECT 122.030 58.100 122.580 58.600 ;
        RECT 86.830 41.400 87.430 41.900 ;
        RECT 87.630 41.400 88.230 41.900 ;
        RECT 88.430 41.400 89.030 41.900 ;
        RECT 89.230 41.400 89.830 41.900 ;
        RECT 90.030 41.400 90.630 41.900 ;
        RECT 98.830 41.400 99.430 41.900 ;
        RECT 99.630 41.400 100.230 41.900 ;
        RECT 100.430 41.400 101.030 41.900 ;
        RECT 101.230 41.400 101.830 41.900 ;
        RECT 102.030 41.400 102.580 41.900 ;
        RECT 106.830 41.400 107.430 41.900 ;
        RECT 107.630 41.400 108.230 41.900 ;
        RECT 108.430 41.400 109.030 41.900 ;
        RECT 109.230 41.400 109.830 41.900 ;
        RECT 110.030 41.400 110.630 41.900 ;
        RECT 118.830 41.400 119.430 41.900 ;
        RECT 119.630 41.400 120.230 41.900 ;
        RECT 120.430 41.400 121.030 41.900 ;
        RECT 121.230 41.400 121.830 41.900 ;
        RECT 122.030 41.400 122.580 41.900 ;
        RECT 6.830 38.100 7.430 38.600 ;
        RECT 7.630 38.100 8.230 38.600 ;
        RECT 8.430 38.100 9.030 38.600 ;
        RECT 9.230 38.100 9.830 38.600 ;
        RECT 10.030 38.100 10.630 38.600 ;
        RECT 18.830 38.100 19.430 38.600 ;
        RECT 19.630 38.100 20.230 38.600 ;
        RECT 20.430 38.100 21.030 38.600 ;
        RECT 21.230 38.100 21.830 38.600 ;
        RECT 22.030 38.100 22.580 38.600 ;
        RECT 2.520 34.925 2.880 35.305 ;
        RECT 3.130 34.925 3.490 35.305 ;
        RECT 3.760 34.925 4.120 35.305 ;
        RECT 2.520 34.190 2.880 34.570 ;
        RECT 3.130 34.190 3.490 34.570 ;
        RECT 3.760 34.190 4.120 34.570 ;
        RECT 2.520 33.505 2.880 33.885 ;
        RECT 3.130 33.505 3.490 33.885 ;
        RECT 3.760 33.505 4.120 33.885 ;
        RECT 2.520 26.115 2.880 26.495 ;
        RECT 3.130 26.115 3.490 26.495 ;
        RECT 3.760 26.115 4.120 26.495 ;
        RECT 2.520 25.380 2.880 25.760 ;
        RECT 3.130 25.380 3.490 25.760 ;
        RECT 3.760 25.380 4.120 25.760 ;
        RECT 2.520 24.695 2.880 25.075 ;
        RECT 3.130 24.695 3.490 25.075 ;
        RECT 3.760 24.695 4.120 25.075 ;
        RECT 26.830 38.100 27.430 38.600 ;
        RECT 27.630 38.100 28.230 38.600 ;
        RECT 28.430 38.100 29.030 38.600 ;
        RECT 29.230 38.100 29.830 38.600 ;
        RECT 30.030 38.100 30.630 38.600 ;
        RECT 38.830 38.100 39.430 38.600 ;
        RECT 39.630 38.100 40.230 38.600 ;
        RECT 40.430 38.100 41.030 38.600 ;
        RECT 41.230 38.100 41.830 38.600 ;
        RECT 42.030 38.100 42.580 38.600 ;
        RECT 6.830 21.400 7.430 21.900 ;
        RECT 7.630 21.400 8.230 21.900 ;
        RECT 8.430 21.400 9.030 21.900 ;
        RECT 9.230 21.400 9.830 21.900 ;
        RECT 10.030 21.400 10.630 21.900 ;
        RECT 18.830 21.400 19.430 21.900 ;
        RECT 19.630 21.400 20.230 21.900 ;
        RECT 20.430 21.400 21.030 21.900 ;
        RECT 21.230 21.400 21.830 21.900 ;
        RECT 22.030 21.400 22.580 21.900 ;
        RECT 46.830 38.100 47.430 38.600 ;
        RECT 47.630 38.100 48.230 38.600 ;
        RECT 48.430 38.100 49.030 38.600 ;
        RECT 49.230 38.100 49.830 38.600 ;
        RECT 50.030 38.100 50.630 38.600 ;
        RECT 58.830 38.100 59.430 38.600 ;
        RECT 59.630 38.100 60.230 38.600 ;
        RECT 60.430 38.100 61.030 38.600 ;
        RECT 61.230 38.100 61.830 38.600 ;
        RECT 62.030 38.100 62.580 38.600 ;
        RECT 26.830 21.400 27.430 21.900 ;
        RECT 27.630 21.400 28.230 21.900 ;
        RECT 28.430 21.400 29.030 21.900 ;
        RECT 29.230 21.400 29.830 21.900 ;
        RECT 30.030 21.400 30.630 21.900 ;
        RECT 38.830 21.400 39.430 21.900 ;
        RECT 39.630 21.400 40.230 21.900 ;
        RECT 40.430 21.400 41.030 21.900 ;
        RECT 41.230 21.400 41.830 21.900 ;
        RECT 42.030 21.400 42.580 21.900 ;
        RECT 66.830 38.100 67.430 38.600 ;
        RECT 67.630 38.100 68.230 38.600 ;
        RECT 68.430 38.100 69.030 38.600 ;
        RECT 69.230 38.100 69.830 38.600 ;
        RECT 70.030 38.100 70.630 38.600 ;
        RECT 78.830 38.100 79.430 38.600 ;
        RECT 79.630 38.100 80.230 38.600 ;
        RECT 80.430 38.100 81.030 38.600 ;
        RECT 81.230 38.100 81.830 38.600 ;
        RECT 82.030 38.100 82.580 38.600 ;
        RECT 46.830 21.400 47.430 21.900 ;
        RECT 47.630 21.400 48.230 21.900 ;
        RECT 48.430 21.400 49.030 21.900 ;
        RECT 49.230 21.400 49.830 21.900 ;
        RECT 50.030 21.400 50.630 21.900 ;
        RECT 58.830 21.400 59.430 21.900 ;
        RECT 59.630 21.400 60.230 21.900 ;
        RECT 60.430 21.400 61.030 21.900 ;
        RECT 61.230 21.400 61.830 21.900 ;
        RECT 62.030 21.400 62.580 21.900 ;
        RECT 86.830 38.100 87.430 38.600 ;
        RECT 87.630 38.100 88.230 38.600 ;
        RECT 88.430 38.100 89.030 38.600 ;
        RECT 89.230 38.100 89.830 38.600 ;
        RECT 90.030 38.100 90.630 38.600 ;
        RECT 98.830 38.100 99.430 38.600 ;
        RECT 99.630 38.100 100.230 38.600 ;
        RECT 100.430 38.100 101.030 38.600 ;
        RECT 101.230 38.100 101.830 38.600 ;
        RECT 102.030 38.100 102.580 38.600 ;
        RECT 66.830 21.400 67.430 21.900 ;
        RECT 67.630 21.400 68.230 21.900 ;
        RECT 68.430 21.400 69.030 21.900 ;
        RECT 69.230 21.400 69.830 21.900 ;
        RECT 70.030 21.400 70.630 21.900 ;
        RECT 78.830 21.400 79.430 21.900 ;
        RECT 79.630 21.400 80.230 21.900 ;
        RECT 80.430 21.400 81.030 21.900 ;
        RECT 81.230 21.400 81.830 21.900 ;
        RECT 82.030 21.400 82.580 21.900 ;
        RECT 106.830 38.100 107.430 38.600 ;
        RECT 107.630 38.100 108.230 38.600 ;
        RECT 108.430 38.100 109.030 38.600 ;
        RECT 109.230 38.100 109.830 38.600 ;
        RECT 110.030 38.100 110.630 38.600 ;
        RECT 118.830 38.100 119.430 38.600 ;
        RECT 119.630 38.100 120.230 38.600 ;
        RECT 120.430 38.100 121.030 38.600 ;
        RECT 121.230 38.100 121.830 38.600 ;
        RECT 122.030 38.100 122.580 38.600 ;
        RECT 86.830 21.400 87.430 21.900 ;
        RECT 87.630 21.400 88.230 21.900 ;
        RECT 88.430 21.400 89.030 21.900 ;
        RECT 89.230 21.400 89.830 21.900 ;
        RECT 90.030 21.400 90.630 21.900 ;
        RECT 98.830 21.400 99.430 21.900 ;
        RECT 99.630 21.400 100.230 21.900 ;
        RECT 100.430 21.400 101.030 21.900 ;
        RECT 101.230 21.400 101.830 21.900 ;
        RECT 102.030 21.400 102.580 21.900 ;
        RECT 106.830 21.400 107.430 21.900 ;
        RECT 107.630 21.400 108.230 21.900 ;
        RECT 108.430 21.400 109.030 21.900 ;
        RECT 109.230 21.400 109.830 21.900 ;
        RECT 110.030 21.400 110.630 21.900 ;
        RECT 118.830 21.400 119.430 21.900 ;
        RECT 119.630 21.400 120.230 21.900 ;
        RECT 120.430 21.400 121.030 21.900 ;
        RECT 121.230 21.400 121.830 21.900 ;
        RECT 122.030 21.400 122.580 21.900 ;
        RECT 6.830 18.100 7.430 18.600 ;
        RECT 7.630 18.100 8.230 18.600 ;
        RECT 8.430 18.100 9.030 18.600 ;
        RECT 9.230 18.100 9.830 18.600 ;
        RECT 10.030 18.100 10.630 18.600 ;
        RECT 18.830 18.100 19.430 18.600 ;
        RECT 19.630 18.100 20.230 18.600 ;
        RECT 20.430 18.100 21.030 18.600 ;
        RECT 21.230 18.100 21.830 18.600 ;
        RECT 22.030 18.100 22.580 18.600 ;
        RECT 2.520 14.925 2.880 15.305 ;
        RECT 3.130 14.925 3.490 15.305 ;
        RECT 3.760 14.925 4.120 15.305 ;
        RECT 2.520 14.190 2.880 14.570 ;
        RECT 3.130 14.190 3.490 14.570 ;
        RECT 3.760 14.190 4.120 14.570 ;
        RECT 2.520 13.505 2.880 13.885 ;
        RECT 3.130 13.505 3.490 13.885 ;
        RECT 3.760 13.505 4.120 13.885 ;
        RECT 2.520 6.120 2.880 6.500 ;
        RECT 3.130 6.120 3.490 6.500 ;
        RECT 3.760 6.120 4.120 6.500 ;
        RECT 2.520 5.385 2.880 5.765 ;
        RECT 3.130 5.385 3.490 5.765 ;
        RECT 3.760 5.385 4.120 5.765 ;
        RECT 2.520 4.700 2.880 5.080 ;
        RECT 3.130 4.700 3.490 5.080 ;
        RECT 3.760 4.700 4.120 5.080 ;
        RECT 26.830 18.100 27.430 18.600 ;
        RECT 27.630 18.100 28.230 18.600 ;
        RECT 28.430 18.100 29.030 18.600 ;
        RECT 29.230 18.100 29.830 18.600 ;
        RECT 30.030 18.100 30.630 18.600 ;
        RECT 38.830 18.100 39.430 18.600 ;
        RECT 39.630 18.100 40.230 18.600 ;
        RECT 40.430 18.100 41.030 18.600 ;
        RECT 41.230 18.100 41.830 18.600 ;
        RECT 42.030 18.100 42.580 18.600 ;
        RECT 6.830 1.400 7.430 1.900 ;
        RECT 7.630 1.400 8.230 1.900 ;
        RECT 8.430 1.400 9.030 1.900 ;
        RECT 9.230 1.400 9.830 1.900 ;
        RECT 10.030 1.400 10.630 1.900 ;
        RECT 18.830 1.400 19.430 1.900 ;
        RECT 19.630 1.400 20.230 1.900 ;
        RECT 20.430 1.400 21.030 1.900 ;
        RECT 21.230 1.400 21.830 1.900 ;
        RECT 22.030 1.400 22.580 1.900 ;
        RECT 46.830 18.100 47.430 18.600 ;
        RECT 47.630 18.100 48.230 18.600 ;
        RECT 48.430 18.100 49.030 18.600 ;
        RECT 49.230 18.100 49.830 18.600 ;
        RECT 50.030 18.100 50.630 18.600 ;
        RECT 58.830 18.100 59.430 18.600 ;
        RECT 59.630 18.100 60.230 18.600 ;
        RECT 60.430 18.100 61.030 18.600 ;
        RECT 61.230 18.100 61.830 18.600 ;
        RECT 62.030 18.100 62.580 18.600 ;
        RECT 26.830 1.400 27.430 1.900 ;
        RECT 27.630 1.400 28.230 1.900 ;
        RECT 28.430 1.400 29.030 1.900 ;
        RECT 29.230 1.400 29.830 1.900 ;
        RECT 30.030 1.400 30.630 1.900 ;
        RECT 38.830 1.400 39.430 1.900 ;
        RECT 39.630 1.400 40.230 1.900 ;
        RECT 40.430 1.400 41.030 1.900 ;
        RECT 41.230 1.400 41.830 1.900 ;
        RECT 42.030 1.400 42.580 1.900 ;
        RECT 66.830 18.100 67.430 18.600 ;
        RECT 67.630 18.100 68.230 18.600 ;
        RECT 68.430 18.100 69.030 18.600 ;
        RECT 69.230 18.100 69.830 18.600 ;
        RECT 70.030 18.100 70.630 18.600 ;
        RECT 78.830 18.100 79.430 18.600 ;
        RECT 79.630 18.100 80.230 18.600 ;
        RECT 80.430 18.100 81.030 18.600 ;
        RECT 81.230 18.100 81.830 18.600 ;
        RECT 82.030 18.100 82.580 18.600 ;
        RECT 46.830 1.400 47.430 1.900 ;
        RECT 47.630 1.400 48.230 1.900 ;
        RECT 48.430 1.400 49.030 1.900 ;
        RECT 49.230 1.400 49.830 1.900 ;
        RECT 50.030 1.400 50.630 1.900 ;
        RECT 58.830 1.400 59.430 1.900 ;
        RECT 59.630 1.400 60.230 1.900 ;
        RECT 60.430 1.400 61.030 1.900 ;
        RECT 61.230 1.400 61.830 1.900 ;
        RECT 62.030 1.400 62.580 1.900 ;
        RECT 86.830 18.100 87.430 18.600 ;
        RECT 87.630 18.100 88.230 18.600 ;
        RECT 88.430 18.100 89.030 18.600 ;
        RECT 89.230 18.100 89.830 18.600 ;
        RECT 90.030 18.100 90.630 18.600 ;
        RECT 98.830 18.100 99.430 18.600 ;
        RECT 99.630 18.100 100.230 18.600 ;
        RECT 100.430 18.100 101.030 18.600 ;
        RECT 101.230 18.100 101.830 18.600 ;
        RECT 102.030 18.100 102.580 18.600 ;
        RECT 66.830 1.400 67.430 1.900 ;
        RECT 67.630 1.400 68.230 1.900 ;
        RECT 68.430 1.400 69.030 1.900 ;
        RECT 69.230 1.400 69.830 1.900 ;
        RECT 70.030 1.400 70.630 1.900 ;
        RECT 78.830 1.400 79.430 1.900 ;
        RECT 79.630 1.400 80.230 1.900 ;
        RECT 80.430 1.400 81.030 1.900 ;
        RECT 81.230 1.400 81.830 1.900 ;
        RECT 82.030 1.400 82.580 1.900 ;
        RECT 106.830 18.100 107.430 18.600 ;
        RECT 107.630 18.100 108.230 18.600 ;
        RECT 108.430 18.100 109.030 18.600 ;
        RECT 109.230 18.100 109.830 18.600 ;
        RECT 110.030 18.100 110.630 18.600 ;
        RECT 118.830 18.100 119.430 18.600 ;
        RECT 119.630 18.100 120.230 18.600 ;
        RECT 120.430 18.100 121.030 18.600 ;
        RECT 121.230 18.100 121.830 18.600 ;
        RECT 122.030 18.100 122.580 18.600 ;
        RECT 86.830 1.400 87.430 1.900 ;
        RECT 87.630 1.400 88.230 1.900 ;
        RECT 88.430 1.400 89.030 1.900 ;
        RECT 89.230 1.400 89.830 1.900 ;
        RECT 90.030 1.400 90.630 1.900 ;
        RECT 98.830 1.400 99.430 1.900 ;
        RECT 99.630 1.400 100.230 1.900 ;
        RECT 100.430 1.400 101.030 1.900 ;
        RECT 101.230 1.400 101.830 1.900 ;
        RECT 102.030 1.400 102.580 1.900 ;
        RECT 106.830 1.400 107.430 1.900 ;
        RECT 107.630 1.400 108.230 1.900 ;
        RECT 108.430 1.400 109.030 1.900 ;
        RECT 109.230 1.400 109.830 1.900 ;
        RECT 110.030 1.400 110.630 1.900 ;
        RECT 118.830 1.400 119.430 1.900 ;
        RECT 119.630 1.400 120.230 1.900 ;
        RECT 120.430 1.400 121.030 1.900 ;
        RECT 121.230 1.400 121.830 1.900 ;
        RECT 122.030 1.400 122.580 1.900 ;
      LAYER met1 ;
        RECT 4.730 339.850 9.130 340.000 ;
        RECT 20.330 339.850 29.130 340.000 ;
        RECT 40.330 339.850 49.130 340.000 ;
        RECT 60.330 339.850 69.130 340.000 ;
        RECT 80.330 339.850 89.130 340.000 ;
        RECT 100.330 339.850 109.130 340.000 ;
        RECT 4.730 338.950 10.730 339.850 ;
        RECT 20.330 339.800 30.730 339.850 ;
        RECT 40.330 339.800 50.730 339.850 ;
        RECT 60.330 339.800 70.730 339.850 ;
        RECT 80.330 339.800 90.730 339.850 ;
        RECT 100.330 339.800 110.730 339.850 ;
        RECT 120.330 339.800 124.730 340.000 ;
        RECT 4.730 338.800 9.130 338.950 ;
        RECT 4.730 337.385 5.930 338.800 ;
        RECT 9.280 338.650 10.730 338.950 ;
        RECT 2.315 336.110 5.930 337.385 ;
        RECT 4.730 335.600 5.930 336.110 ;
        RECT 6.530 338.450 10.730 338.650 ;
        RECT 18.730 338.950 30.730 339.800 ;
        RECT 18.730 338.900 29.130 338.950 ;
        RECT 18.730 338.650 20.180 338.900 ;
        RECT 20.330 338.800 29.130 338.900 ;
        RECT 18.730 338.450 22.930 338.650 ;
        RECT 6.530 338.300 14.080 338.450 ;
        RECT 15.430 338.300 22.930 338.450 ;
        RECT 6.530 338.000 10.730 338.300 ;
        RECT 2.315 333.250 4.315 335.545 ;
        RECT 6.530 335.150 6.680 338.000 ;
        RECT 7.130 330.450 7.280 338.000 ;
        RECT 7.730 330.450 7.880 338.000 ;
        RECT 8.330 330.450 8.480 338.000 ;
        RECT 8.930 330.450 9.080 338.000 ;
        RECT 9.530 330.450 9.680 338.000 ;
        RECT 10.130 337.850 10.730 338.000 ;
        RECT 18.730 338.000 22.930 338.300 ;
        RECT 18.730 337.850 19.330 338.000 ;
        RECT 10.130 337.700 14.080 337.850 ;
        RECT 15.380 337.700 19.330 337.850 ;
        RECT 10.130 337.250 10.730 337.700 ;
        RECT 18.730 337.250 19.330 337.700 ;
        RECT 10.130 337.100 14.080 337.250 ;
        RECT 15.380 337.100 19.330 337.250 ;
        RECT 10.130 336.650 10.730 337.100 ;
        RECT 18.730 336.650 19.330 337.100 ;
        RECT 10.130 336.500 14.080 336.650 ;
        RECT 15.380 336.500 19.330 336.650 ;
        RECT 10.130 336.050 10.730 336.500 ;
        RECT 18.730 336.050 19.330 336.500 ;
        RECT 10.130 335.900 14.080 336.050 ;
        RECT 15.380 335.900 19.330 336.050 ;
        RECT 10.130 335.450 10.730 335.900 ;
        RECT 18.730 335.450 19.330 335.900 ;
        RECT 10.130 335.300 14.080 335.450 ;
        RECT 15.380 335.300 19.330 335.450 ;
        RECT 10.130 334.850 10.730 335.300 ;
        RECT 18.730 334.850 19.330 335.300 ;
        RECT 10.130 334.700 14.080 334.850 ;
        RECT 15.380 334.700 19.330 334.850 ;
        RECT 10.130 334.250 10.730 334.700 ;
        RECT 18.730 334.250 19.330 334.700 ;
        RECT 10.130 334.100 14.080 334.250 ;
        RECT 15.380 334.100 19.330 334.250 ;
        RECT 10.130 333.650 10.730 334.100 ;
        RECT 18.730 333.650 19.330 334.100 ;
        RECT 10.130 333.500 14.080 333.650 ;
        RECT 15.380 333.500 19.330 333.650 ;
        RECT 10.130 333.050 10.730 333.500 ;
        RECT 18.730 333.050 19.330 333.500 ;
        RECT 10.130 332.900 14.080 333.050 ;
        RECT 15.380 332.900 19.330 333.050 ;
        RECT 10.130 332.450 10.730 332.900 ;
        RECT 18.730 332.450 19.330 332.900 ;
        RECT 10.130 332.300 14.080 332.450 ;
        RECT 15.380 332.300 19.330 332.450 ;
        RECT 10.130 331.850 10.730 332.300 ;
        RECT 18.730 331.850 19.330 332.300 ;
        RECT 10.130 331.700 14.080 331.850 ;
        RECT 15.380 331.700 19.330 331.850 ;
        RECT 10.130 331.250 10.730 331.700 ;
        RECT 18.730 331.250 19.330 331.700 ;
        RECT 10.130 331.100 14.080 331.250 ;
        RECT 15.380 331.100 19.330 331.250 ;
        RECT 10.130 330.650 10.730 331.100 ;
        RECT 18.730 330.650 19.330 331.100 ;
        RECT 10.130 330.450 14.080 330.650 ;
        RECT 15.380 330.450 19.330 330.650 ;
        RECT 19.780 330.450 19.930 338.000 ;
        RECT 20.380 330.450 20.530 338.000 ;
        RECT 20.980 330.450 21.130 338.000 ;
        RECT 21.580 330.450 21.730 338.000 ;
        RECT 22.180 330.450 22.330 338.000 ;
        RECT 22.780 335.150 22.930 338.000 ;
        RECT 23.530 335.600 25.930 338.800 ;
        RECT 29.280 338.650 30.730 338.950 ;
        RECT 26.530 338.450 30.730 338.650 ;
        RECT 38.730 338.950 50.730 339.800 ;
        RECT 38.730 338.900 49.130 338.950 ;
        RECT 38.730 338.650 40.180 338.900 ;
        RECT 40.330 338.800 49.130 338.900 ;
        RECT 38.730 338.450 42.930 338.650 ;
        RECT 26.530 338.300 34.080 338.450 ;
        RECT 35.430 338.300 42.930 338.450 ;
        RECT 26.530 338.000 30.730 338.300 ;
        RECT 26.530 335.150 26.680 338.000 ;
        RECT 27.130 330.450 27.280 338.000 ;
        RECT 27.730 330.450 27.880 338.000 ;
        RECT 28.330 330.450 28.480 338.000 ;
        RECT 28.930 330.450 29.080 338.000 ;
        RECT 29.530 330.450 29.680 338.000 ;
        RECT 30.130 337.850 30.730 338.000 ;
        RECT 38.730 338.000 42.930 338.300 ;
        RECT 38.730 337.850 39.330 338.000 ;
        RECT 30.130 337.700 34.080 337.850 ;
        RECT 35.380 337.700 39.330 337.850 ;
        RECT 30.130 337.250 30.730 337.700 ;
        RECT 38.730 337.250 39.330 337.700 ;
        RECT 30.130 337.100 34.080 337.250 ;
        RECT 35.380 337.100 39.330 337.250 ;
        RECT 30.130 336.650 30.730 337.100 ;
        RECT 38.730 336.650 39.330 337.100 ;
        RECT 30.130 336.500 34.080 336.650 ;
        RECT 35.380 336.500 39.330 336.650 ;
        RECT 30.130 336.050 30.730 336.500 ;
        RECT 38.730 336.050 39.330 336.500 ;
        RECT 30.130 335.900 34.080 336.050 ;
        RECT 35.380 335.900 39.330 336.050 ;
        RECT 30.130 335.450 30.730 335.900 ;
        RECT 38.730 335.450 39.330 335.900 ;
        RECT 30.130 335.300 34.080 335.450 ;
        RECT 35.380 335.300 39.330 335.450 ;
        RECT 30.130 334.850 30.730 335.300 ;
        RECT 38.730 334.850 39.330 335.300 ;
        RECT 30.130 334.700 34.080 334.850 ;
        RECT 35.380 334.700 39.330 334.850 ;
        RECT 30.130 334.250 30.730 334.700 ;
        RECT 38.730 334.250 39.330 334.700 ;
        RECT 30.130 334.100 34.080 334.250 ;
        RECT 35.380 334.100 39.330 334.250 ;
        RECT 30.130 333.650 30.730 334.100 ;
        RECT 38.730 333.650 39.330 334.100 ;
        RECT 30.130 333.500 34.080 333.650 ;
        RECT 35.380 333.500 39.330 333.650 ;
        RECT 30.130 333.050 30.730 333.500 ;
        RECT 38.730 333.050 39.330 333.500 ;
        RECT 30.130 332.900 34.080 333.050 ;
        RECT 35.380 332.900 39.330 333.050 ;
        RECT 30.130 332.450 30.730 332.900 ;
        RECT 38.730 332.450 39.330 332.900 ;
        RECT 30.130 332.300 34.080 332.450 ;
        RECT 35.380 332.300 39.330 332.450 ;
        RECT 30.130 331.850 30.730 332.300 ;
        RECT 38.730 331.850 39.330 332.300 ;
        RECT 30.130 331.700 34.080 331.850 ;
        RECT 35.380 331.700 39.330 331.850 ;
        RECT 30.130 331.250 30.730 331.700 ;
        RECT 38.730 331.250 39.330 331.700 ;
        RECT 30.130 331.100 34.080 331.250 ;
        RECT 35.380 331.100 39.330 331.250 ;
        RECT 30.130 330.650 30.730 331.100 ;
        RECT 38.730 330.650 39.330 331.100 ;
        RECT 30.130 330.450 34.080 330.650 ;
        RECT 35.380 330.450 39.330 330.650 ;
        RECT 39.780 330.450 39.930 338.000 ;
        RECT 40.380 330.450 40.530 338.000 ;
        RECT 40.980 330.450 41.130 338.000 ;
        RECT 41.580 330.450 41.730 338.000 ;
        RECT 42.180 330.450 42.330 338.000 ;
        RECT 42.780 335.150 42.930 338.000 ;
        RECT 43.530 335.600 45.930 338.800 ;
        RECT 49.280 338.650 50.730 338.950 ;
        RECT 46.530 338.450 50.730 338.650 ;
        RECT 58.730 338.950 70.730 339.800 ;
        RECT 58.730 338.900 69.130 338.950 ;
        RECT 58.730 338.650 60.180 338.900 ;
        RECT 60.330 338.800 69.130 338.900 ;
        RECT 58.730 338.450 62.930 338.650 ;
        RECT 46.530 338.300 54.080 338.450 ;
        RECT 55.430 338.300 62.930 338.450 ;
        RECT 46.530 338.000 50.730 338.300 ;
        RECT 46.530 335.150 46.680 338.000 ;
        RECT 47.130 330.450 47.280 338.000 ;
        RECT 47.730 330.450 47.880 338.000 ;
        RECT 48.330 330.450 48.480 338.000 ;
        RECT 48.930 330.450 49.080 338.000 ;
        RECT 49.530 330.450 49.680 338.000 ;
        RECT 50.130 337.850 50.730 338.000 ;
        RECT 58.730 338.000 62.930 338.300 ;
        RECT 58.730 337.850 59.330 338.000 ;
        RECT 50.130 337.700 54.080 337.850 ;
        RECT 55.380 337.700 59.330 337.850 ;
        RECT 50.130 337.250 50.730 337.700 ;
        RECT 58.730 337.250 59.330 337.700 ;
        RECT 50.130 337.100 54.080 337.250 ;
        RECT 55.380 337.100 59.330 337.250 ;
        RECT 50.130 336.650 50.730 337.100 ;
        RECT 58.730 336.650 59.330 337.100 ;
        RECT 50.130 336.500 54.080 336.650 ;
        RECT 55.380 336.500 59.330 336.650 ;
        RECT 50.130 336.050 50.730 336.500 ;
        RECT 58.730 336.050 59.330 336.500 ;
        RECT 50.130 335.900 54.080 336.050 ;
        RECT 55.380 335.900 59.330 336.050 ;
        RECT 50.130 335.450 50.730 335.900 ;
        RECT 58.730 335.450 59.330 335.900 ;
        RECT 50.130 335.300 54.080 335.450 ;
        RECT 55.380 335.300 59.330 335.450 ;
        RECT 50.130 334.850 50.730 335.300 ;
        RECT 58.730 334.850 59.330 335.300 ;
        RECT 50.130 334.700 54.080 334.850 ;
        RECT 55.380 334.700 59.330 334.850 ;
        RECT 50.130 334.250 50.730 334.700 ;
        RECT 58.730 334.250 59.330 334.700 ;
        RECT 50.130 334.100 54.080 334.250 ;
        RECT 55.380 334.100 59.330 334.250 ;
        RECT 50.130 333.650 50.730 334.100 ;
        RECT 58.730 333.650 59.330 334.100 ;
        RECT 50.130 333.500 54.080 333.650 ;
        RECT 55.380 333.500 59.330 333.650 ;
        RECT 50.130 333.050 50.730 333.500 ;
        RECT 58.730 333.050 59.330 333.500 ;
        RECT 50.130 332.900 54.080 333.050 ;
        RECT 55.380 332.900 59.330 333.050 ;
        RECT 50.130 332.450 50.730 332.900 ;
        RECT 58.730 332.450 59.330 332.900 ;
        RECT 50.130 332.300 54.080 332.450 ;
        RECT 55.380 332.300 59.330 332.450 ;
        RECT 50.130 331.850 50.730 332.300 ;
        RECT 58.730 331.850 59.330 332.300 ;
        RECT 50.130 331.700 54.080 331.850 ;
        RECT 55.380 331.700 59.330 331.850 ;
        RECT 50.130 331.250 50.730 331.700 ;
        RECT 58.730 331.250 59.330 331.700 ;
        RECT 50.130 331.100 54.080 331.250 ;
        RECT 55.380 331.100 59.330 331.250 ;
        RECT 50.130 330.650 50.730 331.100 ;
        RECT 58.730 330.650 59.330 331.100 ;
        RECT 50.130 330.450 54.080 330.650 ;
        RECT 55.380 330.450 59.330 330.650 ;
        RECT 59.780 330.450 59.930 338.000 ;
        RECT 60.380 330.450 60.530 338.000 ;
        RECT 60.980 330.450 61.130 338.000 ;
        RECT 61.580 330.450 61.730 338.000 ;
        RECT 62.180 330.450 62.330 338.000 ;
        RECT 62.780 335.150 62.930 338.000 ;
        RECT 63.530 335.600 65.930 338.800 ;
        RECT 69.280 338.650 70.730 338.950 ;
        RECT 66.530 338.450 70.730 338.650 ;
        RECT 78.730 338.950 90.730 339.800 ;
        RECT 78.730 338.900 89.130 338.950 ;
        RECT 78.730 338.650 80.180 338.900 ;
        RECT 80.330 338.800 89.130 338.900 ;
        RECT 78.730 338.450 82.930 338.650 ;
        RECT 66.530 338.300 74.080 338.450 ;
        RECT 75.430 338.300 82.930 338.450 ;
        RECT 66.530 338.000 70.730 338.300 ;
        RECT 66.530 335.150 66.680 338.000 ;
        RECT 67.130 330.450 67.280 338.000 ;
        RECT 67.730 330.450 67.880 338.000 ;
        RECT 68.330 330.450 68.480 338.000 ;
        RECT 68.930 330.450 69.080 338.000 ;
        RECT 69.530 330.450 69.680 338.000 ;
        RECT 70.130 337.850 70.730 338.000 ;
        RECT 78.730 338.000 82.930 338.300 ;
        RECT 78.730 337.850 79.330 338.000 ;
        RECT 70.130 337.700 74.080 337.850 ;
        RECT 75.380 337.700 79.330 337.850 ;
        RECT 70.130 337.250 70.730 337.700 ;
        RECT 78.730 337.250 79.330 337.700 ;
        RECT 70.130 337.100 74.080 337.250 ;
        RECT 75.380 337.100 79.330 337.250 ;
        RECT 70.130 336.650 70.730 337.100 ;
        RECT 78.730 336.650 79.330 337.100 ;
        RECT 70.130 336.500 74.080 336.650 ;
        RECT 75.380 336.500 79.330 336.650 ;
        RECT 70.130 336.050 70.730 336.500 ;
        RECT 78.730 336.050 79.330 336.500 ;
        RECT 70.130 335.900 74.080 336.050 ;
        RECT 75.380 335.900 79.330 336.050 ;
        RECT 70.130 335.450 70.730 335.900 ;
        RECT 78.730 335.450 79.330 335.900 ;
        RECT 70.130 335.300 74.080 335.450 ;
        RECT 75.380 335.300 79.330 335.450 ;
        RECT 70.130 334.850 70.730 335.300 ;
        RECT 78.730 334.850 79.330 335.300 ;
        RECT 70.130 334.700 74.080 334.850 ;
        RECT 75.380 334.700 79.330 334.850 ;
        RECT 70.130 334.250 70.730 334.700 ;
        RECT 78.730 334.250 79.330 334.700 ;
        RECT 70.130 334.100 74.080 334.250 ;
        RECT 75.380 334.100 79.330 334.250 ;
        RECT 70.130 333.650 70.730 334.100 ;
        RECT 78.730 333.650 79.330 334.100 ;
        RECT 70.130 333.500 74.080 333.650 ;
        RECT 75.380 333.500 79.330 333.650 ;
        RECT 70.130 333.050 70.730 333.500 ;
        RECT 78.730 333.050 79.330 333.500 ;
        RECT 70.130 332.900 74.080 333.050 ;
        RECT 75.380 332.900 79.330 333.050 ;
        RECT 70.130 332.450 70.730 332.900 ;
        RECT 78.730 332.450 79.330 332.900 ;
        RECT 70.130 332.300 74.080 332.450 ;
        RECT 75.380 332.300 79.330 332.450 ;
        RECT 70.130 331.850 70.730 332.300 ;
        RECT 78.730 331.850 79.330 332.300 ;
        RECT 70.130 331.700 74.080 331.850 ;
        RECT 75.380 331.700 79.330 331.850 ;
        RECT 70.130 331.250 70.730 331.700 ;
        RECT 78.730 331.250 79.330 331.700 ;
        RECT 70.130 331.100 74.080 331.250 ;
        RECT 75.380 331.100 79.330 331.250 ;
        RECT 70.130 330.650 70.730 331.100 ;
        RECT 78.730 330.650 79.330 331.100 ;
        RECT 70.130 330.450 74.080 330.650 ;
        RECT 75.380 330.450 79.330 330.650 ;
        RECT 79.780 330.450 79.930 338.000 ;
        RECT 80.380 330.450 80.530 338.000 ;
        RECT 80.980 330.450 81.130 338.000 ;
        RECT 81.580 330.450 81.730 338.000 ;
        RECT 82.180 330.450 82.330 338.000 ;
        RECT 82.780 335.150 82.930 338.000 ;
        RECT 83.530 335.600 85.930 338.800 ;
        RECT 89.280 338.650 90.730 338.950 ;
        RECT 86.530 338.450 90.730 338.650 ;
        RECT 98.730 338.950 110.730 339.800 ;
        RECT 98.730 338.900 109.130 338.950 ;
        RECT 98.730 338.650 100.180 338.900 ;
        RECT 100.330 338.800 109.130 338.900 ;
        RECT 98.730 338.450 102.930 338.650 ;
        RECT 86.530 338.300 94.080 338.450 ;
        RECT 95.430 338.300 102.930 338.450 ;
        RECT 86.530 338.000 90.730 338.300 ;
        RECT 86.530 335.150 86.680 338.000 ;
        RECT 87.130 330.450 87.280 338.000 ;
        RECT 87.730 330.450 87.880 338.000 ;
        RECT 88.330 330.450 88.480 338.000 ;
        RECT 88.930 330.450 89.080 338.000 ;
        RECT 89.530 330.450 89.680 338.000 ;
        RECT 90.130 337.850 90.730 338.000 ;
        RECT 98.730 338.000 102.930 338.300 ;
        RECT 98.730 337.850 99.330 338.000 ;
        RECT 90.130 337.700 94.080 337.850 ;
        RECT 95.380 337.700 99.330 337.850 ;
        RECT 90.130 337.250 90.730 337.700 ;
        RECT 98.730 337.250 99.330 337.700 ;
        RECT 90.130 337.100 94.080 337.250 ;
        RECT 95.380 337.100 99.330 337.250 ;
        RECT 90.130 336.650 90.730 337.100 ;
        RECT 98.730 336.650 99.330 337.100 ;
        RECT 90.130 336.500 94.080 336.650 ;
        RECT 95.380 336.500 99.330 336.650 ;
        RECT 90.130 336.050 90.730 336.500 ;
        RECT 98.730 336.050 99.330 336.500 ;
        RECT 90.130 335.900 94.080 336.050 ;
        RECT 95.380 335.900 99.330 336.050 ;
        RECT 90.130 335.450 90.730 335.900 ;
        RECT 98.730 335.450 99.330 335.900 ;
        RECT 90.130 335.300 94.080 335.450 ;
        RECT 95.380 335.300 99.330 335.450 ;
        RECT 90.130 334.850 90.730 335.300 ;
        RECT 98.730 334.850 99.330 335.300 ;
        RECT 90.130 334.700 94.080 334.850 ;
        RECT 95.380 334.700 99.330 334.850 ;
        RECT 90.130 334.250 90.730 334.700 ;
        RECT 98.730 334.250 99.330 334.700 ;
        RECT 90.130 334.100 94.080 334.250 ;
        RECT 95.380 334.100 99.330 334.250 ;
        RECT 90.130 333.650 90.730 334.100 ;
        RECT 98.730 333.650 99.330 334.100 ;
        RECT 90.130 333.500 94.080 333.650 ;
        RECT 95.380 333.500 99.330 333.650 ;
        RECT 90.130 333.050 90.730 333.500 ;
        RECT 98.730 333.050 99.330 333.500 ;
        RECT 90.130 332.900 94.080 333.050 ;
        RECT 95.380 332.900 99.330 333.050 ;
        RECT 90.130 332.450 90.730 332.900 ;
        RECT 98.730 332.450 99.330 332.900 ;
        RECT 90.130 332.300 94.080 332.450 ;
        RECT 95.380 332.300 99.330 332.450 ;
        RECT 90.130 331.850 90.730 332.300 ;
        RECT 98.730 331.850 99.330 332.300 ;
        RECT 90.130 331.700 94.080 331.850 ;
        RECT 95.380 331.700 99.330 331.850 ;
        RECT 90.130 331.250 90.730 331.700 ;
        RECT 98.730 331.250 99.330 331.700 ;
        RECT 90.130 331.100 94.080 331.250 ;
        RECT 95.380 331.100 99.330 331.250 ;
        RECT 90.130 330.650 90.730 331.100 ;
        RECT 98.730 330.650 99.330 331.100 ;
        RECT 90.130 330.450 94.080 330.650 ;
        RECT 95.380 330.450 99.330 330.650 ;
        RECT 99.780 330.450 99.930 338.000 ;
        RECT 100.380 330.450 100.530 338.000 ;
        RECT 100.980 330.450 101.130 338.000 ;
        RECT 101.580 330.450 101.730 338.000 ;
        RECT 102.180 330.450 102.330 338.000 ;
        RECT 102.780 335.150 102.930 338.000 ;
        RECT 103.530 335.600 105.930 338.800 ;
        RECT 109.280 338.650 110.730 338.950 ;
        RECT 106.530 338.450 110.730 338.650 ;
        RECT 118.730 338.900 124.730 339.800 ;
        RECT 118.730 338.650 120.180 338.900 ;
        RECT 120.330 338.800 124.730 338.900 ;
        RECT 118.730 338.450 122.930 338.650 ;
        RECT 106.530 338.300 114.080 338.450 ;
        RECT 115.430 338.300 122.930 338.450 ;
        RECT 106.530 338.000 110.730 338.300 ;
        RECT 106.530 335.150 106.680 338.000 ;
        RECT 107.130 330.450 107.280 338.000 ;
        RECT 107.730 330.450 107.880 338.000 ;
        RECT 108.330 330.450 108.480 338.000 ;
        RECT 108.930 330.450 109.080 338.000 ;
        RECT 109.530 330.450 109.680 338.000 ;
        RECT 110.130 337.850 110.730 338.000 ;
        RECT 118.730 338.000 122.930 338.300 ;
        RECT 118.730 337.850 119.330 338.000 ;
        RECT 110.130 337.700 114.080 337.850 ;
        RECT 115.380 337.700 119.330 337.850 ;
        RECT 110.130 337.250 110.730 337.700 ;
        RECT 118.730 337.250 119.330 337.700 ;
        RECT 110.130 337.100 114.080 337.250 ;
        RECT 115.380 337.100 119.330 337.250 ;
        RECT 110.130 336.650 110.730 337.100 ;
        RECT 118.730 336.650 119.330 337.100 ;
        RECT 110.130 336.500 114.080 336.650 ;
        RECT 115.380 336.500 119.330 336.650 ;
        RECT 110.130 336.050 110.730 336.500 ;
        RECT 118.730 336.050 119.330 336.500 ;
        RECT 110.130 335.900 114.080 336.050 ;
        RECT 115.380 335.900 119.330 336.050 ;
        RECT 110.130 335.450 110.730 335.900 ;
        RECT 118.730 335.450 119.330 335.900 ;
        RECT 110.130 335.300 114.080 335.450 ;
        RECT 115.380 335.300 119.330 335.450 ;
        RECT 110.130 334.850 110.730 335.300 ;
        RECT 118.730 334.850 119.330 335.300 ;
        RECT 110.130 334.700 114.080 334.850 ;
        RECT 115.380 334.700 119.330 334.850 ;
        RECT 110.130 334.250 110.730 334.700 ;
        RECT 118.730 334.250 119.330 334.700 ;
        RECT 110.130 334.100 114.080 334.250 ;
        RECT 115.380 334.100 119.330 334.250 ;
        RECT 110.130 333.650 110.730 334.100 ;
        RECT 118.730 333.650 119.330 334.100 ;
        RECT 110.130 333.500 114.080 333.650 ;
        RECT 115.380 333.500 119.330 333.650 ;
        RECT 110.130 333.050 110.730 333.500 ;
        RECT 118.730 333.050 119.330 333.500 ;
        RECT 110.130 332.900 114.080 333.050 ;
        RECT 115.380 332.900 119.330 333.050 ;
        RECT 110.130 332.450 110.730 332.900 ;
        RECT 118.730 332.450 119.330 332.900 ;
        RECT 110.130 332.300 114.080 332.450 ;
        RECT 115.380 332.300 119.330 332.450 ;
        RECT 110.130 331.850 110.730 332.300 ;
        RECT 118.730 331.850 119.330 332.300 ;
        RECT 110.130 331.700 114.080 331.850 ;
        RECT 115.380 331.700 119.330 331.850 ;
        RECT 110.130 331.250 110.730 331.700 ;
        RECT 118.730 331.250 119.330 331.700 ;
        RECT 110.130 331.100 114.080 331.250 ;
        RECT 115.380 331.100 119.330 331.250 ;
        RECT 110.130 330.650 110.730 331.100 ;
        RECT 118.730 330.650 119.330 331.100 ;
        RECT 110.130 330.450 114.080 330.650 ;
        RECT 115.380 330.450 119.330 330.650 ;
        RECT 119.780 330.450 119.930 338.000 ;
        RECT 120.380 330.450 120.530 338.000 ;
        RECT 120.980 330.450 121.130 338.000 ;
        RECT 121.580 330.450 121.730 338.000 ;
        RECT 122.180 330.450 122.330 338.000 ;
        RECT 122.780 335.150 122.930 338.000 ;
        RECT 123.530 337.585 124.730 338.800 ;
        RECT 123.530 336.310 127.130 337.585 ;
        RECT 123.530 335.600 124.730 336.310 ;
        RECT 2.315 324.450 4.315 326.745 ;
        RECT 4.730 324.020 5.930 324.400 ;
        RECT 2.315 322.745 5.930 324.020 ;
        RECT 4.730 321.200 5.930 322.745 ;
        RECT 6.530 322.000 6.680 324.900 ;
        RECT 7.130 322.000 7.280 329.550 ;
        RECT 7.730 322.000 7.880 329.550 ;
        RECT 8.330 322.000 8.480 329.550 ;
        RECT 8.930 322.000 9.080 329.550 ;
        RECT 9.530 322.000 9.680 329.550 ;
        RECT 10.130 329.350 14.080 329.550 ;
        RECT 15.380 329.350 19.330 329.550 ;
        RECT 10.130 328.900 10.730 329.350 ;
        RECT 18.730 328.900 19.330 329.350 ;
        RECT 10.130 328.750 14.080 328.900 ;
        RECT 15.380 328.750 19.330 328.900 ;
        RECT 10.130 328.300 10.730 328.750 ;
        RECT 18.730 328.300 19.330 328.750 ;
        RECT 10.130 328.150 14.080 328.300 ;
        RECT 15.380 328.150 19.330 328.300 ;
        RECT 10.130 327.700 10.730 328.150 ;
        RECT 18.730 327.700 19.330 328.150 ;
        RECT 10.130 327.550 14.080 327.700 ;
        RECT 15.380 327.550 19.330 327.700 ;
        RECT 10.130 327.100 10.730 327.550 ;
        RECT 18.730 327.100 19.330 327.550 ;
        RECT 10.130 326.950 14.080 327.100 ;
        RECT 15.380 326.950 19.330 327.100 ;
        RECT 10.130 326.500 10.730 326.950 ;
        RECT 18.730 326.500 19.330 326.950 ;
        RECT 10.130 326.350 14.080 326.500 ;
        RECT 15.380 326.350 19.330 326.500 ;
        RECT 10.130 325.900 10.730 326.350 ;
        RECT 18.730 325.900 19.330 326.350 ;
        RECT 10.130 325.750 14.080 325.900 ;
        RECT 15.380 325.750 19.330 325.900 ;
        RECT 10.130 325.300 10.730 325.750 ;
        RECT 18.730 325.300 19.330 325.750 ;
        RECT 10.130 325.150 14.080 325.300 ;
        RECT 15.380 325.150 19.330 325.300 ;
        RECT 10.130 324.700 10.730 325.150 ;
        RECT 18.730 324.700 19.330 325.150 ;
        RECT 10.130 324.550 14.080 324.700 ;
        RECT 15.380 324.550 19.330 324.700 ;
        RECT 10.130 324.100 10.730 324.550 ;
        RECT 18.730 324.100 19.330 324.550 ;
        RECT 10.130 323.950 14.080 324.100 ;
        RECT 15.380 323.950 19.330 324.100 ;
        RECT 10.130 323.500 10.730 323.950 ;
        RECT 18.730 323.500 19.330 323.950 ;
        RECT 10.130 323.350 14.080 323.500 ;
        RECT 15.380 323.350 19.330 323.500 ;
        RECT 10.130 322.900 10.730 323.350 ;
        RECT 18.730 322.900 19.330 323.350 ;
        RECT 10.130 322.750 14.080 322.900 ;
        RECT 15.380 322.750 19.330 322.900 ;
        RECT 10.130 322.300 10.730 322.750 ;
        RECT 18.730 322.300 19.330 322.750 ;
        RECT 10.130 322.150 14.080 322.300 ;
        RECT 15.380 322.150 19.330 322.300 ;
        RECT 10.130 322.000 10.730 322.150 ;
        RECT 6.530 321.700 10.730 322.000 ;
        RECT 18.730 322.000 19.330 322.150 ;
        RECT 19.780 322.000 19.930 329.550 ;
        RECT 20.380 322.000 20.530 329.550 ;
        RECT 20.980 322.000 21.130 329.550 ;
        RECT 21.580 322.000 21.730 329.550 ;
        RECT 22.180 322.000 22.330 329.550 ;
        RECT 22.780 322.000 22.930 324.900 ;
        RECT 18.730 321.700 22.930 322.000 ;
        RECT 6.530 321.550 14.080 321.700 ;
        RECT 15.380 321.550 22.930 321.700 ;
        RECT 6.530 321.350 10.730 321.550 ;
        RECT 4.730 321.050 9.130 321.200 ;
        RECT 9.280 321.050 10.730 321.350 ;
        RECT 4.730 320.150 10.730 321.050 ;
        RECT 18.730 321.350 22.930 321.550 ;
        RECT 18.730 321.050 20.180 321.350 ;
        RECT 23.530 321.200 25.930 324.400 ;
        RECT 26.530 322.000 26.680 324.900 ;
        RECT 27.130 322.000 27.280 329.550 ;
        RECT 27.730 322.000 27.880 329.550 ;
        RECT 28.330 322.000 28.480 329.550 ;
        RECT 28.930 322.000 29.080 329.550 ;
        RECT 29.530 322.000 29.680 329.550 ;
        RECT 30.130 329.350 34.080 329.550 ;
        RECT 35.380 329.350 39.330 329.550 ;
        RECT 30.130 328.900 30.730 329.350 ;
        RECT 38.730 328.900 39.330 329.350 ;
        RECT 30.130 328.750 34.080 328.900 ;
        RECT 35.380 328.750 39.330 328.900 ;
        RECT 30.130 328.300 30.730 328.750 ;
        RECT 38.730 328.300 39.330 328.750 ;
        RECT 30.130 328.150 34.080 328.300 ;
        RECT 35.380 328.150 39.330 328.300 ;
        RECT 30.130 327.700 30.730 328.150 ;
        RECT 38.730 327.700 39.330 328.150 ;
        RECT 30.130 327.550 34.080 327.700 ;
        RECT 35.380 327.550 39.330 327.700 ;
        RECT 30.130 327.100 30.730 327.550 ;
        RECT 38.730 327.100 39.330 327.550 ;
        RECT 30.130 326.950 34.080 327.100 ;
        RECT 35.380 326.950 39.330 327.100 ;
        RECT 30.130 326.500 30.730 326.950 ;
        RECT 38.730 326.500 39.330 326.950 ;
        RECT 30.130 326.350 34.080 326.500 ;
        RECT 35.380 326.350 39.330 326.500 ;
        RECT 30.130 325.900 30.730 326.350 ;
        RECT 38.730 325.900 39.330 326.350 ;
        RECT 30.130 325.750 34.080 325.900 ;
        RECT 35.380 325.750 39.330 325.900 ;
        RECT 30.130 325.300 30.730 325.750 ;
        RECT 38.730 325.300 39.330 325.750 ;
        RECT 30.130 325.150 34.080 325.300 ;
        RECT 35.380 325.150 39.330 325.300 ;
        RECT 30.130 324.700 30.730 325.150 ;
        RECT 38.730 324.700 39.330 325.150 ;
        RECT 30.130 324.550 34.080 324.700 ;
        RECT 35.380 324.550 39.330 324.700 ;
        RECT 30.130 324.100 30.730 324.550 ;
        RECT 38.730 324.100 39.330 324.550 ;
        RECT 30.130 323.950 34.080 324.100 ;
        RECT 35.380 323.950 39.330 324.100 ;
        RECT 30.130 323.500 30.730 323.950 ;
        RECT 38.730 323.500 39.330 323.950 ;
        RECT 30.130 323.350 34.080 323.500 ;
        RECT 35.380 323.350 39.330 323.500 ;
        RECT 30.130 322.900 30.730 323.350 ;
        RECT 38.730 322.900 39.330 323.350 ;
        RECT 30.130 322.750 34.080 322.900 ;
        RECT 35.380 322.750 39.330 322.900 ;
        RECT 30.130 322.300 30.730 322.750 ;
        RECT 38.730 322.300 39.330 322.750 ;
        RECT 30.130 322.150 34.080 322.300 ;
        RECT 35.380 322.150 39.330 322.300 ;
        RECT 30.130 322.000 30.730 322.150 ;
        RECT 26.530 321.700 30.730 322.000 ;
        RECT 38.730 322.000 39.330 322.150 ;
        RECT 39.780 322.000 39.930 329.550 ;
        RECT 40.380 322.000 40.530 329.550 ;
        RECT 40.980 322.000 41.130 329.550 ;
        RECT 41.580 322.000 41.730 329.550 ;
        RECT 42.180 322.000 42.330 329.550 ;
        RECT 42.780 322.000 42.930 324.900 ;
        RECT 38.730 321.700 42.930 322.000 ;
        RECT 26.530 321.550 34.080 321.700 ;
        RECT 35.380 321.550 42.930 321.700 ;
        RECT 26.530 321.350 30.730 321.550 ;
        RECT 20.330 321.050 29.130 321.200 ;
        RECT 29.280 321.050 30.730 321.350 ;
        RECT 18.730 320.150 30.730 321.050 ;
        RECT 38.730 321.350 42.930 321.550 ;
        RECT 38.730 321.050 40.180 321.350 ;
        RECT 43.530 321.200 45.930 324.400 ;
        RECT 46.530 322.000 46.680 324.900 ;
        RECT 47.130 322.000 47.280 329.550 ;
        RECT 47.730 322.000 47.880 329.550 ;
        RECT 48.330 322.000 48.480 329.550 ;
        RECT 48.930 322.000 49.080 329.550 ;
        RECT 49.530 322.000 49.680 329.550 ;
        RECT 50.130 329.350 54.080 329.550 ;
        RECT 55.380 329.350 59.330 329.550 ;
        RECT 50.130 328.900 50.730 329.350 ;
        RECT 58.730 328.900 59.330 329.350 ;
        RECT 50.130 328.750 54.080 328.900 ;
        RECT 55.380 328.750 59.330 328.900 ;
        RECT 50.130 328.300 50.730 328.750 ;
        RECT 58.730 328.300 59.330 328.750 ;
        RECT 50.130 328.150 54.080 328.300 ;
        RECT 55.380 328.150 59.330 328.300 ;
        RECT 50.130 327.700 50.730 328.150 ;
        RECT 58.730 327.700 59.330 328.150 ;
        RECT 50.130 327.550 54.080 327.700 ;
        RECT 55.380 327.550 59.330 327.700 ;
        RECT 50.130 327.100 50.730 327.550 ;
        RECT 58.730 327.100 59.330 327.550 ;
        RECT 50.130 326.950 54.080 327.100 ;
        RECT 55.380 326.950 59.330 327.100 ;
        RECT 50.130 326.500 50.730 326.950 ;
        RECT 58.730 326.500 59.330 326.950 ;
        RECT 50.130 326.350 54.080 326.500 ;
        RECT 55.380 326.350 59.330 326.500 ;
        RECT 50.130 325.900 50.730 326.350 ;
        RECT 58.730 325.900 59.330 326.350 ;
        RECT 50.130 325.750 54.080 325.900 ;
        RECT 55.380 325.750 59.330 325.900 ;
        RECT 50.130 325.300 50.730 325.750 ;
        RECT 58.730 325.300 59.330 325.750 ;
        RECT 50.130 325.150 54.080 325.300 ;
        RECT 55.380 325.150 59.330 325.300 ;
        RECT 50.130 324.700 50.730 325.150 ;
        RECT 58.730 324.700 59.330 325.150 ;
        RECT 50.130 324.550 54.080 324.700 ;
        RECT 55.380 324.550 59.330 324.700 ;
        RECT 50.130 324.100 50.730 324.550 ;
        RECT 58.730 324.100 59.330 324.550 ;
        RECT 50.130 323.950 54.080 324.100 ;
        RECT 55.380 323.950 59.330 324.100 ;
        RECT 50.130 323.500 50.730 323.950 ;
        RECT 58.730 323.500 59.330 323.950 ;
        RECT 50.130 323.350 54.080 323.500 ;
        RECT 55.380 323.350 59.330 323.500 ;
        RECT 50.130 322.900 50.730 323.350 ;
        RECT 58.730 322.900 59.330 323.350 ;
        RECT 50.130 322.750 54.080 322.900 ;
        RECT 55.380 322.750 59.330 322.900 ;
        RECT 50.130 322.300 50.730 322.750 ;
        RECT 58.730 322.300 59.330 322.750 ;
        RECT 50.130 322.150 54.080 322.300 ;
        RECT 55.380 322.150 59.330 322.300 ;
        RECT 50.130 322.000 50.730 322.150 ;
        RECT 46.530 321.700 50.730 322.000 ;
        RECT 58.730 322.000 59.330 322.150 ;
        RECT 59.780 322.000 59.930 329.550 ;
        RECT 60.380 322.000 60.530 329.550 ;
        RECT 60.980 322.000 61.130 329.550 ;
        RECT 61.580 322.000 61.730 329.550 ;
        RECT 62.180 322.000 62.330 329.550 ;
        RECT 62.780 322.000 62.930 324.900 ;
        RECT 58.730 321.700 62.930 322.000 ;
        RECT 46.530 321.550 54.080 321.700 ;
        RECT 55.380 321.550 62.930 321.700 ;
        RECT 46.530 321.350 50.730 321.550 ;
        RECT 40.330 321.050 49.130 321.200 ;
        RECT 49.280 321.050 50.730 321.350 ;
        RECT 38.730 320.150 50.730 321.050 ;
        RECT 58.730 321.350 62.930 321.550 ;
        RECT 58.730 321.050 60.180 321.350 ;
        RECT 63.530 321.200 65.930 324.400 ;
        RECT 66.530 322.000 66.680 324.900 ;
        RECT 67.130 322.000 67.280 329.550 ;
        RECT 67.730 322.000 67.880 329.550 ;
        RECT 68.330 322.000 68.480 329.550 ;
        RECT 68.930 322.000 69.080 329.550 ;
        RECT 69.530 322.000 69.680 329.550 ;
        RECT 70.130 329.350 74.080 329.550 ;
        RECT 75.380 329.350 79.330 329.550 ;
        RECT 70.130 328.900 70.730 329.350 ;
        RECT 78.730 328.900 79.330 329.350 ;
        RECT 70.130 328.750 74.080 328.900 ;
        RECT 75.380 328.750 79.330 328.900 ;
        RECT 70.130 328.300 70.730 328.750 ;
        RECT 78.730 328.300 79.330 328.750 ;
        RECT 70.130 328.150 74.080 328.300 ;
        RECT 75.380 328.150 79.330 328.300 ;
        RECT 70.130 327.700 70.730 328.150 ;
        RECT 78.730 327.700 79.330 328.150 ;
        RECT 70.130 327.550 74.080 327.700 ;
        RECT 75.380 327.550 79.330 327.700 ;
        RECT 70.130 327.100 70.730 327.550 ;
        RECT 78.730 327.100 79.330 327.550 ;
        RECT 70.130 326.950 74.080 327.100 ;
        RECT 75.380 326.950 79.330 327.100 ;
        RECT 70.130 326.500 70.730 326.950 ;
        RECT 78.730 326.500 79.330 326.950 ;
        RECT 70.130 326.350 74.080 326.500 ;
        RECT 75.380 326.350 79.330 326.500 ;
        RECT 70.130 325.900 70.730 326.350 ;
        RECT 78.730 325.900 79.330 326.350 ;
        RECT 70.130 325.750 74.080 325.900 ;
        RECT 75.380 325.750 79.330 325.900 ;
        RECT 70.130 325.300 70.730 325.750 ;
        RECT 78.730 325.300 79.330 325.750 ;
        RECT 70.130 325.150 74.080 325.300 ;
        RECT 75.380 325.150 79.330 325.300 ;
        RECT 70.130 324.700 70.730 325.150 ;
        RECT 78.730 324.700 79.330 325.150 ;
        RECT 70.130 324.550 74.080 324.700 ;
        RECT 75.380 324.550 79.330 324.700 ;
        RECT 70.130 324.100 70.730 324.550 ;
        RECT 78.730 324.100 79.330 324.550 ;
        RECT 70.130 323.950 74.080 324.100 ;
        RECT 75.380 323.950 79.330 324.100 ;
        RECT 70.130 323.500 70.730 323.950 ;
        RECT 78.730 323.500 79.330 323.950 ;
        RECT 70.130 323.350 74.080 323.500 ;
        RECT 75.380 323.350 79.330 323.500 ;
        RECT 70.130 322.900 70.730 323.350 ;
        RECT 78.730 322.900 79.330 323.350 ;
        RECT 70.130 322.750 74.080 322.900 ;
        RECT 75.380 322.750 79.330 322.900 ;
        RECT 70.130 322.300 70.730 322.750 ;
        RECT 78.730 322.300 79.330 322.750 ;
        RECT 70.130 322.150 74.080 322.300 ;
        RECT 75.380 322.150 79.330 322.300 ;
        RECT 70.130 322.000 70.730 322.150 ;
        RECT 66.530 321.700 70.730 322.000 ;
        RECT 78.730 322.000 79.330 322.150 ;
        RECT 79.780 322.000 79.930 329.550 ;
        RECT 80.380 322.000 80.530 329.550 ;
        RECT 80.980 322.000 81.130 329.550 ;
        RECT 81.580 322.000 81.730 329.550 ;
        RECT 82.180 322.000 82.330 329.550 ;
        RECT 82.780 322.000 82.930 324.900 ;
        RECT 78.730 321.700 82.930 322.000 ;
        RECT 66.530 321.550 74.080 321.700 ;
        RECT 75.380 321.550 82.930 321.700 ;
        RECT 66.530 321.350 70.730 321.550 ;
        RECT 60.330 321.050 69.130 321.200 ;
        RECT 69.280 321.050 70.730 321.350 ;
        RECT 58.730 320.150 70.730 321.050 ;
        RECT 78.730 321.350 82.930 321.550 ;
        RECT 78.730 321.050 80.180 321.350 ;
        RECT 83.530 321.200 85.930 324.400 ;
        RECT 86.530 322.000 86.680 324.900 ;
        RECT 87.130 322.000 87.280 329.550 ;
        RECT 87.730 322.000 87.880 329.550 ;
        RECT 88.330 322.000 88.480 329.550 ;
        RECT 88.930 322.000 89.080 329.550 ;
        RECT 89.530 322.000 89.680 329.550 ;
        RECT 90.130 329.350 94.080 329.550 ;
        RECT 95.380 329.350 99.330 329.550 ;
        RECT 90.130 328.900 90.730 329.350 ;
        RECT 98.730 328.900 99.330 329.350 ;
        RECT 90.130 328.750 94.080 328.900 ;
        RECT 95.380 328.750 99.330 328.900 ;
        RECT 90.130 328.300 90.730 328.750 ;
        RECT 98.730 328.300 99.330 328.750 ;
        RECT 90.130 328.150 94.080 328.300 ;
        RECT 95.380 328.150 99.330 328.300 ;
        RECT 90.130 327.700 90.730 328.150 ;
        RECT 98.730 327.700 99.330 328.150 ;
        RECT 90.130 327.550 94.080 327.700 ;
        RECT 95.380 327.550 99.330 327.700 ;
        RECT 90.130 327.100 90.730 327.550 ;
        RECT 98.730 327.100 99.330 327.550 ;
        RECT 90.130 326.950 94.080 327.100 ;
        RECT 95.380 326.950 99.330 327.100 ;
        RECT 90.130 326.500 90.730 326.950 ;
        RECT 98.730 326.500 99.330 326.950 ;
        RECT 90.130 326.350 94.080 326.500 ;
        RECT 95.380 326.350 99.330 326.500 ;
        RECT 90.130 325.900 90.730 326.350 ;
        RECT 98.730 325.900 99.330 326.350 ;
        RECT 90.130 325.750 94.080 325.900 ;
        RECT 95.380 325.750 99.330 325.900 ;
        RECT 90.130 325.300 90.730 325.750 ;
        RECT 98.730 325.300 99.330 325.750 ;
        RECT 90.130 325.150 94.080 325.300 ;
        RECT 95.380 325.150 99.330 325.300 ;
        RECT 90.130 324.700 90.730 325.150 ;
        RECT 98.730 324.700 99.330 325.150 ;
        RECT 90.130 324.550 94.080 324.700 ;
        RECT 95.380 324.550 99.330 324.700 ;
        RECT 90.130 324.100 90.730 324.550 ;
        RECT 98.730 324.100 99.330 324.550 ;
        RECT 90.130 323.950 94.080 324.100 ;
        RECT 95.380 323.950 99.330 324.100 ;
        RECT 90.130 323.500 90.730 323.950 ;
        RECT 98.730 323.500 99.330 323.950 ;
        RECT 90.130 323.350 94.080 323.500 ;
        RECT 95.380 323.350 99.330 323.500 ;
        RECT 90.130 322.900 90.730 323.350 ;
        RECT 98.730 322.900 99.330 323.350 ;
        RECT 90.130 322.750 94.080 322.900 ;
        RECT 95.380 322.750 99.330 322.900 ;
        RECT 90.130 322.300 90.730 322.750 ;
        RECT 98.730 322.300 99.330 322.750 ;
        RECT 90.130 322.150 94.080 322.300 ;
        RECT 95.380 322.150 99.330 322.300 ;
        RECT 90.130 322.000 90.730 322.150 ;
        RECT 86.530 321.700 90.730 322.000 ;
        RECT 98.730 322.000 99.330 322.150 ;
        RECT 99.780 322.000 99.930 329.550 ;
        RECT 100.380 322.000 100.530 329.550 ;
        RECT 100.980 322.000 101.130 329.550 ;
        RECT 101.580 322.000 101.730 329.550 ;
        RECT 102.180 322.000 102.330 329.550 ;
        RECT 102.780 322.000 102.930 324.900 ;
        RECT 98.730 321.700 102.930 322.000 ;
        RECT 86.530 321.550 94.080 321.700 ;
        RECT 95.380 321.550 102.930 321.700 ;
        RECT 86.530 321.350 90.730 321.550 ;
        RECT 80.330 321.050 89.130 321.200 ;
        RECT 89.280 321.050 90.730 321.350 ;
        RECT 78.730 320.150 90.730 321.050 ;
        RECT 98.730 321.350 102.930 321.550 ;
        RECT 98.730 321.050 100.180 321.350 ;
        RECT 103.530 321.200 105.930 324.400 ;
        RECT 106.530 322.000 106.680 324.900 ;
        RECT 107.130 322.000 107.280 329.550 ;
        RECT 107.730 322.000 107.880 329.550 ;
        RECT 108.330 322.000 108.480 329.550 ;
        RECT 108.930 322.000 109.080 329.550 ;
        RECT 109.530 322.000 109.680 329.550 ;
        RECT 110.130 329.350 114.080 329.550 ;
        RECT 115.380 329.350 119.330 329.550 ;
        RECT 110.130 328.900 110.730 329.350 ;
        RECT 118.730 328.900 119.330 329.350 ;
        RECT 110.130 328.750 114.080 328.900 ;
        RECT 115.380 328.750 119.330 328.900 ;
        RECT 110.130 328.300 110.730 328.750 ;
        RECT 118.730 328.300 119.330 328.750 ;
        RECT 110.130 328.150 114.080 328.300 ;
        RECT 115.380 328.150 119.330 328.300 ;
        RECT 110.130 327.700 110.730 328.150 ;
        RECT 118.730 327.700 119.330 328.150 ;
        RECT 110.130 327.550 114.080 327.700 ;
        RECT 115.380 327.550 119.330 327.700 ;
        RECT 110.130 327.100 110.730 327.550 ;
        RECT 118.730 327.100 119.330 327.550 ;
        RECT 110.130 326.950 114.080 327.100 ;
        RECT 115.380 326.950 119.330 327.100 ;
        RECT 110.130 326.500 110.730 326.950 ;
        RECT 118.730 326.500 119.330 326.950 ;
        RECT 110.130 326.350 114.080 326.500 ;
        RECT 115.380 326.350 119.330 326.500 ;
        RECT 110.130 325.900 110.730 326.350 ;
        RECT 118.730 325.900 119.330 326.350 ;
        RECT 110.130 325.750 114.080 325.900 ;
        RECT 115.380 325.750 119.330 325.900 ;
        RECT 110.130 325.300 110.730 325.750 ;
        RECT 118.730 325.300 119.330 325.750 ;
        RECT 110.130 325.150 114.080 325.300 ;
        RECT 115.380 325.150 119.330 325.300 ;
        RECT 110.130 324.700 110.730 325.150 ;
        RECT 118.730 324.700 119.330 325.150 ;
        RECT 110.130 324.550 114.080 324.700 ;
        RECT 115.380 324.550 119.330 324.700 ;
        RECT 110.130 324.100 110.730 324.550 ;
        RECT 118.730 324.100 119.330 324.550 ;
        RECT 110.130 323.950 114.080 324.100 ;
        RECT 115.380 323.950 119.330 324.100 ;
        RECT 110.130 323.500 110.730 323.950 ;
        RECT 118.730 323.500 119.330 323.950 ;
        RECT 110.130 323.350 114.080 323.500 ;
        RECT 115.380 323.350 119.330 323.500 ;
        RECT 110.130 322.900 110.730 323.350 ;
        RECT 118.730 322.900 119.330 323.350 ;
        RECT 110.130 322.750 114.080 322.900 ;
        RECT 115.380 322.750 119.330 322.900 ;
        RECT 110.130 322.300 110.730 322.750 ;
        RECT 118.730 322.300 119.330 322.750 ;
        RECT 110.130 322.150 114.080 322.300 ;
        RECT 115.380 322.150 119.330 322.300 ;
        RECT 110.130 322.000 110.730 322.150 ;
        RECT 106.530 321.700 110.730 322.000 ;
        RECT 118.730 322.000 119.330 322.150 ;
        RECT 119.780 322.000 119.930 329.550 ;
        RECT 120.380 322.000 120.530 329.550 ;
        RECT 120.980 322.000 121.130 329.550 ;
        RECT 121.580 322.000 121.730 329.550 ;
        RECT 122.180 322.000 122.330 329.550 ;
        RECT 122.780 322.000 122.930 324.900 ;
        RECT 118.730 321.700 122.930 322.000 ;
        RECT 106.530 321.550 114.080 321.700 ;
        RECT 115.380 321.550 122.930 321.700 ;
        RECT 106.530 321.350 110.730 321.550 ;
        RECT 100.330 321.050 109.130 321.200 ;
        RECT 109.280 321.050 110.730 321.350 ;
        RECT 98.730 320.150 110.730 321.050 ;
        RECT 118.730 321.350 122.930 321.550 ;
        RECT 123.530 323.600 124.730 324.400 ;
        RECT 123.530 322.325 127.140 323.600 ;
        RECT 118.730 321.050 120.180 321.350 ;
        RECT 123.530 321.200 124.730 322.325 ;
        RECT 120.330 321.050 124.730 321.200 ;
        RECT 118.730 320.150 124.730 321.050 ;
        RECT 4.730 319.850 9.130 320.150 ;
        RECT 20.330 319.850 29.130 320.150 ;
        RECT 40.330 319.850 49.130 320.150 ;
        RECT 60.330 319.850 69.130 320.150 ;
        RECT 80.330 319.850 89.130 320.150 ;
        RECT 100.330 319.850 109.130 320.150 ;
        RECT 4.730 318.950 10.730 319.850 ;
        RECT 20.330 319.800 30.730 319.850 ;
        RECT 40.330 319.800 50.730 319.850 ;
        RECT 60.330 319.800 70.730 319.850 ;
        RECT 80.330 319.800 90.730 319.850 ;
        RECT 100.330 319.800 110.730 319.850 ;
        RECT 120.330 319.800 124.730 320.150 ;
        RECT 4.730 318.800 9.130 318.950 ;
        RECT 4.730 317.375 5.930 318.800 ;
        RECT 9.280 318.650 10.730 318.950 ;
        RECT 2.315 316.100 5.930 317.375 ;
        RECT 4.730 315.600 5.930 316.100 ;
        RECT 6.530 318.450 10.730 318.650 ;
        RECT 18.730 318.950 30.730 319.800 ;
        RECT 18.730 318.900 29.130 318.950 ;
        RECT 18.730 318.650 20.180 318.900 ;
        RECT 20.330 318.800 29.130 318.900 ;
        RECT 18.730 318.450 22.930 318.650 ;
        RECT 6.530 318.300 14.080 318.450 ;
        RECT 15.430 318.300 22.930 318.450 ;
        RECT 6.530 318.000 10.730 318.300 ;
        RECT 2.315 313.250 4.315 315.545 ;
        RECT 6.530 315.150 6.680 318.000 ;
        RECT 7.130 310.450 7.280 318.000 ;
        RECT 7.730 310.450 7.880 318.000 ;
        RECT 8.330 310.450 8.480 318.000 ;
        RECT 8.930 310.450 9.080 318.000 ;
        RECT 9.530 310.450 9.680 318.000 ;
        RECT 10.130 317.850 10.730 318.000 ;
        RECT 18.730 318.000 22.930 318.300 ;
        RECT 18.730 317.850 19.330 318.000 ;
        RECT 10.130 317.700 14.080 317.850 ;
        RECT 15.380 317.700 19.330 317.850 ;
        RECT 10.130 317.250 10.730 317.700 ;
        RECT 18.730 317.250 19.330 317.700 ;
        RECT 10.130 317.100 14.080 317.250 ;
        RECT 15.380 317.100 19.330 317.250 ;
        RECT 10.130 316.650 10.730 317.100 ;
        RECT 18.730 316.650 19.330 317.100 ;
        RECT 10.130 316.500 14.080 316.650 ;
        RECT 15.380 316.500 19.330 316.650 ;
        RECT 10.130 316.050 10.730 316.500 ;
        RECT 18.730 316.050 19.330 316.500 ;
        RECT 10.130 315.900 14.080 316.050 ;
        RECT 15.380 315.900 19.330 316.050 ;
        RECT 10.130 315.450 10.730 315.900 ;
        RECT 18.730 315.450 19.330 315.900 ;
        RECT 10.130 315.300 14.080 315.450 ;
        RECT 15.380 315.300 19.330 315.450 ;
        RECT 10.130 314.850 10.730 315.300 ;
        RECT 18.730 314.850 19.330 315.300 ;
        RECT 10.130 314.700 14.080 314.850 ;
        RECT 15.380 314.700 19.330 314.850 ;
        RECT 10.130 314.250 10.730 314.700 ;
        RECT 18.730 314.250 19.330 314.700 ;
        RECT 10.130 314.100 14.080 314.250 ;
        RECT 15.380 314.100 19.330 314.250 ;
        RECT 10.130 313.650 10.730 314.100 ;
        RECT 18.730 313.650 19.330 314.100 ;
        RECT 10.130 313.500 14.080 313.650 ;
        RECT 15.380 313.500 19.330 313.650 ;
        RECT 10.130 313.050 10.730 313.500 ;
        RECT 18.730 313.050 19.330 313.500 ;
        RECT 10.130 312.900 14.080 313.050 ;
        RECT 15.380 312.900 19.330 313.050 ;
        RECT 10.130 312.450 10.730 312.900 ;
        RECT 18.730 312.450 19.330 312.900 ;
        RECT 10.130 312.300 14.080 312.450 ;
        RECT 15.380 312.300 19.330 312.450 ;
        RECT 10.130 311.850 10.730 312.300 ;
        RECT 18.730 311.850 19.330 312.300 ;
        RECT 10.130 311.700 14.080 311.850 ;
        RECT 15.380 311.700 19.330 311.850 ;
        RECT 10.130 311.250 10.730 311.700 ;
        RECT 18.730 311.250 19.330 311.700 ;
        RECT 10.130 311.100 14.080 311.250 ;
        RECT 15.380 311.100 19.330 311.250 ;
        RECT 10.130 310.650 10.730 311.100 ;
        RECT 18.730 310.650 19.330 311.100 ;
        RECT 10.130 310.450 14.080 310.650 ;
        RECT 15.380 310.450 19.330 310.650 ;
        RECT 19.780 310.450 19.930 318.000 ;
        RECT 20.380 310.450 20.530 318.000 ;
        RECT 20.980 310.450 21.130 318.000 ;
        RECT 21.580 310.450 21.730 318.000 ;
        RECT 22.180 310.450 22.330 318.000 ;
        RECT 22.780 315.150 22.930 318.000 ;
        RECT 23.530 315.600 25.930 318.800 ;
        RECT 29.280 318.650 30.730 318.950 ;
        RECT 26.530 318.450 30.730 318.650 ;
        RECT 38.730 318.950 50.730 319.800 ;
        RECT 38.730 318.900 49.130 318.950 ;
        RECT 38.730 318.650 40.180 318.900 ;
        RECT 40.330 318.800 49.130 318.900 ;
        RECT 38.730 318.450 42.930 318.650 ;
        RECT 26.530 318.300 34.080 318.450 ;
        RECT 35.430 318.300 42.930 318.450 ;
        RECT 26.530 318.000 30.730 318.300 ;
        RECT 26.530 315.150 26.680 318.000 ;
        RECT 27.130 310.450 27.280 318.000 ;
        RECT 27.730 310.450 27.880 318.000 ;
        RECT 28.330 310.450 28.480 318.000 ;
        RECT 28.930 310.450 29.080 318.000 ;
        RECT 29.530 310.450 29.680 318.000 ;
        RECT 30.130 317.850 30.730 318.000 ;
        RECT 38.730 318.000 42.930 318.300 ;
        RECT 38.730 317.850 39.330 318.000 ;
        RECT 30.130 317.700 34.080 317.850 ;
        RECT 35.380 317.700 39.330 317.850 ;
        RECT 30.130 317.250 30.730 317.700 ;
        RECT 38.730 317.250 39.330 317.700 ;
        RECT 30.130 317.100 34.080 317.250 ;
        RECT 35.380 317.100 39.330 317.250 ;
        RECT 30.130 316.650 30.730 317.100 ;
        RECT 38.730 316.650 39.330 317.100 ;
        RECT 30.130 316.500 34.080 316.650 ;
        RECT 35.380 316.500 39.330 316.650 ;
        RECT 30.130 316.050 30.730 316.500 ;
        RECT 38.730 316.050 39.330 316.500 ;
        RECT 30.130 315.900 34.080 316.050 ;
        RECT 35.380 315.900 39.330 316.050 ;
        RECT 30.130 315.450 30.730 315.900 ;
        RECT 38.730 315.450 39.330 315.900 ;
        RECT 30.130 315.300 34.080 315.450 ;
        RECT 35.380 315.300 39.330 315.450 ;
        RECT 30.130 314.850 30.730 315.300 ;
        RECT 38.730 314.850 39.330 315.300 ;
        RECT 30.130 314.700 34.080 314.850 ;
        RECT 35.380 314.700 39.330 314.850 ;
        RECT 30.130 314.250 30.730 314.700 ;
        RECT 38.730 314.250 39.330 314.700 ;
        RECT 30.130 314.100 34.080 314.250 ;
        RECT 35.380 314.100 39.330 314.250 ;
        RECT 30.130 313.650 30.730 314.100 ;
        RECT 38.730 313.650 39.330 314.100 ;
        RECT 30.130 313.500 34.080 313.650 ;
        RECT 35.380 313.500 39.330 313.650 ;
        RECT 30.130 313.050 30.730 313.500 ;
        RECT 38.730 313.050 39.330 313.500 ;
        RECT 30.130 312.900 34.080 313.050 ;
        RECT 35.380 312.900 39.330 313.050 ;
        RECT 30.130 312.450 30.730 312.900 ;
        RECT 38.730 312.450 39.330 312.900 ;
        RECT 30.130 312.300 34.080 312.450 ;
        RECT 35.380 312.300 39.330 312.450 ;
        RECT 30.130 311.850 30.730 312.300 ;
        RECT 38.730 311.850 39.330 312.300 ;
        RECT 30.130 311.700 34.080 311.850 ;
        RECT 35.380 311.700 39.330 311.850 ;
        RECT 30.130 311.250 30.730 311.700 ;
        RECT 38.730 311.250 39.330 311.700 ;
        RECT 30.130 311.100 34.080 311.250 ;
        RECT 35.380 311.100 39.330 311.250 ;
        RECT 30.130 310.650 30.730 311.100 ;
        RECT 38.730 310.650 39.330 311.100 ;
        RECT 30.130 310.450 34.080 310.650 ;
        RECT 35.380 310.450 39.330 310.650 ;
        RECT 39.780 310.450 39.930 318.000 ;
        RECT 40.380 310.450 40.530 318.000 ;
        RECT 40.980 310.450 41.130 318.000 ;
        RECT 41.580 310.450 41.730 318.000 ;
        RECT 42.180 310.450 42.330 318.000 ;
        RECT 42.780 315.150 42.930 318.000 ;
        RECT 43.530 315.600 45.930 318.800 ;
        RECT 49.280 318.650 50.730 318.950 ;
        RECT 46.530 318.450 50.730 318.650 ;
        RECT 58.730 318.950 70.730 319.800 ;
        RECT 58.730 318.900 69.130 318.950 ;
        RECT 58.730 318.650 60.180 318.900 ;
        RECT 60.330 318.800 69.130 318.900 ;
        RECT 58.730 318.450 62.930 318.650 ;
        RECT 46.530 318.300 54.080 318.450 ;
        RECT 55.430 318.300 62.930 318.450 ;
        RECT 46.530 318.000 50.730 318.300 ;
        RECT 46.530 315.150 46.680 318.000 ;
        RECT 47.130 310.450 47.280 318.000 ;
        RECT 47.730 310.450 47.880 318.000 ;
        RECT 48.330 310.450 48.480 318.000 ;
        RECT 48.930 310.450 49.080 318.000 ;
        RECT 49.530 310.450 49.680 318.000 ;
        RECT 50.130 317.850 50.730 318.000 ;
        RECT 58.730 318.000 62.930 318.300 ;
        RECT 58.730 317.850 59.330 318.000 ;
        RECT 50.130 317.700 54.080 317.850 ;
        RECT 55.380 317.700 59.330 317.850 ;
        RECT 50.130 317.250 50.730 317.700 ;
        RECT 58.730 317.250 59.330 317.700 ;
        RECT 50.130 317.100 54.080 317.250 ;
        RECT 55.380 317.100 59.330 317.250 ;
        RECT 50.130 316.650 50.730 317.100 ;
        RECT 58.730 316.650 59.330 317.100 ;
        RECT 50.130 316.500 54.080 316.650 ;
        RECT 55.380 316.500 59.330 316.650 ;
        RECT 50.130 316.050 50.730 316.500 ;
        RECT 58.730 316.050 59.330 316.500 ;
        RECT 50.130 315.900 54.080 316.050 ;
        RECT 55.380 315.900 59.330 316.050 ;
        RECT 50.130 315.450 50.730 315.900 ;
        RECT 58.730 315.450 59.330 315.900 ;
        RECT 50.130 315.300 54.080 315.450 ;
        RECT 55.380 315.300 59.330 315.450 ;
        RECT 50.130 314.850 50.730 315.300 ;
        RECT 58.730 314.850 59.330 315.300 ;
        RECT 50.130 314.700 54.080 314.850 ;
        RECT 55.380 314.700 59.330 314.850 ;
        RECT 50.130 314.250 50.730 314.700 ;
        RECT 58.730 314.250 59.330 314.700 ;
        RECT 50.130 314.100 54.080 314.250 ;
        RECT 55.380 314.100 59.330 314.250 ;
        RECT 50.130 313.650 50.730 314.100 ;
        RECT 58.730 313.650 59.330 314.100 ;
        RECT 50.130 313.500 54.080 313.650 ;
        RECT 55.380 313.500 59.330 313.650 ;
        RECT 50.130 313.050 50.730 313.500 ;
        RECT 58.730 313.050 59.330 313.500 ;
        RECT 50.130 312.900 54.080 313.050 ;
        RECT 55.380 312.900 59.330 313.050 ;
        RECT 50.130 312.450 50.730 312.900 ;
        RECT 58.730 312.450 59.330 312.900 ;
        RECT 50.130 312.300 54.080 312.450 ;
        RECT 55.380 312.300 59.330 312.450 ;
        RECT 50.130 311.850 50.730 312.300 ;
        RECT 58.730 311.850 59.330 312.300 ;
        RECT 50.130 311.700 54.080 311.850 ;
        RECT 55.380 311.700 59.330 311.850 ;
        RECT 50.130 311.250 50.730 311.700 ;
        RECT 58.730 311.250 59.330 311.700 ;
        RECT 50.130 311.100 54.080 311.250 ;
        RECT 55.380 311.100 59.330 311.250 ;
        RECT 50.130 310.650 50.730 311.100 ;
        RECT 58.730 310.650 59.330 311.100 ;
        RECT 50.130 310.450 54.080 310.650 ;
        RECT 55.380 310.450 59.330 310.650 ;
        RECT 59.780 310.450 59.930 318.000 ;
        RECT 60.380 310.450 60.530 318.000 ;
        RECT 60.980 310.450 61.130 318.000 ;
        RECT 61.580 310.450 61.730 318.000 ;
        RECT 62.180 310.450 62.330 318.000 ;
        RECT 62.780 315.150 62.930 318.000 ;
        RECT 63.530 315.600 65.930 318.800 ;
        RECT 69.280 318.650 70.730 318.950 ;
        RECT 66.530 318.450 70.730 318.650 ;
        RECT 78.730 318.950 90.730 319.800 ;
        RECT 78.730 318.900 89.130 318.950 ;
        RECT 78.730 318.650 80.180 318.900 ;
        RECT 80.330 318.800 89.130 318.900 ;
        RECT 78.730 318.450 82.930 318.650 ;
        RECT 66.530 318.300 74.080 318.450 ;
        RECT 75.430 318.300 82.930 318.450 ;
        RECT 66.530 318.000 70.730 318.300 ;
        RECT 66.530 315.150 66.680 318.000 ;
        RECT 67.130 310.450 67.280 318.000 ;
        RECT 67.730 310.450 67.880 318.000 ;
        RECT 68.330 310.450 68.480 318.000 ;
        RECT 68.930 310.450 69.080 318.000 ;
        RECT 69.530 310.450 69.680 318.000 ;
        RECT 70.130 317.850 70.730 318.000 ;
        RECT 78.730 318.000 82.930 318.300 ;
        RECT 78.730 317.850 79.330 318.000 ;
        RECT 70.130 317.700 74.080 317.850 ;
        RECT 75.380 317.700 79.330 317.850 ;
        RECT 70.130 317.250 70.730 317.700 ;
        RECT 78.730 317.250 79.330 317.700 ;
        RECT 70.130 317.100 74.080 317.250 ;
        RECT 75.380 317.100 79.330 317.250 ;
        RECT 70.130 316.650 70.730 317.100 ;
        RECT 78.730 316.650 79.330 317.100 ;
        RECT 70.130 316.500 74.080 316.650 ;
        RECT 75.380 316.500 79.330 316.650 ;
        RECT 70.130 316.050 70.730 316.500 ;
        RECT 78.730 316.050 79.330 316.500 ;
        RECT 70.130 315.900 74.080 316.050 ;
        RECT 75.380 315.900 79.330 316.050 ;
        RECT 70.130 315.450 70.730 315.900 ;
        RECT 78.730 315.450 79.330 315.900 ;
        RECT 70.130 315.300 74.080 315.450 ;
        RECT 75.380 315.300 79.330 315.450 ;
        RECT 70.130 314.850 70.730 315.300 ;
        RECT 78.730 314.850 79.330 315.300 ;
        RECT 70.130 314.700 74.080 314.850 ;
        RECT 75.380 314.700 79.330 314.850 ;
        RECT 70.130 314.250 70.730 314.700 ;
        RECT 78.730 314.250 79.330 314.700 ;
        RECT 70.130 314.100 74.080 314.250 ;
        RECT 75.380 314.100 79.330 314.250 ;
        RECT 70.130 313.650 70.730 314.100 ;
        RECT 78.730 313.650 79.330 314.100 ;
        RECT 70.130 313.500 74.080 313.650 ;
        RECT 75.380 313.500 79.330 313.650 ;
        RECT 70.130 313.050 70.730 313.500 ;
        RECT 78.730 313.050 79.330 313.500 ;
        RECT 70.130 312.900 74.080 313.050 ;
        RECT 75.380 312.900 79.330 313.050 ;
        RECT 70.130 312.450 70.730 312.900 ;
        RECT 78.730 312.450 79.330 312.900 ;
        RECT 70.130 312.300 74.080 312.450 ;
        RECT 75.380 312.300 79.330 312.450 ;
        RECT 70.130 311.850 70.730 312.300 ;
        RECT 78.730 311.850 79.330 312.300 ;
        RECT 70.130 311.700 74.080 311.850 ;
        RECT 75.380 311.700 79.330 311.850 ;
        RECT 70.130 311.250 70.730 311.700 ;
        RECT 78.730 311.250 79.330 311.700 ;
        RECT 70.130 311.100 74.080 311.250 ;
        RECT 75.380 311.100 79.330 311.250 ;
        RECT 70.130 310.650 70.730 311.100 ;
        RECT 78.730 310.650 79.330 311.100 ;
        RECT 70.130 310.450 74.080 310.650 ;
        RECT 75.380 310.450 79.330 310.650 ;
        RECT 79.780 310.450 79.930 318.000 ;
        RECT 80.380 310.450 80.530 318.000 ;
        RECT 80.980 310.450 81.130 318.000 ;
        RECT 81.580 310.450 81.730 318.000 ;
        RECT 82.180 310.450 82.330 318.000 ;
        RECT 82.780 315.150 82.930 318.000 ;
        RECT 83.530 315.600 85.930 318.800 ;
        RECT 89.280 318.650 90.730 318.950 ;
        RECT 86.530 318.450 90.730 318.650 ;
        RECT 98.730 318.950 110.730 319.800 ;
        RECT 98.730 318.900 109.130 318.950 ;
        RECT 98.730 318.650 100.180 318.900 ;
        RECT 100.330 318.800 109.130 318.900 ;
        RECT 98.730 318.450 102.930 318.650 ;
        RECT 86.530 318.300 94.080 318.450 ;
        RECT 95.430 318.300 102.930 318.450 ;
        RECT 86.530 318.000 90.730 318.300 ;
        RECT 86.530 315.150 86.680 318.000 ;
        RECT 87.130 310.450 87.280 318.000 ;
        RECT 87.730 310.450 87.880 318.000 ;
        RECT 88.330 310.450 88.480 318.000 ;
        RECT 88.930 310.450 89.080 318.000 ;
        RECT 89.530 310.450 89.680 318.000 ;
        RECT 90.130 317.850 90.730 318.000 ;
        RECT 98.730 318.000 102.930 318.300 ;
        RECT 98.730 317.850 99.330 318.000 ;
        RECT 90.130 317.700 94.080 317.850 ;
        RECT 95.380 317.700 99.330 317.850 ;
        RECT 90.130 317.250 90.730 317.700 ;
        RECT 98.730 317.250 99.330 317.700 ;
        RECT 90.130 317.100 94.080 317.250 ;
        RECT 95.380 317.100 99.330 317.250 ;
        RECT 90.130 316.650 90.730 317.100 ;
        RECT 98.730 316.650 99.330 317.100 ;
        RECT 90.130 316.500 94.080 316.650 ;
        RECT 95.380 316.500 99.330 316.650 ;
        RECT 90.130 316.050 90.730 316.500 ;
        RECT 98.730 316.050 99.330 316.500 ;
        RECT 90.130 315.900 94.080 316.050 ;
        RECT 95.380 315.900 99.330 316.050 ;
        RECT 90.130 315.450 90.730 315.900 ;
        RECT 98.730 315.450 99.330 315.900 ;
        RECT 90.130 315.300 94.080 315.450 ;
        RECT 95.380 315.300 99.330 315.450 ;
        RECT 90.130 314.850 90.730 315.300 ;
        RECT 98.730 314.850 99.330 315.300 ;
        RECT 90.130 314.700 94.080 314.850 ;
        RECT 95.380 314.700 99.330 314.850 ;
        RECT 90.130 314.250 90.730 314.700 ;
        RECT 98.730 314.250 99.330 314.700 ;
        RECT 90.130 314.100 94.080 314.250 ;
        RECT 95.380 314.100 99.330 314.250 ;
        RECT 90.130 313.650 90.730 314.100 ;
        RECT 98.730 313.650 99.330 314.100 ;
        RECT 90.130 313.500 94.080 313.650 ;
        RECT 95.380 313.500 99.330 313.650 ;
        RECT 90.130 313.050 90.730 313.500 ;
        RECT 98.730 313.050 99.330 313.500 ;
        RECT 90.130 312.900 94.080 313.050 ;
        RECT 95.380 312.900 99.330 313.050 ;
        RECT 90.130 312.450 90.730 312.900 ;
        RECT 98.730 312.450 99.330 312.900 ;
        RECT 90.130 312.300 94.080 312.450 ;
        RECT 95.380 312.300 99.330 312.450 ;
        RECT 90.130 311.850 90.730 312.300 ;
        RECT 98.730 311.850 99.330 312.300 ;
        RECT 90.130 311.700 94.080 311.850 ;
        RECT 95.380 311.700 99.330 311.850 ;
        RECT 90.130 311.250 90.730 311.700 ;
        RECT 98.730 311.250 99.330 311.700 ;
        RECT 90.130 311.100 94.080 311.250 ;
        RECT 95.380 311.100 99.330 311.250 ;
        RECT 90.130 310.650 90.730 311.100 ;
        RECT 98.730 310.650 99.330 311.100 ;
        RECT 90.130 310.450 94.080 310.650 ;
        RECT 95.380 310.450 99.330 310.650 ;
        RECT 99.780 310.450 99.930 318.000 ;
        RECT 100.380 310.450 100.530 318.000 ;
        RECT 100.980 310.450 101.130 318.000 ;
        RECT 101.580 310.450 101.730 318.000 ;
        RECT 102.180 310.450 102.330 318.000 ;
        RECT 102.780 315.150 102.930 318.000 ;
        RECT 103.530 315.600 105.930 318.800 ;
        RECT 109.280 318.650 110.730 318.950 ;
        RECT 106.530 318.450 110.730 318.650 ;
        RECT 118.730 318.900 124.730 319.800 ;
        RECT 118.730 318.650 120.180 318.900 ;
        RECT 120.330 318.800 124.730 318.900 ;
        RECT 118.730 318.450 122.930 318.650 ;
        RECT 106.530 318.300 114.080 318.450 ;
        RECT 115.430 318.300 122.930 318.450 ;
        RECT 106.530 318.000 110.730 318.300 ;
        RECT 106.530 315.150 106.680 318.000 ;
        RECT 107.130 310.450 107.280 318.000 ;
        RECT 107.730 310.450 107.880 318.000 ;
        RECT 108.330 310.450 108.480 318.000 ;
        RECT 108.930 310.450 109.080 318.000 ;
        RECT 109.530 310.450 109.680 318.000 ;
        RECT 110.130 317.850 110.730 318.000 ;
        RECT 118.730 318.000 122.930 318.300 ;
        RECT 118.730 317.850 119.330 318.000 ;
        RECT 110.130 317.700 114.080 317.850 ;
        RECT 115.380 317.700 119.330 317.850 ;
        RECT 110.130 317.250 110.730 317.700 ;
        RECT 118.730 317.250 119.330 317.700 ;
        RECT 110.130 317.100 114.080 317.250 ;
        RECT 115.380 317.100 119.330 317.250 ;
        RECT 110.130 316.650 110.730 317.100 ;
        RECT 118.730 316.650 119.330 317.100 ;
        RECT 110.130 316.500 114.080 316.650 ;
        RECT 115.380 316.500 119.330 316.650 ;
        RECT 110.130 316.050 110.730 316.500 ;
        RECT 118.730 316.050 119.330 316.500 ;
        RECT 110.130 315.900 114.080 316.050 ;
        RECT 115.380 315.900 119.330 316.050 ;
        RECT 110.130 315.450 110.730 315.900 ;
        RECT 118.730 315.450 119.330 315.900 ;
        RECT 110.130 315.300 114.080 315.450 ;
        RECT 115.380 315.300 119.330 315.450 ;
        RECT 110.130 314.850 110.730 315.300 ;
        RECT 118.730 314.850 119.330 315.300 ;
        RECT 110.130 314.700 114.080 314.850 ;
        RECT 115.380 314.700 119.330 314.850 ;
        RECT 110.130 314.250 110.730 314.700 ;
        RECT 118.730 314.250 119.330 314.700 ;
        RECT 110.130 314.100 114.080 314.250 ;
        RECT 115.380 314.100 119.330 314.250 ;
        RECT 110.130 313.650 110.730 314.100 ;
        RECT 118.730 313.650 119.330 314.100 ;
        RECT 110.130 313.500 114.080 313.650 ;
        RECT 115.380 313.500 119.330 313.650 ;
        RECT 110.130 313.050 110.730 313.500 ;
        RECT 118.730 313.050 119.330 313.500 ;
        RECT 110.130 312.900 114.080 313.050 ;
        RECT 115.380 312.900 119.330 313.050 ;
        RECT 110.130 312.450 110.730 312.900 ;
        RECT 118.730 312.450 119.330 312.900 ;
        RECT 110.130 312.300 114.080 312.450 ;
        RECT 115.380 312.300 119.330 312.450 ;
        RECT 110.130 311.850 110.730 312.300 ;
        RECT 118.730 311.850 119.330 312.300 ;
        RECT 110.130 311.700 114.080 311.850 ;
        RECT 115.380 311.700 119.330 311.850 ;
        RECT 110.130 311.250 110.730 311.700 ;
        RECT 118.730 311.250 119.330 311.700 ;
        RECT 110.130 311.100 114.080 311.250 ;
        RECT 115.380 311.100 119.330 311.250 ;
        RECT 110.130 310.650 110.730 311.100 ;
        RECT 118.730 310.650 119.330 311.100 ;
        RECT 110.130 310.450 114.080 310.650 ;
        RECT 115.380 310.450 119.330 310.650 ;
        RECT 119.780 310.450 119.930 318.000 ;
        RECT 120.380 310.450 120.530 318.000 ;
        RECT 120.980 310.450 121.130 318.000 ;
        RECT 121.580 310.450 121.730 318.000 ;
        RECT 122.180 310.450 122.330 318.000 ;
        RECT 122.780 315.150 122.930 318.000 ;
        RECT 123.530 317.585 124.730 318.800 ;
        RECT 123.530 316.310 127.130 317.585 ;
        RECT 123.530 315.600 124.730 316.310 ;
        RECT 2.315 304.455 4.315 306.750 ;
        RECT 4.730 303.675 5.930 304.400 ;
        RECT 2.315 302.400 5.930 303.675 ;
        RECT 4.730 301.200 5.930 302.400 ;
        RECT 6.530 302.000 6.680 304.900 ;
        RECT 7.130 302.000 7.280 309.550 ;
        RECT 7.730 302.000 7.880 309.550 ;
        RECT 8.330 302.000 8.480 309.550 ;
        RECT 8.930 302.000 9.080 309.550 ;
        RECT 9.530 302.000 9.680 309.550 ;
        RECT 10.130 309.350 14.080 309.550 ;
        RECT 15.380 309.350 19.330 309.550 ;
        RECT 10.130 308.900 10.730 309.350 ;
        RECT 18.730 308.900 19.330 309.350 ;
        RECT 10.130 308.750 14.080 308.900 ;
        RECT 15.380 308.750 19.330 308.900 ;
        RECT 10.130 308.300 10.730 308.750 ;
        RECT 18.730 308.300 19.330 308.750 ;
        RECT 10.130 308.150 14.080 308.300 ;
        RECT 15.380 308.150 19.330 308.300 ;
        RECT 10.130 307.700 10.730 308.150 ;
        RECT 18.730 307.700 19.330 308.150 ;
        RECT 10.130 307.550 14.080 307.700 ;
        RECT 15.380 307.550 19.330 307.700 ;
        RECT 10.130 307.100 10.730 307.550 ;
        RECT 18.730 307.100 19.330 307.550 ;
        RECT 10.130 306.950 14.080 307.100 ;
        RECT 15.380 306.950 19.330 307.100 ;
        RECT 10.130 306.500 10.730 306.950 ;
        RECT 18.730 306.500 19.330 306.950 ;
        RECT 10.130 306.350 14.080 306.500 ;
        RECT 15.380 306.350 19.330 306.500 ;
        RECT 10.130 305.900 10.730 306.350 ;
        RECT 18.730 305.900 19.330 306.350 ;
        RECT 10.130 305.750 14.080 305.900 ;
        RECT 15.380 305.750 19.330 305.900 ;
        RECT 10.130 305.300 10.730 305.750 ;
        RECT 18.730 305.300 19.330 305.750 ;
        RECT 10.130 305.150 14.080 305.300 ;
        RECT 15.380 305.150 19.330 305.300 ;
        RECT 10.130 304.700 10.730 305.150 ;
        RECT 18.730 304.700 19.330 305.150 ;
        RECT 10.130 304.550 14.080 304.700 ;
        RECT 15.380 304.550 19.330 304.700 ;
        RECT 10.130 304.100 10.730 304.550 ;
        RECT 18.730 304.100 19.330 304.550 ;
        RECT 10.130 303.950 14.080 304.100 ;
        RECT 15.380 303.950 19.330 304.100 ;
        RECT 10.130 303.500 10.730 303.950 ;
        RECT 18.730 303.500 19.330 303.950 ;
        RECT 10.130 303.350 14.080 303.500 ;
        RECT 15.380 303.350 19.330 303.500 ;
        RECT 10.130 302.900 10.730 303.350 ;
        RECT 18.730 302.900 19.330 303.350 ;
        RECT 10.130 302.750 14.080 302.900 ;
        RECT 15.380 302.750 19.330 302.900 ;
        RECT 10.130 302.300 10.730 302.750 ;
        RECT 18.730 302.300 19.330 302.750 ;
        RECT 10.130 302.150 14.080 302.300 ;
        RECT 15.380 302.150 19.330 302.300 ;
        RECT 10.130 302.000 10.730 302.150 ;
        RECT 6.530 301.700 10.730 302.000 ;
        RECT 18.730 302.000 19.330 302.150 ;
        RECT 19.780 302.000 19.930 309.550 ;
        RECT 20.380 302.000 20.530 309.550 ;
        RECT 20.980 302.000 21.130 309.550 ;
        RECT 21.580 302.000 21.730 309.550 ;
        RECT 22.180 302.000 22.330 309.550 ;
        RECT 22.780 302.000 22.930 304.900 ;
        RECT 18.730 301.700 22.930 302.000 ;
        RECT 6.530 301.550 14.080 301.700 ;
        RECT 15.380 301.550 22.930 301.700 ;
        RECT 6.530 301.350 10.730 301.550 ;
        RECT 4.730 301.050 9.130 301.200 ;
        RECT 9.280 301.050 10.730 301.350 ;
        RECT 4.730 300.150 10.730 301.050 ;
        RECT 18.730 301.350 22.930 301.550 ;
        RECT 18.730 301.050 20.180 301.350 ;
        RECT 23.530 301.200 25.930 304.400 ;
        RECT 26.530 302.000 26.680 304.900 ;
        RECT 27.130 302.000 27.280 309.550 ;
        RECT 27.730 302.000 27.880 309.550 ;
        RECT 28.330 302.000 28.480 309.550 ;
        RECT 28.930 302.000 29.080 309.550 ;
        RECT 29.530 302.000 29.680 309.550 ;
        RECT 30.130 309.350 34.080 309.550 ;
        RECT 35.380 309.350 39.330 309.550 ;
        RECT 30.130 308.900 30.730 309.350 ;
        RECT 38.730 308.900 39.330 309.350 ;
        RECT 30.130 308.750 34.080 308.900 ;
        RECT 35.380 308.750 39.330 308.900 ;
        RECT 30.130 308.300 30.730 308.750 ;
        RECT 38.730 308.300 39.330 308.750 ;
        RECT 30.130 308.150 34.080 308.300 ;
        RECT 35.380 308.150 39.330 308.300 ;
        RECT 30.130 307.700 30.730 308.150 ;
        RECT 38.730 307.700 39.330 308.150 ;
        RECT 30.130 307.550 34.080 307.700 ;
        RECT 35.380 307.550 39.330 307.700 ;
        RECT 30.130 307.100 30.730 307.550 ;
        RECT 38.730 307.100 39.330 307.550 ;
        RECT 30.130 306.950 34.080 307.100 ;
        RECT 35.380 306.950 39.330 307.100 ;
        RECT 30.130 306.500 30.730 306.950 ;
        RECT 38.730 306.500 39.330 306.950 ;
        RECT 30.130 306.350 34.080 306.500 ;
        RECT 35.380 306.350 39.330 306.500 ;
        RECT 30.130 305.900 30.730 306.350 ;
        RECT 38.730 305.900 39.330 306.350 ;
        RECT 30.130 305.750 34.080 305.900 ;
        RECT 35.380 305.750 39.330 305.900 ;
        RECT 30.130 305.300 30.730 305.750 ;
        RECT 38.730 305.300 39.330 305.750 ;
        RECT 30.130 305.150 34.080 305.300 ;
        RECT 35.380 305.150 39.330 305.300 ;
        RECT 30.130 304.700 30.730 305.150 ;
        RECT 38.730 304.700 39.330 305.150 ;
        RECT 30.130 304.550 34.080 304.700 ;
        RECT 35.380 304.550 39.330 304.700 ;
        RECT 30.130 304.100 30.730 304.550 ;
        RECT 38.730 304.100 39.330 304.550 ;
        RECT 30.130 303.950 34.080 304.100 ;
        RECT 35.380 303.950 39.330 304.100 ;
        RECT 30.130 303.500 30.730 303.950 ;
        RECT 38.730 303.500 39.330 303.950 ;
        RECT 30.130 303.350 34.080 303.500 ;
        RECT 35.380 303.350 39.330 303.500 ;
        RECT 30.130 302.900 30.730 303.350 ;
        RECT 38.730 302.900 39.330 303.350 ;
        RECT 30.130 302.750 34.080 302.900 ;
        RECT 35.380 302.750 39.330 302.900 ;
        RECT 30.130 302.300 30.730 302.750 ;
        RECT 38.730 302.300 39.330 302.750 ;
        RECT 30.130 302.150 34.080 302.300 ;
        RECT 35.380 302.150 39.330 302.300 ;
        RECT 30.130 302.000 30.730 302.150 ;
        RECT 26.530 301.700 30.730 302.000 ;
        RECT 38.730 302.000 39.330 302.150 ;
        RECT 39.780 302.000 39.930 309.550 ;
        RECT 40.380 302.000 40.530 309.550 ;
        RECT 40.980 302.000 41.130 309.550 ;
        RECT 41.580 302.000 41.730 309.550 ;
        RECT 42.180 302.000 42.330 309.550 ;
        RECT 42.780 302.000 42.930 304.900 ;
        RECT 38.730 301.700 42.930 302.000 ;
        RECT 26.530 301.550 34.080 301.700 ;
        RECT 35.380 301.550 42.930 301.700 ;
        RECT 26.530 301.350 30.730 301.550 ;
        RECT 20.330 301.050 29.130 301.200 ;
        RECT 29.280 301.050 30.730 301.350 ;
        RECT 18.730 300.150 30.730 301.050 ;
        RECT 38.730 301.350 42.930 301.550 ;
        RECT 38.730 301.050 40.180 301.350 ;
        RECT 43.530 301.200 45.930 304.400 ;
        RECT 46.530 302.000 46.680 304.900 ;
        RECT 47.130 302.000 47.280 309.550 ;
        RECT 47.730 302.000 47.880 309.550 ;
        RECT 48.330 302.000 48.480 309.550 ;
        RECT 48.930 302.000 49.080 309.550 ;
        RECT 49.530 302.000 49.680 309.550 ;
        RECT 50.130 309.350 54.080 309.550 ;
        RECT 55.380 309.350 59.330 309.550 ;
        RECT 50.130 308.900 50.730 309.350 ;
        RECT 58.730 308.900 59.330 309.350 ;
        RECT 50.130 308.750 54.080 308.900 ;
        RECT 55.380 308.750 59.330 308.900 ;
        RECT 50.130 308.300 50.730 308.750 ;
        RECT 58.730 308.300 59.330 308.750 ;
        RECT 50.130 308.150 54.080 308.300 ;
        RECT 55.380 308.150 59.330 308.300 ;
        RECT 50.130 307.700 50.730 308.150 ;
        RECT 58.730 307.700 59.330 308.150 ;
        RECT 50.130 307.550 54.080 307.700 ;
        RECT 55.380 307.550 59.330 307.700 ;
        RECT 50.130 307.100 50.730 307.550 ;
        RECT 58.730 307.100 59.330 307.550 ;
        RECT 50.130 306.950 54.080 307.100 ;
        RECT 55.380 306.950 59.330 307.100 ;
        RECT 50.130 306.500 50.730 306.950 ;
        RECT 58.730 306.500 59.330 306.950 ;
        RECT 50.130 306.350 54.080 306.500 ;
        RECT 55.380 306.350 59.330 306.500 ;
        RECT 50.130 305.900 50.730 306.350 ;
        RECT 58.730 305.900 59.330 306.350 ;
        RECT 50.130 305.750 54.080 305.900 ;
        RECT 55.380 305.750 59.330 305.900 ;
        RECT 50.130 305.300 50.730 305.750 ;
        RECT 58.730 305.300 59.330 305.750 ;
        RECT 50.130 305.150 54.080 305.300 ;
        RECT 55.380 305.150 59.330 305.300 ;
        RECT 50.130 304.700 50.730 305.150 ;
        RECT 58.730 304.700 59.330 305.150 ;
        RECT 50.130 304.550 54.080 304.700 ;
        RECT 55.380 304.550 59.330 304.700 ;
        RECT 50.130 304.100 50.730 304.550 ;
        RECT 58.730 304.100 59.330 304.550 ;
        RECT 50.130 303.950 54.080 304.100 ;
        RECT 55.380 303.950 59.330 304.100 ;
        RECT 50.130 303.500 50.730 303.950 ;
        RECT 58.730 303.500 59.330 303.950 ;
        RECT 50.130 303.350 54.080 303.500 ;
        RECT 55.380 303.350 59.330 303.500 ;
        RECT 50.130 302.900 50.730 303.350 ;
        RECT 58.730 302.900 59.330 303.350 ;
        RECT 50.130 302.750 54.080 302.900 ;
        RECT 55.380 302.750 59.330 302.900 ;
        RECT 50.130 302.300 50.730 302.750 ;
        RECT 58.730 302.300 59.330 302.750 ;
        RECT 50.130 302.150 54.080 302.300 ;
        RECT 55.380 302.150 59.330 302.300 ;
        RECT 50.130 302.000 50.730 302.150 ;
        RECT 46.530 301.700 50.730 302.000 ;
        RECT 58.730 302.000 59.330 302.150 ;
        RECT 59.780 302.000 59.930 309.550 ;
        RECT 60.380 302.000 60.530 309.550 ;
        RECT 60.980 302.000 61.130 309.550 ;
        RECT 61.580 302.000 61.730 309.550 ;
        RECT 62.180 302.000 62.330 309.550 ;
        RECT 62.780 302.000 62.930 304.900 ;
        RECT 58.730 301.700 62.930 302.000 ;
        RECT 46.530 301.550 54.080 301.700 ;
        RECT 55.380 301.550 62.930 301.700 ;
        RECT 46.530 301.350 50.730 301.550 ;
        RECT 40.330 301.050 49.130 301.200 ;
        RECT 49.280 301.050 50.730 301.350 ;
        RECT 38.730 300.150 50.730 301.050 ;
        RECT 58.730 301.350 62.930 301.550 ;
        RECT 58.730 301.050 60.180 301.350 ;
        RECT 63.530 301.200 65.930 304.400 ;
        RECT 66.530 302.000 66.680 304.900 ;
        RECT 67.130 302.000 67.280 309.550 ;
        RECT 67.730 302.000 67.880 309.550 ;
        RECT 68.330 302.000 68.480 309.550 ;
        RECT 68.930 302.000 69.080 309.550 ;
        RECT 69.530 302.000 69.680 309.550 ;
        RECT 70.130 309.350 74.080 309.550 ;
        RECT 75.380 309.350 79.330 309.550 ;
        RECT 70.130 308.900 70.730 309.350 ;
        RECT 78.730 308.900 79.330 309.350 ;
        RECT 70.130 308.750 74.080 308.900 ;
        RECT 75.380 308.750 79.330 308.900 ;
        RECT 70.130 308.300 70.730 308.750 ;
        RECT 78.730 308.300 79.330 308.750 ;
        RECT 70.130 308.150 74.080 308.300 ;
        RECT 75.380 308.150 79.330 308.300 ;
        RECT 70.130 307.700 70.730 308.150 ;
        RECT 78.730 307.700 79.330 308.150 ;
        RECT 70.130 307.550 74.080 307.700 ;
        RECT 75.380 307.550 79.330 307.700 ;
        RECT 70.130 307.100 70.730 307.550 ;
        RECT 78.730 307.100 79.330 307.550 ;
        RECT 70.130 306.950 74.080 307.100 ;
        RECT 75.380 306.950 79.330 307.100 ;
        RECT 70.130 306.500 70.730 306.950 ;
        RECT 78.730 306.500 79.330 306.950 ;
        RECT 70.130 306.350 74.080 306.500 ;
        RECT 75.380 306.350 79.330 306.500 ;
        RECT 70.130 305.900 70.730 306.350 ;
        RECT 78.730 305.900 79.330 306.350 ;
        RECT 70.130 305.750 74.080 305.900 ;
        RECT 75.380 305.750 79.330 305.900 ;
        RECT 70.130 305.300 70.730 305.750 ;
        RECT 78.730 305.300 79.330 305.750 ;
        RECT 70.130 305.150 74.080 305.300 ;
        RECT 75.380 305.150 79.330 305.300 ;
        RECT 70.130 304.700 70.730 305.150 ;
        RECT 78.730 304.700 79.330 305.150 ;
        RECT 70.130 304.550 74.080 304.700 ;
        RECT 75.380 304.550 79.330 304.700 ;
        RECT 70.130 304.100 70.730 304.550 ;
        RECT 78.730 304.100 79.330 304.550 ;
        RECT 70.130 303.950 74.080 304.100 ;
        RECT 75.380 303.950 79.330 304.100 ;
        RECT 70.130 303.500 70.730 303.950 ;
        RECT 78.730 303.500 79.330 303.950 ;
        RECT 70.130 303.350 74.080 303.500 ;
        RECT 75.380 303.350 79.330 303.500 ;
        RECT 70.130 302.900 70.730 303.350 ;
        RECT 78.730 302.900 79.330 303.350 ;
        RECT 70.130 302.750 74.080 302.900 ;
        RECT 75.380 302.750 79.330 302.900 ;
        RECT 70.130 302.300 70.730 302.750 ;
        RECT 78.730 302.300 79.330 302.750 ;
        RECT 70.130 302.150 74.080 302.300 ;
        RECT 75.380 302.150 79.330 302.300 ;
        RECT 70.130 302.000 70.730 302.150 ;
        RECT 66.530 301.700 70.730 302.000 ;
        RECT 78.730 302.000 79.330 302.150 ;
        RECT 79.780 302.000 79.930 309.550 ;
        RECT 80.380 302.000 80.530 309.550 ;
        RECT 80.980 302.000 81.130 309.550 ;
        RECT 81.580 302.000 81.730 309.550 ;
        RECT 82.180 302.000 82.330 309.550 ;
        RECT 82.780 302.000 82.930 304.900 ;
        RECT 78.730 301.700 82.930 302.000 ;
        RECT 66.530 301.550 74.080 301.700 ;
        RECT 75.380 301.550 82.930 301.700 ;
        RECT 66.530 301.350 70.730 301.550 ;
        RECT 60.330 301.050 69.130 301.200 ;
        RECT 69.280 301.050 70.730 301.350 ;
        RECT 58.730 300.150 70.730 301.050 ;
        RECT 78.730 301.350 82.930 301.550 ;
        RECT 78.730 301.050 80.180 301.350 ;
        RECT 83.530 301.200 85.930 304.400 ;
        RECT 86.530 302.000 86.680 304.900 ;
        RECT 87.130 302.000 87.280 309.550 ;
        RECT 87.730 302.000 87.880 309.550 ;
        RECT 88.330 302.000 88.480 309.550 ;
        RECT 88.930 302.000 89.080 309.550 ;
        RECT 89.530 302.000 89.680 309.550 ;
        RECT 90.130 309.350 94.080 309.550 ;
        RECT 95.380 309.350 99.330 309.550 ;
        RECT 90.130 308.900 90.730 309.350 ;
        RECT 98.730 308.900 99.330 309.350 ;
        RECT 90.130 308.750 94.080 308.900 ;
        RECT 95.380 308.750 99.330 308.900 ;
        RECT 90.130 308.300 90.730 308.750 ;
        RECT 98.730 308.300 99.330 308.750 ;
        RECT 90.130 308.150 94.080 308.300 ;
        RECT 95.380 308.150 99.330 308.300 ;
        RECT 90.130 307.700 90.730 308.150 ;
        RECT 98.730 307.700 99.330 308.150 ;
        RECT 90.130 307.550 94.080 307.700 ;
        RECT 95.380 307.550 99.330 307.700 ;
        RECT 90.130 307.100 90.730 307.550 ;
        RECT 98.730 307.100 99.330 307.550 ;
        RECT 90.130 306.950 94.080 307.100 ;
        RECT 95.380 306.950 99.330 307.100 ;
        RECT 90.130 306.500 90.730 306.950 ;
        RECT 98.730 306.500 99.330 306.950 ;
        RECT 90.130 306.350 94.080 306.500 ;
        RECT 95.380 306.350 99.330 306.500 ;
        RECT 90.130 305.900 90.730 306.350 ;
        RECT 98.730 305.900 99.330 306.350 ;
        RECT 90.130 305.750 94.080 305.900 ;
        RECT 95.380 305.750 99.330 305.900 ;
        RECT 90.130 305.300 90.730 305.750 ;
        RECT 98.730 305.300 99.330 305.750 ;
        RECT 90.130 305.150 94.080 305.300 ;
        RECT 95.380 305.150 99.330 305.300 ;
        RECT 90.130 304.700 90.730 305.150 ;
        RECT 98.730 304.700 99.330 305.150 ;
        RECT 90.130 304.550 94.080 304.700 ;
        RECT 95.380 304.550 99.330 304.700 ;
        RECT 90.130 304.100 90.730 304.550 ;
        RECT 98.730 304.100 99.330 304.550 ;
        RECT 90.130 303.950 94.080 304.100 ;
        RECT 95.380 303.950 99.330 304.100 ;
        RECT 90.130 303.500 90.730 303.950 ;
        RECT 98.730 303.500 99.330 303.950 ;
        RECT 90.130 303.350 94.080 303.500 ;
        RECT 95.380 303.350 99.330 303.500 ;
        RECT 90.130 302.900 90.730 303.350 ;
        RECT 98.730 302.900 99.330 303.350 ;
        RECT 90.130 302.750 94.080 302.900 ;
        RECT 95.380 302.750 99.330 302.900 ;
        RECT 90.130 302.300 90.730 302.750 ;
        RECT 98.730 302.300 99.330 302.750 ;
        RECT 90.130 302.150 94.080 302.300 ;
        RECT 95.380 302.150 99.330 302.300 ;
        RECT 90.130 302.000 90.730 302.150 ;
        RECT 86.530 301.700 90.730 302.000 ;
        RECT 98.730 302.000 99.330 302.150 ;
        RECT 99.780 302.000 99.930 309.550 ;
        RECT 100.380 302.000 100.530 309.550 ;
        RECT 100.980 302.000 101.130 309.550 ;
        RECT 101.580 302.000 101.730 309.550 ;
        RECT 102.180 302.000 102.330 309.550 ;
        RECT 102.780 302.000 102.930 304.900 ;
        RECT 98.730 301.700 102.930 302.000 ;
        RECT 86.530 301.550 94.080 301.700 ;
        RECT 95.380 301.550 102.930 301.700 ;
        RECT 86.530 301.350 90.730 301.550 ;
        RECT 80.330 301.050 89.130 301.200 ;
        RECT 89.280 301.050 90.730 301.350 ;
        RECT 78.730 300.150 90.730 301.050 ;
        RECT 98.730 301.350 102.930 301.550 ;
        RECT 98.730 301.050 100.180 301.350 ;
        RECT 103.530 301.200 105.930 304.400 ;
        RECT 106.530 302.000 106.680 304.900 ;
        RECT 107.130 302.000 107.280 309.550 ;
        RECT 107.730 302.000 107.880 309.550 ;
        RECT 108.330 302.000 108.480 309.550 ;
        RECT 108.930 302.000 109.080 309.550 ;
        RECT 109.530 302.000 109.680 309.550 ;
        RECT 110.130 309.350 114.080 309.550 ;
        RECT 115.380 309.350 119.330 309.550 ;
        RECT 110.130 308.900 110.730 309.350 ;
        RECT 118.730 308.900 119.330 309.350 ;
        RECT 110.130 308.750 114.080 308.900 ;
        RECT 115.380 308.750 119.330 308.900 ;
        RECT 110.130 308.300 110.730 308.750 ;
        RECT 118.730 308.300 119.330 308.750 ;
        RECT 110.130 308.150 114.080 308.300 ;
        RECT 115.380 308.150 119.330 308.300 ;
        RECT 110.130 307.700 110.730 308.150 ;
        RECT 118.730 307.700 119.330 308.150 ;
        RECT 110.130 307.550 114.080 307.700 ;
        RECT 115.380 307.550 119.330 307.700 ;
        RECT 110.130 307.100 110.730 307.550 ;
        RECT 118.730 307.100 119.330 307.550 ;
        RECT 110.130 306.950 114.080 307.100 ;
        RECT 115.380 306.950 119.330 307.100 ;
        RECT 110.130 306.500 110.730 306.950 ;
        RECT 118.730 306.500 119.330 306.950 ;
        RECT 110.130 306.350 114.080 306.500 ;
        RECT 115.380 306.350 119.330 306.500 ;
        RECT 110.130 305.900 110.730 306.350 ;
        RECT 118.730 305.900 119.330 306.350 ;
        RECT 110.130 305.750 114.080 305.900 ;
        RECT 115.380 305.750 119.330 305.900 ;
        RECT 110.130 305.300 110.730 305.750 ;
        RECT 118.730 305.300 119.330 305.750 ;
        RECT 110.130 305.150 114.080 305.300 ;
        RECT 115.380 305.150 119.330 305.300 ;
        RECT 110.130 304.700 110.730 305.150 ;
        RECT 118.730 304.700 119.330 305.150 ;
        RECT 110.130 304.550 114.080 304.700 ;
        RECT 115.380 304.550 119.330 304.700 ;
        RECT 110.130 304.100 110.730 304.550 ;
        RECT 118.730 304.100 119.330 304.550 ;
        RECT 110.130 303.950 114.080 304.100 ;
        RECT 115.380 303.950 119.330 304.100 ;
        RECT 110.130 303.500 110.730 303.950 ;
        RECT 118.730 303.500 119.330 303.950 ;
        RECT 110.130 303.350 114.080 303.500 ;
        RECT 115.380 303.350 119.330 303.500 ;
        RECT 110.130 302.900 110.730 303.350 ;
        RECT 118.730 302.900 119.330 303.350 ;
        RECT 110.130 302.750 114.080 302.900 ;
        RECT 115.380 302.750 119.330 302.900 ;
        RECT 110.130 302.300 110.730 302.750 ;
        RECT 118.730 302.300 119.330 302.750 ;
        RECT 110.130 302.150 114.080 302.300 ;
        RECT 115.380 302.150 119.330 302.300 ;
        RECT 110.130 302.000 110.730 302.150 ;
        RECT 106.530 301.700 110.730 302.000 ;
        RECT 118.730 302.000 119.330 302.150 ;
        RECT 119.780 302.000 119.930 309.550 ;
        RECT 120.380 302.000 120.530 309.550 ;
        RECT 120.980 302.000 121.130 309.550 ;
        RECT 121.580 302.000 121.730 309.550 ;
        RECT 122.180 302.000 122.330 309.550 ;
        RECT 122.780 302.000 122.930 304.900 ;
        RECT 118.730 301.700 122.930 302.000 ;
        RECT 106.530 301.550 114.080 301.700 ;
        RECT 115.380 301.550 122.930 301.700 ;
        RECT 106.530 301.350 110.730 301.550 ;
        RECT 100.330 301.050 109.130 301.200 ;
        RECT 109.280 301.050 110.730 301.350 ;
        RECT 98.730 300.150 110.730 301.050 ;
        RECT 118.730 301.350 122.930 301.550 ;
        RECT 123.530 303.600 124.730 304.400 ;
        RECT 123.530 302.325 127.140 303.600 ;
        RECT 118.730 301.050 120.180 301.350 ;
        RECT 123.530 301.200 124.730 302.325 ;
        RECT 120.330 301.050 124.730 301.200 ;
        RECT 118.730 300.150 124.730 301.050 ;
        RECT 4.730 299.850 9.130 300.150 ;
        RECT 20.330 299.850 29.130 300.150 ;
        RECT 40.330 299.850 49.130 300.150 ;
        RECT 60.330 299.850 69.130 300.150 ;
        RECT 80.330 299.850 89.130 300.150 ;
        RECT 100.330 299.850 109.130 300.150 ;
        RECT 4.730 298.950 10.730 299.850 ;
        RECT 20.330 299.800 30.730 299.850 ;
        RECT 40.330 299.800 50.730 299.850 ;
        RECT 60.330 299.800 70.730 299.850 ;
        RECT 80.330 299.800 90.730 299.850 ;
        RECT 100.330 299.800 110.730 299.850 ;
        RECT 120.330 299.800 124.730 300.150 ;
        RECT 4.730 298.800 9.130 298.950 ;
        RECT 4.730 297.785 5.930 298.800 ;
        RECT 9.280 298.650 10.730 298.950 ;
        RECT 2.315 296.510 5.930 297.785 ;
        RECT 4.730 295.600 5.930 296.510 ;
        RECT 6.530 298.450 10.730 298.650 ;
        RECT 18.730 298.950 30.730 299.800 ;
        RECT 18.730 298.900 29.130 298.950 ;
        RECT 18.730 298.650 20.180 298.900 ;
        RECT 20.330 298.800 29.130 298.900 ;
        RECT 18.730 298.450 22.930 298.650 ;
        RECT 6.530 298.300 14.080 298.450 ;
        RECT 15.430 298.300 22.930 298.450 ;
        RECT 6.530 298.000 10.730 298.300 ;
        RECT 2.320 295.340 4.320 295.545 ;
        RECT 2.315 293.250 4.320 295.340 ;
        RECT 6.530 295.150 6.680 298.000 ;
        RECT 7.130 290.450 7.280 298.000 ;
        RECT 7.730 290.450 7.880 298.000 ;
        RECT 8.330 290.450 8.480 298.000 ;
        RECT 8.930 290.450 9.080 298.000 ;
        RECT 9.530 290.450 9.680 298.000 ;
        RECT 10.130 297.850 10.730 298.000 ;
        RECT 18.730 298.000 22.930 298.300 ;
        RECT 18.730 297.850 19.330 298.000 ;
        RECT 10.130 297.700 14.080 297.850 ;
        RECT 15.380 297.700 19.330 297.850 ;
        RECT 10.130 297.250 10.730 297.700 ;
        RECT 18.730 297.250 19.330 297.700 ;
        RECT 10.130 297.100 14.080 297.250 ;
        RECT 15.380 297.100 19.330 297.250 ;
        RECT 10.130 296.650 10.730 297.100 ;
        RECT 18.730 296.650 19.330 297.100 ;
        RECT 10.130 296.500 14.080 296.650 ;
        RECT 15.380 296.500 19.330 296.650 ;
        RECT 10.130 296.050 10.730 296.500 ;
        RECT 18.730 296.050 19.330 296.500 ;
        RECT 10.130 295.900 14.080 296.050 ;
        RECT 15.380 295.900 19.330 296.050 ;
        RECT 10.130 295.450 10.730 295.900 ;
        RECT 18.730 295.450 19.330 295.900 ;
        RECT 10.130 295.300 14.080 295.450 ;
        RECT 15.380 295.300 19.330 295.450 ;
        RECT 10.130 294.850 10.730 295.300 ;
        RECT 18.730 294.850 19.330 295.300 ;
        RECT 10.130 294.700 14.080 294.850 ;
        RECT 15.380 294.700 19.330 294.850 ;
        RECT 10.130 294.250 10.730 294.700 ;
        RECT 18.730 294.250 19.330 294.700 ;
        RECT 10.130 294.100 14.080 294.250 ;
        RECT 15.380 294.100 19.330 294.250 ;
        RECT 10.130 293.650 10.730 294.100 ;
        RECT 18.730 293.650 19.330 294.100 ;
        RECT 10.130 293.500 14.080 293.650 ;
        RECT 15.380 293.500 19.330 293.650 ;
        RECT 10.130 293.050 10.730 293.500 ;
        RECT 18.730 293.050 19.330 293.500 ;
        RECT 10.130 292.900 14.080 293.050 ;
        RECT 15.380 292.900 19.330 293.050 ;
        RECT 10.130 292.450 10.730 292.900 ;
        RECT 18.730 292.450 19.330 292.900 ;
        RECT 10.130 292.300 14.080 292.450 ;
        RECT 15.380 292.300 19.330 292.450 ;
        RECT 10.130 291.850 10.730 292.300 ;
        RECT 18.730 291.850 19.330 292.300 ;
        RECT 10.130 291.700 14.080 291.850 ;
        RECT 15.380 291.700 19.330 291.850 ;
        RECT 10.130 291.250 10.730 291.700 ;
        RECT 18.730 291.250 19.330 291.700 ;
        RECT 10.130 291.100 14.080 291.250 ;
        RECT 15.380 291.100 19.330 291.250 ;
        RECT 10.130 290.650 10.730 291.100 ;
        RECT 18.730 290.650 19.330 291.100 ;
        RECT 10.130 290.450 14.080 290.650 ;
        RECT 15.380 290.450 19.330 290.650 ;
        RECT 19.780 290.450 19.930 298.000 ;
        RECT 20.380 290.450 20.530 298.000 ;
        RECT 20.980 290.450 21.130 298.000 ;
        RECT 21.580 290.450 21.730 298.000 ;
        RECT 22.180 290.450 22.330 298.000 ;
        RECT 22.780 295.150 22.930 298.000 ;
        RECT 23.530 295.600 25.930 298.800 ;
        RECT 29.280 298.650 30.730 298.950 ;
        RECT 26.530 298.450 30.730 298.650 ;
        RECT 38.730 298.950 50.730 299.800 ;
        RECT 38.730 298.900 49.130 298.950 ;
        RECT 38.730 298.650 40.180 298.900 ;
        RECT 40.330 298.800 49.130 298.900 ;
        RECT 38.730 298.450 42.930 298.650 ;
        RECT 26.530 298.300 34.080 298.450 ;
        RECT 35.430 298.300 42.930 298.450 ;
        RECT 26.530 298.000 30.730 298.300 ;
        RECT 26.530 295.150 26.680 298.000 ;
        RECT 27.130 290.450 27.280 298.000 ;
        RECT 27.730 290.450 27.880 298.000 ;
        RECT 28.330 290.450 28.480 298.000 ;
        RECT 28.930 290.450 29.080 298.000 ;
        RECT 29.530 290.450 29.680 298.000 ;
        RECT 30.130 297.850 30.730 298.000 ;
        RECT 38.730 298.000 42.930 298.300 ;
        RECT 38.730 297.850 39.330 298.000 ;
        RECT 30.130 297.700 34.080 297.850 ;
        RECT 35.380 297.700 39.330 297.850 ;
        RECT 30.130 297.250 30.730 297.700 ;
        RECT 38.730 297.250 39.330 297.700 ;
        RECT 30.130 297.100 34.080 297.250 ;
        RECT 35.380 297.100 39.330 297.250 ;
        RECT 30.130 296.650 30.730 297.100 ;
        RECT 38.730 296.650 39.330 297.100 ;
        RECT 30.130 296.500 34.080 296.650 ;
        RECT 35.380 296.500 39.330 296.650 ;
        RECT 30.130 296.050 30.730 296.500 ;
        RECT 38.730 296.050 39.330 296.500 ;
        RECT 30.130 295.900 34.080 296.050 ;
        RECT 35.380 295.900 39.330 296.050 ;
        RECT 30.130 295.450 30.730 295.900 ;
        RECT 38.730 295.450 39.330 295.900 ;
        RECT 30.130 295.300 34.080 295.450 ;
        RECT 35.380 295.300 39.330 295.450 ;
        RECT 30.130 294.850 30.730 295.300 ;
        RECT 38.730 294.850 39.330 295.300 ;
        RECT 30.130 294.700 34.080 294.850 ;
        RECT 35.380 294.700 39.330 294.850 ;
        RECT 30.130 294.250 30.730 294.700 ;
        RECT 38.730 294.250 39.330 294.700 ;
        RECT 30.130 294.100 34.080 294.250 ;
        RECT 35.380 294.100 39.330 294.250 ;
        RECT 30.130 293.650 30.730 294.100 ;
        RECT 38.730 293.650 39.330 294.100 ;
        RECT 30.130 293.500 34.080 293.650 ;
        RECT 35.380 293.500 39.330 293.650 ;
        RECT 30.130 293.050 30.730 293.500 ;
        RECT 38.730 293.050 39.330 293.500 ;
        RECT 30.130 292.900 34.080 293.050 ;
        RECT 35.380 292.900 39.330 293.050 ;
        RECT 30.130 292.450 30.730 292.900 ;
        RECT 38.730 292.450 39.330 292.900 ;
        RECT 30.130 292.300 34.080 292.450 ;
        RECT 35.380 292.300 39.330 292.450 ;
        RECT 30.130 291.850 30.730 292.300 ;
        RECT 38.730 291.850 39.330 292.300 ;
        RECT 30.130 291.700 34.080 291.850 ;
        RECT 35.380 291.700 39.330 291.850 ;
        RECT 30.130 291.250 30.730 291.700 ;
        RECT 38.730 291.250 39.330 291.700 ;
        RECT 30.130 291.100 34.080 291.250 ;
        RECT 35.380 291.100 39.330 291.250 ;
        RECT 30.130 290.650 30.730 291.100 ;
        RECT 38.730 290.650 39.330 291.100 ;
        RECT 30.130 290.450 34.080 290.650 ;
        RECT 35.380 290.450 39.330 290.650 ;
        RECT 39.780 290.450 39.930 298.000 ;
        RECT 40.380 290.450 40.530 298.000 ;
        RECT 40.980 290.450 41.130 298.000 ;
        RECT 41.580 290.450 41.730 298.000 ;
        RECT 42.180 290.450 42.330 298.000 ;
        RECT 42.780 295.150 42.930 298.000 ;
        RECT 43.530 295.600 45.930 298.800 ;
        RECT 49.280 298.650 50.730 298.950 ;
        RECT 46.530 298.450 50.730 298.650 ;
        RECT 58.730 298.950 70.730 299.800 ;
        RECT 58.730 298.900 69.130 298.950 ;
        RECT 58.730 298.650 60.180 298.900 ;
        RECT 60.330 298.800 69.130 298.900 ;
        RECT 58.730 298.450 62.930 298.650 ;
        RECT 46.530 298.300 54.080 298.450 ;
        RECT 55.430 298.300 62.930 298.450 ;
        RECT 46.530 298.000 50.730 298.300 ;
        RECT 46.530 295.150 46.680 298.000 ;
        RECT 47.130 290.450 47.280 298.000 ;
        RECT 47.730 290.450 47.880 298.000 ;
        RECT 48.330 290.450 48.480 298.000 ;
        RECT 48.930 290.450 49.080 298.000 ;
        RECT 49.530 290.450 49.680 298.000 ;
        RECT 50.130 297.850 50.730 298.000 ;
        RECT 58.730 298.000 62.930 298.300 ;
        RECT 58.730 297.850 59.330 298.000 ;
        RECT 50.130 297.700 54.080 297.850 ;
        RECT 55.380 297.700 59.330 297.850 ;
        RECT 50.130 297.250 50.730 297.700 ;
        RECT 58.730 297.250 59.330 297.700 ;
        RECT 50.130 297.100 54.080 297.250 ;
        RECT 55.380 297.100 59.330 297.250 ;
        RECT 50.130 296.650 50.730 297.100 ;
        RECT 58.730 296.650 59.330 297.100 ;
        RECT 50.130 296.500 54.080 296.650 ;
        RECT 55.380 296.500 59.330 296.650 ;
        RECT 50.130 296.050 50.730 296.500 ;
        RECT 58.730 296.050 59.330 296.500 ;
        RECT 50.130 295.900 54.080 296.050 ;
        RECT 55.380 295.900 59.330 296.050 ;
        RECT 50.130 295.450 50.730 295.900 ;
        RECT 58.730 295.450 59.330 295.900 ;
        RECT 50.130 295.300 54.080 295.450 ;
        RECT 55.380 295.300 59.330 295.450 ;
        RECT 50.130 294.850 50.730 295.300 ;
        RECT 58.730 294.850 59.330 295.300 ;
        RECT 50.130 294.700 54.080 294.850 ;
        RECT 55.380 294.700 59.330 294.850 ;
        RECT 50.130 294.250 50.730 294.700 ;
        RECT 58.730 294.250 59.330 294.700 ;
        RECT 50.130 294.100 54.080 294.250 ;
        RECT 55.380 294.100 59.330 294.250 ;
        RECT 50.130 293.650 50.730 294.100 ;
        RECT 58.730 293.650 59.330 294.100 ;
        RECT 50.130 293.500 54.080 293.650 ;
        RECT 55.380 293.500 59.330 293.650 ;
        RECT 50.130 293.050 50.730 293.500 ;
        RECT 58.730 293.050 59.330 293.500 ;
        RECT 50.130 292.900 54.080 293.050 ;
        RECT 55.380 292.900 59.330 293.050 ;
        RECT 50.130 292.450 50.730 292.900 ;
        RECT 58.730 292.450 59.330 292.900 ;
        RECT 50.130 292.300 54.080 292.450 ;
        RECT 55.380 292.300 59.330 292.450 ;
        RECT 50.130 291.850 50.730 292.300 ;
        RECT 58.730 291.850 59.330 292.300 ;
        RECT 50.130 291.700 54.080 291.850 ;
        RECT 55.380 291.700 59.330 291.850 ;
        RECT 50.130 291.250 50.730 291.700 ;
        RECT 58.730 291.250 59.330 291.700 ;
        RECT 50.130 291.100 54.080 291.250 ;
        RECT 55.380 291.100 59.330 291.250 ;
        RECT 50.130 290.650 50.730 291.100 ;
        RECT 58.730 290.650 59.330 291.100 ;
        RECT 50.130 290.450 54.080 290.650 ;
        RECT 55.380 290.450 59.330 290.650 ;
        RECT 59.780 290.450 59.930 298.000 ;
        RECT 60.380 290.450 60.530 298.000 ;
        RECT 60.980 290.450 61.130 298.000 ;
        RECT 61.580 290.450 61.730 298.000 ;
        RECT 62.180 290.450 62.330 298.000 ;
        RECT 62.780 295.150 62.930 298.000 ;
        RECT 63.530 295.600 65.930 298.800 ;
        RECT 69.280 298.650 70.730 298.950 ;
        RECT 66.530 298.450 70.730 298.650 ;
        RECT 78.730 298.950 90.730 299.800 ;
        RECT 78.730 298.900 89.130 298.950 ;
        RECT 78.730 298.650 80.180 298.900 ;
        RECT 80.330 298.800 89.130 298.900 ;
        RECT 78.730 298.450 82.930 298.650 ;
        RECT 66.530 298.300 74.080 298.450 ;
        RECT 75.430 298.300 82.930 298.450 ;
        RECT 66.530 298.000 70.730 298.300 ;
        RECT 66.530 295.150 66.680 298.000 ;
        RECT 67.130 290.450 67.280 298.000 ;
        RECT 67.730 290.450 67.880 298.000 ;
        RECT 68.330 290.450 68.480 298.000 ;
        RECT 68.930 290.450 69.080 298.000 ;
        RECT 69.530 290.450 69.680 298.000 ;
        RECT 70.130 297.850 70.730 298.000 ;
        RECT 78.730 298.000 82.930 298.300 ;
        RECT 78.730 297.850 79.330 298.000 ;
        RECT 70.130 297.700 74.080 297.850 ;
        RECT 75.380 297.700 79.330 297.850 ;
        RECT 70.130 297.250 70.730 297.700 ;
        RECT 78.730 297.250 79.330 297.700 ;
        RECT 70.130 297.100 74.080 297.250 ;
        RECT 75.380 297.100 79.330 297.250 ;
        RECT 70.130 296.650 70.730 297.100 ;
        RECT 78.730 296.650 79.330 297.100 ;
        RECT 70.130 296.500 74.080 296.650 ;
        RECT 75.380 296.500 79.330 296.650 ;
        RECT 70.130 296.050 70.730 296.500 ;
        RECT 78.730 296.050 79.330 296.500 ;
        RECT 70.130 295.900 74.080 296.050 ;
        RECT 75.380 295.900 79.330 296.050 ;
        RECT 70.130 295.450 70.730 295.900 ;
        RECT 78.730 295.450 79.330 295.900 ;
        RECT 70.130 295.300 74.080 295.450 ;
        RECT 75.380 295.300 79.330 295.450 ;
        RECT 70.130 294.850 70.730 295.300 ;
        RECT 78.730 294.850 79.330 295.300 ;
        RECT 70.130 294.700 74.080 294.850 ;
        RECT 75.380 294.700 79.330 294.850 ;
        RECT 70.130 294.250 70.730 294.700 ;
        RECT 78.730 294.250 79.330 294.700 ;
        RECT 70.130 294.100 74.080 294.250 ;
        RECT 75.380 294.100 79.330 294.250 ;
        RECT 70.130 293.650 70.730 294.100 ;
        RECT 78.730 293.650 79.330 294.100 ;
        RECT 70.130 293.500 74.080 293.650 ;
        RECT 75.380 293.500 79.330 293.650 ;
        RECT 70.130 293.050 70.730 293.500 ;
        RECT 78.730 293.050 79.330 293.500 ;
        RECT 70.130 292.900 74.080 293.050 ;
        RECT 75.380 292.900 79.330 293.050 ;
        RECT 70.130 292.450 70.730 292.900 ;
        RECT 78.730 292.450 79.330 292.900 ;
        RECT 70.130 292.300 74.080 292.450 ;
        RECT 75.380 292.300 79.330 292.450 ;
        RECT 70.130 291.850 70.730 292.300 ;
        RECT 78.730 291.850 79.330 292.300 ;
        RECT 70.130 291.700 74.080 291.850 ;
        RECT 75.380 291.700 79.330 291.850 ;
        RECT 70.130 291.250 70.730 291.700 ;
        RECT 78.730 291.250 79.330 291.700 ;
        RECT 70.130 291.100 74.080 291.250 ;
        RECT 75.380 291.100 79.330 291.250 ;
        RECT 70.130 290.650 70.730 291.100 ;
        RECT 78.730 290.650 79.330 291.100 ;
        RECT 70.130 290.450 74.080 290.650 ;
        RECT 75.380 290.450 79.330 290.650 ;
        RECT 79.780 290.450 79.930 298.000 ;
        RECT 80.380 290.450 80.530 298.000 ;
        RECT 80.980 290.450 81.130 298.000 ;
        RECT 81.580 290.450 81.730 298.000 ;
        RECT 82.180 290.450 82.330 298.000 ;
        RECT 82.780 295.150 82.930 298.000 ;
        RECT 83.530 295.600 85.930 298.800 ;
        RECT 89.280 298.650 90.730 298.950 ;
        RECT 86.530 298.450 90.730 298.650 ;
        RECT 98.730 298.950 110.730 299.800 ;
        RECT 98.730 298.900 109.130 298.950 ;
        RECT 98.730 298.650 100.180 298.900 ;
        RECT 100.330 298.800 109.130 298.900 ;
        RECT 98.730 298.450 102.930 298.650 ;
        RECT 86.530 298.300 94.080 298.450 ;
        RECT 95.430 298.300 102.930 298.450 ;
        RECT 86.530 298.000 90.730 298.300 ;
        RECT 86.530 295.150 86.680 298.000 ;
        RECT 87.130 290.450 87.280 298.000 ;
        RECT 87.730 290.450 87.880 298.000 ;
        RECT 88.330 290.450 88.480 298.000 ;
        RECT 88.930 290.450 89.080 298.000 ;
        RECT 89.530 290.450 89.680 298.000 ;
        RECT 90.130 297.850 90.730 298.000 ;
        RECT 98.730 298.000 102.930 298.300 ;
        RECT 98.730 297.850 99.330 298.000 ;
        RECT 90.130 297.700 94.080 297.850 ;
        RECT 95.380 297.700 99.330 297.850 ;
        RECT 90.130 297.250 90.730 297.700 ;
        RECT 98.730 297.250 99.330 297.700 ;
        RECT 90.130 297.100 94.080 297.250 ;
        RECT 95.380 297.100 99.330 297.250 ;
        RECT 90.130 296.650 90.730 297.100 ;
        RECT 98.730 296.650 99.330 297.100 ;
        RECT 90.130 296.500 94.080 296.650 ;
        RECT 95.380 296.500 99.330 296.650 ;
        RECT 90.130 296.050 90.730 296.500 ;
        RECT 98.730 296.050 99.330 296.500 ;
        RECT 90.130 295.900 94.080 296.050 ;
        RECT 95.380 295.900 99.330 296.050 ;
        RECT 90.130 295.450 90.730 295.900 ;
        RECT 98.730 295.450 99.330 295.900 ;
        RECT 90.130 295.300 94.080 295.450 ;
        RECT 95.380 295.300 99.330 295.450 ;
        RECT 90.130 294.850 90.730 295.300 ;
        RECT 98.730 294.850 99.330 295.300 ;
        RECT 90.130 294.700 94.080 294.850 ;
        RECT 95.380 294.700 99.330 294.850 ;
        RECT 90.130 294.250 90.730 294.700 ;
        RECT 98.730 294.250 99.330 294.700 ;
        RECT 90.130 294.100 94.080 294.250 ;
        RECT 95.380 294.100 99.330 294.250 ;
        RECT 90.130 293.650 90.730 294.100 ;
        RECT 98.730 293.650 99.330 294.100 ;
        RECT 90.130 293.500 94.080 293.650 ;
        RECT 95.380 293.500 99.330 293.650 ;
        RECT 90.130 293.050 90.730 293.500 ;
        RECT 98.730 293.050 99.330 293.500 ;
        RECT 90.130 292.900 94.080 293.050 ;
        RECT 95.380 292.900 99.330 293.050 ;
        RECT 90.130 292.450 90.730 292.900 ;
        RECT 98.730 292.450 99.330 292.900 ;
        RECT 90.130 292.300 94.080 292.450 ;
        RECT 95.380 292.300 99.330 292.450 ;
        RECT 90.130 291.850 90.730 292.300 ;
        RECT 98.730 291.850 99.330 292.300 ;
        RECT 90.130 291.700 94.080 291.850 ;
        RECT 95.380 291.700 99.330 291.850 ;
        RECT 90.130 291.250 90.730 291.700 ;
        RECT 98.730 291.250 99.330 291.700 ;
        RECT 90.130 291.100 94.080 291.250 ;
        RECT 95.380 291.100 99.330 291.250 ;
        RECT 90.130 290.650 90.730 291.100 ;
        RECT 98.730 290.650 99.330 291.100 ;
        RECT 90.130 290.450 94.080 290.650 ;
        RECT 95.380 290.450 99.330 290.650 ;
        RECT 99.780 290.450 99.930 298.000 ;
        RECT 100.380 290.450 100.530 298.000 ;
        RECT 100.980 290.450 101.130 298.000 ;
        RECT 101.580 290.450 101.730 298.000 ;
        RECT 102.180 290.450 102.330 298.000 ;
        RECT 102.780 295.150 102.930 298.000 ;
        RECT 103.530 295.600 105.930 298.800 ;
        RECT 109.280 298.650 110.730 298.950 ;
        RECT 106.530 298.450 110.730 298.650 ;
        RECT 118.730 298.900 124.730 299.800 ;
        RECT 118.730 298.650 120.180 298.900 ;
        RECT 120.330 298.800 124.730 298.900 ;
        RECT 118.730 298.450 122.930 298.650 ;
        RECT 106.530 298.300 114.080 298.450 ;
        RECT 115.430 298.300 122.930 298.450 ;
        RECT 106.530 298.000 110.730 298.300 ;
        RECT 106.530 295.150 106.680 298.000 ;
        RECT 107.130 290.450 107.280 298.000 ;
        RECT 107.730 290.450 107.880 298.000 ;
        RECT 108.330 290.450 108.480 298.000 ;
        RECT 108.930 290.450 109.080 298.000 ;
        RECT 109.530 290.450 109.680 298.000 ;
        RECT 110.130 297.850 110.730 298.000 ;
        RECT 118.730 298.000 122.930 298.300 ;
        RECT 118.730 297.850 119.330 298.000 ;
        RECT 110.130 297.700 114.080 297.850 ;
        RECT 115.380 297.700 119.330 297.850 ;
        RECT 110.130 297.250 110.730 297.700 ;
        RECT 118.730 297.250 119.330 297.700 ;
        RECT 110.130 297.100 114.080 297.250 ;
        RECT 115.380 297.100 119.330 297.250 ;
        RECT 110.130 296.650 110.730 297.100 ;
        RECT 118.730 296.650 119.330 297.100 ;
        RECT 110.130 296.500 114.080 296.650 ;
        RECT 115.380 296.500 119.330 296.650 ;
        RECT 110.130 296.050 110.730 296.500 ;
        RECT 118.730 296.050 119.330 296.500 ;
        RECT 110.130 295.900 114.080 296.050 ;
        RECT 115.380 295.900 119.330 296.050 ;
        RECT 110.130 295.450 110.730 295.900 ;
        RECT 118.730 295.450 119.330 295.900 ;
        RECT 110.130 295.300 114.080 295.450 ;
        RECT 115.380 295.300 119.330 295.450 ;
        RECT 110.130 294.850 110.730 295.300 ;
        RECT 118.730 294.850 119.330 295.300 ;
        RECT 110.130 294.700 114.080 294.850 ;
        RECT 115.380 294.700 119.330 294.850 ;
        RECT 110.130 294.250 110.730 294.700 ;
        RECT 118.730 294.250 119.330 294.700 ;
        RECT 110.130 294.100 114.080 294.250 ;
        RECT 115.380 294.100 119.330 294.250 ;
        RECT 110.130 293.650 110.730 294.100 ;
        RECT 118.730 293.650 119.330 294.100 ;
        RECT 110.130 293.500 114.080 293.650 ;
        RECT 115.380 293.500 119.330 293.650 ;
        RECT 110.130 293.050 110.730 293.500 ;
        RECT 118.730 293.050 119.330 293.500 ;
        RECT 110.130 292.900 114.080 293.050 ;
        RECT 115.380 292.900 119.330 293.050 ;
        RECT 110.130 292.450 110.730 292.900 ;
        RECT 118.730 292.450 119.330 292.900 ;
        RECT 110.130 292.300 114.080 292.450 ;
        RECT 115.380 292.300 119.330 292.450 ;
        RECT 110.130 291.850 110.730 292.300 ;
        RECT 118.730 291.850 119.330 292.300 ;
        RECT 110.130 291.700 114.080 291.850 ;
        RECT 115.380 291.700 119.330 291.850 ;
        RECT 110.130 291.250 110.730 291.700 ;
        RECT 118.730 291.250 119.330 291.700 ;
        RECT 110.130 291.100 114.080 291.250 ;
        RECT 115.380 291.100 119.330 291.250 ;
        RECT 110.130 290.650 110.730 291.100 ;
        RECT 118.730 290.650 119.330 291.100 ;
        RECT 110.130 290.450 114.080 290.650 ;
        RECT 115.380 290.450 119.330 290.650 ;
        RECT 119.780 290.450 119.930 298.000 ;
        RECT 120.380 290.450 120.530 298.000 ;
        RECT 120.980 290.450 121.130 298.000 ;
        RECT 121.580 290.450 121.730 298.000 ;
        RECT 122.180 290.450 122.330 298.000 ;
        RECT 122.780 295.150 122.930 298.000 ;
        RECT 123.530 297.585 124.730 298.800 ;
        RECT 123.530 296.310 127.130 297.585 ;
        RECT 123.530 295.600 124.730 296.310 ;
        RECT 2.315 284.455 4.315 286.750 ;
        RECT 4.730 283.545 5.930 284.400 ;
        RECT 2.315 282.270 5.930 283.545 ;
        RECT 4.730 281.200 5.930 282.270 ;
        RECT 6.530 282.000 6.680 284.900 ;
        RECT 7.130 282.000 7.280 289.550 ;
        RECT 7.730 282.000 7.880 289.550 ;
        RECT 8.330 282.000 8.480 289.550 ;
        RECT 8.930 282.000 9.080 289.550 ;
        RECT 9.530 282.000 9.680 289.550 ;
        RECT 10.130 289.350 14.080 289.550 ;
        RECT 15.380 289.350 19.330 289.550 ;
        RECT 10.130 288.900 10.730 289.350 ;
        RECT 18.730 288.900 19.330 289.350 ;
        RECT 10.130 288.750 14.080 288.900 ;
        RECT 15.380 288.750 19.330 288.900 ;
        RECT 10.130 288.300 10.730 288.750 ;
        RECT 18.730 288.300 19.330 288.750 ;
        RECT 10.130 288.150 14.080 288.300 ;
        RECT 15.380 288.150 19.330 288.300 ;
        RECT 10.130 287.700 10.730 288.150 ;
        RECT 18.730 287.700 19.330 288.150 ;
        RECT 10.130 287.550 14.080 287.700 ;
        RECT 15.380 287.550 19.330 287.700 ;
        RECT 10.130 287.100 10.730 287.550 ;
        RECT 18.730 287.100 19.330 287.550 ;
        RECT 10.130 286.950 14.080 287.100 ;
        RECT 15.380 286.950 19.330 287.100 ;
        RECT 10.130 286.500 10.730 286.950 ;
        RECT 18.730 286.500 19.330 286.950 ;
        RECT 10.130 286.350 14.080 286.500 ;
        RECT 15.380 286.350 19.330 286.500 ;
        RECT 10.130 285.900 10.730 286.350 ;
        RECT 18.730 285.900 19.330 286.350 ;
        RECT 10.130 285.750 14.080 285.900 ;
        RECT 15.380 285.750 19.330 285.900 ;
        RECT 10.130 285.300 10.730 285.750 ;
        RECT 18.730 285.300 19.330 285.750 ;
        RECT 10.130 285.150 14.080 285.300 ;
        RECT 15.380 285.150 19.330 285.300 ;
        RECT 10.130 284.700 10.730 285.150 ;
        RECT 18.730 284.700 19.330 285.150 ;
        RECT 10.130 284.550 14.080 284.700 ;
        RECT 15.380 284.550 19.330 284.700 ;
        RECT 10.130 284.100 10.730 284.550 ;
        RECT 18.730 284.100 19.330 284.550 ;
        RECT 10.130 283.950 14.080 284.100 ;
        RECT 15.380 283.950 19.330 284.100 ;
        RECT 10.130 283.500 10.730 283.950 ;
        RECT 18.730 283.500 19.330 283.950 ;
        RECT 10.130 283.350 14.080 283.500 ;
        RECT 15.380 283.350 19.330 283.500 ;
        RECT 10.130 282.900 10.730 283.350 ;
        RECT 18.730 282.900 19.330 283.350 ;
        RECT 10.130 282.750 14.080 282.900 ;
        RECT 15.380 282.750 19.330 282.900 ;
        RECT 10.130 282.300 10.730 282.750 ;
        RECT 18.730 282.300 19.330 282.750 ;
        RECT 10.130 282.150 14.080 282.300 ;
        RECT 15.380 282.150 19.330 282.300 ;
        RECT 10.130 282.000 10.730 282.150 ;
        RECT 6.530 281.700 10.730 282.000 ;
        RECT 18.730 282.000 19.330 282.150 ;
        RECT 19.780 282.000 19.930 289.550 ;
        RECT 20.380 282.000 20.530 289.550 ;
        RECT 20.980 282.000 21.130 289.550 ;
        RECT 21.580 282.000 21.730 289.550 ;
        RECT 22.180 282.000 22.330 289.550 ;
        RECT 22.780 282.000 22.930 284.900 ;
        RECT 18.730 281.700 22.930 282.000 ;
        RECT 6.530 281.550 14.080 281.700 ;
        RECT 15.380 281.550 22.930 281.700 ;
        RECT 6.530 281.350 10.730 281.550 ;
        RECT 4.730 281.050 9.130 281.200 ;
        RECT 9.280 281.050 10.730 281.350 ;
        RECT 4.730 280.150 10.730 281.050 ;
        RECT 18.730 281.350 22.930 281.550 ;
        RECT 18.730 281.050 20.180 281.350 ;
        RECT 23.530 281.200 25.930 284.400 ;
        RECT 26.530 282.000 26.680 284.900 ;
        RECT 27.130 282.000 27.280 289.550 ;
        RECT 27.730 282.000 27.880 289.550 ;
        RECT 28.330 282.000 28.480 289.550 ;
        RECT 28.930 282.000 29.080 289.550 ;
        RECT 29.530 282.000 29.680 289.550 ;
        RECT 30.130 289.350 34.080 289.550 ;
        RECT 35.380 289.350 39.330 289.550 ;
        RECT 30.130 288.900 30.730 289.350 ;
        RECT 38.730 288.900 39.330 289.350 ;
        RECT 30.130 288.750 34.080 288.900 ;
        RECT 35.380 288.750 39.330 288.900 ;
        RECT 30.130 288.300 30.730 288.750 ;
        RECT 38.730 288.300 39.330 288.750 ;
        RECT 30.130 288.150 34.080 288.300 ;
        RECT 35.380 288.150 39.330 288.300 ;
        RECT 30.130 287.700 30.730 288.150 ;
        RECT 38.730 287.700 39.330 288.150 ;
        RECT 30.130 287.550 34.080 287.700 ;
        RECT 35.380 287.550 39.330 287.700 ;
        RECT 30.130 287.100 30.730 287.550 ;
        RECT 38.730 287.100 39.330 287.550 ;
        RECT 30.130 286.950 34.080 287.100 ;
        RECT 35.380 286.950 39.330 287.100 ;
        RECT 30.130 286.500 30.730 286.950 ;
        RECT 38.730 286.500 39.330 286.950 ;
        RECT 30.130 286.350 34.080 286.500 ;
        RECT 35.380 286.350 39.330 286.500 ;
        RECT 30.130 285.900 30.730 286.350 ;
        RECT 38.730 285.900 39.330 286.350 ;
        RECT 30.130 285.750 34.080 285.900 ;
        RECT 35.380 285.750 39.330 285.900 ;
        RECT 30.130 285.300 30.730 285.750 ;
        RECT 38.730 285.300 39.330 285.750 ;
        RECT 30.130 285.150 34.080 285.300 ;
        RECT 35.380 285.150 39.330 285.300 ;
        RECT 30.130 284.700 30.730 285.150 ;
        RECT 38.730 284.700 39.330 285.150 ;
        RECT 30.130 284.550 34.080 284.700 ;
        RECT 35.380 284.550 39.330 284.700 ;
        RECT 30.130 284.100 30.730 284.550 ;
        RECT 38.730 284.100 39.330 284.550 ;
        RECT 30.130 283.950 34.080 284.100 ;
        RECT 35.380 283.950 39.330 284.100 ;
        RECT 30.130 283.500 30.730 283.950 ;
        RECT 38.730 283.500 39.330 283.950 ;
        RECT 30.130 283.350 34.080 283.500 ;
        RECT 35.380 283.350 39.330 283.500 ;
        RECT 30.130 282.900 30.730 283.350 ;
        RECT 38.730 282.900 39.330 283.350 ;
        RECT 30.130 282.750 34.080 282.900 ;
        RECT 35.380 282.750 39.330 282.900 ;
        RECT 30.130 282.300 30.730 282.750 ;
        RECT 38.730 282.300 39.330 282.750 ;
        RECT 30.130 282.150 34.080 282.300 ;
        RECT 35.380 282.150 39.330 282.300 ;
        RECT 30.130 282.000 30.730 282.150 ;
        RECT 26.530 281.700 30.730 282.000 ;
        RECT 38.730 282.000 39.330 282.150 ;
        RECT 39.780 282.000 39.930 289.550 ;
        RECT 40.380 282.000 40.530 289.550 ;
        RECT 40.980 282.000 41.130 289.550 ;
        RECT 41.580 282.000 41.730 289.550 ;
        RECT 42.180 282.000 42.330 289.550 ;
        RECT 42.780 282.000 42.930 284.900 ;
        RECT 38.730 281.700 42.930 282.000 ;
        RECT 26.530 281.550 34.080 281.700 ;
        RECT 35.380 281.550 42.930 281.700 ;
        RECT 26.530 281.350 30.730 281.550 ;
        RECT 20.330 281.050 29.130 281.200 ;
        RECT 29.280 281.050 30.730 281.350 ;
        RECT 18.730 280.150 30.730 281.050 ;
        RECT 38.730 281.350 42.930 281.550 ;
        RECT 38.730 281.050 40.180 281.350 ;
        RECT 43.530 281.200 45.930 284.400 ;
        RECT 46.530 282.000 46.680 284.900 ;
        RECT 47.130 282.000 47.280 289.550 ;
        RECT 47.730 282.000 47.880 289.550 ;
        RECT 48.330 282.000 48.480 289.550 ;
        RECT 48.930 282.000 49.080 289.550 ;
        RECT 49.530 282.000 49.680 289.550 ;
        RECT 50.130 289.350 54.080 289.550 ;
        RECT 55.380 289.350 59.330 289.550 ;
        RECT 50.130 288.900 50.730 289.350 ;
        RECT 58.730 288.900 59.330 289.350 ;
        RECT 50.130 288.750 54.080 288.900 ;
        RECT 55.380 288.750 59.330 288.900 ;
        RECT 50.130 288.300 50.730 288.750 ;
        RECT 58.730 288.300 59.330 288.750 ;
        RECT 50.130 288.150 54.080 288.300 ;
        RECT 55.380 288.150 59.330 288.300 ;
        RECT 50.130 287.700 50.730 288.150 ;
        RECT 58.730 287.700 59.330 288.150 ;
        RECT 50.130 287.550 54.080 287.700 ;
        RECT 55.380 287.550 59.330 287.700 ;
        RECT 50.130 287.100 50.730 287.550 ;
        RECT 58.730 287.100 59.330 287.550 ;
        RECT 50.130 286.950 54.080 287.100 ;
        RECT 55.380 286.950 59.330 287.100 ;
        RECT 50.130 286.500 50.730 286.950 ;
        RECT 58.730 286.500 59.330 286.950 ;
        RECT 50.130 286.350 54.080 286.500 ;
        RECT 55.380 286.350 59.330 286.500 ;
        RECT 50.130 285.900 50.730 286.350 ;
        RECT 58.730 285.900 59.330 286.350 ;
        RECT 50.130 285.750 54.080 285.900 ;
        RECT 55.380 285.750 59.330 285.900 ;
        RECT 50.130 285.300 50.730 285.750 ;
        RECT 58.730 285.300 59.330 285.750 ;
        RECT 50.130 285.150 54.080 285.300 ;
        RECT 55.380 285.150 59.330 285.300 ;
        RECT 50.130 284.700 50.730 285.150 ;
        RECT 58.730 284.700 59.330 285.150 ;
        RECT 50.130 284.550 54.080 284.700 ;
        RECT 55.380 284.550 59.330 284.700 ;
        RECT 50.130 284.100 50.730 284.550 ;
        RECT 58.730 284.100 59.330 284.550 ;
        RECT 50.130 283.950 54.080 284.100 ;
        RECT 55.380 283.950 59.330 284.100 ;
        RECT 50.130 283.500 50.730 283.950 ;
        RECT 58.730 283.500 59.330 283.950 ;
        RECT 50.130 283.350 54.080 283.500 ;
        RECT 55.380 283.350 59.330 283.500 ;
        RECT 50.130 282.900 50.730 283.350 ;
        RECT 58.730 282.900 59.330 283.350 ;
        RECT 50.130 282.750 54.080 282.900 ;
        RECT 55.380 282.750 59.330 282.900 ;
        RECT 50.130 282.300 50.730 282.750 ;
        RECT 58.730 282.300 59.330 282.750 ;
        RECT 50.130 282.150 54.080 282.300 ;
        RECT 55.380 282.150 59.330 282.300 ;
        RECT 50.130 282.000 50.730 282.150 ;
        RECT 46.530 281.700 50.730 282.000 ;
        RECT 58.730 282.000 59.330 282.150 ;
        RECT 59.780 282.000 59.930 289.550 ;
        RECT 60.380 282.000 60.530 289.550 ;
        RECT 60.980 282.000 61.130 289.550 ;
        RECT 61.580 282.000 61.730 289.550 ;
        RECT 62.180 282.000 62.330 289.550 ;
        RECT 62.780 282.000 62.930 284.900 ;
        RECT 58.730 281.700 62.930 282.000 ;
        RECT 46.530 281.550 54.080 281.700 ;
        RECT 55.380 281.550 62.930 281.700 ;
        RECT 46.530 281.350 50.730 281.550 ;
        RECT 40.330 281.050 49.130 281.200 ;
        RECT 49.280 281.050 50.730 281.350 ;
        RECT 38.730 280.150 50.730 281.050 ;
        RECT 58.730 281.350 62.930 281.550 ;
        RECT 58.730 281.050 60.180 281.350 ;
        RECT 63.530 281.200 65.930 284.400 ;
        RECT 66.530 282.000 66.680 284.900 ;
        RECT 67.130 282.000 67.280 289.550 ;
        RECT 67.730 282.000 67.880 289.550 ;
        RECT 68.330 282.000 68.480 289.550 ;
        RECT 68.930 282.000 69.080 289.550 ;
        RECT 69.530 282.000 69.680 289.550 ;
        RECT 70.130 289.350 74.080 289.550 ;
        RECT 75.380 289.350 79.330 289.550 ;
        RECT 70.130 288.900 70.730 289.350 ;
        RECT 78.730 288.900 79.330 289.350 ;
        RECT 70.130 288.750 74.080 288.900 ;
        RECT 75.380 288.750 79.330 288.900 ;
        RECT 70.130 288.300 70.730 288.750 ;
        RECT 78.730 288.300 79.330 288.750 ;
        RECT 70.130 288.150 74.080 288.300 ;
        RECT 75.380 288.150 79.330 288.300 ;
        RECT 70.130 287.700 70.730 288.150 ;
        RECT 78.730 287.700 79.330 288.150 ;
        RECT 70.130 287.550 74.080 287.700 ;
        RECT 75.380 287.550 79.330 287.700 ;
        RECT 70.130 287.100 70.730 287.550 ;
        RECT 78.730 287.100 79.330 287.550 ;
        RECT 70.130 286.950 74.080 287.100 ;
        RECT 75.380 286.950 79.330 287.100 ;
        RECT 70.130 286.500 70.730 286.950 ;
        RECT 78.730 286.500 79.330 286.950 ;
        RECT 70.130 286.350 74.080 286.500 ;
        RECT 75.380 286.350 79.330 286.500 ;
        RECT 70.130 285.900 70.730 286.350 ;
        RECT 78.730 285.900 79.330 286.350 ;
        RECT 70.130 285.750 74.080 285.900 ;
        RECT 75.380 285.750 79.330 285.900 ;
        RECT 70.130 285.300 70.730 285.750 ;
        RECT 78.730 285.300 79.330 285.750 ;
        RECT 70.130 285.150 74.080 285.300 ;
        RECT 75.380 285.150 79.330 285.300 ;
        RECT 70.130 284.700 70.730 285.150 ;
        RECT 78.730 284.700 79.330 285.150 ;
        RECT 70.130 284.550 74.080 284.700 ;
        RECT 75.380 284.550 79.330 284.700 ;
        RECT 70.130 284.100 70.730 284.550 ;
        RECT 78.730 284.100 79.330 284.550 ;
        RECT 70.130 283.950 74.080 284.100 ;
        RECT 75.380 283.950 79.330 284.100 ;
        RECT 70.130 283.500 70.730 283.950 ;
        RECT 78.730 283.500 79.330 283.950 ;
        RECT 70.130 283.350 74.080 283.500 ;
        RECT 75.380 283.350 79.330 283.500 ;
        RECT 70.130 282.900 70.730 283.350 ;
        RECT 78.730 282.900 79.330 283.350 ;
        RECT 70.130 282.750 74.080 282.900 ;
        RECT 75.380 282.750 79.330 282.900 ;
        RECT 70.130 282.300 70.730 282.750 ;
        RECT 78.730 282.300 79.330 282.750 ;
        RECT 70.130 282.150 74.080 282.300 ;
        RECT 75.380 282.150 79.330 282.300 ;
        RECT 70.130 282.000 70.730 282.150 ;
        RECT 66.530 281.700 70.730 282.000 ;
        RECT 78.730 282.000 79.330 282.150 ;
        RECT 79.780 282.000 79.930 289.550 ;
        RECT 80.380 282.000 80.530 289.550 ;
        RECT 80.980 282.000 81.130 289.550 ;
        RECT 81.580 282.000 81.730 289.550 ;
        RECT 82.180 282.000 82.330 289.550 ;
        RECT 82.780 282.000 82.930 284.900 ;
        RECT 78.730 281.700 82.930 282.000 ;
        RECT 66.530 281.550 74.080 281.700 ;
        RECT 75.380 281.550 82.930 281.700 ;
        RECT 66.530 281.350 70.730 281.550 ;
        RECT 60.330 281.050 69.130 281.200 ;
        RECT 69.280 281.050 70.730 281.350 ;
        RECT 58.730 280.150 70.730 281.050 ;
        RECT 78.730 281.350 82.930 281.550 ;
        RECT 78.730 281.050 80.180 281.350 ;
        RECT 83.530 281.200 85.930 284.400 ;
        RECT 86.530 282.000 86.680 284.900 ;
        RECT 87.130 282.000 87.280 289.550 ;
        RECT 87.730 282.000 87.880 289.550 ;
        RECT 88.330 282.000 88.480 289.550 ;
        RECT 88.930 282.000 89.080 289.550 ;
        RECT 89.530 282.000 89.680 289.550 ;
        RECT 90.130 289.350 94.080 289.550 ;
        RECT 95.380 289.350 99.330 289.550 ;
        RECT 90.130 288.900 90.730 289.350 ;
        RECT 98.730 288.900 99.330 289.350 ;
        RECT 90.130 288.750 94.080 288.900 ;
        RECT 95.380 288.750 99.330 288.900 ;
        RECT 90.130 288.300 90.730 288.750 ;
        RECT 98.730 288.300 99.330 288.750 ;
        RECT 90.130 288.150 94.080 288.300 ;
        RECT 95.380 288.150 99.330 288.300 ;
        RECT 90.130 287.700 90.730 288.150 ;
        RECT 98.730 287.700 99.330 288.150 ;
        RECT 90.130 287.550 94.080 287.700 ;
        RECT 95.380 287.550 99.330 287.700 ;
        RECT 90.130 287.100 90.730 287.550 ;
        RECT 98.730 287.100 99.330 287.550 ;
        RECT 90.130 286.950 94.080 287.100 ;
        RECT 95.380 286.950 99.330 287.100 ;
        RECT 90.130 286.500 90.730 286.950 ;
        RECT 98.730 286.500 99.330 286.950 ;
        RECT 90.130 286.350 94.080 286.500 ;
        RECT 95.380 286.350 99.330 286.500 ;
        RECT 90.130 285.900 90.730 286.350 ;
        RECT 98.730 285.900 99.330 286.350 ;
        RECT 90.130 285.750 94.080 285.900 ;
        RECT 95.380 285.750 99.330 285.900 ;
        RECT 90.130 285.300 90.730 285.750 ;
        RECT 98.730 285.300 99.330 285.750 ;
        RECT 90.130 285.150 94.080 285.300 ;
        RECT 95.380 285.150 99.330 285.300 ;
        RECT 90.130 284.700 90.730 285.150 ;
        RECT 98.730 284.700 99.330 285.150 ;
        RECT 90.130 284.550 94.080 284.700 ;
        RECT 95.380 284.550 99.330 284.700 ;
        RECT 90.130 284.100 90.730 284.550 ;
        RECT 98.730 284.100 99.330 284.550 ;
        RECT 90.130 283.950 94.080 284.100 ;
        RECT 95.380 283.950 99.330 284.100 ;
        RECT 90.130 283.500 90.730 283.950 ;
        RECT 98.730 283.500 99.330 283.950 ;
        RECT 90.130 283.350 94.080 283.500 ;
        RECT 95.380 283.350 99.330 283.500 ;
        RECT 90.130 282.900 90.730 283.350 ;
        RECT 98.730 282.900 99.330 283.350 ;
        RECT 90.130 282.750 94.080 282.900 ;
        RECT 95.380 282.750 99.330 282.900 ;
        RECT 90.130 282.300 90.730 282.750 ;
        RECT 98.730 282.300 99.330 282.750 ;
        RECT 90.130 282.150 94.080 282.300 ;
        RECT 95.380 282.150 99.330 282.300 ;
        RECT 90.130 282.000 90.730 282.150 ;
        RECT 86.530 281.700 90.730 282.000 ;
        RECT 98.730 282.000 99.330 282.150 ;
        RECT 99.780 282.000 99.930 289.550 ;
        RECT 100.380 282.000 100.530 289.550 ;
        RECT 100.980 282.000 101.130 289.550 ;
        RECT 101.580 282.000 101.730 289.550 ;
        RECT 102.180 282.000 102.330 289.550 ;
        RECT 102.780 282.000 102.930 284.900 ;
        RECT 98.730 281.700 102.930 282.000 ;
        RECT 86.530 281.550 94.080 281.700 ;
        RECT 95.380 281.550 102.930 281.700 ;
        RECT 86.530 281.350 90.730 281.550 ;
        RECT 80.330 281.050 89.130 281.200 ;
        RECT 89.280 281.050 90.730 281.350 ;
        RECT 78.730 280.150 90.730 281.050 ;
        RECT 98.730 281.350 102.930 281.550 ;
        RECT 98.730 281.050 100.180 281.350 ;
        RECT 103.530 281.200 105.930 284.400 ;
        RECT 106.530 282.000 106.680 284.900 ;
        RECT 107.130 282.000 107.280 289.550 ;
        RECT 107.730 282.000 107.880 289.550 ;
        RECT 108.330 282.000 108.480 289.550 ;
        RECT 108.930 282.000 109.080 289.550 ;
        RECT 109.530 282.000 109.680 289.550 ;
        RECT 110.130 289.350 114.080 289.550 ;
        RECT 115.380 289.350 119.330 289.550 ;
        RECT 110.130 288.900 110.730 289.350 ;
        RECT 118.730 288.900 119.330 289.350 ;
        RECT 110.130 288.750 114.080 288.900 ;
        RECT 115.380 288.750 119.330 288.900 ;
        RECT 110.130 288.300 110.730 288.750 ;
        RECT 118.730 288.300 119.330 288.750 ;
        RECT 110.130 288.150 114.080 288.300 ;
        RECT 115.380 288.150 119.330 288.300 ;
        RECT 110.130 287.700 110.730 288.150 ;
        RECT 118.730 287.700 119.330 288.150 ;
        RECT 110.130 287.550 114.080 287.700 ;
        RECT 115.380 287.550 119.330 287.700 ;
        RECT 110.130 287.100 110.730 287.550 ;
        RECT 118.730 287.100 119.330 287.550 ;
        RECT 110.130 286.950 114.080 287.100 ;
        RECT 115.380 286.950 119.330 287.100 ;
        RECT 110.130 286.500 110.730 286.950 ;
        RECT 118.730 286.500 119.330 286.950 ;
        RECT 110.130 286.350 114.080 286.500 ;
        RECT 115.380 286.350 119.330 286.500 ;
        RECT 110.130 285.900 110.730 286.350 ;
        RECT 118.730 285.900 119.330 286.350 ;
        RECT 110.130 285.750 114.080 285.900 ;
        RECT 115.380 285.750 119.330 285.900 ;
        RECT 110.130 285.300 110.730 285.750 ;
        RECT 118.730 285.300 119.330 285.750 ;
        RECT 110.130 285.150 114.080 285.300 ;
        RECT 115.380 285.150 119.330 285.300 ;
        RECT 110.130 284.700 110.730 285.150 ;
        RECT 118.730 284.700 119.330 285.150 ;
        RECT 110.130 284.550 114.080 284.700 ;
        RECT 115.380 284.550 119.330 284.700 ;
        RECT 110.130 284.100 110.730 284.550 ;
        RECT 118.730 284.100 119.330 284.550 ;
        RECT 110.130 283.950 114.080 284.100 ;
        RECT 115.380 283.950 119.330 284.100 ;
        RECT 110.130 283.500 110.730 283.950 ;
        RECT 118.730 283.500 119.330 283.950 ;
        RECT 110.130 283.350 114.080 283.500 ;
        RECT 115.380 283.350 119.330 283.500 ;
        RECT 110.130 282.900 110.730 283.350 ;
        RECT 118.730 282.900 119.330 283.350 ;
        RECT 110.130 282.750 114.080 282.900 ;
        RECT 115.380 282.750 119.330 282.900 ;
        RECT 110.130 282.300 110.730 282.750 ;
        RECT 118.730 282.300 119.330 282.750 ;
        RECT 110.130 282.150 114.080 282.300 ;
        RECT 115.380 282.150 119.330 282.300 ;
        RECT 110.130 282.000 110.730 282.150 ;
        RECT 106.530 281.700 110.730 282.000 ;
        RECT 118.730 282.000 119.330 282.150 ;
        RECT 119.780 282.000 119.930 289.550 ;
        RECT 120.380 282.000 120.530 289.550 ;
        RECT 120.980 282.000 121.130 289.550 ;
        RECT 121.580 282.000 121.730 289.550 ;
        RECT 122.180 282.000 122.330 289.550 ;
        RECT 122.780 282.000 122.930 284.900 ;
        RECT 118.730 281.700 122.930 282.000 ;
        RECT 106.530 281.550 114.080 281.700 ;
        RECT 115.380 281.550 122.930 281.700 ;
        RECT 106.530 281.350 110.730 281.550 ;
        RECT 100.330 281.050 109.130 281.200 ;
        RECT 109.280 281.050 110.730 281.350 ;
        RECT 98.730 280.150 110.730 281.050 ;
        RECT 118.730 281.350 122.930 281.550 ;
        RECT 123.530 283.600 124.730 284.400 ;
        RECT 123.530 282.325 127.140 283.600 ;
        RECT 118.730 281.050 120.180 281.350 ;
        RECT 123.530 281.200 124.730 282.325 ;
        RECT 120.330 281.050 124.730 281.200 ;
        RECT 118.730 280.150 124.730 281.050 ;
        RECT 4.730 279.850 9.130 280.150 ;
        RECT 20.330 279.850 29.130 280.150 ;
        RECT 40.330 279.850 49.130 280.150 ;
        RECT 60.330 279.850 69.130 280.150 ;
        RECT 80.330 279.850 89.130 280.150 ;
        RECT 100.330 279.850 109.130 280.150 ;
        RECT 4.730 278.950 10.730 279.850 ;
        RECT 20.330 279.800 30.730 279.850 ;
        RECT 40.330 279.800 50.730 279.850 ;
        RECT 60.330 279.800 70.730 279.850 ;
        RECT 80.330 279.800 90.730 279.850 ;
        RECT 100.330 279.800 110.730 279.850 ;
        RECT 120.330 279.800 124.730 280.150 ;
        RECT 4.730 278.800 9.130 278.950 ;
        RECT 4.730 277.530 5.930 278.800 ;
        RECT 9.280 278.650 10.730 278.950 ;
        RECT 2.315 276.255 5.930 277.530 ;
        RECT 4.730 275.600 5.930 276.255 ;
        RECT 6.530 278.450 10.730 278.650 ;
        RECT 18.730 278.950 30.730 279.800 ;
        RECT 18.730 278.900 29.130 278.950 ;
        RECT 18.730 278.650 20.180 278.900 ;
        RECT 20.330 278.800 29.130 278.900 ;
        RECT 18.730 278.450 22.930 278.650 ;
        RECT 6.530 278.300 14.080 278.450 ;
        RECT 15.430 278.300 22.930 278.450 ;
        RECT 6.530 278.000 10.730 278.300 ;
        RECT 2.320 275.340 4.320 275.545 ;
        RECT 2.315 273.250 4.320 275.340 ;
        RECT 6.530 275.150 6.680 278.000 ;
        RECT 7.130 270.450 7.280 278.000 ;
        RECT 7.730 270.450 7.880 278.000 ;
        RECT 8.330 270.450 8.480 278.000 ;
        RECT 8.930 270.450 9.080 278.000 ;
        RECT 9.530 270.450 9.680 278.000 ;
        RECT 10.130 277.850 10.730 278.000 ;
        RECT 18.730 278.000 22.930 278.300 ;
        RECT 18.730 277.850 19.330 278.000 ;
        RECT 10.130 277.700 14.080 277.850 ;
        RECT 15.380 277.700 19.330 277.850 ;
        RECT 10.130 277.250 10.730 277.700 ;
        RECT 18.730 277.250 19.330 277.700 ;
        RECT 10.130 277.100 14.080 277.250 ;
        RECT 15.380 277.100 19.330 277.250 ;
        RECT 10.130 276.650 10.730 277.100 ;
        RECT 18.730 276.650 19.330 277.100 ;
        RECT 10.130 276.500 14.080 276.650 ;
        RECT 15.380 276.500 19.330 276.650 ;
        RECT 10.130 276.050 10.730 276.500 ;
        RECT 18.730 276.050 19.330 276.500 ;
        RECT 10.130 275.900 14.080 276.050 ;
        RECT 15.380 275.900 19.330 276.050 ;
        RECT 10.130 275.450 10.730 275.900 ;
        RECT 18.730 275.450 19.330 275.900 ;
        RECT 10.130 275.300 14.080 275.450 ;
        RECT 15.380 275.300 19.330 275.450 ;
        RECT 10.130 274.850 10.730 275.300 ;
        RECT 18.730 274.850 19.330 275.300 ;
        RECT 10.130 274.700 14.080 274.850 ;
        RECT 15.380 274.700 19.330 274.850 ;
        RECT 10.130 274.250 10.730 274.700 ;
        RECT 18.730 274.250 19.330 274.700 ;
        RECT 10.130 274.100 14.080 274.250 ;
        RECT 15.380 274.100 19.330 274.250 ;
        RECT 10.130 273.650 10.730 274.100 ;
        RECT 18.730 273.650 19.330 274.100 ;
        RECT 10.130 273.500 14.080 273.650 ;
        RECT 15.380 273.500 19.330 273.650 ;
        RECT 10.130 273.050 10.730 273.500 ;
        RECT 18.730 273.050 19.330 273.500 ;
        RECT 10.130 272.900 14.080 273.050 ;
        RECT 15.380 272.900 19.330 273.050 ;
        RECT 10.130 272.450 10.730 272.900 ;
        RECT 18.730 272.450 19.330 272.900 ;
        RECT 10.130 272.300 14.080 272.450 ;
        RECT 15.380 272.300 19.330 272.450 ;
        RECT 10.130 271.850 10.730 272.300 ;
        RECT 18.730 271.850 19.330 272.300 ;
        RECT 10.130 271.700 14.080 271.850 ;
        RECT 15.380 271.700 19.330 271.850 ;
        RECT 10.130 271.250 10.730 271.700 ;
        RECT 18.730 271.250 19.330 271.700 ;
        RECT 10.130 271.100 14.080 271.250 ;
        RECT 15.380 271.100 19.330 271.250 ;
        RECT 10.130 270.650 10.730 271.100 ;
        RECT 18.730 270.650 19.330 271.100 ;
        RECT 10.130 270.450 14.080 270.650 ;
        RECT 15.380 270.450 19.330 270.650 ;
        RECT 19.780 270.450 19.930 278.000 ;
        RECT 20.380 270.450 20.530 278.000 ;
        RECT 20.980 270.450 21.130 278.000 ;
        RECT 21.580 270.450 21.730 278.000 ;
        RECT 22.180 270.450 22.330 278.000 ;
        RECT 22.780 275.150 22.930 278.000 ;
        RECT 23.530 275.600 25.930 278.800 ;
        RECT 29.280 278.650 30.730 278.950 ;
        RECT 26.530 278.450 30.730 278.650 ;
        RECT 38.730 278.950 50.730 279.800 ;
        RECT 38.730 278.900 49.130 278.950 ;
        RECT 38.730 278.650 40.180 278.900 ;
        RECT 40.330 278.800 49.130 278.900 ;
        RECT 38.730 278.450 42.930 278.650 ;
        RECT 26.530 278.300 34.080 278.450 ;
        RECT 35.430 278.300 42.930 278.450 ;
        RECT 26.530 278.000 30.730 278.300 ;
        RECT 26.530 275.150 26.680 278.000 ;
        RECT 27.130 270.450 27.280 278.000 ;
        RECT 27.730 270.450 27.880 278.000 ;
        RECT 28.330 270.450 28.480 278.000 ;
        RECT 28.930 270.450 29.080 278.000 ;
        RECT 29.530 270.450 29.680 278.000 ;
        RECT 30.130 277.850 30.730 278.000 ;
        RECT 38.730 278.000 42.930 278.300 ;
        RECT 38.730 277.850 39.330 278.000 ;
        RECT 30.130 277.700 34.080 277.850 ;
        RECT 35.380 277.700 39.330 277.850 ;
        RECT 30.130 277.250 30.730 277.700 ;
        RECT 38.730 277.250 39.330 277.700 ;
        RECT 30.130 277.100 34.080 277.250 ;
        RECT 35.380 277.100 39.330 277.250 ;
        RECT 30.130 276.650 30.730 277.100 ;
        RECT 38.730 276.650 39.330 277.100 ;
        RECT 30.130 276.500 34.080 276.650 ;
        RECT 35.380 276.500 39.330 276.650 ;
        RECT 30.130 276.050 30.730 276.500 ;
        RECT 38.730 276.050 39.330 276.500 ;
        RECT 30.130 275.900 34.080 276.050 ;
        RECT 35.380 275.900 39.330 276.050 ;
        RECT 30.130 275.450 30.730 275.900 ;
        RECT 38.730 275.450 39.330 275.900 ;
        RECT 30.130 275.300 34.080 275.450 ;
        RECT 35.380 275.300 39.330 275.450 ;
        RECT 30.130 274.850 30.730 275.300 ;
        RECT 38.730 274.850 39.330 275.300 ;
        RECT 30.130 274.700 34.080 274.850 ;
        RECT 35.380 274.700 39.330 274.850 ;
        RECT 30.130 274.250 30.730 274.700 ;
        RECT 38.730 274.250 39.330 274.700 ;
        RECT 30.130 274.100 34.080 274.250 ;
        RECT 35.380 274.100 39.330 274.250 ;
        RECT 30.130 273.650 30.730 274.100 ;
        RECT 38.730 273.650 39.330 274.100 ;
        RECT 30.130 273.500 34.080 273.650 ;
        RECT 35.380 273.500 39.330 273.650 ;
        RECT 30.130 273.050 30.730 273.500 ;
        RECT 38.730 273.050 39.330 273.500 ;
        RECT 30.130 272.900 34.080 273.050 ;
        RECT 35.380 272.900 39.330 273.050 ;
        RECT 30.130 272.450 30.730 272.900 ;
        RECT 38.730 272.450 39.330 272.900 ;
        RECT 30.130 272.300 34.080 272.450 ;
        RECT 35.380 272.300 39.330 272.450 ;
        RECT 30.130 271.850 30.730 272.300 ;
        RECT 38.730 271.850 39.330 272.300 ;
        RECT 30.130 271.700 34.080 271.850 ;
        RECT 35.380 271.700 39.330 271.850 ;
        RECT 30.130 271.250 30.730 271.700 ;
        RECT 38.730 271.250 39.330 271.700 ;
        RECT 30.130 271.100 34.080 271.250 ;
        RECT 35.380 271.100 39.330 271.250 ;
        RECT 30.130 270.650 30.730 271.100 ;
        RECT 38.730 270.650 39.330 271.100 ;
        RECT 30.130 270.450 34.080 270.650 ;
        RECT 35.380 270.450 39.330 270.650 ;
        RECT 39.780 270.450 39.930 278.000 ;
        RECT 40.380 270.450 40.530 278.000 ;
        RECT 40.980 270.450 41.130 278.000 ;
        RECT 41.580 270.450 41.730 278.000 ;
        RECT 42.180 270.450 42.330 278.000 ;
        RECT 42.780 275.150 42.930 278.000 ;
        RECT 43.530 275.600 45.930 278.800 ;
        RECT 49.280 278.650 50.730 278.950 ;
        RECT 46.530 278.450 50.730 278.650 ;
        RECT 58.730 278.950 70.730 279.800 ;
        RECT 58.730 278.900 69.130 278.950 ;
        RECT 58.730 278.650 60.180 278.900 ;
        RECT 60.330 278.800 69.130 278.900 ;
        RECT 58.730 278.450 62.930 278.650 ;
        RECT 46.530 278.300 54.080 278.450 ;
        RECT 55.430 278.300 62.930 278.450 ;
        RECT 46.530 278.000 50.730 278.300 ;
        RECT 46.530 275.150 46.680 278.000 ;
        RECT 47.130 270.450 47.280 278.000 ;
        RECT 47.730 270.450 47.880 278.000 ;
        RECT 48.330 270.450 48.480 278.000 ;
        RECT 48.930 270.450 49.080 278.000 ;
        RECT 49.530 270.450 49.680 278.000 ;
        RECT 50.130 277.850 50.730 278.000 ;
        RECT 58.730 278.000 62.930 278.300 ;
        RECT 58.730 277.850 59.330 278.000 ;
        RECT 50.130 277.700 54.080 277.850 ;
        RECT 55.380 277.700 59.330 277.850 ;
        RECT 50.130 277.250 50.730 277.700 ;
        RECT 58.730 277.250 59.330 277.700 ;
        RECT 50.130 277.100 54.080 277.250 ;
        RECT 55.380 277.100 59.330 277.250 ;
        RECT 50.130 276.650 50.730 277.100 ;
        RECT 58.730 276.650 59.330 277.100 ;
        RECT 50.130 276.500 54.080 276.650 ;
        RECT 55.380 276.500 59.330 276.650 ;
        RECT 50.130 276.050 50.730 276.500 ;
        RECT 58.730 276.050 59.330 276.500 ;
        RECT 50.130 275.900 54.080 276.050 ;
        RECT 55.380 275.900 59.330 276.050 ;
        RECT 50.130 275.450 50.730 275.900 ;
        RECT 58.730 275.450 59.330 275.900 ;
        RECT 50.130 275.300 54.080 275.450 ;
        RECT 55.380 275.300 59.330 275.450 ;
        RECT 50.130 274.850 50.730 275.300 ;
        RECT 58.730 274.850 59.330 275.300 ;
        RECT 50.130 274.700 54.080 274.850 ;
        RECT 55.380 274.700 59.330 274.850 ;
        RECT 50.130 274.250 50.730 274.700 ;
        RECT 58.730 274.250 59.330 274.700 ;
        RECT 50.130 274.100 54.080 274.250 ;
        RECT 55.380 274.100 59.330 274.250 ;
        RECT 50.130 273.650 50.730 274.100 ;
        RECT 58.730 273.650 59.330 274.100 ;
        RECT 50.130 273.500 54.080 273.650 ;
        RECT 55.380 273.500 59.330 273.650 ;
        RECT 50.130 273.050 50.730 273.500 ;
        RECT 58.730 273.050 59.330 273.500 ;
        RECT 50.130 272.900 54.080 273.050 ;
        RECT 55.380 272.900 59.330 273.050 ;
        RECT 50.130 272.450 50.730 272.900 ;
        RECT 58.730 272.450 59.330 272.900 ;
        RECT 50.130 272.300 54.080 272.450 ;
        RECT 55.380 272.300 59.330 272.450 ;
        RECT 50.130 271.850 50.730 272.300 ;
        RECT 58.730 271.850 59.330 272.300 ;
        RECT 50.130 271.700 54.080 271.850 ;
        RECT 55.380 271.700 59.330 271.850 ;
        RECT 50.130 271.250 50.730 271.700 ;
        RECT 58.730 271.250 59.330 271.700 ;
        RECT 50.130 271.100 54.080 271.250 ;
        RECT 55.380 271.100 59.330 271.250 ;
        RECT 50.130 270.650 50.730 271.100 ;
        RECT 58.730 270.650 59.330 271.100 ;
        RECT 50.130 270.450 54.080 270.650 ;
        RECT 55.380 270.450 59.330 270.650 ;
        RECT 59.780 270.450 59.930 278.000 ;
        RECT 60.380 270.450 60.530 278.000 ;
        RECT 60.980 270.450 61.130 278.000 ;
        RECT 61.580 270.450 61.730 278.000 ;
        RECT 62.180 270.450 62.330 278.000 ;
        RECT 62.780 275.150 62.930 278.000 ;
        RECT 63.530 275.600 65.930 278.800 ;
        RECT 69.280 278.650 70.730 278.950 ;
        RECT 66.530 278.450 70.730 278.650 ;
        RECT 78.730 278.950 90.730 279.800 ;
        RECT 78.730 278.900 89.130 278.950 ;
        RECT 78.730 278.650 80.180 278.900 ;
        RECT 80.330 278.800 89.130 278.900 ;
        RECT 78.730 278.450 82.930 278.650 ;
        RECT 66.530 278.300 74.080 278.450 ;
        RECT 75.430 278.300 82.930 278.450 ;
        RECT 66.530 278.000 70.730 278.300 ;
        RECT 66.530 275.150 66.680 278.000 ;
        RECT 67.130 270.450 67.280 278.000 ;
        RECT 67.730 270.450 67.880 278.000 ;
        RECT 68.330 270.450 68.480 278.000 ;
        RECT 68.930 270.450 69.080 278.000 ;
        RECT 69.530 270.450 69.680 278.000 ;
        RECT 70.130 277.850 70.730 278.000 ;
        RECT 78.730 278.000 82.930 278.300 ;
        RECT 78.730 277.850 79.330 278.000 ;
        RECT 70.130 277.700 74.080 277.850 ;
        RECT 75.380 277.700 79.330 277.850 ;
        RECT 70.130 277.250 70.730 277.700 ;
        RECT 78.730 277.250 79.330 277.700 ;
        RECT 70.130 277.100 74.080 277.250 ;
        RECT 75.380 277.100 79.330 277.250 ;
        RECT 70.130 276.650 70.730 277.100 ;
        RECT 78.730 276.650 79.330 277.100 ;
        RECT 70.130 276.500 74.080 276.650 ;
        RECT 75.380 276.500 79.330 276.650 ;
        RECT 70.130 276.050 70.730 276.500 ;
        RECT 78.730 276.050 79.330 276.500 ;
        RECT 70.130 275.900 74.080 276.050 ;
        RECT 75.380 275.900 79.330 276.050 ;
        RECT 70.130 275.450 70.730 275.900 ;
        RECT 78.730 275.450 79.330 275.900 ;
        RECT 70.130 275.300 74.080 275.450 ;
        RECT 75.380 275.300 79.330 275.450 ;
        RECT 70.130 274.850 70.730 275.300 ;
        RECT 78.730 274.850 79.330 275.300 ;
        RECT 70.130 274.700 74.080 274.850 ;
        RECT 75.380 274.700 79.330 274.850 ;
        RECT 70.130 274.250 70.730 274.700 ;
        RECT 78.730 274.250 79.330 274.700 ;
        RECT 70.130 274.100 74.080 274.250 ;
        RECT 75.380 274.100 79.330 274.250 ;
        RECT 70.130 273.650 70.730 274.100 ;
        RECT 78.730 273.650 79.330 274.100 ;
        RECT 70.130 273.500 74.080 273.650 ;
        RECT 75.380 273.500 79.330 273.650 ;
        RECT 70.130 273.050 70.730 273.500 ;
        RECT 78.730 273.050 79.330 273.500 ;
        RECT 70.130 272.900 74.080 273.050 ;
        RECT 75.380 272.900 79.330 273.050 ;
        RECT 70.130 272.450 70.730 272.900 ;
        RECT 78.730 272.450 79.330 272.900 ;
        RECT 70.130 272.300 74.080 272.450 ;
        RECT 75.380 272.300 79.330 272.450 ;
        RECT 70.130 271.850 70.730 272.300 ;
        RECT 78.730 271.850 79.330 272.300 ;
        RECT 70.130 271.700 74.080 271.850 ;
        RECT 75.380 271.700 79.330 271.850 ;
        RECT 70.130 271.250 70.730 271.700 ;
        RECT 78.730 271.250 79.330 271.700 ;
        RECT 70.130 271.100 74.080 271.250 ;
        RECT 75.380 271.100 79.330 271.250 ;
        RECT 70.130 270.650 70.730 271.100 ;
        RECT 78.730 270.650 79.330 271.100 ;
        RECT 70.130 270.450 74.080 270.650 ;
        RECT 75.380 270.450 79.330 270.650 ;
        RECT 79.780 270.450 79.930 278.000 ;
        RECT 80.380 270.450 80.530 278.000 ;
        RECT 80.980 270.450 81.130 278.000 ;
        RECT 81.580 270.450 81.730 278.000 ;
        RECT 82.180 270.450 82.330 278.000 ;
        RECT 82.780 275.150 82.930 278.000 ;
        RECT 83.530 275.600 85.930 278.800 ;
        RECT 89.280 278.650 90.730 278.950 ;
        RECT 86.530 278.450 90.730 278.650 ;
        RECT 98.730 278.950 110.730 279.800 ;
        RECT 98.730 278.900 109.130 278.950 ;
        RECT 98.730 278.650 100.180 278.900 ;
        RECT 100.330 278.800 109.130 278.900 ;
        RECT 98.730 278.450 102.930 278.650 ;
        RECT 86.530 278.300 94.080 278.450 ;
        RECT 95.430 278.300 102.930 278.450 ;
        RECT 86.530 278.000 90.730 278.300 ;
        RECT 86.530 275.150 86.680 278.000 ;
        RECT 87.130 270.450 87.280 278.000 ;
        RECT 87.730 270.450 87.880 278.000 ;
        RECT 88.330 270.450 88.480 278.000 ;
        RECT 88.930 270.450 89.080 278.000 ;
        RECT 89.530 270.450 89.680 278.000 ;
        RECT 90.130 277.850 90.730 278.000 ;
        RECT 98.730 278.000 102.930 278.300 ;
        RECT 98.730 277.850 99.330 278.000 ;
        RECT 90.130 277.700 94.080 277.850 ;
        RECT 95.380 277.700 99.330 277.850 ;
        RECT 90.130 277.250 90.730 277.700 ;
        RECT 98.730 277.250 99.330 277.700 ;
        RECT 90.130 277.100 94.080 277.250 ;
        RECT 95.380 277.100 99.330 277.250 ;
        RECT 90.130 276.650 90.730 277.100 ;
        RECT 98.730 276.650 99.330 277.100 ;
        RECT 90.130 276.500 94.080 276.650 ;
        RECT 95.380 276.500 99.330 276.650 ;
        RECT 90.130 276.050 90.730 276.500 ;
        RECT 98.730 276.050 99.330 276.500 ;
        RECT 90.130 275.900 94.080 276.050 ;
        RECT 95.380 275.900 99.330 276.050 ;
        RECT 90.130 275.450 90.730 275.900 ;
        RECT 98.730 275.450 99.330 275.900 ;
        RECT 90.130 275.300 94.080 275.450 ;
        RECT 95.380 275.300 99.330 275.450 ;
        RECT 90.130 274.850 90.730 275.300 ;
        RECT 98.730 274.850 99.330 275.300 ;
        RECT 90.130 274.700 94.080 274.850 ;
        RECT 95.380 274.700 99.330 274.850 ;
        RECT 90.130 274.250 90.730 274.700 ;
        RECT 98.730 274.250 99.330 274.700 ;
        RECT 90.130 274.100 94.080 274.250 ;
        RECT 95.380 274.100 99.330 274.250 ;
        RECT 90.130 273.650 90.730 274.100 ;
        RECT 98.730 273.650 99.330 274.100 ;
        RECT 90.130 273.500 94.080 273.650 ;
        RECT 95.380 273.500 99.330 273.650 ;
        RECT 90.130 273.050 90.730 273.500 ;
        RECT 98.730 273.050 99.330 273.500 ;
        RECT 90.130 272.900 94.080 273.050 ;
        RECT 95.380 272.900 99.330 273.050 ;
        RECT 90.130 272.450 90.730 272.900 ;
        RECT 98.730 272.450 99.330 272.900 ;
        RECT 90.130 272.300 94.080 272.450 ;
        RECT 95.380 272.300 99.330 272.450 ;
        RECT 90.130 271.850 90.730 272.300 ;
        RECT 98.730 271.850 99.330 272.300 ;
        RECT 90.130 271.700 94.080 271.850 ;
        RECT 95.380 271.700 99.330 271.850 ;
        RECT 90.130 271.250 90.730 271.700 ;
        RECT 98.730 271.250 99.330 271.700 ;
        RECT 90.130 271.100 94.080 271.250 ;
        RECT 95.380 271.100 99.330 271.250 ;
        RECT 90.130 270.650 90.730 271.100 ;
        RECT 98.730 270.650 99.330 271.100 ;
        RECT 90.130 270.450 94.080 270.650 ;
        RECT 95.380 270.450 99.330 270.650 ;
        RECT 99.780 270.450 99.930 278.000 ;
        RECT 100.380 270.450 100.530 278.000 ;
        RECT 100.980 270.450 101.130 278.000 ;
        RECT 101.580 270.450 101.730 278.000 ;
        RECT 102.180 270.450 102.330 278.000 ;
        RECT 102.780 275.150 102.930 278.000 ;
        RECT 103.530 275.600 105.930 278.800 ;
        RECT 109.280 278.650 110.730 278.950 ;
        RECT 106.530 278.450 110.730 278.650 ;
        RECT 118.730 278.900 124.730 279.800 ;
        RECT 118.730 278.650 120.180 278.900 ;
        RECT 120.330 278.800 124.730 278.900 ;
        RECT 118.730 278.450 122.930 278.650 ;
        RECT 106.530 278.300 114.080 278.450 ;
        RECT 115.430 278.300 122.930 278.450 ;
        RECT 106.530 278.000 110.730 278.300 ;
        RECT 106.530 275.150 106.680 278.000 ;
        RECT 107.130 270.450 107.280 278.000 ;
        RECT 107.730 270.450 107.880 278.000 ;
        RECT 108.330 270.450 108.480 278.000 ;
        RECT 108.930 270.450 109.080 278.000 ;
        RECT 109.530 270.450 109.680 278.000 ;
        RECT 110.130 277.850 110.730 278.000 ;
        RECT 118.730 278.000 122.930 278.300 ;
        RECT 118.730 277.850 119.330 278.000 ;
        RECT 110.130 277.700 114.080 277.850 ;
        RECT 115.380 277.700 119.330 277.850 ;
        RECT 110.130 277.250 110.730 277.700 ;
        RECT 118.730 277.250 119.330 277.700 ;
        RECT 110.130 277.100 114.080 277.250 ;
        RECT 115.380 277.100 119.330 277.250 ;
        RECT 110.130 276.650 110.730 277.100 ;
        RECT 118.730 276.650 119.330 277.100 ;
        RECT 110.130 276.500 114.080 276.650 ;
        RECT 115.380 276.500 119.330 276.650 ;
        RECT 110.130 276.050 110.730 276.500 ;
        RECT 118.730 276.050 119.330 276.500 ;
        RECT 110.130 275.900 114.080 276.050 ;
        RECT 115.380 275.900 119.330 276.050 ;
        RECT 110.130 275.450 110.730 275.900 ;
        RECT 118.730 275.450 119.330 275.900 ;
        RECT 110.130 275.300 114.080 275.450 ;
        RECT 115.380 275.300 119.330 275.450 ;
        RECT 110.130 274.850 110.730 275.300 ;
        RECT 118.730 274.850 119.330 275.300 ;
        RECT 110.130 274.700 114.080 274.850 ;
        RECT 115.380 274.700 119.330 274.850 ;
        RECT 110.130 274.250 110.730 274.700 ;
        RECT 118.730 274.250 119.330 274.700 ;
        RECT 110.130 274.100 114.080 274.250 ;
        RECT 115.380 274.100 119.330 274.250 ;
        RECT 110.130 273.650 110.730 274.100 ;
        RECT 118.730 273.650 119.330 274.100 ;
        RECT 110.130 273.500 114.080 273.650 ;
        RECT 115.380 273.500 119.330 273.650 ;
        RECT 110.130 273.050 110.730 273.500 ;
        RECT 118.730 273.050 119.330 273.500 ;
        RECT 110.130 272.900 114.080 273.050 ;
        RECT 115.380 272.900 119.330 273.050 ;
        RECT 110.130 272.450 110.730 272.900 ;
        RECT 118.730 272.450 119.330 272.900 ;
        RECT 110.130 272.300 114.080 272.450 ;
        RECT 115.380 272.300 119.330 272.450 ;
        RECT 110.130 271.850 110.730 272.300 ;
        RECT 118.730 271.850 119.330 272.300 ;
        RECT 110.130 271.700 114.080 271.850 ;
        RECT 115.380 271.700 119.330 271.850 ;
        RECT 110.130 271.250 110.730 271.700 ;
        RECT 118.730 271.250 119.330 271.700 ;
        RECT 110.130 271.100 114.080 271.250 ;
        RECT 115.380 271.100 119.330 271.250 ;
        RECT 110.130 270.650 110.730 271.100 ;
        RECT 118.730 270.650 119.330 271.100 ;
        RECT 110.130 270.450 114.080 270.650 ;
        RECT 115.380 270.450 119.330 270.650 ;
        RECT 119.780 270.450 119.930 278.000 ;
        RECT 120.380 270.450 120.530 278.000 ;
        RECT 120.980 270.450 121.130 278.000 ;
        RECT 121.580 270.450 121.730 278.000 ;
        RECT 122.180 270.450 122.330 278.000 ;
        RECT 122.780 275.150 122.930 278.000 ;
        RECT 123.530 277.855 124.730 278.800 ;
        RECT 123.530 276.580 127.135 277.855 ;
        RECT 123.530 275.600 124.730 276.580 ;
        RECT 2.315 264.445 4.315 266.740 ;
        RECT 4.730 263.645 5.930 264.400 ;
        RECT 2.315 262.370 5.930 263.645 ;
        RECT 4.730 261.200 5.930 262.370 ;
        RECT 6.530 262.000 6.680 264.900 ;
        RECT 7.130 262.000 7.280 269.550 ;
        RECT 7.730 262.000 7.880 269.550 ;
        RECT 8.330 262.000 8.480 269.550 ;
        RECT 8.930 262.000 9.080 269.550 ;
        RECT 9.530 262.000 9.680 269.550 ;
        RECT 10.130 269.350 14.080 269.550 ;
        RECT 15.380 269.350 19.330 269.550 ;
        RECT 10.130 268.900 10.730 269.350 ;
        RECT 18.730 268.900 19.330 269.350 ;
        RECT 10.130 268.750 14.080 268.900 ;
        RECT 15.380 268.750 19.330 268.900 ;
        RECT 10.130 268.300 10.730 268.750 ;
        RECT 18.730 268.300 19.330 268.750 ;
        RECT 10.130 268.150 14.080 268.300 ;
        RECT 15.380 268.150 19.330 268.300 ;
        RECT 10.130 267.700 10.730 268.150 ;
        RECT 18.730 267.700 19.330 268.150 ;
        RECT 10.130 267.550 14.080 267.700 ;
        RECT 15.380 267.550 19.330 267.700 ;
        RECT 10.130 267.100 10.730 267.550 ;
        RECT 18.730 267.100 19.330 267.550 ;
        RECT 10.130 266.950 14.080 267.100 ;
        RECT 15.380 266.950 19.330 267.100 ;
        RECT 10.130 266.500 10.730 266.950 ;
        RECT 18.730 266.500 19.330 266.950 ;
        RECT 10.130 266.350 14.080 266.500 ;
        RECT 15.380 266.350 19.330 266.500 ;
        RECT 10.130 265.900 10.730 266.350 ;
        RECT 18.730 265.900 19.330 266.350 ;
        RECT 10.130 265.750 14.080 265.900 ;
        RECT 15.380 265.750 19.330 265.900 ;
        RECT 10.130 265.300 10.730 265.750 ;
        RECT 18.730 265.300 19.330 265.750 ;
        RECT 10.130 265.150 14.080 265.300 ;
        RECT 15.380 265.150 19.330 265.300 ;
        RECT 10.130 264.700 10.730 265.150 ;
        RECT 18.730 264.700 19.330 265.150 ;
        RECT 10.130 264.550 14.080 264.700 ;
        RECT 15.380 264.550 19.330 264.700 ;
        RECT 10.130 264.100 10.730 264.550 ;
        RECT 18.730 264.100 19.330 264.550 ;
        RECT 10.130 263.950 14.080 264.100 ;
        RECT 15.380 263.950 19.330 264.100 ;
        RECT 10.130 263.500 10.730 263.950 ;
        RECT 18.730 263.500 19.330 263.950 ;
        RECT 10.130 263.350 14.080 263.500 ;
        RECT 15.380 263.350 19.330 263.500 ;
        RECT 10.130 262.900 10.730 263.350 ;
        RECT 18.730 262.900 19.330 263.350 ;
        RECT 10.130 262.750 14.080 262.900 ;
        RECT 15.380 262.750 19.330 262.900 ;
        RECT 10.130 262.300 10.730 262.750 ;
        RECT 18.730 262.300 19.330 262.750 ;
        RECT 10.130 262.150 14.080 262.300 ;
        RECT 15.380 262.150 19.330 262.300 ;
        RECT 10.130 262.000 10.730 262.150 ;
        RECT 6.530 261.700 10.730 262.000 ;
        RECT 18.730 262.000 19.330 262.150 ;
        RECT 19.780 262.000 19.930 269.550 ;
        RECT 20.380 262.000 20.530 269.550 ;
        RECT 20.980 262.000 21.130 269.550 ;
        RECT 21.580 262.000 21.730 269.550 ;
        RECT 22.180 262.000 22.330 269.550 ;
        RECT 22.780 262.000 22.930 264.900 ;
        RECT 18.730 261.700 22.930 262.000 ;
        RECT 6.530 261.550 14.080 261.700 ;
        RECT 15.380 261.550 22.930 261.700 ;
        RECT 6.530 261.350 10.730 261.550 ;
        RECT 4.730 261.050 9.130 261.200 ;
        RECT 9.280 261.050 10.730 261.350 ;
        RECT 4.730 260.150 10.730 261.050 ;
        RECT 18.730 261.350 22.930 261.550 ;
        RECT 18.730 261.050 20.180 261.350 ;
        RECT 23.530 261.200 25.930 264.400 ;
        RECT 26.530 262.000 26.680 264.900 ;
        RECT 27.130 262.000 27.280 269.550 ;
        RECT 27.730 262.000 27.880 269.550 ;
        RECT 28.330 262.000 28.480 269.550 ;
        RECT 28.930 262.000 29.080 269.550 ;
        RECT 29.530 262.000 29.680 269.550 ;
        RECT 30.130 269.350 34.080 269.550 ;
        RECT 35.380 269.350 39.330 269.550 ;
        RECT 30.130 268.900 30.730 269.350 ;
        RECT 38.730 268.900 39.330 269.350 ;
        RECT 30.130 268.750 34.080 268.900 ;
        RECT 35.380 268.750 39.330 268.900 ;
        RECT 30.130 268.300 30.730 268.750 ;
        RECT 38.730 268.300 39.330 268.750 ;
        RECT 30.130 268.150 34.080 268.300 ;
        RECT 35.380 268.150 39.330 268.300 ;
        RECT 30.130 267.700 30.730 268.150 ;
        RECT 38.730 267.700 39.330 268.150 ;
        RECT 30.130 267.550 34.080 267.700 ;
        RECT 35.380 267.550 39.330 267.700 ;
        RECT 30.130 267.100 30.730 267.550 ;
        RECT 38.730 267.100 39.330 267.550 ;
        RECT 30.130 266.950 34.080 267.100 ;
        RECT 35.380 266.950 39.330 267.100 ;
        RECT 30.130 266.500 30.730 266.950 ;
        RECT 38.730 266.500 39.330 266.950 ;
        RECT 30.130 266.350 34.080 266.500 ;
        RECT 35.380 266.350 39.330 266.500 ;
        RECT 30.130 265.900 30.730 266.350 ;
        RECT 38.730 265.900 39.330 266.350 ;
        RECT 30.130 265.750 34.080 265.900 ;
        RECT 35.380 265.750 39.330 265.900 ;
        RECT 30.130 265.300 30.730 265.750 ;
        RECT 38.730 265.300 39.330 265.750 ;
        RECT 30.130 265.150 34.080 265.300 ;
        RECT 35.380 265.150 39.330 265.300 ;
        RECT 30.130 264.700 30.730 265.150 ;
        RECT 38.730 264.700 39.330 265.150 ;
        RECT 30.130 264.550 34.080 264.700 ;
        RECT 35.380 264.550 39.330 264.700 ;
        RECT 30.130 264.100 30.730 264.550 ;
        RECT 38.730 264.100 39.330 264.550 ;
        RECT 30.130 263.950 34.080 264.100 ;
        RECT 35.380 263.950 39.330 264.100 ;
        RECT 30.130 263.500 30.730 263.950 ;
        RECT 38.730 263.500 39.330 263.950 ;
        RECT 30.130 263.350 34.080 263.500 ;
        RECT 35.380 263.350 39.330 263.500 ;
        RECT 30.130 262.900 30.730 263.350 ;
        RECT 38.730 262.900 39.330 263.350 ;
        RECT 30.130 262.750 34.080 262.900 ;
        RECT 35.380 262.750 39.330 262.900 ;
        RECT 30.130 262.300 30.730 262.750 ;
        RECT 38.730 262.300 39.330 262.750 ;
        RECT 30.130 262.150 34.080 262.300 ;
        RECT 35.380 262.150 39.330 262.300 ;
        RECT 30.130 262.000 30.730 262.150 ;
        RECT 26.530 261.700 30.730 262.000 ;
        RECT 38.730 262.000 39.330 262.150 ;
        RECT 39.780 262.000 39.930 269.550 ;
        RECT 40.380 262.000 40.530 269.550 ;
        RECT 40.980 262.000 41.130 269.550 ;
        RECT 41.580 262.000 41.730 269.550 ;
        RECT 42.180 262.000 42.330 269.550 ;
        RECT 42.780 262.000 42.930 264.900 ;
        RECT 38.730 261.700 42.930 262.000 ;
        RECT 26.530 261.550 34.080 261.700 ;
        RECT 35.380 261.550 42.930 261.700 ;
        RECT 26.530 261.350 30.730 261.550 ;
        RECT 20.330 261.050 29.130 261.200 ;
        RECT 29.280 261.050 30.730 261.350 ;
        RECT 18.730 260.150 30.730 261.050 ;
        RECT 38.730 261.350 42.930 261.550 ;
        RECT 38.730 261.050 40.180 261.350 ;
        RECT 43.530 261.200 45.930 264.400 ;
        RECT 46.530 262.000 46.680 264.900 ;
        RECT 47.130 262.000 47.280 269.550 ;
        RECT 47.730 262.000 47.880 269.550 ;
        RECT 48.330 262.000 48.480 269.550 ;
        RECT 48.930 262.000 49.080 269.550 ;
        RECT 49.530 262.000 49.680 269.550 ;
        RECT 50.130 269.350 54.080 269.550 ;
        RECT 55.380 269.350 59.330 269.550 ;
        RECT 50.130 268.900 50.730 269.350 ;
        RECT 58.730 268.900 59.330 269.350 ;
        RECT 50.130 268.750 54.080 268.900 ;
        RECT 55.380 268.750 59.330 268.900 ;
        RECT 50.130 268.300 50.730 268.750 ;
        RECT 58.730 268.300 59.330 268.750 ;
        RECT 50.130 268.150 54.080 268.300 ;
        RECT 55.380 268.150 59.330 268.300 ;
        RECT 50.130 267.700 50.730 268.150 ;
        RECT 58.730 267.700 59.330 268.150 ;
        RECT 50.130 267.550 54.080 267.700 ;
        RECT 55.380 267.550 59.330 267.700 ;
        RECT 50.130 267.100 50.730 267.550 ;
        RECT 58.730 267.100 59.330 267.550 ;
        RECT 50.130 266.950 54.080 267.100 ;
        RECT 55.380 266.950 59.330 267.100 ;
        RECT 50.130 266.500 50.730 266.950 ;
        RECT 58.730 266.500 59.330 266.950 ;
        RECT 50.130 266.350 54.080 266.500 ;
        RECT 55.380 266.350 59.330 266.500 ;
        RECT 50.130 265.900 50.730 266.350 ;
        RECT 58.730 265.900 59.330 266.350 ;
        RECT 50.130 265.750 54.080 265.900 ;
        RECT 55.380 265.750 59.330 265.900 ;
        RECT 50.130 265.300 50.730 265.750 ;
        RECT 58.730 265.300 59.330 265.750 ;
        RECT 50.130 265.150 54.080 265.300 ;
        RECT 55.380 265.150 59.330 265.300 ;
        RECT 50.130 264.700 50.730 265.150 ;
        RECT 58.730 264.700 59.330 265.150 ;
        RECT 50.130 264.550 54.080 264.700 ;
        RECT 55.380 264.550 59.330 264.700 ;
        RECT 50.130 264.100 50.730 264.550 ;
        RECT 58.730 264.100 59.330 264.550 ;
        RECT 50.130 263.950 54.080 264.100 ;
        RECT 55.380 263.950 59.330 264.100 ;
        RECT 50.130 263.500 50.730 263.950 ;
        RECT 58.730 263.500 59.330 263.950 ;
        RECT 50.130 263.350 54.080 263.500 ;
        RECT 55.380 263.350 59.330 263.500 ;
        RECT 50.130 262.900 50.730 263.350 ;
        RECT 58.730 262.900 59.330 263.350 ;
        RECT 50.130 262.750 54.080 262.900 ;
        RECT 55.380 262.750 59.330 262.900 ;
        RECT 50.130 262.300 50.730 262.750 ;
        RECT 58.730 262.300 59.330 262.750 ;
        RECT 50.130 262.150 54.080 262.300 ;
        RECT 55.380 262.150 59.330 262.300 ;
        RECT 50.130 262.000 50.730 262.150 ;
        RECT 46.530 261.700 50.730 262.000 ;
        RECT 58.730 262.000 59.330 262.150 ;
        RECT 59.780 262.000 59.930 269.550 ;
        RECT 60.380 262.000 60.530 269.550 ;
        RECT 60.980 262.000 61.130 269.550 ;
        RECT 61.580 262.000 61.730 269.550 ;
        RECT 62.180 262.000 62.330 269.550 ;
        RECT 62.780 262.000 62.930 264.900 ;
        RECT 58.730 261.700 62.930 262.000 ;
        RECT 46.530 261.550 54.080 261.700 ;
        RECT 55.380 261.550 62.930 261.700 ;
        RECT 46.530 261.350 50.730 261.550 ;
        RECT 40.330 261.050 49.130 261.200 ;
        RECT 49.280 261.050 50.730 261.350 ;
        RECT 38.730 260.150 50.730 261.050 ;
        RECT 58.730 261.350 62.930 261.550 ;
        RECT 58.730 261.050 60.180 261.350 ;
        RECT 63.530 261.200 65.930 264.400 ;
        RECT 66.530 262.000 66.680 264.900 ;
        RECT 67.130 262.000 67.280 269.550 ;
        RECT 67.730 262.000 67.880 269.550 ;
        RECT 68.330 262.000 68.480 269.550 ;
        RECT 68.930 262.000 69.080 269.550 ;
        RECT 69.530 262.000 69.680 269.550 ;
        RECT 70.130 269.350 74.080 269.550 ;
        RECT 75.380 269.350 79.330 269.550 ;
        RECT 70.130 268.900 70.730 269.350 ;
        RECT 78.730 268.900 79.330 269.350 ;
        RECT 70.130 268.750 74.080 268.900 ;
        RECT 75.380 268.750 79.330 268.900 ;
        RECT 70.130 268.300 70.730 268.750 ;
        RECT 78.730 268.300 79.330 268.750 ;
        RECT 70.130 268.150 74.080 268.300 ;
        RECT 75.380 268.150 79.330 268.300 ;
        RECT 70.130 267.700 70.730 268.150 ;
        RECT 78.730 267.700 79.330 268.150 ;
        RECT 70.130 267.550 74.080 267.700 ;
        RECT 75.380 267.550 79.330 267.700 ;
        RECT 70.130 267.100 70.730 267.550 ;
        RECT 78.730 267.100 79.330 267.550 ;
        RECT 70.130 266.950 74.080 267.100 ;
        RECT 75.380 266.950 79.330 267.100 ;
        RECT 70.130 266.500 70.730 266.950 ;
        RECT 78.730 266.500 79.330 266.950 ;
        RECT 70.130 266.350 74.080 266.500 ;
        RECT 75.380 266.350 79.330 266.500 ;
        RECT 70.130 265.900 70.730 266.350 ;
        RECT 78.730 265.900 79.330 266.350 ;
        RECT 70.130 265.750 74.080 265.900 ;
        RECT 75.380 265.750 79.330 265.900 ;
        RECT 70.130 265.300 70.730 265.750 ;
        RECT 78.730 265.300 79.330 265.750 ;
        RECT 70.130 265.150 74.080 265.300 ;
        RECT 75.380 265.150 79.330 265.300 ;
        RECT 70.130 264.700 70.730 265.150 ;
        RECT 78.730 264.700 79.330 265.150 ;
        RECT 70.130 264.550 74.080 264.700 ;
        RECT 75.380 264.550 79.330 264.700 ;
        RECT 70.130 264.100 70.730 264.550 ;
        RECT 78.730 264.100 79.330 264.550 ;
        RECT 70.130 263.950 74.080 264.100 ;
        RECT 75.380 263.950 79.330 264.100 ;
        RECT 70.130 263.500 70.730 263.950 ;
        RECT 78.730 263.500 79.330 263.950 ;
        RECT 70.130 263.350 74.080 263.500 ;
        RECT 75.380 263.350 79.330 263.500 ;
        RECT 70.130 262.900 70.730 263.350 ;
        RECT 78.730 262.900 79.330 263.350 ;
        RECT 70.130 262.750 74.080 262.900 ;
        RECT 75.380 262.750 79.330 262.900 ;
        RECT 70.130 262.300 70.730 262.750 ;
        RECT 78.730 262.300 79.330 262.750 ;
        RECT 70.130 262.150 74.080 262.300 ;
        RECT 75.380 262.150 79.330 262.300 ;
        RECT 70.130 262.000 70.730 262.150 ;
        RECT 66.530 261.700 70.730 262.000 ;
        RECT 78.730 262.000 79.330 262.150 ;
        RECT 79.780 262.000 79.930 269.550 ;
        RECT 80.380 262.000 80.530 269.550 ;
        RECT 80.980 262.000 81.130 269.550 ;
        RECT 81.580 262.000 81.730 269.550 ;
        RECT 82.180 262.000 82.330 269.550 ;
        RECT 82.780 262.000 82.930 264.900 ;
        RECT 78.730 261.700 82.930 262.000 ;
        RECT 66.530 261.550 74.080 261.700 ;
        RECT 75.380 261.550 82.930 261.700 ;
        RECT 66.530 261.350 70.730 261.550 ;
        RECT 60.330 261.050 69.130 261.200 ;
        RECT 69.280 261.050 70.730 261.350 ;
        RECT 58.730 260.150 70.730 261.050 ;
        RECT 78.730 261.350 82.930 261.550 ;
        RECT 78.730 261.050 80.180 261.350 ;
        RECT 83.530 261.200 85.930 264.400 ;
        RECT 86.530 262.000 86.680 264.900 ;
        RECT 87.130 262.000 87.280 269.550 ;
        RECT 87.730 262.000 87.880 269.550 ;
        RECT 88.330 262.000 88.480 269.550 ;
        RECT 88.930 262.000 89.080 269.550 ;
        RECT 89.530 262.000 89.680 269.550 ;
        RECT 90.130 269.350 94.080 269.550 ;
        RECT 95.380 269.350 99.330 269.550 ;
        RECT 90.130 268.900 90.730 269.350 ;
        RECT 98.730 268.900 99.330 269.350 ;
        RECT 90.130 268.750 94.080 268.900 ;
        RECT 95.380 268.750 99.330 268.900 ;
        RECT 90.130 268.300 90.730 268.750 ;
        RECT 98.730 268.300 99.330 268.750 ;
        RECT 90.130 268.150 94.080 268.300 ;
        RECT 95.380 268.150 99.330 268.300 ;
        RECT 90.130 267.700 90.730 268.150 ;
        RECT 98.730 267.700 99.330 268.150 ;
        RECT 90.130 267.550 94.080 267.700 ;
        RECT 95.380 267.550 99.330 267.700 ;
        RECT 90.130 267.100 90.730 267.550 ;
        RECT 98.730 267.100 99.330 267.550 ;
        RECT 90.130 266.950 94.080 267.100 ;
        RECT 95.380 266.950 99.330 267.100 ;
        RECT 90.130 266.500 90.730 266.950 ;
        RECT 98.730 266.500 99.330 266.950 ;
        RECT 90.130 266.350 94.080 266.500 ;
        RECT 95.380 266.350 99.330 266.500 ;
        RECT 90.130 265.900 90.730 266.350 ;
        RECT 98.730 265.900 99.330 266.350 ;
        RECT 90.130 265.750 94.080 265.900 ;
        RECT 95.380 265.750 99.330 265.900 ;
        RECT 90.130 265.300 90.730 265.750 ;
        RECT 98.730 265.300 99.330 265.750 ;
        RECT 90.130 265.150 94.080 265.300 ;
        RECT 95.380 265.150 99.330 265.300 ;
        RECT 90.130 264.700 90.730 265.150 ;
        RECT 98.730 264.700 99.330 265.150 ;
        RECT 90.130 264.550 94.080 264.700 ;
        RECT 95.380 264.550 99.330 264.700 ;
        RECT 90.130 264.100 90.730 264.550 ;
        RECT 98.730 264.100 99.330 264.550 ;
        RECT 90.130 263.950 94.080 264.100 ;
        RECT 95.380 263.950 99.330 264.100 ;
        RECT 90.130 263.500 90.730 263.950 ;
        RECT 98.730 263.500 99.330 263.950 ;
        RECT 90.130 263.350 94.080 263.500 ;
        RECT 95.380 263.350 99.330 263.500 ;
        RECT 90.130 262.900 90.730 263.350 ;
        RECT 98.730 262.900 99.330 263.350 ;
        RECT 90.130 262.750 94.080 262.900 ;
        RECT 95.380 262.750 99.330 262.900 ;
        RECT 90.130 262.300 90.730 262.750 ;
        RECT 98.730 262.300 99.330 262.750 ;
        RECT 90.130 262.150 94.080 262.300 ;
        RECT 95.380 262.150 99.330 262.300 ;
        RECT 90.130 262.000 90.730 262.150 ;
        RECT 86.530 261.700 90.730 262.000 ;
        RECT 98.730 262.000 99.330 262.150 ;
        RECT 99.780 262.000 99.930 269.550 ;
        RECT 100.380 262.000 100.530 269.550 ;
        RECT 100.980 262.000 101.130 269.550 ;
        RECT 101.580 262.000 101.730 269.550 ;
        RECT 102.180 262.000 102.330 269.550 ;
        RECT 102.780 262.000 102.930 264.900 ;
        RECT 98.730 261.700 102.930 262.000 ;
        RECT 86.530 261.550 94.080 261.700 ;
        RECT 95.380 261.550 102.930 261.700 ;
        RECT 86.530 261.350 90.730 261.550 ;
        RECT 80.330 261.050 89.130 261.200 ;
        RECT 89.280 261.050 90.730 261.350 ;
        RECT 78.730 260.150 90.730 261.050 ;
        RECT 98.730 261.350 102.930 261.550 ;
        RECT 98.730 261.050 100.180 261.350 ;
        RECT 103.530 261.200 105.930 264.400 ;
        RECT 106.530 262.000 106.680 264.900 ;
        RECT 107.130 262.000 107.280 269.550 ;
        RECT 107.730 262.000 107.880 269.550 ;
        RECT 108.330 262.000 108.480 269.550 ;
        RECT 108.930 262.000 109.080 269.550 ;
        RECT 109.530 262.000 109.680 269.550 ;
        RECT 110.130 269.350 114.080 269.550 ;
        RECT 115.380 269.350 119.330 269.550 ;
        RECT 110.130 268.900 110.730 269.350 ;
        RECT 118.730 268.900 119.330 269.350 ;
        RECT 110.130 268.750 114.080 268.900 ;
        RECT 115.380 268.750 119.330 268.900 ;
        RECT 110.130 268.300 110.730 268.750 ;
        RECT 118.730 268.300 119.330 268.750 ;
        RECT 110.130 268.150 114.080 268.300 ;
        RECT 115.380 268.150 119.330 268.300 ;
        RECT 110.130 267.700 110.730 268.150 ;
        RECT 118.730 267.700 119.330 268.150 ;
        RECT 110.130 267.550 114.080 267.700 ;
        RECT 115.380 267.550 119.330 267.700 ;
        RECT 110.130 267.100 110.730 267.550 ;
        RECT 118.730 267.100 119.330 267.550 ;
        RECT 110.130 266.950 114.080 267.100 ;
        RECT 115.380 266.950 119.330 267.100 ;
        RECT 110.130 266.500 110.730 266.950 ;
        RECT 118.730 266.500 119.330 266.950 ;
        RECT 110.130 266.350 114.080 266.500 ;
        RECT 115.380 266.350 119.330 266.500 ;
        RECT 110.130 265.900 110.730 266.350 ;
        RECT 118.730 265.900 119.330 266.350 ;
        RECT 110.130 265.750 114.080 265.900 ;
        RECT 115.380 265.750 119.330 265.900 ;
        RECT 110.130 265.300 110.730 265.750 ;
        RECT 118.730 265.300 119.330 265.750 ;
        RECT 110.130 265.150 114.080 265.300 ;
        RECT 115.380 265.150 119.330 265.300 ;
        RECT 110.130 264.700 110.730 265.150 ;
        RECT 118.730 264.700 119.330 265.150 ;
        RECT 110.130 264.550 114.080 264.700 ;
        RECT 115.380 264.550 119.330 264.700 ;
        RECT 110.130 264.100 110.730 264.550 ;
        RECT 118.730 264.100 119.330 264.550 ;
        RECT 110.130 263.950 114.080 264.100 ;
        RECT 115.380 263.950 119.330 264.100 ;
        RECT 110.130 263.500 110.730 263.950 ;
        RECT 118.730 263.500 119.330 263.950 ;
        RECT 110.130 263.350 114.080 263.500 ;
        RECT 115.380 263.350 119.330 263.500 ;
        RECT 110.130 262.900 110.730 263.350 ;
        RECT 118.730 262.900 119.330 263.350 ;
        RECT 110.130 262.750 114.080 262.900 ;
        RECT 115.380 262.750 119.330 262.900 ;
        RECT 110.130 262.300 110.730 262.750 ;
        RECT 118.730 262.300 119.330 262.750 ;
        RECT 110.130 262.150 114.080 262.300 ;
        RECT 115.380 262.150 119.330 262.300 ;
        RECT 110.130 262.000 110.730 262.150 ;
        RECT 106.530 261.700 110.730 262.000 ;
        RECT 118.730 262.000 119.330 262.150 ;
        RECT 119.780 262.000 119.930 269.550 ;
        RECT 120.380 262.000 120.530 269.550 ;
        RECT 120.980 262.000 121.130 269.550 ;
        RECT 121.580 262.000 121.730 269.550 ;
        RECT 122.180 262.000 122.330 269.550 ;
        RECT 122.780 262.000 122.930 264.900 ;
        RECT 118.730 261.700 122.930 262.000 ;
        RECT 106.530 261.550 114.080 261.700 ;
        RECT 115.380 261.550 122.930 261.700 ;
        RECT 106.530 261.350 110.730 261.550 ;
        RECT 100.330 261.050 109.130 261.200 ;
        RECT 109.280 261.050 110.730 261.350 ;
        RECT 98.730 260.150 110.730 261.050 ;
        RECT 118.730 261.350 122.930 261.550 ;
        RECT 123.530 263.275 124.730 264.400 ;
        RECT 123.530 262.000 127.140 263.275 ;
        RECT 118.730 261.050 120.180 261.350 ;
        RECT 123.530 261.200 124.730 262.000 ;
        RECT 120.330 261.050 124.730 261.200 ;
        RECT 118.730 260.150 124.730 261.050 ;
        RECT 4.730 259.850 9.130 260.150 ;
        RECT 20.330 259.850 29.130 260.150 ;
        RECT 40.330 259.850 49.130 260.150 ;
        RECT 60.330 259.850 69.130 260.150 ;
        RECT 80.330 259.850 89.130 260.150 ;
        RECT 100.330 259.850 109.130 260.150 ;
        RECT 4.730 258.950 10.730 259.850 ;
        RECT 20.330 259.800 30.730 259.850 ;
        RECT 40.330 259.800 50.730 259.850 ;
        RECT 60.330 259.800 70.730 259.850 ;
        RECT 80.330 259.800 90.730 259.850 ;
        RECT 100.330 259.800 110.730 259.850 ;
        RECT 120.330 259.800 124.730 260.150 ;
        RECT 4.730 258.800 9.130 258.950 ;
        RECT 4.730 257.610 5.930 258.800 ;
        RECT 9.280 258.650 10.730 258.950 ;
        RECT 2.315 256.335 5.930 257.610 ;
        RECT 4.730 255.600 5.930 256.335 ;
        RECT 6.530 258.450 10.730 258.650 ;
        RECT 18.730 258.950 30.730 259.800 ;
        RECT 18.730 258.900 29.130 258.950 ;
        RECT 18.730 258.650 20.180 258.900 ;
        RECT 20.330 258.800 29.130 258.900 ;
        RECT 18.730 258.450 22.930 258.650 ;
        RECT 6.530 258.300 14.080 258.450 ;
        RECT 15.430 258.300 22.930 258.450 ;
        RECT 6.530 258.000 10.730 258.300 ;
        RECT 2.315 253.250 4.315 255.545 ;
        RECT 6.530 255.150 6.680 258.000 ;
        RECT 7.130 250.450 7.280 258.000 ;
        RECT 7.730 250.450 7.880 258.000 ;
        RECT 8.330 250.450 8.480 258.000 ;
        RECT 8.930 250.450 9.080 258.000 ;
        RECT 9.530 250.450 9.680 258.000 ;
        RECT 10.130 257.850 10.730 258.000 ;
        RECT 18.730 258.000 22.930 258.300 ;
        RECT 18.730 257.850 19.330 258.000 ;
        RECT 10.130 257.700 14.080 257.850 ;
        RECT 15.380 257.700 19.330 257.850 ;
        RECT 10.130 257.250 10.730 257.700 ;
        RECT 18.730 257.250 19.330 257.700 ;
        RECT 10.130 257.100 14.080 257.250 ;
        RECT 15.380 257.100 19.330 257.250 ;
        RECT 10.130 256.650 10.730 257.100 ;
        RECT 18.730 256.650 19.330 257.100 ;
        RECT 10.130 256.500 14.080 256.650 ;
        RECT 15.380 256.500 19.330 256.650 ;
        RECT 10.130 256.050 10.730 256.500 ;
        RECT 18.730 256.050 19.330 256.500 ;
        RECT 10.130 255.900 14.080 256.050 ;
        RECT 15.380 255.900 19.330 256.050 ;
        RECT 10.130 255.450 10.730 255.900 ;
        RECT 18.730 255.450 19.330 255.900 ;
        RECT 10.130 255.300 14.080 255.450 ;
        RECT 15.380 255.300 19.330 255.450 ;
        RECT 10.130 254.850 10.730 255.300 ;
        RECT 18.730 254.850 19.330 255.300 ;
        RECT 10.130 254.700 14.080 254.850 ;
        RECT 15.380 254.700 19.330 254.850 ;
        RECT 10.130 254.250 10.730 254.700 ;
        RECT 18.730 254.250 19.330 254.700 ;
        RECT 10.130 254.100 14.080 254.250 ;
        RECT 15.380 254.100 19.330 254.250 ;
        RECT 10.130 253.650 10.730 254.100 ;
        RECT 18.730 253.650 19.330 254.100 ;
        RECT 10.130 253.500 14.080 253.650 ;
        RECT 15.380 253.500 19.330 253.650 ;
        RECT 10.130 253.050 10.730 253.500 ;
        RECT 18.730 253.050 19.330 253.500 ;
        RECT 10.130 252.900 14.080 253.050 ;
        RECT 15.380 252.900 19.330 253.050 ;
        RECT 10.130 252.450 10.730 252.900 ;
        RECT 18.730 252.450 19.330 252.900 ;
        RECT 10.130 252.300 14.080 252.450 ;
        RECT 15.380 252.300 19.330 252.450 ;
        RECT 10.130 251.850 10.730 252.300 ;
        RECT 18.730 251.850 19.330 252.300 ;
        RECT 10.130 251.700 14.080 251.850 ;
        RECT 15.380 251.700 19.330 251.850 ;
        RECT 10.130 251.250 10.730 251.700 ;
        RECT 18.730 251.250 19.330 251.700 ;
        RECT 10.130 251.100 14.080 251.250 ;
        RECT 15.380 251.100 19.330 251.250 ;
        RECT 10.130 250.650 10.730 251.100 ;
        RECT 18.730 250.650 19.330 251.100 ;
        RECT 10.130 250.450 14.080 250.650 ;
        RECT 15.380 250.450 19.330 250.650 ;
        RECT 19.780 250.450 19.930 258.000 ;
        RECT 20.380 250.450 20.530 258.000 ;
        RECT 20.980 250.450 21.130 258.000 ;
        RECT 21.580 250.450 21.730 258.000 ;
        RECT 22.180 250.450 22.330 258.000 ;
        RECT 22.780 255.150 22.930 258.000 ;
        RECT 23.530 255.600 25.930 258.800 ;
        RECT 29.280 258.650 30.730 258.950 ;
        RECT 26.530 258.450 30.730 258.650 ;
        RECT 38.730 258.950 50.730 259.800 ;
        RECT 38.730 258.900 49.130 258.950 ;
        RECT 38.730 258.650 40.180 258.900 ;
        RECT 40.330 258.800 49.130 258.900 ;
        RECT 38.730 258.450 42.930 258.650 ;
        RECT 26.530 258.300 34.080 258.450 ;
        RECT 35.430 258.300 42.930 258.450 ;
        RECT 26.530 258.000 30.730 258.300 ;
        RECT 26.530 255.150 26.680 258.000 ;
        RECT 27.130 250.450 27.280 258.000 ;
        RECT 27.730 250.450 27.880 258.000 ;
        RECT 28.330 250.450 28.480 258.000 ;
        RECT 28.930 250.450 29.080 258.000 ;
        RECT 29.530 250.450 29.680 258.000 ;
        RECT 30.130 257.850 30.730 258.000 ;
        RECT 38.730 258.000 42.930 258.300 ;
        RECT 38.730 257.850 39.330 258.000 ;
        RECT 30.130 257.700 34.080 257.850 ;
        RECT 35.380 257.700 39.330 257.850 ;
        RECT 30.130 257.250 30.730 257.700 ;
        RECT 38.730 257.250 39.330 257.700 ;
        RECT 30.130 257.100 34.080 257.250 ;
        RECT 35.380 257.100 39.330 257.250 ;
        RECT 30.130 256.650 30.730 257.100 ;
        RECT 38.730 256.650 39.330 257.100 ;
        RECT 30.130 256.500 34.080 256.650 ;
        RECT 35.380 256.500 39.330 256.650 ;
        RECT 30.130 256.050 30.730 256.500 ;
        RECT 38.730 256.050 39.330 256.500 ;
        RECT 30.130 255.900 34.080 256.050 ;
        RECT 35.380 255.900 39.330 256.050 ;
        RECT 30.130 255.450 30.730 255.900 ;
        RECT 38.730 255.450 39.330 255.900 ;
        RECT 30.130 255.300 34.080 255.450 ;
        RECT 35.380 255.300 39.330 255.450 ;
        RECT 30.130 254.850 30.730 255.300 ;
        RECT 38.730 254.850 39.330 255.300 ;
        RECT 30.130 254.700 34.080 254.850 ;
        RECT 35.380 254.700 39.330 254.850 ;
        RECT 30.130 254.250 30.730 254.700 ;
        RECT 38.730 254.250 39.330 254.700 ;
        RECT 30.130 254.100 34.080 254.250 ;
        RECT 35.380 254.100 39.330 254.250 ;
        RECT 30.130 253.650 30.730 254.100 ;
        RECT 38.730 253.650 39.330 254.100 ;
        RECT 30.130 253.500 34.080 253.650 ;
        RECT 35.380 253.500 39.330 253.650 ;
        RECT 30.130 253.050 30.730 253.500 ;
        RECT 38.730 253.050 39.330 253.500 ;
        RECT 30.130 252.900 34.080 253.050 ;
        RECT 35.380 252.900 39.330 253.050 ;
        RECT 30.130 252.450 30.730 252.900 ;
        RECT 38.730 252.450 39.330 252.900 ;
        RECT 30.130 252.300 34.080 252.450 ;
        RECT 35.380 252.300 39.330 252.450 ;
        RECT 30.130 251.850 30.730 252.300 ;
        RECT 38.730 251.850 39.330 252.300 ;
        RECT 30.130 251.700 34.080 251.850 ;
        RECT 35.380 251.700 39.330 251.850 ;
        RECT 30.130 251.250 30.730 251.700 ;
        RECT 38.730 251.250 39.330 251.700 ;
        RECT 30.130 251.100 34.080 251.250 ;
        RECT 35.380 251.100 39.330 251.250 ;
        RECT 30.130 250.650 30.730 251.100 ;
        RECT 38.730 250.650 39.330 251.100 ;
        RECT 30.130 250.450 34.080 250.650 ;
        RECT 35.380 250.450 39.330 250.650 ;
        RECT 39.780 250.450 39.930 258.000 ;
        RECT 40.380 250.450 40.530 258.000 ;
        RECT 40.980 250.450 41.130 258.000 ;
        RECT 41.580 250.450 41.730 258.000 ;
        RECT 42.180 250.450 42.330 258.000 ;
        RECT 42.780 255.150 42.930 258.000 ;
        RECT 43.530 255.600 45.930 258.800 ;
        RECT 49.280 258.650 50.730 258.950 ;
        RECT 46.530 258.450 50.730 258.650 ;
        RECT 58.730 258.950 70.730 259.800 ;
        RECT 58.730 258.900 69.130 258.950 ;
        RECT 58.730 258.650 60.180 258.900 ;
        RECT 60.330 258.800 69.130 258.900 ;
        RECT 58.730 258.450 62.930 258.650 ;
        RECT 46.530 258.300 54.080 258.450 ;
        RECT 55.430 258.300 62.930 258.450 ;
        RECT 46.530 258.000 50.730 258.300 ;
        RECT 46.530 255.150 46.680 258.000 ;
        RECT 47.130 250.450 47.280 258.000 ;
        RECT 47.730 250.450 47.880 258.000 ;
        RECT 48.330 250.450 48.480 258.000 ;
        RECT 48.930 250.450 49.080 258.000 ;
        RECT 49.530 250.450 49.680 258.000 ;
        RECT 50.130 257.850 50.730 258.000 ;
        RECT 58.730 258.000 62.930 258.300 ;
        RECT 58.730 257.850 59.330 258.000 ;
        RECT 50.130 257.700 54.080 257.850 ;
        RECT 55.380 257.700 59.330 257.850 ;
        RECT 50.130 257.250 50.730 257.700 ;
        RECT 58.730 257.250 59.330 257.700 ;
        RECT 50.130 257.100 54.080 257.250 ;
        RECT 55.380 257.100 59.330 257.250 ;
        RECT 50.130 256.650 50.730 257.100 ;
        RECT 58.730 256.650 59.330 257.100 ;
        RECT 50.130 256.500 54.080 256.650 ;
        RECT 55.380 256.500 59.330 256.650 ;
        RECT 50.130 256.050 50.730 256.500 ;
        RECT 58.730 256.050 59.330 256.500 ;
        RECT 50.130 255.900 54.080 256.050 ;
        RECT 55.380 255.900 59.330 256.050 ;
        RECT 50.130 255.450 50.730 255.900 ;
        RECT 58.730 255.450 59.330 255.900 ;
        RECT 50.130 255.300 54.080 255.450 ;
        RECT 55.380 255.300 59.330 255.450 ;
        RECT 50.130 254.850 50.730 255.300 ;
        RECT 58.730 254.850 59.330 255.300 ;
        RECT 50.130 254.700 54.080 254.850 ;
        RECT 55.380 254.700 59.330 254.850 ;
        RECT 50.130 254.250 50.730 254.700 ;
        RECT 58.730 254.250 59.330 254.700 ;
        RECT 50.130 254.100 54.080 254.250 ;
        RECT 55.380 254.100 59.330 254.250 ;
        RECT 50.130 253.650 50.730 254.100 ;
        RECT 58.730 253.650 59.330 254.100 ;
        RECT 50.130 253.500 54.080 253.650 ;
        RECT 55.380 253.500 59.330 253.650 ;
        RECT 50.130 253.050 50.730 253.500 ;
        RECT 58.730 253.050 59.330 253.500 ;
        RECT 50.130 252.900 54.080 253.050 ;
        RECT 55.380 252.900 59.330 253.050 ;
        RECT 50.130 252.450 50.730 252.900 ;
        RECT 58.730 252.450 59.330 252.900 ;
        RECT 50.130 252.300 54.080 252.450 ;
        RECT 55.380 252.300 59.330 252.450 ;
        RECT 50.130 251.850 50.730 252.300 ;
        RECT 58.730 251.850 59.330 252.300 ;
        RECT 50.130 251.700 54.080 251.850 ;
        RECT 55.380 251.700 59.330 251.850 ;
        RECT 50.130 251.250 50.730 251.700 ;
        RECT 58.730 251.250 59.330 251.700 ;
        RECT 50.130 251.100 54.080 251.250 ;
        RECT 55.380 251.100 59.330 251.250 ;
        RECT 50.130 250.650 50.730 251.100 ;
        RECT 58.730 250.650 59.330 251.100 ;
        RECT 50.130 250.450 54.080 250.650 ;
        RECT 55.380 250.450 59.330 250.650 ;
        RECT 59.780 250.450 59.930 258.000 ;
        RECT 60.380 250.450 60.530 258.000 ;
        RECT 60.980 250.450 61.130 258.000 ;
        RECT 61.580 250.450 61.730 258.000 ;
        RECT 62.180 250.450 62.330 258.000 ;
        RECT 62.780 255.150 62.930 258.000 ;
        RECT 63.530 255.600 65.930 258.800 ;
        RECT 69.280 258.650 70.730 258.950 ;
        RECT 66.530 258.450 70.730 258.650 ;
        RECT 78.730 258.950 90.730 259.800 ;
        RECT 78.730 258.900 89.130 258.950 ;
        RECT 78.730 258.650 80.180 258.900 ;
        RECT 80.330 258.800 89.130 258.900 ;
        RECT 78.730 258.450 82.930 258.650 ;
        RECT 66.530 258.300 74.080 258.450 ;
        RECT 75.430 258.300 82.930 258.450 ;
        RECT 66.530 258.000 70.730 258.300 ;
        RECT 66.530 255.150 66.680 258.000 ;
        RECT 67.130 250.450 67.280 258.000 ;
        RECT 67.730 250.450 67.880 258.000 ;
        RECT 68.330 250.450 68.480 258.000 ;
        RECT 68.930 250.450 69.080 258.000 ;
        RECT 69.530 250.450 69.680 258.000 ;
        RECT 70.130 257.850 70.730 258.000 ;
        RECT 78.730 258.000 82.930 258.300 ;
        RECT 78.730 257.850 79.330 258.000 ;
        RECT 70.130 257.700 74.080 257.850 ;
        RECT 75.380 257.700 79.330 257.850 ;
        RECT 70.130 257.250 70.730 257.700 ;
        RECT 78.730 257.250 79.330 257.700 ;
        RECT 70.130 257.100 74.080 257.250 ;
        RECT 75.380 257.100 79.330 257.250 ;
        RECT 70.130 256.650 70.730 257.100 ;
        RECT 78.730 256.650 79.330 257.100 ;
        RECT 70.130 256.500 74.080 256.650 ;
        RECT 75.380 256.500 79.330 256.650 ;
        RECT 70.130 256.050 70.730 256.500 ;
        RECT 78.730 256.050 79.330 256.500 ;
        RECT 70.130 255.900 74.080 256.050 ;
        RECT 75.380 255.900 79.330 256.050 ;
        RECT 70.130 255.450 70.730 255.900 ;
        RECT 78.730 255.450 79.330 255.900 ;
        RECT 70.130 255.300 74.080 255.450 ;
        RECT 75.380 255.300 79.330 255.450 ;
        RECT 70.130 254.850 70.730 255.300 ;
        RECT 78.730 254.850 79.330 255.300 ;
        RECT 70.130 254.700 74.080 254.850 ;
        RECT 75.380 254.700 79.330 254.850 ;
        RECT 70.130 254.250 70.730 254.700 ;
        RECT 78.730 254.250 79.330 254.700 ;
        RECT 70.130 254.100 74.080 254.250 ;
        RECT 75.380 254.100 79.330 254.250 ;
        RECT 70.130 253.650 70.730 254.100 ;
        RECT 78.730 253.650 79.330 254.100 ;
        RECT 70.130 253.500 74.080 253.650 ;
        RECT 75.380 253.500 79.330 253.650 ;
        RECT 70.130 253.050 70.730 253.500 ;
        RECT 78.730 253.050 79.330 253.500 ;
        RECT 70.130 252.900 74.080 253.050 ;
        RECT 75.380 252.900 79.330 253.050 ;
        RECT 70.130 252.450 70.730 252.900 ;
        RECT 78.730 252.450 79.330 252.900 ;
        RECT 70.130 252.300 74.080 252.450 ;
        RECT 75.380 252.300 79.330 252.450 ;
        RECT 70.130 251.850 70.730 252.300 ;
        RECT 78.730 251.850 79.330 252.300 ;
        RECT 70.130 251.700 74.080 251.850 ;
        RECT 75.380 251.700 79.330 251.850 ;
        RECT 70.130 251.250 70.730 251.700 ;
        RECT 78.730 251.250 79.330 251.700 ;
        RECT 70.130 251.100 74.080 251.250 ;
        RECT 75.380 251.100 79.330 251.250 ;
        RECT 70.130 250.650 70.730 251.100 ;
        RECT 78.730 250.650 79.330 251.100 ;
        RECT 70.130 250.450 74.080 250.650 ;
        RECT 75.380 250.450 79.330 250.650 ;
        RECT 79.780 250.450 79.930 258.000 ;
        RECT 80.380 250.450 80.530 258.000 ;
        RECT 80.980 250.450 81.130 258.000 ;
        RECT 81.580 250.450 81.730 258.000 ;
        RECT 82.180 250.450 82.330 258.000 ;
        RECT 82.780 255.150 82.930 258.000 ;
        RECT 83.530 255.600 85.930 258.800 ;
        RECT 89.280 258.650 90.730 258.950 ;
        RECT 86.530 258.450 90.730 258.650 ;
        RECT 98.730 258.950 110.730 259.800 ;
        RECT 98.730 258.900 109.130 258.950 ;
        RECT 98.730 258.650 100.180 258.900 ;
        RECT 100.330 258.800 109.130 258.900 ;
        RECT 98.730 258.450 102.930 258.650 ;
        RECT 86.530 258.300 94.080 258.450 ;
        RECT 95.430 258.300 102.930 258.450 ;
        RECT 86.530 258.000 90.730 258.300 ;
        RECT 86.530 255.150 86.680 258.000 ;
        RECT 87.130 250.450 87.280 258.000 ;
        RECT 87.730 250.450 87.880 258.000 ;
        RECT 88.330 250.450 88.480 258.000 ;
        RECT 88.930 250.450 89.080 258.000 ;
        RECT 89.530 250.450 89.680 258.000 ;
        RECT 90.130 257.850 90.730 258.000 ;
        RECT 98.730 258.000 102.930 258.300 ;
        RECT 98.730 257.850 99.330 258.000 ;
        RECT 90.130 257.700 94.080 257.850 ;
        RECT 95.380 257.700 99.330 257.850 ;
        RECT 90.130 257.250 90.730 257.700 ;
        RECT 98.730 257.250 99.330 257.700 ;
        RECT 90.130 257.100 94.080 257.250 ;
        RECT 95.380 257.100 99.330 257.250 ;
        RECT 90.130 256.650 90.730 257.100 ;
        RECT 98.730 256.650 99.330 257.100 ;
        RECT 90.130 256.500 94.080 256.650 ;
        RECT 95.380 256.500 99.330 256.650 ;
        RECT 90.130 256.050 90.730 256.500 ;
        RECT 98.730 256.050 99.330 256.500 ;
        RECT 90.130 255.900 94.080 256.050 ;
        RECT 95.380 255.900 99.330 256.050 ;
        RECT 90.130 255.450 90.730 255.900 ;
        RECT 98.730 255.450 99.330 255.900 ;
        RECT 90.130 255.300 94.080 255.450 ;
        RECT 95.380 255.300 99.330 255.450 ;
        RECT 90.130 254.850 90.730 255.300 ;
        RECT 98.730 254.850 99.330 255.300 ;
        RECT 90.130 254.700 94.080 254.850 ;
        RECT 95.380 254.700 99.330 254.850 ;
        RECT 90.130 254.250 90.730 254.700 ;
        RECT 98.730 254.250 99.330 254.700 ;
        RECT 90.130 254.100 94.080 254.250 ;
        RECT 95.380 254.100 99.330 254.250 ;
        RECT 90.130 253.650 90.730 254.100 ;
        RECT 98.730 253.650 99.330 254.100 ;
        RECT 90.130 253.500 94.080 253.650 ;
        RECT 95.380 253.500 99.330 253.650 ;
        RECT 90.130 253.050 90.730 253.500 ;
        RECT 98.730 253.050 99.330 253.500 ;
        RECT 90.130 252.900 94.080 253.050 ;
        RECT 95.380 252.900 99.330 253.050 ;
        RECT 90.130 252.450 90.730 252.900 ;
        RECT 98.730 252.450 99.330 252.900 ;
        RECT 90.130 252.300 94.080 252.450 ;
        RECT 95.380 252.300 99.330 252.450 ;
        RECT 90.130 251.850 90.730 252.300 ;
        RECT 98.730 251.850 99.330 252.300 ;
        RECT 90.130 251.700 94.080 251.850 ;
        RECT 95.380 251.700 99.330 251.850 ;
        RECT 90.130 251.250 90.730 251.700 ;
        RECT 98.730 251.250 99.330 251.700 ;
        RECT 90.130 251.100 94.080 251.250 ;
        RECT 95.380 251.100 99.330 251.250 ;
        RECT 90.130 250.650 90.730 251.100 ;
        RECT 98.730 250.650 99.330 251.100 ;
        RECT 90.130 250.450 94.080 250.650 ;
        RECT 95.380 250.450 99.330 250.650 ;
        RECT 99.780 250.450 99.930 258.000 ;
        RECT 100.380 250.450 100.530 258.000 ;
        RECT 100.980 250.450 101.130 258.000 ;
        RECT 101.580 250.450 101.730 258.000 ;
        RECT 102.180 250.450 102.330 258.000 ;
        RECT 102.780 255.150 102.930 258.000 ;
        RECT 103.530 255.600 105.930 258.800 ;
        RECT 109.280 258.650 110.730 258.950 ;
        RECT 106.530 258.450 110.730 258.650 ;
        RECT 118.730 258.900 124.730 259.800 ;
        RECT 118.730 258.650 120.180 258.900 ;
        RECT 120.330 258.800 124.730 258.900 ;
        RECT 118.730 258.450 122.930 258.650 ;
        RECT 106.530 258.300 114.080 258.450 ;
        RECT 115.430 258.300 122.930 258.450 ;
        RECT 106.530 258.000 110.730 258.300 ;
        RECT 106.530 255.150 106.680 258.000 ;
        RECT 107.130 250.450 107.280 258.000 ;
        RECT 107.730 250.450 107.880 258.000 ;
        RECT 108.330 250.450 108.480 258.000 ;
        RECT 108.930 250.450 109.080 258.000 ;
        RECT 109.530 250.450 109.680 258.000 ;
        RECT 110.130 257.850 110.730 258.000 ;
        RECT 118.730 258.000 122.930 258.300 ;
        RECT 118.730 257.850 119.330 258.000 ;
        RECT 110.130 257.700 114.080 257.850 ;
        RECT 115.380 257.700 119.330 257.850 ;
        RECT 110.130 257.250 110.730 257.700 ;
        RECT 118.730 257.250 119.330 257.700 ;
        RECT 110.130 257.100 114.080 257.250 ;
        RECT 115.380 257.100 119.330 257.250 ;
        RECT 110.130 256.650 110.730 257.100 ;
        RECT 118.730 256.650 119.330 257.100 ;
        RECT 110.130 256.500 114.080 256.650 ;
        RECT 115.380 256.500 119.330 256.650 ;
        RECT 110.130 256.050 110.730 256.500 ;
        RECT 118.730 256.050 119.330 256.500 ;
        RECT 110.130 255.900 114.080 256.050 ;
        RECT 115.380 255.900 119.330 256.050 ;
        RECT 110.130 255.450 110.730 255.900 ;
        RECT 118.730 255.450 119.330 255.900 ;
        RECT 110.130 255.300 114.080 255.450 ;
        RECT 115.380 255.300 119.330 255.450 ;
        RECT 110.130 254.850 110.730 255.300 ;
        RECT 118.730 254.850 119.330 255.300 ;
        RECT 110.130 254.700 114.080 254.850 ;
        RECT 115.380 254.700 119.330 254.850 ;
        RECT 110.130 254.250 110.730 254.700 ;
        RECT 118.730 254.250 119.330 254.700 ;
        RECT 110.130 254.100 114.080 254.250 ;
        RECT 115.380 254.100 119.330 254.250 ;
        RECT 110.130 253.650 110.730 254.100 ;
        RECT 118.730 253.650 119.330 254.100 ;
        RECT 110.130 253.500 114.080 253.650 ;
        RECT 115.380 253.500 119.330 253.650 ;
        RECT 110.130 253.050 110.730 253.500 ;
        RECT 118.730 253.050 119.330 253.500 ;
        RECT 110.130 252.900 114.080 253.050 ;
        RECT 115.380 252.900 119.330 253.050 ;
        RECT 110.130 252.450 110.730 252.900 ;
        RECT 118.730 252.450 119.330 252.900 ;
        RECT 110.130 252.300 114.080 252.450 ;
        RECT 115.380 252.300 119.330 252.450 ;
        RECT 110.130 251.850 110.730 252.300 ;
        RECT 118.730 251.850 119.330 252.300 ;
        RECT 110.130 251.700 114.080 251.850 ;
        RECT 115.380 251.700 119.330 251.850 ;
        RECT 110.130 251.250 110.730 251.700 ;
        RECT 118.730 251.250 119.330 251.700 ;
        RECT 110.130 251.100 114.080 251.250 ;
        RECT 115.380 251.100 119.330 251.250 ;
        RECT 110.130 250.650 110.730 251.100 ;
        RECT 118.730 250.650 119.330 251.100 ;
        RECT 110.130 250.450 114.080 250.650 ;
        RECT 115.380 250.450 119.330 250.650 ;
        RECT 119.780 250.450 119.930 258.000 ;
        RECT 120.380 250.450 120.530 258.000 ;
        RECT 120.980 250.450 121.130 258.000 ;
        RECT 121.580 250.450 121.730 258.000 ;
        RECT 122.180 250.450 122.330 258.000 ;
        RECT 122.780 255.150 122.930 258.000 ;
        RECT 123.530 257.360 124.730 258.800 ;
        RECT 123.530 256.085 127.135 257.360 ;
        RECT 123.530 255.600 124.730 256.085 ;
        RECT 2.315 244.455 4.315 246.750 ;
        RECT 4.730 243.780 5.930 244.400 ;
        RECT 2.315 242.505 5.930 243.780 ;
        RECT 4.730 241.200 5.930 242.505 ;
        RECT 6.530 242.000 6.680 244.900 ;
        RECT 7.130 242.000 7.280 249.550 ;
        RECT 7.730 242.000 7.880 249.550 ;
        RECT 8.330 242.000 8.480 249.550 ;
        RECT 8.930 242.000 9.080 249.550 ;
        RECT 9.530 242.000 9.680 249.550 ;
        RECT 10.130 249.350 14.080 249.550 ;
        RECT 15.380 249.350 19.330 249.550 ;
        RECT 10.130 248.900 10.730 249.350 ;
        RECT 18.730 248.900 19.330 249.350 ;
        RECT 10.130 248.750 14.080 248.900 ;
        RECT 15.380 248.750 19.330 248.900 ;
        RECT 10.130 248.300 10.730 248.750 ;
        RECT 18.730 248.300 19.330 248.750 ;
        RECT 10.130 248.150 14.080 248.300 ;
        RECT 15.380 248.150 19.330 248.300 ;
        RECT 10.130 247.700 10.730 248.150 ;
        RECT 18.730 247.700 19.330 248.150 ;
        RECT 10.130 247.550 14.080 247.700 ;
        RECT 15.380 247.550 19.330 247.700 ;
        RECT 10.130 247.100 10.730 247.550 ;
        RECT 18.730 247.100 19.330 247.550 ;
        RECT 10.130 246.950 14.080 247.100 ;
        RECT 15.380 246.950 19.330 247.100 ;
        RECT 10.130 246.500 10.730 246.950 ;
        RECT 18.730 246.500 19.330 246.950 ;
        RECT 10.130 246.350 14.080 246.500 ;
        RECT 15.380 246.350 19.330 246.500 ;
        RECT 10.130 245.900 10.730 246.350 ;
        RECT 18.730 245.900 19.330 246.350 ;
        RECT 10.130 245.750 14.080 245.900 ;
        RECT 15.380 245.750 19.330 245.900 ;
        RECT 10.130 245.300 10.730 245.750 ;
        RECT 18.730 245.300 19.330 245.750 ;
        RECT 10.130 245.150 14.080 245.300 ;
        RECT 15.380 245.150 19.330 245.300 ;
        RECT 10.130 244.700 10.730 245.150 ;
        RECT 18.730 244.700 19.330 245.150 ;
        RECT 10.130 244.550 14.080 244.700 ;
        RECT 15.380 244.550 19.330 244.700 ;
        RECT 10.130 244.100 10.730 244.550 ;
        RECT 18.730 244.100 19.330 244.550 ;
        RECT 10.130 243.950 14.080 244.100 ;
        RECT 15.380 243.950 19.330 244.100 ;
        RECT 10.130 243.500 10.730 243.950 ;
        RECT 18.730 243.500 19.330 243.950 ;
        RECT 10.130 243.350 14.080 243.500 ;
        RECT 15.380 243.350 19.330 243.500 ;
        RECT 10.130 242.900 10.730 243.350 ;
        RECT 18.730 242.900 19.330 243.350 ;
        RECT 10.130 242.750 14.080 242.900 ;
        RECT 15.380 242.750 19.330 242.900 ;
        RECT 10.130 242.300 10.730 242.750 ;
        RECT 18.730 242.300 19.330 242.750 ;
        RECT 10.130 242.150 14.080 242.300 ;
        RECT 15.380 242.150 19.330 242.300 ;
        RECT 10.130 242.000 10.730 242.150 ;
        RECT 6.530 241.700 10.730 242.000 ;
        RECT 18.730 242.000 19.330 242.150 ;
        RECT 19.780 242.000 19.930 249.550 ;
        RECT 20.380 242.000 20.530 249.550 ;
        RECT 20.980 242.000 21.130 249.550 ;
        RECT 21.580 242.000 21.730 249.550 ;
        RECT 22.180 242.000 22.330 249.550 ;
        RECT 22.780 242.000 22.930 244.900 ;
        RECT 18.730 241.700 22.930 242.000 ;
        RECT 6.530 241.550 14.080 241.700 ;
        RECT 15.380 241.550 22.930 241.700 ;
        RECT 6.530 241.350 10.730 241.550 ;
        RECT 4.730 241.050 9.130 241.200 ;
        RECT 9.280 241.050 10.730 241.350 ;
        RECT 4.730 240.150 10.730 241.050 ;
        RECT 18.730 241.350 22.930 241.550 ;
        RECT 18.730 241.050 20.180 241.350 ;
        RECT 23.530 241.200 25.930 244.400 ;
        RECT 26.530 242.000 26.680 244.900 ;
        RECT 27.130 242.000 27.280 249.550 ;
        RECT 27.730 242.000 27.880 249.550 ;
        RECT 28.330 242.000 28.480 249.550 ;
        RECT 28.930 242.000 29.080 249.550 ;
        RECT 29.530 242.000 29.680 249.550 ;
        RECT 30.130 249.350 34.080 249.550 ;
        RECT 35.380 249.350 39.330 249.550 ;
        RECT 30.130 248.900 30.730 249.350 ;
        RECT 38.730 248.900 39.330 249.350 ;
        RECT 30.130 248.750 34.080 248.900 ;
        RECT 35.380 248.750 39.330 248.900 ;
        RECT 30.130 248.300 30.730 248.750 ;
        RECT 38.730 248.300 39.330 248.750 ;
        RECT 30.130 248.150 34.080 248.300 ;
        RECT 35.380 248.150 39.330 248.300 ;
        RECT 30.130 247.700 30.730 248.150 ;
        RECT 38.730 247.700 39.330 248.150 ;
        RECT 30.130 247.550 34.080 247.700 ;
        RECT 35.380 247.550 39.330 247.700 ;
        RECT 30.130 247.100 30.730 247.550 ;
        RECT 38.730 247.100 39.330 247.550 ;
        RECT 30.130 246.950 34.080 247.100 ;
        RECT 35.380 246.950 39.330 247.100 ;
        RECT 30.130 246.500 30.730 246.950 ;
        RECT 38.730 246.500 39.330 246.950 ;
        RECT 30.130 246.350 34.080 246.500 ;
        RECT 35.380 246.350 39.330 246.500 ;
        RECT 30.130 245.900 30.730 246.350 ;
        RECT 38.730 245.900 39.330 246.350 ;
        RECT 30.130 245.750 34.080 245.900 ;
        RECT 35.380 245.750 39.330 245.900 ;
        RECT 30.130 245.300 30.730 245.750 ;
        RECT 38.730 245.300 39.330 245.750 ;
        RECT 30.130 245.150 34.080 245.300 ;
        RECT 35.380 245.150 39.330 245.300 ;
        RECT 30.130 244.700 30.730 245.150 ;
        RECT 38.730 244.700 39.330 245.150 ;
        RECT 30.130 244.550 34.080 244.700 ;
        RECT 35.380 244.550 39.330 244.700 ;
        RECT 30.130 244.100 30.730 244.550 ;
        RECT 38.730 244.100 39.330 244.550 ;
        RECT 30.130 243.950 34.080 244.100 ;
        RECT 35.380 243.950 39.330 244.100 ;
        RECT 30.130 243.500 30.730 243.950 ;
        RECT 38.730 243.500 39.330 243.950 ;
        RECT 30.130 243.350 34.080 243.500 ;
        RECT 35.380 243.350 39.330 243.500 ;
        RECT 30.130 242.900 30.730 243.350 ;
        RECT 38.730 242.900 39.330 243.350 ;
        RECT 30.130 242.750 34.080 242.900 ;
        RECT 35.380 242.750 39.330 242.900 ;
        RECT 30.130 242.300 30.730 242.750 ;
        RECT 38.730 242.300 39.330 242.750 ;
        RECT 30.130 242.150 34.080 242.300 ;
        RECT 35.380 242.150 39.330 242.300 ;
        RECT 30.130 242.000 30.730 242.150 ;
        RECT 26.530 241.700 30.730 242.000 ;
        RECT 38.730 242.000 39.330 242.150 ;
        RECT 39.780 242.000 39.930 249.550 ;
        RECT 40.380 242.000 40.530 249.550 ;
        RECT 40.980 242.000 41.130 249.550 ;
        RECT 41.580 242.000 41.730 249.550 ;
        RECT 42.180 242.000 42.330 249.550 ;
        RECT 42.780 242.000 42.930 244.900 ;
        RECT 38.730 241.700 42.930 242.000 ;
        RECT 26.530 241.550 34.080 241.700 ;
        RECT 35.380 241.550 42.930 241.700 ;
        RECT 26.530 241.350 30.730 241.550 ;
        RECT 20.330 241.050 29.130 241.200 ;
        RECT 29.280 241.050 30.730 241.350 ;
        RECT 18.730 240.150 30.730 241.050 ;
        RECT 38.730 241.350 42.930 241.550 ;
        RECT 38.730 241.050 40.180 241.350 ;
        RECT 43.530 241.200 45.930 244.400 ;
        RECT 46.530 242.000 46.680 244.900 ;
        RECT 47.130 242.000 47.280 249.550 ;
        RECT 47.730 242.000 47.880 249.550 ;
        RECT 48.330 242.000 48.480 249.550 ;
        RECT 48.930 242.000 49.080 249.550 ;
        RECT 49.530 242.000 49.680 249.550 ;
        RECT 50.130 249.350 54.080 249.550 ;
        RECT 55.380 249.350 59.330 249.550 ;
        RECT 50.130 248.900 50.730 249.350 ;
        RECT 58.730 248.900 59.330 249.350 ;
        RECT 50.130 248.750 54.080 248.900 ;
        RECT 55.380 248.750 59.330 248.900 ;
        RECT 50.130 248.300 50.730 248.750 ;
        RECT 58.730 248.300 59.330 248.750 ;
        RECT 50.130 248.150 54.080 248.300 ;
        RECT 55.380 248.150 59.330 248.300 ;
        RECT 50.130 247.700 50.730 248.150 ;
        RECT 58.730 247.700 59.330 248.150 ;
        RECT 50.130 247.550 54.080 247.700 ;
        RECT 55.380 247.550 59.330 247.700 ;
        RECT 50.130 247.100 50.730 247.550 ;
        RECT 58.730 247.100 59.330 247.550 ;
        RECT 50.130 246.950 54.080 247.100 ;
        RECT 55.380 246.950 59.330 247.100 ;
        RECT 50.130 246.500 50.730 246.950 ;
        RECT 58.730 246.500 59.330 246.950 ;
        RECT 50.130 246.350 54.080 246.500 ;
        RECT 55.380 246.350 59.330 246.500 ;
        RECT 50.130 245.900 50.730 246.350 ;
        RECT 58.730 245.900 59.330 246.350 ;
        RECT 50.130 245.750 54.080 245.900 ;
        RECT 55.380 245.750 59.330 245.900 ;
        RECT 50.130 245.300 50.730 245.750 ;
        RECT 58.730 245.300 59.330 245.750 ;
        RECT 50.130 245.150 54.080 245.300 ;
        RECT 55.380 245.150 59.330 245.300 ;
        RECT 50.130 244.700 50.730 245.150 ;
        RECT 58.730 244.700 59.330 245.150 ;
        RECT 50.130 244.550 54.080 244.700 ;
        RECT 55.380 244.550 59.330 244.700 ;
        RECT 50.130 244.100 50.730 244.550 ;
        RECT 58.730 244.100 59.330 244.550 ;
        RECT 50.130 243.950 54.080 244.100 ;
        RECT 55.380 243.950 59.330 244.100 ;
        RECT 50.130 243.500 50.730 243.950 ;
        RECT 58.730 243.500 59.330 243.950 ;
        RECT 50.130 243.350 54.080 243.500 ;
        RECT 55.380 243.350 59.330 243.500 ;
        RECT 50.130 242.900 50.730 243.350 ;
        RECT 58.730 242.900 59.330 243.350 ;
        RECT 50.130 242.750 54.080 242.900 ;
        RECT 55.380 242.750 59.330 242.900 ;
        RECT 50.130 242.300 50.730 242.750 ;
        RECT 58.730 242.300 59.330 242.750 ;
        RECT 50.130 242.150 54.080 242.300 ;
        RECT 55.380 242.150 59.330 242.300 ;
        RECT 50.130 242.000 50.730 242.150 ;
        RECT 46.530 241.700 50.730 242.000 ;
        RECT 58.730 242.000 59.330 242.150 ;
        RECT 59.780 242.000 59.930 249.550 ;
        RECT 60.380 242.000 60.530 249.550 ;
        RECT 60.980 242.000 61.130 249.550 ;
        RECT 61.580 242.000 61.730 249.550 ;
        RECT 62.180 242.000 62.330 249.550 ;
        RECT 62.780 242.000 62.930 244.900 ;
        RECT 58.730 241.700 62.930 242.000 ;
        RECT 46.530 241.550 54.080 241.700 ;
        RECT 55.380 241.550 62.930 241.700 ;
        RECT 46.530 241.350 50.730 241.550 ;
        RECT 40.330 241.050 49.130 241.200 ;
        RECT 49.280 241.050 50.730 241.350 ;
        RECT 38.730 240.150 50.730 241.050 ;
        RECT 58.730 241.350 62.930 241.550 ;
        RECT 58.730 241.050 60.180 241.350 ;
        RECT 63.530 241.200 65.930 244.400 ;
        RECT 66.530 242.000 66.680 244.900 ;
        RECT 67.130 242.000 67.280 249.550 ;
        RECT 67.730 242.000 67.880 249.550 ;
        RECT 68.330 242.000 68.480 249.550 ;
        RECT 68.930 242.000 69.080 249.550 ;
        RECT 69.530 242.000 69.680 249.550 ;
        RECT 70.130 249.350 74.080 249.550 ;
        RECT 75.380 249.350 79.330 249.550 ;
        RECT 70.130 248.900 70.730 249.350 ;
        RECT 78.730 248.900 79.330 249.350 ;
        RECT 70.130 248.750 74.080 248.900 ;
        RECT 75.380 248.750 79.330 248.900 ;
        RECT 70.130 248.300 70.730 248.750 ;
        RECT 78.730 248.300 79.330 248.750 ;
        RECT 70.130 248.150 74.080 248.300 ;
        RECT 75.380 248.150 79.330 248.300 ;
        RECT 70.130 247.700 70.730 248.150 ;
        RECT 78.730 247.700 79.330 248.150 ;
        RECT 70.130 247.550 74.080 247.700 ;
        RECT 75.380 247.550 79.330 247.700 ;
        RECT 70.130 247.100 70.730 247.550 ;
        RECT 78.730 247.100 79.330 247.550 ;
        RECT 70.130 246.950 74.080 247.100 ;
        RECT 75.380 246.950 79.330 247.100 ;
        RECT 70.130 246.500 70.730 246.950 ;
        RECT 78.730 246.500 79.330 246.950 ;
        RECT 70.130 246.350 74.080 246.500 ;
        RECT 75.380 246.350 79.330 246.500 ;
        RECT 70.130 245.900 70.730 246.350 ;
        RECT 78.730 245.900 79.330 246.350 ;
        RECT 70.130 245.750 74.080 245.900 ;
        RECT 75.380 245.750 79.330 245.900 ;
        RECT 70.130 245.300 70.730 245.750 ;
        RECT 78.730 245.300 79.330 245.750 ;
        RECT 70.130 245.150 74.080 245.300 ;
        RECT 75.380 245.150 79.330 245.300 ;
        RECT 70.130 244.700 70.730 245.150 ;
        RECT 78.730 244.700 79.330 245.150 ;
        RECT 70.130 244.550 74.080 244.700 ;
        RECT 75.380 244.550 79.330 244.700 ;
        RECT 70.130 244.100 70.730 244.550 ;
        RECT 78.730 244.100 79.330 244.550 ;
        RECT 70.130 243.950 74.080 244.100 ;
        RECT 75.380 243.950 79.330 244.100 ;
        RECT 70.130 243.500 70.730 243.950 ;
        RECT 78.730 243.500 79.330 243.950 ;
        RECT 70.130 243.350 74.080 243.500 ;
        RECT 75.380 243.350 79.330 243.500 ;
        RECT 70.130 242.900 70.730 243.350 ;
        RECT 78.730 242.900 79.330 243.350 ;
        RECT 70.130 242.750 74.080 242.900 ;
        RECT 75.380 242.750 79.330 242.900 ;
        RECT 70.130 242.300 70.730 242.750 ;
        RECT 78.730 242.300 79.330 242.750 ;
        RECT 70.130 242.150 74.080 242.300 ;
        RECT 75.380 242.150 79.330 242.300 ;
        RECT 70.130 242.000 70.730 242.150 ;
        RECT 66.530 241.700 70.730 242.000 ;
        RECT 78.730 242.000 79.330 242.150 ;
        RECT 79.780 242.000 79.930 249.550 ;
        RECT 80.380 242.000 80.530 249.550 ;
        RECT 80.980 242.000 81.130 249.550 ;
        RECT 81.580 242.000 81.730 249.550 ;
        RECT 82.180 242.000 82.330 249.550 ;
        RECT 82.780 242.000 82.930 244.900 ;
        RECT 78.730 241.700 82.930 242.000 ;
        RECT 66.530 241.550 74.080 241.700 ;
        RECT 75.380 241.550 82.930 241.700 ;
        RECT 66.530 241.350 70.730 241.550 ;
        RECT 60.330 241.050 69.130 241.200 ;
        RECT 69.280 241.050 70.730 241.350 ;
        RECT 58.730 240.150 70.730 241.050 ;
        RECT 78.730 241.350 82.930 241.550 ;
        RECT 78.730 241.050 80.180 241.350 ;
        RECT 83.530 241.200 85.930 244.400 ;
        RECT 86.530 242.000 86.680 244.900 ;
        RECT 87.130 242.000 87.280 249.550 ;
        RECT 87.730 242.000 87.880 249.550 ;
        RECT 88.330 242.000 88.480 249.550 ;
        RECT 88.930 242.000 89.080 249.550 ;
        RECT 89.530 242.000 89.680 249.550 ;
        RECT 90.130 249.350 94.080 249.550 ;
        RECT 95.380 249.350 99.330 249.550 ;
        RECT 90.130 248.900 90.730 249.350 ;
        RECT 98.730 248.900 99.330 249.350 ;
        RECT 90.130 248.750 94.080 248.900 ;
        RECT 95.380 248.750 99.330 248.900 ;
        RECT 90.130 248.300 90.730 248.750 ;
        RECT 98.730 248.300 99.330 248.750 ;
        RECT 90.130 248.150 94.080 248.300 ;
        RECT 95.380 248.150 99.330 248.300 ;
        RECT 90.130 247.700 90.730 248.150 ;
        RECT 98.730 247.700 99.330 248.150 ;
        RECT 90.130 247.550 94.080 247.700 ;
        RECT 95.380 247.550 99.330 247.700 ;
        RECT 90.130 247.100 90.730 247.550 ;
        RECT 98.730 247.100 99.330 247.550 ;
        RECT 90.130 246.950 94.080 247.100 ;
        RECT 95.380 246.950 99.330 247.100 ;
        RECT 90.130 246.500 90.730 246.950 ;
        RECT 98.730 246.500 99.330 246.950 ;
        RECT 90.130 246.350 94.080 246.500 ;
        RECT 95.380 246.350 99.330 246.500 ;
        RECT 90.130 245.900 90.730 246.350 ;
        RECT 98.730 245.900 99.330 246.350 ;
        RECT 90.130 245.750 94.080 245.900 ;
        RECT 95.380 245.750 99.330 245.900 ;
        RECT 90.130 245.300 90.730 245.750 ;
        RECT 98.730 245.300 99.330 245.750 ;
        RECT 90.130 245.150 94.080 245.300 ;
        RECT 95.380 245.150 99.330 245.300 ;
        RECT 90.130 244.700 90.730 245.150 ;
        RECT 98.730 244.700 99.330 245.150 ;
        RECT 90.130 244.550 94.080 244.700 ;
        RECT 95.380 244.550 99.330 244.700 ;
        RECT 90.130 244.100 90.730 244.550 ;
        RECT 98.730 244.100 99.330 244.550 ;
        RECT 90.130 243.950 94.080 244.100 ;
        RECT 95.380 243.950 99.330 244.100 ;
        RECT 90.130 243.500 90.730 243.950 ;
        RECT 98.730 243.500 99.330 243.950 ;
        RECT 90.130 243.350 94.080 243.500 ;
        RECT 95.380 243.350 99.330 243.500 ;
        RECT 90.130 242.900 90.730 243.350 ;
        RECT 98.730 242.900 99.330 243.350 ;
        RECT 90.130 242.750 94.080 242.900 ;
        RECT 95.380 242.750 99.330 242.900 ;
        RECT 90.130 242.300 90.730 242.750 ;
        RECT 98.730 242.300 99.330 242.750 ;
        RECT 90.130 242.150 94.080 242.300 ;
        RECT 95.380 242.150 99.330 242.300 ;
        RECT 90.130 242.000 90.730 242.150 ;
        RECT 86.530 241.700 90.730 242.000 ;
        RECT 98.730 242.000 99.330 242.150 ;
        RECT 99.780 242.000 99.930 249.550 ;
        RECT 100.380 242.000 100.530 249.550 ;
        RECT 100.980 242.000 101.130 249.550 ;
        RECT 101.580 242.000 101.730 249.550 ;
        RECT 102.180 242.000 102.330 249.550 ;
        RECT 102.780 242.000 102.930 244.900 ;
        RECT 98.730 241.700 102.930 242.000 ;
        RECT 86.530 241.550 94.080 241.700 ;
        RECT 95.380 241.550 102.930 241.700 ;
        RECT 86.530 241.350 90.730 241.550 ;
        RECT 80.330 241.050 89.130 241.200 ;
        RECT 89.280 241.050 90.730 241.350 ;
        RECT 78.730 240.150 90.730 241.050 ;
        RECT 98.730 241.350 102.930 241.550 ;
        RECT 98.730 241.050 100.180 241.350 ;
        RECT 103.530 241.200 105.930 244.400 ;
        RECT 106.530 242.000 106.680 244.900 ;
        RECT 107.130 242.000 107.280 249.550 ;
        RECT 107.730 242.000 107.880 249.550 ;
        RECT 108.330 242.000 108.480 249.550 ;
        RECT 108.930 242.000 109.080 249.550 ;
        RECT 109.530 242.000 109.680 249.550 ;
        RECT 110.130 249.350 114.080 249.550 ;
        RECT 115.380 249.350 119.330 249.550 ;
        RECT 110.130 248.900 110.730 249.350 ;
        RECT 118.730 248.900 119.330 249.350 ;
        RECT 110.130 248.750 114.080 248.900 ;
        RECT 115.380 248.750 119.330 248.900 ;
        RECT 110.130 248.300 110.730 248.750 ;
        RECT 118.730 248.300 119.330 248.750 ;
        RECT 110.130 248.150 114.080 248.300 ;
        RECT 115.380 248.150 119.330 248.300 ;
        RECT 110.130 247.700 110.730 248.150 ;
        RECT 118.730 247.700 119.330 248.150 ;
        RECT 110.130 247.550 114.080 247.700 ;
        RECT 115.380 247.550 119.330 247.700 ;
        RECT 110.130 247.100 110.730 247.550 ;
        RECT 118.730 247.100 119.330 247.550 ;
        RECT 110.130 246.950 114.080 247.100 ;
        RECT 115.380 246.950 119.330 247.100 ;
        RECT 110.130 246.500 110.730 246.950 ;
        RECT 118.730 246.500 119.330 246.950 ;
        RECT 110.130 246.350 114.080 246.500 ;
        RECT 115.380 246.350 119.330 246.500 ;
        RECT 110.130 245.900 110.730 246.350 ;
        RECT 118.730 245.900 119.330 246.350 ;
        RECT 110.130 245.750 114.080 245.900 ;
        RECT 115.380 245.750 119.330 245.900 ;
        RECT 110.130 245.300 110.730 245.750 ;
        RECT 118.730 245.300 119.330 245.750 ;
        RECT 110.130 245.150 114.080 245.300 ;
        RECT 115.380 245.150 119.330 245.300 ;
        RECT 110.130 244.700 110.730 245.150 ;
        RECT 118.730 244.700 119.330 245.150 ;
        RECT 110.130 244.550 114.080 244.700 ;
        RECT 115.380 244.550 119.330 244.700 ;
        RECT 110.130 244.100 110.730 244.550 ;
        RECT 118.730 244.100 119.330 244.550 ;
        RECT 110.130 243.950 114.080 244.100 ;
        RECT 115.380 243.950 119.330 244.100 ;
        RECT 110.130 243.500 110.730 243.950 ;
        RECT 118.730 243.500 119.330 243.950 ;
        RECT 110.130 243.350 114.080 243.500 ;
        RECT 115.380 243.350 119.330 243.500 ;
        RECT 110.130 242.900 110.730 243.350 ;
        RECT 118.730 242.900 119.330 243.350 ;
        RECT 110.130 242.750 114.080 242.900 ;
        RECT 115.380 242.750 119.330 242.900 ;
        RECT 110.130 242.300 110.730 242.750 ;
        RECT 118.730 242.300 119.330 242.750 ;
        RECT 110.130 242.150 114.080 242.300 ;
        RECT 115.380 242.150 119.330 242.300 ;
        RECT 110.130 242.000 110.730 242.150 ;
        RECT 106.530 241.700 110.730 242.000 ;
        RECT 118.730 242.000 119.330 242.150 ;
        RECT 119.780 242.000 119.930 249.550 ;
        RECT 120.380 242.000 120.530 249.550 ;
        RECT 120.980 242.000 121.130 249.550 ;
        RECT 121.580 242.000 121.730 249.550 ;
        RECT 122.180 242.000 122.330 249.550 ;
        RECT 122.780 242.000 122.930 244.900 ;
        RECT 118.730 241.700 122.930 242.000 ;
        RECT 106.530 241.550 114.080 241.700 ;
        RECT 115.380 241.550 122.930 241.700 ;
        RECT 106.530 241.350 110.730 241.550 ;
        RECT 100.330 241.050 109.130 241.200 ;
        RECT 109.280 241.050 110.730 241.350 ;
        RECT 98.730 240.150 110.730 241.050 ;
        RECT 118.730 241.350 122.930 241.550 ;
        RECT 123.530 243.000 124.730 244.400 ;
        RECT 123.530 241.725 127.140 243.000 ;
        RECT 118.730 241.050 120.180 241.350 ;
        RECT 123.530 241.200 124.730 241.725 ;
        RECT 120.330 241.050 124.730 241.200 ;
        RECT 118.730 240.150 124.730 241.050 ;
        RECT 4.730 239.850 9.130 240.150 ;
        RECT 20.330 239.850 29.130 240.150 ;
        RECT 40.330 239.850 49.130 240.150 ;
        RECT 60.330 239.850 69.130 240.150 ;
        RECT 80.330 239.850 89.130 240.150 ;
        RECT 100.330 239.850 109.130 240.150 ;
        RECT 4.730 238.950 10.730 239.850 ;
        RECT 20.330 239.800 30.730 239.850 ;
        RECT 40.330 239.800 50.730 239.850 ;
        RECT 60.330 239.800 70.730 239.850 ;
        RECT 80.330 239.800 90.730 239.850 ;
        RECT 100.330 239.800 110.730 239.850 ;
        RECT 120.330 239.800 124.730 240.150 ;
        RECT 4.730 238.800 9.130 238.950 ;
        RECT 4.730 237.845 5.930 238.800 ;
        RECT 9.280 238.650 10.730 238.950 ;
        RECT 2.315 236.570 5.930 237.845 ;
        RECT 4.730 235.600 5.930 236.570 ;
        RECT 6.530 238.450 10.730 238.650 ;
        RECT 18.730 238.950 30.730 239.800 ;
        RECT 18.730 238.900 29.130 238.950 ;
        RECT 18.730 238.650 20.180 238.900 ;
        RECT 20.330 238.800 29.130 238.900 ;
        RECT 18.730 238.450 22.930 238.650 ;
        RECT 6.530 238.300 14.080 238.450 ;
        RECT 15.430 238.300 22.930 238.450 ;
        RECT 6.530 238.000 10.730 238.300 ;
        RECT 2.315 233.250 4.315 235.545 ;
        RECT 6.530 235.150 6.680 238.000 ;
        RECT 7.130 230.450 7.280 238.000 ;
        RECT 7.730 230.450 7.880 238.000 ;
        RECT 8.330 230.450 8.480 238.000 ;
        RECT 8.930 230.450 9.080 238.000 ;
        RECT 9.530 230.450 9.680 238.000 ;
        RECT 10.130 237.850 10.730 238.000 ;
        RECT 18.730 238.000 22.930 238.300 ;
        RECT 18.730 237.850 19.330 238.000 ;
        RECT 10.130 237.700 14.080 237.850 ;
        RECT 15.380 237.700 19.330 237.850 ;
        RECT 10.130 237.250 10.730 237.700 ;
        RECT 18.730 237.250 19.330 237.700 ;
        RECT 10.130 237.100 14.080 237.250 ;
        RECT 15.380 237.100 19.330 237.250 ;
        RECT 10.130 236.650 10.730 237.100 ;
        RECT 18.730 236.650 19.330 237.100 ;
        RECT 10.130 236.500 14.080 236.650 ;
        RECT 15.380 236.500 19.330 236.650 ;
        RECT 10.130 236.050 10.730 236.500 ;
        RECT 18.730 236.050 19.330 236.500 ;
        RECT 10.130 235.900 14.080 236.050 ;
        RECT 15.380 235.900 19.330 236.050 ;
        RECT 10.130 235.450 10.730 235.900 ;
        RECT 18.730 235.450 19.330 235.900 ;
        RECT 10.130 235.300 14.080 235.450 ;
        RECT 15.380 235.300 19.330 235.450 ;
        RECT 10.130 234.850 10.730 235.300 ;
        RECT 18.730 234.850 19.330 235.300 ;
        RECT 10.130 234.700 14.080 234.850 ;
        RECT 15.380 234.700 19.330 234.850 ;
        RECT 10.130 234.250 10.730 234.700 ;
        RECT 18.730 234.250 19.330 234.700 ;
        RECT 10.130 234.100 14.080 234.250 ;
        RECT 15.380 234.100 19.330 234.250 ;
        RECT 10.130 233.650 10.730 234.100 ;
        RECT 18.730 233.650 19.330 234.100 ;
        RECT 10.130 233.500 14.080 233.650 ;
        RECT 15.380 233.500 19.330 233.650 ;
        RECT 10.130 233.050 10.730 233.500 ;
        RECT 18.730 233.050 19.330 233.500 ;
        RECT 10.130 232.900 14.080 233.050 ;
        RECT 15.380 232.900 19.330 233.050 ;
        RECT 10.130 232.450 10.730 232.900 ;
        RECT 18.730 232.450 19.330 232.900 ;
        RECT 10.130 232.300 14.080 232.450 ;
        RECT 15.380 232.300 19.330 232.450 ;
        RECT 10.130 231.850 10.730 232.300 ;
        RECT 18.730 231.850 19.330 232.300 ;
        RECT 10.130 231.700 14.080 231.850 ;
        RECT 15.380 231.700 19.330 231.850 ;
        RECT 10.130 231.250 10.730 231.700 ;
        RECT 18.730 231.250 19.330 231.700 ;
        RECT 10.130 231.100 14.080 231.250 ;
        RECT 15.380 231.100 19.330 231.250 ;
        RECT 10.130 230.650 10.730 231.100 ;
        RECT 18.730 230.650 19.330 231.100 ;
        RECT 10.130 230.450 14.080 230.650 ;
        RECT 15.380 230.450 19.330 230.650 ;
        RECT 19.780 230.450 19.930 238.000 ;
        RECT 20.380 230.450 20.530 238.000 ;
        RECT 20.980 230.450 21.130 238.000 ;
        RECT 21.580 230.450 21.730 238.000 ;
        RECT 22.180 230.450 22.330 238.000 ;
        RECT 22.780 235.150 22.930 238.000 ;
        RECT 23.530 235.600 25.930 238.800 ;
        RECT 29.280 238.650 30.730 238.950 ;
        RECT 26.530 238.450 30.730 238.650 ;
        RECT 38.730 238.950 50.730 239.800 ;
        RECT 38.730 238.900 49.130 238.950 ;
        RECT 38.730 238.650 40.180 238.900 ;
        RECT 40.330 238.800 49.130 238.900 ;
        RECT 38.730 238.450 42.930 238.650 ;
        RECT 26.530 238.300 34.080 238.450 ;
        RECT 35.430 238.300 42.930 238.450 ;
        RECT 26.530 238.000 30.730 238.300 ;
        RECT 26.530 235.150 26.680 238.000 ;
        RECT 27.130 230.450 27.280 238.000 ;
        RECT 27.730 230.450 27.880 238.000 ;
        RECT 28.330 230.450 28.480 238.000 ;
        RECT 28.930 230.450 29.080 238.000 ;
        RECT 29.530 230.450 29.680 238.000 ;
        RECT 30.130 237.850 30.730 238.000 ;
        RECT 38.730 238.000 42.930 238.300 ;
        RECT 38.730 237.850 39.330 238.000 ;
        RECT 30.130 237.700 34.080 237.850 ;
        RECT 35.380 237.700 39.330 237.850 ;
        RECT 30.130 237.250 30.730 237.700 ;
        RECT 38.730 237.250 39.330 237.700 ;
        RECT 30.130 237.100 34.080 237.250 ;
        RECT 35.380 237.100 39.330 237.250 ;
        RECT 30.130 236.650 30.730 237.100 ;
        RECT 38.730 236.650 39.330 237.100 ;
        RECT 30.130 236.500 34.080 236.650 ;
        RECT 35.380 236.500 39.330 236.650 ;
        RECT 30.130 236.050 30.730 236.500 ;
        RECT 38.730 236.050 39.330 236.500 ;
        RECT 30.130 235.900 34.080 236.050 ;
        RECT 35.380 235.900 39.330 236.050 ;
        RECT 30.130 235.450 30.730 235.900 ;
        RECT 38.730 235.450 39.330 235.900 ;
        RECT 30.130 235.300 34.080 235.450 ;
        RECT 35.380 235.300 39.330 235.450 ;
        RECT 30.130 234.850 30.730 235.300 ;
        RECT 38.730 234.850 39.330 235.300 ;
        RECT 30.130 234.700 34.080 234.850 ;
        RECT 35.380 234.700 39.330 234.850 ;
        RECT 30.130 234.250 30.730 234.700 ;
        RECT 38.730 234.250 39.330 234.700 ;
        RECT 30.130 234.100 34.080 234.250 ;
        RECT 35.380 234.100 39.330 234.250 ;
        RECT 30.130 233.650 30.730 234.100 ;
        RECT 38.730 233.650 39.330 234.100 ;
        RECT 30.130 233.500 34.080 233.650 ;
        RECT 35.380 233.500 39.330 233.650 ;
        RECT 30.130 233.050 30.730 233.500 ;
        RECT 38.730 233.050 39.330 233.500 ;
        RECT 30.130 232.900 34.080 233.050 ;
        RECT 35.380 232.900 39.330 233.050 ;
        RECT 30.130 232.450 30.730 232.900 ;
        RECT 38.730 232.450 39.330 232.900 ;
        RECT 30.130 232.300 34.080 232.450 ;
        RECT 35.380 232.300 39.330 232.450 ;
        RECT 30.130 231.850 30.730 232.300 ;
        RECT 38.730 231.850 39.330 232.300 ;
        RECT 30.130 231.700 34.080 231.850 ;
        RECT 35.380 231.700 39.330 231.850 ;
        RECT 30.130 231.250 30.730 231.700 ;
        RECT 38.730 231.250 39.330 231.700 ;
        RECT 30.130 231.100 34.080 231.250 ;
        RECT 35.380 231.100 39.330 231.250 ;
        RECT 30.130 230.650 30.730 231.100 ;
        RECT 38.730 230.650 39.330 231.100 ;
        RECT 30.130 230.450 34.080 230.650 ;
        RECT 35.380 230.450 39.330 230.650 ;
        RECT 39.780 230.450 39.930 238.000 ;
        RECT 40.380 230.450 40.530 238.000 ;
        RECT 40.980 230.450 41.130 238.000 ;
        RECT 41.580 230.450 41.730 238.000 ;
        RECT 42.180 230.450 42.330 238.000 ;
        RECT 42.780 235.150 42.930 238.000 ;
        RECT 43.530 235.600 45.930 238.800 ;
        RECT 49.280 238.650 50.730 238.950 ;
        RECT 46.530 238.450 50.730 238.650 ;
        RECT 58.730 238.950 70.730 239.800 ;
        RECT 58.730 238.900 69.130 238.950 ;
        RECT 58.730 238.650 60.180 238.900 ;
        RECT 60.330 238.800 69.130 238.900 ;
        RECT 58.730 238.450 62.930 238.650 ;
        RECT 46.530 238.300 54.080 238.450 ;
        RECT 55.430 238.300 62.930 238.450 ;
        RECT 46.530 238.000 50.730 238.300 ;
        RECT 46.530 235.150 46.680 238.000 ;
        RECT 47.130 230.450 47.280 238.000 ;
        RECT 47.730 230.450 47.880 238.000 ;
        RECT 48.330 230.450 48.480 238.000 ;
        RECT 48.930 230.450 49.080 238.000 ;
        RECT 49.530 230.450 49.680 238.000 ;
        RECT 50.130 237.850 50.730 238.000 ;
        RECT 58.730 238.000 62.930 238.300 ;
        RECT 58.730 237.850 59.330 238.000 ;
        RECT 50.130 237.700 54.080 237.850 ;
        RECT 55.380 237.700 59.330 237.850 ;
        RECT 50.130 237.250 50.730 237.700 ;
        RECT 58.730 237.250 59.330 237.700 ;
        RECT 50.130 237.100 54.080 237.250 ;
        RECT 55.380 237.100 59.330 237.250 ;
        RECT 50.130 236.650 50.730 237.100 ;
        RECT 58.730 236.650 59.330 237.100 ;
        RECT 50.130 236.500 54.080 236.650 ;
        RECT 55.380 236.500 59.330 236.650 ;
        RECT 50.130 236.050 50.730 236.500 ;
        RECT 58.730 236.050 59.330 236.500 ;
        RECT 50.130 235.900 54.080 236.050 ;
        RECT 55.380 235.900 59.330 236.050 ;
        RECT 50.130 235.450 50.730 235.900 ;
        RECT 58.730 235.450 59.330 235.900 ;
        RECT 50.130 235.300 54.080 235.450 ;
        RECT 55.380 235.300 59.330 235.450 ;
        RECT 50.130 234.850 50.730 235.300 ;
        RECT 58.730 234.850 59.330 235.300 ;
        RECT 50.130 234.700 54.080 234.850 ;
        RECT 55.380 234.700 59.330 234.850 ;
        RECT 50.130 234.250 50.730 234.700 ;
        RECT 58.730 234.250 59.330 234.700 ;
        RECT 50.130 234.100 54.080 234.250 ;
        RECT 55.380 234.100 59.330 234.250 ;
        RECT 50.130 233.650 50.730 234.100 ;
        RECT 58.730 233.650 59.330 234.100 ;
        RECT 50.130 233.500 54.080 233.650 ;
        RECT 55.380 233.500 59.330 233.650 ;
        RECT 50.130 233.050 50.730 233.500 ;
        RECT 58.730 233.050 59.330 233.500 ;
        RECT 50.130 232.900 54.080 233.050 ;
        RECT 55.380 232.900 59.330 233.050 ;
        RECT 50.130 232.450 50.730 232.900 ;
        RECT 58.730 232.450 59.330 232.900 ;
        RECT 50.130 232.300 54.080 232.450 ;
        RECT 55.380 232.300 59.330 232.450 ;
        RECT 50.130 231.850 50.730 232.300 ;
        RECT 58.730 231.850 59.330 232.300 ;
        RECT 50.130 231.700 54.080 231.850 ;
        RECT 55.380 231.700 59.330 231.850 ;
        RECT 50.130 231.250 50.730 231.700 ;
        RECT 58.730 231.250 59.330 231.700 ;
        RECT 50.130 231.100 54.080 231.250 ;
        RECT 55.380 231.100 59.330 231.250 ;
        RECT 50.130 230.650 50.730 231.100 ;
        RECT 58.730 230.650 59.330 231.100 ;
        RECT 50.130 230.450 54.080 230.650 ;
        RECT 55.380 230.450 59.330 230.650 ;
        RECT 59.780 230.450 59.930 238.000 ;
        RECT 60.380 230.450 60.530 238.000 ;
        RECT 60.980 230.450 61.130 238.000 ;
        RECT 61.580 230.450 61.730 238.000 ;
        RECT 62.180 230.450 62.330 238.000 ;
        RECT 62.780 235.150 62.930 238.000 ;
        RECT 63.530 235.600 65.930 238.800 ;
        RECT 69.280 238.650 70.730 238.950 ;
        RECT 66.530 238.450 70.730 238.650 ;
        RECT 78.730 238.950 90.730 239.800 ;
        RECT 78.730 238.900 89.130 238.950 ;
        RECT 78.730 238.650 80.180 238.900 ;
        RECT 80.330 238.800 89.130 238.900 ;
        RECT 78.730 238.450 82.930 238.650 ;
        RECT 66.530 238.300 74.080 238.450 ;
        RECT 75.430 238.300 82.930 238.450 ;
        RECT 66.530 238.000 70.730 238.300 ;
        RECT 66.530 235.150 66.680 238.000 ;
        RECT 67.130 230.450 67.280 238.000 ;
        RECT 67.730 230.450 67.880 238.000 ;
        RECT 68.330 230.450 68.480 238.000 ;
        RECT 68.930 230.450 69.080 238.000 ;
        RECT 69.530 230.450 69.680 238.000 ;
        RECT 70.130 237.850 70.730 238.000 ;
        RECT 78.730 238.000 82.930 238.300 ;
        RECT 78.730 237.850 79.330 238.000 ;
        RECT 70.130 237.700 74.080 237.850 ;
        RECT 75.380 237.700 79.330 237.850 ;
        RECT 70.130 237.250 70.730 237.700 ;
        RECT 78.730 237.250 79.330 237.700 ;
        RECT 70.130 237.100 74.080 237.250 ;
        RECT 75.380 237.100 79.330 237.250 ;
        RECT 70.130 236.650 70.730 237.100 ;
        RECT 78.730 236.650 79.330 237.100 ;
        RECT 70.130 236.500 74.080 236.650 ;
        RECT 75.380 236.500 79.330 236.650 ;
        RECT 70.130 236.050 70.730 236.500 ;
        RECT 78.730 236.050 79.330 236.500 ;
        RECT 70.130 235.900 74.080 236.050 ;
        RECT 75.380 235.900 79.330 236.050 ;
        RECT 70.130 235.450 70.730 235.900 ;
        RECT 78.730 235.450 79.330 235.900 ;
        RECT 70.130 235.300 74.080 235.450 ;
        RECT 75.380 235.300 79.330 235.450 ;
        RECT 70.130 234.850 70.730 235.300 ;
        RECT 78.730 234.850 79.330 235.300 ;
        RECT 70.130 234.700 74.080 234.850 ;
        RECT 75.380 234.700 79.330 234.850 ;
        RECT 70.130 234.250 70.730 234.700 ;
        RECT 78.730 234.250 79.330 234.700 ;
        RECT 70.130 234.100 74.080 234.250 ;
        RECT 75.380 234.100 79.330 234.250 ;
        RECT 70.130 233.650 70.730 234.100 ;
        RECT 78.730 233.650 79.330 234.100 ;
        RECT 70.130 233.500 74.080 233.650 ;
        RECT 75.380 233.500 79.330 233.650 ;
        RECT 70.130 233.050 70.730 233.500 ;
        RECT 78.730 233.050 79.330 233.500 ;
        RECT 70.130 232.900 74.080 233.050 ;
        RECT 75.380 232.900 79.330 233.050 ;
        RECT 70.130 232.450 70.730 232.900 ;
        RECT 78.730 232.450 79.330 232.900 ;
        RECT 70.130 232.300 74.080 232.450 ;
        RECT 75.380 232.300 79.330 232.450 ;
        RECT 70.130 231.850 70.730 232.300 ;
        RECT 78.730 231.850 79.330 232.300 ;
        RECT 70.130 231.700 74.080 231.850 ;
        RECT 75.380 231.700 79.330 231.850 ;
        RECT 70.130 231.250 70.730 231.700 ;
        RECT 78.730 231.250 79.330 231.700 ;
        RECT 70.130 231.100 74.080 231.250 ;
        RECT 75.380 231.100 79.330 231.250 ;
        RECT 70.130 230.650 70.730 231.100 ;
        RECT 78.730 230.650 79.330 231.100 ;
        RECT 70.130 230.450 74.080 230.650 ;
        RECT 75.380 230.450 79.330 230.650 ;
        RECT 79.780 230.450 79.930 238.000 ;
        RECT 80.380 230.450 80.530 238.000 ;
        RECT 80.980 230.450 81.130 238.000 ;
        RECT 81.580 230.450 81.730 238.000 ;
        RECT 82.180 230.450 82.330 238.000 ;
        RECT 82.780 235.150 82.930 238.000 ;
        RECT 83.530 235.600 85.930 238.800 ;
        RECT 89.280 238.650 90.730 238.950 ;
        RECT 86.530 238.450 90.730 238.650 ;
        RECT 98.730 238.950 110.730 239.800 ;
        RECT 98.730 238.900 109.130 238.950 ;
        RECT 98.730 238.650 100.180 238.900 ;
        RECT 100.330 238.800 109.130 238.900 ;
        RECT 98.730 238.450 102.930 238.650 ;
        RECT 86.530 238.300 94.080 238.450 ;
        RECT 95.430 238.300 102.930 238.450 ;
        RECT 86.530 238.000 90.730 238.300 ;
        RECT 86.530 235.150 86.680 238.000 ;
        RECT 87.130 230.450 87.280 238.000 ;
        RECT 87.730 230.450 87.880 238.000 ;
        RECT 88.330 230.450 88.480 238.000 ;
        RECT 88.930 230.450 89.080 238.000 ;
        RECT 89.530 230.450 89.680 238.000 ;
        RECT 90.130 237.850 90.730 238.000 ;
        RECT 98.730 238.000 102.930 238.300 ;
        RECT 98.730 237.850 99.330 238.000 ;
        RECT 90.130 237.700 94.080 237.850 ;
        RECT 95.380 237.700 99.330 237.850 ;
        RECT 90.130 237.250 90.730 237.700 ;
        RECT 98.730 237.250 99.330 237.700 ;
        RECT 90.130 237.100 94.080 237.250 ;
        RECT 95.380 237.100 99.330 237.250 ;
        RECT 90.130 236.650 90.730 237.100 ;
        RECT 98.730 236.650 99.330 237.100 ;
        RECT 90.130 236.500 94.080 236.650 ;
        RECT 95.380 236.500 99.330 236.650 ;
        RECT 90.130 236.050 90.730 236.500 ;
        RECT 98.730 236.050 99.330 236.500 ;
        RECT 90.130 235.900 94.080 236.050 ;
        RECT 95.380 235.900 99.330 236.050 ;
        RECT 90.130 235.450 90.730 235.900 ;
        RECT 98.730 235.450 99.330 235.900 ;
        RECT 90.130 235.300 94.080 235.450 ;
        RECT 95.380 235.300 99.330 235.450 ;
        RECT 90.130 234.850 90.730 235.300 ;
        RECT 98.730 234.850 99.330 235.300 ;
        RECT 90.130 234.700 94.080 234.850 ;
        RECT 95.380 234.700 99.330 234.850 ;
        RECT 90.130 234.250 90.730 234.700 ;
        RECT 98.730 234.250 99.330 234.700 ;
        RECT 90.130 234.100 94.080 234.250 ;
        RECT 95.380 234.100 99.330 234.250 ;
        RECT 90.130 233.650 90.730 234.100 ;
        RECT 98.730 233.650 99.330 234.100 ;
        RECT 90.130 233.500 94.080 233.650 ;
        RECT 95.380 233.500 99.330 233.650 ;
        RECT 90.130 233.050 90.730 233.500 ;
        RECT 98.730 233.050 99.330 233.500 ;
        RECT 90.130 232.900 94.080 233.050 ;
        RECT 95.380 232.900 99.330 233.050 ;
        RECT 90.130 232.450 90.730 232.900 ;
        RECT 98.730 232.450 99.330 232.900 ;
        RECT 90.130 232.300 94.080 232.450 ;
        RECT 95.380 232.300 99.330 232.450 ;
        RECT 90.130 231.850 90.730 232.300 ;
        RECT 98.730 231.850 99.330 232.300 ;
        RECT 90.130 231.700 94.080 231.850 ;
        RECT 95.380 231.700 99.330 231.850 ;
        RECT 90.130 231.250 90.730 231.700 ;
        RECT 98.730 231.250 99.330 231.700 ;
        RECT 90.130 231.100 94.080 231.250 ;
        RECT 95.380 231.100 99.330 231.250 ;
        RECT 90.130 230.650 90.730 231.100 ;
        RECT 98.730 230.650 99.330 231.100 ;
        RECT 90.130 230.450 94.080 230.650 ;
        RECT 95.380 230.450 99.330 230.650 ;
        RECT 99.780 230.450 99.930 238.000 ;
        RECT 100.380 230.450 100.530 238.000 ;
        RECT 100.980 230.450 101.130 238.000 ;
        RECT 101.580 230.450 101.730 238.000 ;
        RECT 102.180 230.450 102.330 238.000 ;
        RECT 102.780 235.150 102.930 238.000 ;
        RECT 103.530 235.600 105.930 238.800 ;
        RECT 109.280 238.650 110.730 238.950 ;
        RECT 106.530 238.450 110.730 238.650 ;
        RECT 118.730 238.900 124.730 239.800 ;
        RECT 118.730 238.650 120.180 238.900 ;
        RECT 120.330 238.800 124.730 238.900 ;
        RECT 118.730 238.450 122.930 238.650 ;
        RECT 106.530 238.300 114.080 238.450 ;
        RECT 115.430 238.300 122.930 238.450 ;
        RECT 106.530 238.000 110.730 238.300 ;
        RECT 106.530 235.150 106.680 238.000 ;
        RECT 107.130 230.450 107.280 238.000 ;
        RECT 107.730 230.450 107.880 238.000 ;
        RECT 108.330 230.450 108.480 238.000 ;
        RECT 108.930 230.450 109.080 238.000 ;
        RECT 109.530 230.450 109.680 238.000 ;
        RECT 110.130 237.850 110.730 238.000 ;
        RECT 118.730 238.000 122.930 238.300 ;
        RECT 118.730 237.850 119.330 238.000 ;
        RECT 110.130 237.700 114.080 237.850 ;
        RECT 115.380 237.700 119.330 237.850 ;
        RECT 110.130 237.250 110.730 237.700 ;
        RECT 118.730 237.250 119.330 237.700 ;
        RECT 110.130 237.100 114.080 237.250 ;
        RECT 115.380 237.100 119.330 237.250 ;
        RECT 110.130 236.650 110.730 237.100 ;
        RECT 118.730 236.650 119.330 237.100 ;
        RECT 110.130 236.500 114.080 236.650 ;
        RECT 115.380 236.500 119.330 236.650 ;
        RECT 110.130 236.050 110.730 236.500 ;
        RECT 118.730 236.050 119.330 236.500 ;
        RECT 110.130 235.900 114.080 236.050 ;
        RECT 115.380 235.900 119.330 236.050 ;
        RECT 110.130 235.450 110.730 235.900 ;
        RECT 118.730 235.450 119.330 235.900 ;
        RECT 110.130 235.300 114.080 235.450 ;
        RECT 115.380 235.300 119.330 235.450 ;
        RECT 110.130 234.850 110.730 235.300 ;
        RECT 118.730 234.850 119.330 235.300 ;
        RECT 110.130 234.700 114.080 234.850 ;
        RECT 115.380 234.700 119.330 234.850 ;
        RECT 110.130 234.250 110.730 234.700 ;
        RECT 118.730 234.250 119.330 234.700 ;
        RECT 110.130 234.100 114.080 234.250 ;
        RECT 115.380 234.100 119.330 234.250 ;
        RECT 110.130 233.650 110.730 234.100 ;
        RECT 118.730 233.650 119.330 234.100 ;
        RECT 110.130 233.500 114.080 233.650 ;
        RECT 115.380 233.500 119.330 233.650 ;
        RECT 110.130 233.050 110.730 233.500 ;
        RECT 118.730 233.050 119.330 233.500 ;
        RECT 110.130 232.900 114.080 233.050 ;
        RECT 115.380 232.900 119.330 233.050 ;
        RECT 110.130 232.450 110.730 232.900 ;
        RECT 118.730 232.450 119.330 232.900 ;
        RECT 110.130 232.300 114.080 232.450 ;
        RECT 115.380 232.300 119.330 232.450 ;
        RECT 110.130 231.850 110.730 232.300 ;
        RECT 118.730 231.850 119.330 232.300 ;
        RECT 110.130 231.700 114.080 231.850 ;
        RECT 115.380 231.700 119.330 231.850 ;
        RECT 110.130 231.250 110.730 231.700 ;
        RECT 118.730 231.250 119.330 231.700 ;
        RECT 110.130 231.100 114.080 231.250 ;
        RECT 115.380 231.100 119.330 231.250 ;
        RECT 110.130 230.650 110.730 231.100 ;
        RECT 118.730 230.650 119.330 231.100 ;
        RECT 110.130 230.450 114.080 230.650 ;
        RECT 115.380 230.450 119.330 230.650 ;
        RECT 119.780 230.450 119.930 238.000 ;
        RECT 120.380 230.450 120.530 238.000 ;
        RECT 120.980 230.450 121.130 238.000 ;
        RECT 121.580 230.450 121.730 238.000 ;
        RECT 122.180 230.450 122.330 238.000 ;
        RECT 122.780 235.150 122.930 238.000 ;
        RECT 123.530 237.325 124.730 238.800 ;
        RECT 123.530 236.050 127.140 237.325 ;
        RECT 123.530 235.600 124.730 236.050 ;
        RECT 2.315 224.455 4.315 226.750 ;
        RECT 4.730 223.735 5.930 224.400 ;
        RECT 2.315 222.460 5.930 223.735 ;
        RECT 4.730 221.200 5.930 222.460 ;
        RECT 6.530 222.000 6.680 224.900 ;
        RECT 7.130 222.000 7.280 229.550 ;
        RECT 7.730 222.000 7.880 229.550 ;
        RECT 8.330 222.000 8.480 229.550 ;
        RECT 8.930 222.000 9.080 229.550 ;
        RECT 9.530 222.000 9.680 229.550 ;
        RECT 10.130 229.350 14.080 229.550 ;
        RECT 15.380 229.350 19.330 229.550 ;
        RECT 10.130 228.900 10.730 229.350 ;
        RECT 18.730 228.900 19.330 229.350 ;
        RECT 10.130 228.750 14.080 228.900 ;
        RECT 15.380 228.750 19.330 228.900 ;
        RECT 10.130 228.300 10.730 228.750 ;
        RECT 18.730 228.300 19.330 228.750 ;
        RECT 10.130 228.150 14.080 228.300 ;
        RECT 15.380 228.150 19.330 228.300 ;
        RECT 10.130 227.700 10.730 228.150 ;
        RECT 18.730 227.700 19.330 228.150 ;
        RECT 10.130 227.550 14.080 227.700 ;
        RECT 15.380 227.550 19.330 227.700 ;
        RECT 10.130 227.100 10.730 227.550 ;
        RECT 18.730 227.100 19.330 227.550 ;
        RECT 10.130 226.950 14.080 227.100 ;
        RECT 15.380 226.950 19.330 227.100 ;
        RECT 10.130 226.500 10.730 226.950 ;
        RECT 18.730 226.500 19.330 226.950 ;
        RECT 10.130 226.350 14.080 226.500 ;
        RECT 15.380 226.350 19.330 226.500 ;
        RECT 10.130 225.900 10.730 226.350 ;
        RECT 18.730 225.900 19.330 226.350 ;
        RECT 10.130 225.750 14.080 225.900 ;
        RECT 15.380 225.750 19.330 225.900 ;
        RECT 10.130 225.300 10.730 225.750 ;
        RECT 18.730 225.300 19.330 225.750 ;
        RECT 10.130 225.150 14.080 225.300 ;
        RECT 15.380 225.150 19.330 225.300 ;
        RECT 10.130 224.700 10.730 225.150 ;
        RECT 18.730 224.700 19.330 225.150 ;
        RECT 10.130 224.550 14.080 224.700 ;
        RECT 15.380 224.550 19.330 224.700 ;
        RECT 10.130 224.100 10.730 224.550 ;
        RECT 18.730 224.100 19.330 224.550 ;
        RECT 10.130 223.950 14.080 224.100 ;
        RECT 15.380 223.950 19.330 224.100 ;
        RECT 10.130 223.500 10.730 223.950 ;
        RECT 18.730 223.500 19.330 223.950 ;
        RECT 10.130 223.350 14.080 223.500 ;
        RECT 15.380 223.350 19.330 223.500 ;
        RECT 10.130 222.900 10.730 223.350 ;
        RECT 18.730 222.900 19.330 223.350 ;
        RECT 10.130 222.750 14.080 222.900 ;
        RECT 15.380 222.750 19.330 222.900 ;
        RECT 10.130 222.300 10.730 222.750 ;
        RECT 18.730 222.300 19.330 222.750 ;
        RECT 10.130 222.150 14.080 222.300 ;
        RECT 15.380 222.150 19.330 222.300 ;
        RECT 10.130 222.000 10.730 222.150 ;
        RECT 6.530 221.700 10.730 222.000 ;
        RECT 18.730 222.000 19.330 222.150 ;
        RECT 19.780 222.000 19.930 229.550 ;
        RECT 20.380 222.000 20.530 229.550 ;
        RECT 20.980 222.000 21.130 229.550 ;
        RECT 21.580 222.000 21.730 229.550 ;
        RECT 22.180 222.000 22.330 229.550 ;
        RECT 22.780 222.000 22.930 224.900 ;
        RECT 18.730 221.700 22.930 222.000 ;
        RECT 6.530 221.550 14.080 221.700 ;
        RECT 15.380 221.550 22.930 221.700 ;
        RECT 6.530 221.350 10.730 221.550 ;
        RECT 4.730 221.050 9.130 221.200 ;
        RECT 9.280 221.050 10.730 221.350 ;
        RECT 4.730 220.150 10.730 221.050 ;
        RECT 18.730 221.350 22.930 221.550 ;
        RECT 18.730 221.050 20.180 221.350 ;
        RECT 23.530 221.200 25.930 224.400 ;
        RECT 26.530 222.000 26.680 224.900 ;
        RECT 27.130 222.000 27.280 229.550 ;
        RECT 27.730 222.000 27.880 229.550 ;
        RECT 28.330 222.000 28.480 229.550 ;
        RECT 28.930 222.000 29.080 229.550 ;
        RECT 29.530 222.000 29.680 229.550 ;
        RECT 30.130 229.350 34.080 229.550 ;
        RECT 35.380 229.350 39.330 229.550 ;
        RECT 30.130 228.900 30.730 229.350 ;
        RECT 38.730 228.900 39.330 229.350 ;
        RECT 30.130 228.750 34.080 228.900 ;
        RECT 35.380 228.750 39.330 228.900 ;
        RECT 30.130 228.300 30.730 228.750 ;
        RECT 38.730 228.300 39.330 228.750 ;
        RECT 30.130 228.150 34.080 228.300 ;
        RECT 35.380 228.150 39.330 228.300 ;
        RECT 30.130 227.700 30.730 228.150 ;
        RECT 38.730 227.700 39.330 228.150 ;
        RECT 30.130 227.550 34.080 227.700 ;
        RECT 35.380 227.550 39.330 227.700 ;
        RECT 30.130 227.100 30.730 227.550 ;
        RECT 38.730 227.100 39.330 227.550 ;
        RECT 30.130 226.950 34.080 227.100 ;
        RECT 35.380 226.950 39.330 227.100 ;
        RECT 30.130 226.500 30.730 226.950 ;
        RECT 38.730 226.500 39.330 226.950 ;
        RECT 30.130 226.350 34.080 226.500 ;
        RECT 35.380 226.350 39.330 226.500 ;
        RECT 30.130 225.900 30.730 226.350 ;
        RECT 38.730 225.900 39.330 226.350 ;
        RECT 30.130 225.750 34.080 225.900 ;
        RECT 35.380 225.750 39.330 225.900 ;
        RECT 30.130 225.300 30.730 225.750 ;
        RECT 38.730 225.300 39.330 225.750 ;
        RECT 30.130 225.150 34.080 225.300 ;
        RECT 35.380 225.150 39.330 225.300 ;
        RECT 30.130 224.700 30.730 225.150 ;
        RECT 38.730 224.700 39.330 225.150 ;
        RECT 30.130 224.550 34.080 224.700 ;
        RECT 35.380 224.550 39.330 224.700 ;
        RECT 30.130 224.100 30.730 224.550 ;
        RECT 38.730 224.100 39.330 224.550 ;
        RECT 30.130 223.950 34.080 224.100 ;
        RECT 35.380 223.950 39.330 224.100 ;
        RECT 30.130 223.500 30.730 223.950 ;
        RECT 38.730 223.500 39.330 223.950 ;
        RECT 30.130 223.350 34.080 223.500 ;
        RECT 35.380 223.350 39.330 223.500 ;
        RECT 30.130 222.900 30.730 223.350 ;
        RECT 38.730 222.900 39.330 223.350 ;
        RECT 30.130 222.750 34.080 222.900 ;
        RECT 35.380 222.750 39.330 222.900 ;
        RECT 30.130 222.300 30.730 222.750 ;
        RECT 38.730 222.300 39.330 222.750 ;
        RECT 30.130 222.150 34.080 222.300 ;
        RECT 35.380 222.150 39.330 222.300 ;
        RECT 30.130 222.000 30.730 222.150 ;
        RECT 26.530 221.700 30.730 222.000 ;
        RECT 38.730 222.000 39.330 222.150 ;
        RECT 39.780 222.000 39.930 229.550 ;
        RECT 40.380 222.000 40.530 229.550 ;
        RECT 40.980 222.000 41.130 229.550 ;
        RECT 41.580 222.000 41.730 229.550 ;
        RECT 42.180 222.000 42.330 229.550 ;
        RECT 42.780 222.000 42.930 224.900 ;
        RECT 38.730 221.700 42.930 222.000 ;
        RECT 26.530 221.550 34.080 221.700 ;
        RECT 35.380 221.550 42.930 221.700 ;
        RECT 26.530 221.350 30.730 221.550 ;
        RECT 20.330 221.050 29.130 221.200 ;
        RECT 29.280 221.050 30.730 221.350 ;
        RECT 18.730 220.150 30.730 221.050 ;
        RECT 38.730 221.350 42.930 221.550 ;
        RECT 38.730 221.050 40.180 221.350 ;
        RECT 43.530 221.200 45.930 224.400 ;
        RECT 46.530 222.000 46.680 224.900 ;
        RECT 47.130 222.000 47.280 229.550 ;
        RECT 47.730 222.000 47.880 229.550 ;
        RECT 48.330 222.000 48.480 229.550 ;
        RECT 48.930 222.000 49.080 229.550 ;
        RECT 49.530 222.000 49.680 229.550 ;
        RECT 50.130 229.350 54.080 229.550 ;
        RECT 55.380 229.350 59.330 229.550 ;
        RECT 50.130 228.900 50.730 229.350 ;
        RECT 58.730 228.900 59.330 229.350 ;
        RECT 50.130 228.750 54.080 228.900 ;
        RECT 55.380 228.750 59.330 228.900 ;
        RECT 50.130 228.300 50.730 228.750 ;
        RECT 58.730 228.300 59.330 228.750 ;
        RECT 50.130 228.150 54.080 228.300 ;
        RECT 55.380 228.150 59.330 228.300 ;
        RECT 50.130 227.700 50.730 228.150 ;
        RECT 58.730 227.700 59.330 228.150 ;
        RECT 50.130 227.550 54.080 227.700 ;
        RECT 55.380 227.550 59.330 227.700 ;
        RECT 50.130 227.100 50.730 227.550 ;
        RECT 58.730 227.100 59.330 227.550 ;
        RECT 50.130 226.950 54.080 227.100 ;
        RECT 55.380 226.950 59.330 227.100 ;
        RECT 50.130 226.500 50.730 226.950 ;
        RECT 58.730 226.500 59.330 226.950 ;
        RECT 50.130 226.350 54.080 226.500 ;
        RECT 55.380 226.350 59.330 226.500 ;
        RECT 50.130 225.900 50.730 226.350 ;
        RECT 58.730 225.900 59.330 226.350 ;
        RECT 50.130 225.750 54.080 225.900 ;
        RECT 55.380 225.750 59.330 225.900 ;
        RECT 50.130 225.300 50.730 225.750 ;
        RECT 58.730 225.300 59.330 225.750 ;
        RECT 50.130 225.150 54.080 225.300 ;
        RECT 55.380 225.150 59.330 225.300 ;
        RECT 50.130 224.700 50.730 225.150 ;
        RECT 58.730 224.700 59.330 225.150 ;
        RECT 50.130 224.550 54.080 224.700 ;
        RECT 55.380 224.550 59.330 224.700 ;
        RECT 50.130 224.100 50.730 224.550 ;
        RECT 58.730 224.100 59.330 224.550 ;
        RECT 50.130 223.950 54.080 224.100 ;
        RECT 55.380 223.950 59.330 224.100 ;
        RECT 50.130 223.500 50.730 223.950 ;
        RECT 58.730 223.500 59.330 223.950 ;
        RECT 50.130 223.350 54.080 223.500 ;
        RECT 55.380 223.350 59.330 223.500 ;
        RECT 50.130 222.900 50.730 223.350 ;
        RECT 58.730 222.900 59.330 223.350 ;
        RECT 50.130 222.750 54.080 222.900 ;
        RECT 55.380 222.750 59.330 222.900 ;
        RECT 50.130 222.300 50.730 222.750 ;
        RECT 58.730 222.300 59.330 222.750 ;
        RECT 50.130 222.150 54.080 222.300 ;
        RECT 55.380 222.150 59.330 222.300 ;
        RECT 50.130 222.000 50.730 222.150 ;
        RECT 46.530 221.700 50.730 222.000 ;
        RECT 58.730 222.000 59.330 222.150 ;
        RECT 59.780 222.000 59.930 229.550 ;
        RECT 60.380 222.000 60.530 229.550 ;
        RECT 60.980 222.000 61.130 229.550 ;
        RECT 61.580 222.000 61.730 229.550 ;
        RECT 62.180 222.000 62.330 229.550 ;
        RECT 62.780 222.000 62.930 224.900 ;
        RECT 58.730 221.700 62.930 222.000 ;
        RECT 46.530 221.550 54.080 221.700 ;
        RECT 55.380 221.550 62.930 221.700 ;
        RECT 46.530 221.350 50.730 221.550 ;
        RECT 40.330 221.050 49.130 221.200 ;
        RECT 49.280 221.050 50.730 221.350 ;
        RECT 38.730 220.150 50.730 221.050 ;
        RECT 58.730 221.350 62.930 221.550 ;
        RECT 58.730 221.050 60.180 221.350 ;
        RECT 63.530 221.200 65.930 224.400 ;
        RECT 66.530 222.000 66.680 224.900 ;
        RECT 67.130 222.000 67.280 229.550 ;
        RECT 67.730 222.000 67.880 229.550 ;
        RECT 68.330 222.000 68.480 229.550 ;
        RECT 68.930 222.000 69.080 229.550 ;
        RECT 69.530 222.000 69.680 229.550 ;
        RECT 70.130 229.350 74.080 229.550 ;
        RECT 75.380 229.350 79.330 229.550 ;
        RECT 70.130 228.900 70.730 229.350 ;
        RECT 78.730 228.900 79.330 229.350 ;
        RECT 70.130 228.750 74.080 228.900 ;
        RECT 75.380 228.750 79.330 228.900 ;
        RECT 70.130 228.300 70.730 228.750 ;
        RECT 78.730 228.300 79.330 228.750 ;
        RECT 70.130 228.150 74.080 228.300 ;
        RECT 75.380 228.150 79.330 228.300 ;
        RECT 70.130 227.700 70.730 228.150 ;
        RECT 78.730 227.700 79.330 228.150 ;
        RECT 70.130 227.550 74.080 227.700 ;
        RECT 75.380 227.550 79.330 227.700 ;
        RECT 70.130 227.100 70.730 227.550 ;
        RECT 78.730 227.100 79.330 227.550 ;
        RECT 70.130 226.950 74.080 227.100 ;
        RECT 75.380 226.950 79.330 227.100 ;
        RECT 70.130 226.500 70.730 226.950 ;
        RECT 78.730 226.500 79.330 226.950 ;
        RECT 70.130 226.350 74.080 226.500 ;
        RECT 75.380 226.350 79.330 226.500 ;
        RECT 70.130 225.900 70.730 226.350 ;
        RECT 78.730 225.900 79.330 226.350 ;
        RECT 70.130 225.750 74.080 225.900 ;
        RECT 75.380 225.750 79.330 225.900 ;
        RECT 70.130 225.300 70.730 225.750 ;
        RECT 78.730 225.300 79.330 225.750 ;
        RECT 70.130 225.150 74.080 225.300 ;
        RECT 75.380 225.150 79.330 225.300 ;
        RECT 70.130 224.700 70.730 225.150 ;
        RECT 78.730 224.700 79.330 225.150 ;
        RECT 70.130 224.550 74.080 224.700 ;
        RECT 75.380 224.550 79.330 224.700 ;
        RECT 70.130 224.100 70.730 224.550 ;
        RECT 78.730 224.100 79.330 224.550 ;
        RECT 70.130 223.950 74.080 224.100 ;
        RECT 75.380 223.950 79.330 224.100 ;
        RECT 70.130 223.500 70.730 223.950 ;
        RECT 78.730 223.500 79.330 223.950 ;
        RECT 70.130 223.350 74.080 223.500 ;
        RECT 75.380 223.350 79.330 223.500 ;
        RECT 70.130 222.900 70.730 223.350 ;
        RECT 78.730 222.900 79.330 223.350 ;
        RECT 70.130 222.750 74.080 222.900 ;
        RECT 75.380 222.750 79.330 222.900 ;
        RECT 70.130 222.300 70.730 222.750 ;
        RECT 78.730 222.300 79.330 222.750 ;
        RECT 70.130 222.150 74.080 222.300 ;
        RECT 75.380 222.150 79.330 222.300 ;
        RECT 70.130 222.000 70.730 222.150 ;
        RECT 66.530 221.700 70.730 222.000 ;
        RECT 78.730 222.000 79.330 222.150 ;
        RECT 79.780 222.000 79.930 229.550 ;
        RECT 80.380 222.000 80.530 229.550 ;
        RECT 80.980 222.000 81.130 229.550 ;
        RECT 81.580 222.000 81.730 229.550 ;
        RECT 82.180 222.000 82.330 229.550 ;
        RECT 82.780 222.000 82.930 224.900 ;
        RECT 78.730 221.700 82.930 222.000 ;
        RECT 66.530 221.550 74.080 221.700 ;
        RECT 75.380 221.550 82.930 221.700 ;
        RECT 66.530 221.350 70.730 221.550 ;
        RECT 60.330 221.050 69.130 221.200 ;
        RECT 69.280 221.050 70.730 221.350 ;
        RECT 58.730 220.150 70.730 221.050 ;
        RECT 78.730 221.350 82.930 221.550 ;
        RECT 78.730 221.050 80.180 221.350 ;
        RECT 83.530 221.200 85.930 224.400 ;
        RECT 86.530 222.000 86.680 224.900 ;
        RECT 87.130 222.000 87.280 229.550 ;
        RECT 87.730 222.000 87.880 229.550 ;
        RECT 88.330 222.000 88.480 229.550 ;
        RECT 88.930 222.000 89.080 229.550 ;
        RECT 89.530 222.000 89.680 229.550 ;
        RECT 90.130 229.350 94.080 229.550 ;
        RECT 95.380 229.350 99.330 229.550 ;
        RECT 90.130 228.900 90.730 229.350 ;
        RECT 98.730 228.900 99.330 229.350 ;
        RECT 90.130 228.750 94.080 228.900 ;
        RECT 95.380 228.750 99.330 228.900 ;
        RECT 90.130 228.300 90.730 228.750 ;
        RECT 98.730 228.300 99.330 228.750 ;
        RECT 90.130 228.150 94.080 228.300 ;
        RECT 95.380 228.150 99.330 228.300 ;
        RECT 90.130 227.700 90.730 228.150 ;
        RECT 98.730 227.700 99.330 228.150 ;
        RECT 90.130 227.550 94.080 227.700 ;
        RECT 95.380 227.550 99.330 227.700 ;
        RECT 90.130 227.100 90.730 227.550 ;
        RECT 98.730 227.100 99.330 227.550 ;
        RECT 90.130 226.950 94.080 227.100 ;
        RECT 95.380 226.950 99.330 227.100 ;
        RECT 90.130 226.500 90.730 226.950 ;
        RECT 98.730 226.500 99.330 226.950 ;
        RECT 90.130 226.350 94.080 226.500 ;
        RECT 95.380 226.350 99.330 226.500 ;
        RECT 90.130 225.900 90.730 226.350 ;
        RECT 98.730 225.900 99.330 226.350 ;
        RECT 90.130 225.750 94.080 225.900 ;
        RECT 95.380 225.750 99.330 225.900 ;
        RECT 90.130 225.300 90.730 225.750 ;
        RECT 98.730 225.300 99.330 225.750 ;
        RECT 90.130 225.150 94.080 225.300 ;
        RECT 95.380 225.150 99.330 225.300 ;
        RECT 90.130 224.700 90.730 225.150 ;
        RECT 98.730 224.700 99.330 225.150 ;
        RECT 90.130 224.550 94.080 224.700 ;
        RECT 95.380 224.550 99.330 224.700 ;
        RECT 90.130 224.100 90.730 224.550 ;
        RECT 98.730 224.100 99.330 224.550 ;
        RECT 90.130 223.950 94.080 224.100 ;
        RECT 95.380 223.950 99.330 224.100 ;
        RECT 90.130 223.500 90.730 223.950 ;
        RECT 98.730 223.500 99.330 223.950 ;
        RECT 90.130 223.350 94.080 223.500 ;
        RECT 95.380 223.350 99.330 223.500 ;
        RECT 90.130 222.900 90.730 223.350 ;
        RECT 98.730 222.900 99.330 223.350 ;
        RECT 90.130 222.750 94.080 222.900 ;
        RECT 95.380 222.750 99.330 222.900 ;
        RECT 90.130 222.300 90.730 222.750 ;
        RECT 98.730 222.300 99.330 222.750 ;
        RECT 90.130 222.150 94.080 222.300 ;
        RECT 95.380 222.150 99.330 222.300 ;
        RECT 90.130 222.000 90.730 222.150 ;
        RECT 86.530 221.700 90.730 222.000 ;
        RECT 98.730 222.000 99.330 222.150 ;
        RECT 99.780 222.000 99.930 229.550 ;
        RECT 100.380 222.000 100.530 229.550 ;
        RECT 100.980 222.000 101.130 229.550 ;
        RECT 101.580 222.000 101.730 229.550 ;
        RECT 102.180 222.000 102.330 229.550 ;
        RECT 102.780 222.000 102.930 224.900 ;
        RECT 98.730 221.700 102.930 222.000 ;
        RECT 86.530 221.550 94.080 221.700 ;
        RECT 95.380 221.550 102.930 221.700 ;
        RECT 86.530 221.350 90.730 221.550 ;
        RECT 80.330 221.050 89.130 221.200 ;
        RECT 89.280 221.050 90.730 221.350 ;
        RECT 78.730 220.150 90.730 221.050 ;
        RECT 98.730 221.350 102.930 221.550 ;
        RECT 98.730 221.050 100.180 221.350 ;
        RECT 103.530 221.200 105.930 224.400 ;
        RECT 106.530 222.000 106.680 224.900 ;
        RECT 107.130 222.000 107.280 229.550 ;
        RECT 107.730 222.000 107.880 229.550 ;
        RECT 108.330 222.000 108.480 229.550 ;
        RECT 108.930 222.000 109.080 229.550 ;
        RECT 109.530 222.000 109.680 229.550 ;
        RECT 110.130 229.350 114.080 229.550 ;
        RECT 115.380 229.350 119.330 229.550 ;
        RECT 110.130 228.900 110.730 229.350 ;
        RECT 118.730 228.900 119.330 229.350 ;
        RECT 110.130 228.750 114.080 228.900 ;
        RECT 115.380 228.750 119.330 228.900 ;
        RECT 110.130 228.300 110.730 228.750 ;
        RECT 118.730 228.300 119.330 228.750 ;
        RECT 110.130 228.150 114.080 228.300 ;
        RECT 115.380 228.150 119.330 228.300 ;
        RECT 110.130 227.700 110.730 228.150 ;
        RECT 118.730 227.700 119.330 228.150 ;
        RECT 110.130 227.550 114.080 227.700 ;
        RECT 115.380 227.550 119.330 227.700 ;
        RECT 110.130 227.100 110.730 227.550 ;
        RECT 118.730 227.100 119.330 227.550 ;
        RECT 110.130 226.950 114.080 227.100 ;
        RECT 115.380 226.950 119.330 227.100 ;
        RECT 110.130 226.500 110.730 226.950 ;
        RECT 118.730 226.500 119.330 226.950 ;
        RECT 110.130 226.350 114.080 226.500 ;
        RECT 115.380 226.350 119.330 226.500 ;
        RECT 110.130 225.900 110.730 226.350 ;
        RECT 118.730 225.900 119.330 226.350 ;
        RECT 110.130 225.750 114.080 225.900 ;
        RECT 115.380 225.750 119.330 225.900 ;
        RECT 110.130 225.300 110.730 225.750 ;
        RECT 118.730 225.300 119.330 225.750 ;
        RECT 110.130 225.150 114.080 225.300 ;
        RECT 115.380 225.150 119.330 225.300 ;
        RECT 110.130 224.700 110.730 225.150 ;
        RECT 118.730 224.700 119.330 225.150 ;
        RECT 110.130 224.550 114.080 224.700 ;
        RECT 115.380 224.550 119.330 224.700 ;
        RECT 110.130 224.100 110.730 224.550 ;
        RECT 118.730 224.100 119.330 224.550 ;
        RECT 110.130 223.950 114.080 224.100 ;
        RECT 115.380 223.950 119.330 224.100 ;
        RECT 110.130 223.500 110.730 223.950 ;
        RECT 118.730 223.500 119.330 223.950 ;
        RECT 110.130 223.350 114.080 223.500 ;
        RECT 115.380 223.350 119.330 223.500 ;
        RECT 110.130 222.900 110.730 223.350 ;
        RECT 118.730 222.900 119.330 223.350 ;
        RECT 110.130 222.750 114.080 222.900 ;
        RECT 115.380 222.750 119.330 222.900 ;
        RECT 110.130 222.300 110.730 222.750 ;
        RECT 118.730 222.300 119.330 222.750 ;
        RECT 110.130 222.150 114.080 222.300 ;
        RECT 115.380 222.150 119.330 222.300 ;
        RECT 110.130 222.000 110.730 222.150 ;
        RECT 106.530 221.700 110.730 222.000 ;
        RECT 118.730 222.000 119.330 222.150 ;
        RECT 119.780 222.000 119.930 229.550 ;
        RECT 120.380 222.000 120.530 229.550 ;
        RECT 120.980 222.000 121.130 229.550 ;
        RECT 121.580 222.000 121.730 229.550 ;
        RECT 122.180 222.000 122.330 229.550 ;
        RECT 122.780 222.000 122.930 224.900 ;
        RECT 118.730 221.700 122.930 222.000 ;
        RECT 106.530 221.550 114.080 221.700 ;
        RECT 115.380 221.550 122.930 221.700 ;
        RECT 106.530 221.350 110.730 221.550 ;
        RECT 100.330 221.050 109.130 221.200 ;
        RECT 109.280 221.050 110.730 221.350 ;
        RECT 98.730 220.150 110.730 221.050 ;
        RECT 118.730 221.350 122.930 221.550 ;
        RECT 123.530 223.530 124.730 224.400 ;
        RECT 123.530 222.255 127.140 223.530 ;
        RECT 118.730 221.050 120.180 221.350 ;
        RECT 123.530 221.200 124.730 222.255 ;
        RECT 120.330 221.050 124.730 221.200 ;
        RECT 118.730 220.150 124.730 221.050 ;
        RECT 4.730 219.850 9.130 220.150 ;
        RECT 20.330 219.850 29.130 220.150 ;
        RECT 40.330 219.850 49.130 220.150 ;
        RECT 60.330 219.850 69.130 220.150 ;
        RECT 80.330 219.850 89.130 220.150 ;
        RECT 100.330 219.850 109.130 220.150 ;
        RECT 4.730 218.950 10.730 219.850 ;
        RECT 20.330 219.800 30.730 219.850 ;
        RECT 40.330 219.800 50.730 219.850 ;
        RECT 60.330 219.800 70.730 219.850 ;
        RECT 80.330 219.800 90.730 219.850 ;
        RECT 100.330 219.800 110.730 219.850 ;
        RECT 120.330 219.800 124.730 220.150 ;
        RECT 4.730 218.800 9.130 218.950 ;
        RECT 4.730 217.970 5.930 218.800 ;
        RECT 9.280 218.650 10.730 218.950 ;
        RECT 2.315 216.695 5.930 217.970 ;
        RECT 4.730 215.600 5.930 216.695 ;
        RECT 6.530 218.450 10.730 218.650 ;
        RECT 18.730 218.950 30.730 219.800 ;
        RECT 18.730 218.900 29.130 218.950 ;
        RECT 18.730 218.650 20.180 218.900 ;
        RECT 20.330 218.800 29.130 218.900 ;
        RECT 18.730 218.450 22.930 218.650 ;
        RECT 6.530 218.300 14.080 218.450 ;
        RECT 15.430 218.300 22.930 218.450 ;
        RECT 6.530 218.000 10.730 218.300 ;
        RECT 2.315 213.250 4.315 215.545 ;
        RECT 6.530 215.150 6.680 218.000 ;
        RECT 7.130 210.450 7.280 218.000 ;
        RECT 7.730 210.450 7.880 218.000 ;
        RECT 8.330 210.450 8.480 218.000 ;
        RECT 8.930 210.450 9.080 218.000 ;
        RECT 9.530 210.450 9.680 218.000 ;
        RECT 10.130 217.850 10.730 218.000 ;
        RECT 18.730 218.000 22.930 218.300 ;
        RECT 18.730 217.850 19.330 218.000 ;
        RECT 10.130 217.700 14.080 217.850 ;
        RECT 15.380 217.700 19.330 217.850 ;
        RECT 10.130 217.250 10.730 217.700 ;
        RECT 18.730 217.250 19.330 217.700 ;
        RECT 10.130 217.100 14.080 217.250 ;
        RECT 15.380 217.100 19.330 217.250 ;
        RECT 10.130 216.650 10.730 217.100 ;
        RECT 18.730 216.650 19.330 217.100 ;
        RECT 10.130 216.500 14.080 216.650 ;
        RECT 15.380 216.500 19.330 216.650 ;
        RECT 10.130 216.050 10.730 216.500 ;
        RECT 18.730 216.050 19.330 216.500 ;
        RECT 10.130 215.900 14.080 216.050 ;
        RECT 15.380 215.900 19.330 216.050 ;
        RECT 10.130 215.450 10.730 215.900 ;
        RECT 18.730 215.450 19.330 215.900 ;
        RECT 10.130 215.300 14.080 215.450 ;
        RECT 15.380 215.300 19.330 215.450 ;
        RECT 10.130 214.850 10.730 215.300 ;
        RECT 18.730 214.850 19.330 215.300 ;
        RECT 10.130 214.700 14.080 214.850 ;
        RECT 15.380 214.700 19.330 214.850 ;
        RECT 10.130 214.250 10.730 214.700 ;
        RECT 18.730 214.250 19.330 214.700 ;
        RECT 10.130 214.100 14.080 214.250 ;
        RECT 15.380 214.100 19.330 214.250 ;
        RECT 10.130 213.650 10.730 214.100 ;
        RECT 18.730 213.650 19.330 214.100 ;
        RECT 10.130 213.500 14.080 213.650 ;
        RECT 15.380 213.500 19.330 213.650 ;
        RECT 10.130 213.050 10.730 213.500 ;
        RECT 18.730 213.050 19.330 213.500 ;
        RECT 10.130 212.900 14.080 213.050 ;
        RECT 15.380 212.900 19.330 213.050 ;
        RECT 10.130 212.450 10.730 212.900 ;
        RECT 18.730 212.450 19.330 212.900 ;
        RECT 10.130 212.300 14.080 212.450 ;
        RECT 15.380 212.300 19.330 212.450 ;
        RECT 10.130 211.850 10.730 212.300 ;
        RECT 18.730 211.850 19.330 212.300 ;
        RECT 10.130 211.700 14.080 211.850 ;
        RECT 15.380 211.700 19.330 211.850 ;
        RECT 10.130 211.250 10.730 211.700 ;
        RECT 18.730 211.250 19.330 211.700 ;
        RECT 10.130 211.100 14.080 211.250 ;
        RECT 15.380 211.100 19.330 211.250 ;
        RECT 10.130 210.650 10.730 211.100 ;
        RECT 18.730 210.650 19.330 211.100 ;
        RECT 10.130 210.450 14.080 210.650 ;
        RECT 15.380 210.450 19.330 210.650 ;
        RECT 19.780 210.450 19.930 218.000 ;
        RECT 20.380 210.450 20.530 218.000 ;
        RECT 20.980 210.450 21.130 218.000 ;
        RECT 21.580 210.450 21.730 218.000 ;
        RECT 22.180 210.450 22.330 218.000 ;
        RECT 22.780 215.150 22.930 218.000 ;
        RECT 23.530 215.600 25.930 218.800 ;
        RECT 29.280 218.650 30.730 218.950 ;
        RECT 26.530 218.450 30.730 218.650 ;
        RECT 38.730 218.950 50.730 219.800 ;
        RECT 38.730 218.900 49.130 218.950 ;
        RECT 38.730 218.650 40.180 218.900 ;
        RECT 40.330 218.800 49.130 218.900 ;
        RECT 38.730 218.450 42.930 218.650 ;
        RECT 26.530 218.300 34.080 218.450 ;
        RECT 35.430 218.300 42.930 218.450 ;
        RECT 26.530 218.000 30.730 218.300 ;
        RECT 26.530 215.150 26.680 218.000 ;
        RECT 27.130 210.450 27.280 218.000 ;
        RECT 27.730 210.450 27.880 218.000 ;
        RECT 28.330 210.450 28.480 218.000 ;
        RECT 28.930 210.450 29.080 218.000 ;
        RECT 29.530 210.450 29.680 218.000 ;
        RECT 30.130 217.850 30.730 218.000 ;
        RECT 38.730 218.000 42.930 218.300 ;
        RECT 38.730 217.850 39.330 218.000 ;
        RECT 30.130 217.700 34.080 217.850 ;
        RECT 35.380 217.700 39.330 217.850 ;
        RECT 30.130 217.250 30.730 217.700 ;
        RECT 38.730 217.250 39.330 217.700 ;
        RECT 30.130 217.100 34.080 217.250 ;
        RECT 35.380 217.100 39.330 217.250 ;
        RECT 30.130 216.650 30.730 217.100 ;
        RECT 38.730 216.650 39.330 217.100 ;
        RECT 30.130 216.500 34.080 216.650 ;
        RECT 35.380 216.500 39.330 216.650 ;
        RECT 30.130 216.050 30.730 216.500 ;
        RECT 38.730 216.050 39.330 216.500 ;
        RECT 30.130 215.900 34.080 216.050 ;
        RECT 35.380 215.900 39.330 216.050 ;
        RECT 30.130 215.450 30.730 215.900 ;
        RECT 38.730 215.450 39.330 215.900 ;
        RECT 30.130 215.300 34.080 215.450 ;
        RECT 35.380 215.300 39.330 215.450 ;
        RECT 30.130 214.850 30.730 215.300 ;
        RECT 38.730 214.850 39.330 215.300 ;
        RECT 30.130 214.700 34.080 214.850 ;
        RECT 35.380 214.700 39.330 214.850 ;
        RECT 30.130 214.250 30.730 214.700 ;
        RECT 38.730 214.250 39.330 214.700 ;
        RECT 30.130 214.100 34.080 214.250 ;
        RECT 35.380 214.100 39.330 214.250 ;
        RECT 30.130 213.650 30.730 214.100 ;
        RECT 38.730 213.650 39.330 214.100 ;
        RECT 30.130 213.500 34.080 213.650 ;
        RECT 35.380 213.500 39.330 213.650 ;
        RECT 30.130 213.050 30.730 213.500 ;
        RECT 38.730 213.050 39.330 213.500 ;
        RECT 30.130 212.900 34.080 213.050 ;
        RECT 35.380 212.900 39.330 213.050 ;
        RECT 30.130 212.450 30.730 212.900 ;
        RECT 38.730 212.450 39.330 212.900 ;
        RECT 30.130 212.300 34.080 212.450 ;
        RECT 35.380 212.300 39.330 212.450 ;
        RECT 30.130 211.850 30.730 212.300 ;
        RECT 38.730 211.850 39.330 212.300 ;
        RECT 30.130 211.700 34.080 211.850 ;
        RECT 35.380 211.700 39.330 211.850 ;
        RECT 30.130 211.250 30.730 211.700 ;
        RECT 38.730 211.250 39.330 211.700 ;
        RECT 30.130 211.100 34.080 211.250 ;
        RECT 35.380 211.100 39.330 211.250 ;
        RECT 30.130 210.650 30.730 211.100 ;
        RECT 38.730 210.650 39.330 211.100 ;
        RECT 30.130 210.450 34.080 210.650 ;
        RECT 35.380 210.450 39.330 210.650 ;
        RECT 39.780 210.450 39.930 218.000 ;
        RECT 40.380 210.450 40.530 218.000 ;
        RECT 40.980 210.450 41.130 218.000 ;
        RECT 41.580 210.450 41.730 218.000 ;
        RECT 42.180 210.450 42.330 218.000 ;
        RECT 42.780 215.150 42.930 218.000 ;
        RECT 43.530 215.600 45.930 218.800 ;
        RECT 49.280 218.650 50.730 218.950 ;
        RECT 46.530 218.450 50.730 218.650 ;
        RECT 58.730 218.950 70.730 219.800 ;
        RECT 58.730 218.900 69.130 218.950 ;
        RECT 58.730 218.650 60.180 218.900 ;
        RECT 60.330 218.800 69.130 218.900 ;
        RECT 58.730 218.450 62.930 218.650 ;
        RECT 46.530 218.300 54.080 218.450 ;
        RECT 55.430 218.300 62.930 218.450 ;
        RECT 46.530 218.000 50.730 218.300 ;
        RECT 46.530 215.150 46.680 218.000 ;
        RECT 47.130 210.450 47.280 218.000 ;
        RECT 47.730 210.450 47.880 218.000 ;
        RECT 48.330 210.450 48.480 218.000 ;
        RECT 48.930 210.450 49.080 218.000 ;
        RECT 49.530 210.450 49.680 218.000 ;
        RECT 50.130 217.850 50.730 218.000 ;
        RECT 58.730 218.000 62.930 218.300 ;
        RECT 58.730 217.850 59.330 218.000 ;
        RECT 50.130 217.700 54.080 217.850 ;
        RECT 55.380 217.700 59.330 217.850 ;
        RECT 50.130 217.250 50.730 217.700 ;
        RECT 58.730 217.250 59.330 217.700 ;
        RECT 50.130 217.100 54.080 217.250 ;
        RECT 55.380 217.100 59.330 217.250 ;
        RECT 50.130 216.650 50.730 217.100 ;
        RECT 58.730 216.650 59.330 217.100 ;
        RECT 50.130 216.500 54.080 216.650 ;
        RECT 55.380 216.500 59.330 216.650 ;
        RECT 50.130 216.050 50.730 216.500 ;
        RECT 58.730 216.050 59.330 216.500 ;
        RECT 50.130 215.900 54.080 216.050 ;
        RECT 55.380 215.900 59.330 216.050 ;
        RECT 50.130 215.450 50.730 215.900 ;
        RECT 58.730 215.450 59.330 215.900 ;
        RECT 50.130 215.300 54.080 215.450 ;
        RECT 55.380 215.300 59.330 215.450 ;
        RECT 50.130 214.850 50.730 215.300 ;
        RECT 58.730 214.850 59.330 215.300 ;
        RECT 50.130 214.700 54.080 214.850 ;
        RECT 55.380 214.700 59.330 214.850 ;
        RECT 50.130 214.250 50.730 214.700 ;
        RECT 58.730 214.250 59.330 214.700 ;
        RECT 50.130 214.100 54.080 214.250 ;
        RECT 55.380 214.100 59.330 214.250 ;
        RECT 50.130 213.650 50.730 214.100 ;
        RECT 58.730 213.650 59.330 214.100 ;
        RECT 50.130 213.500 54.080 213.650 ;
        RECT 55.380 213.500 59.330 213.650 ;
        RECT 50.130 213.050 50.730 213.500 ;
        RECT 58.730 213.050 59.330 213.500 ;
        RECT 50.130 212.900 54.080 213.050 ;
        RECT 55.380 212.900 59.330 213.050 ;
        RECT 50.130 212.450 50.730 212.900 ;
        RECT 58.730 212.450 59.330 212.900 ;
        RECT 50.130 212.300 54.080 212.450 ;
        RECT 55.380 212.300 59.330 212.450 ;
        RECT 50.130 211.850 50.730 212.300 ;
        RECT 58.730 211.850 59.330 212.300 ;
        RECT 50.130 211.700 54.080 211.850 ;
        RECT 55.380 211.700 59.330 211.850 ;
        RECT 50.130 211.250 50.730 211.700 ;
        RECT 58.730 211.250 59.330 211.700 ;
        RECT 50.130 211.100 54.080 211.250 ;
        RECT 55.380 211.100 59.330 211.250 ;
        RECT 50.130 210.650 50.730 211.100 ;
        RECT 58.730 210.650 59.330 211.100 ;
        RECT 50.130 210.450 54.080 210.650 ;
        RECT 55.380 210.450 59.330 210.650 ;
        RECT 59.780 210.450 59.930 218.000 ;
        RECT 60.380 210.450 60.530 218.000 ;
        RECT 60.980 210.450 61.130 218.000 ;
        RECT 61.580 210.450 61.730 218.000 ;
        RECT 62.180 210.450 62.330 218.000 ;
        RECT 62.780 215.150 62.930 218.000 ;
        RECT 63.530 215.600 65.930 218.800 ;
        RECT 69.280 218.650 70.730 218.950 ;
        RECT 66.530 218.450 70.730 218.650 ;
        RECT 78.730 218.950 90.730 219.800 ;
        RECT 78.730 218.900 89.130 218.950 ;
        RECT 78.730 218.650 80.180 218.900 ;
        RECT 80.330 218.800 89.130 218.900 ;
        RECT 78.730 218.450 82.930 218.650 ;
        RECT 66.530 218.300 74.080 218.450 ;
        RECT 75.430 218.300 82.930 218.450 ;
        RECT 66.530 218.000 70.730 218.300 ;
        RECT 66.530 215.150 66.680 218.000 ;
        RECT 67.130 210.450 67.280 218.000 ;
        RECT 67.730 210.450 67.880 218.000 ;
        RECT 68.330 210.450 68.480 218.000 ;
        RECT 68.930 210.450 69.080 218.000 ;
        RECT 69.530 210.450 69.680 218.000 ;
        RECT 70.130 217.850 70.730 218.000 ;
        RECT 78.730 218.000 82.930 218.300 ;
        RECT 78.730 217.850 79.330 218.000 ;
        RECT 70.130 217.700 74.080 217.850 ;
        RECT 75.380 217.700 79.330 217.850 ;
        RECT 70.130 217.250 70.730 217.700 ;
        RECT 78.730 217.250 79.330 217.700 ;
        RECT 70.130 217.100 74.080 217.250 ;
        RECT 75.380 217.100 79.330 217.250 ;
        RECT 70.130 216.650 70.730 217.100 ;
        RECT 78.730 216.650 79.330 217.100 ;
        RECT 70.130 216.500 74.080 216.650 ;
        RECT 75.380 216.500 79.330 216.650 ;
        RECT 70.130 216.050 70.730 216.500 ;
        RECT 78.730 216.050 79.330 216.500 ;
        RECT 70.130 215.900 74.080 216.050 ;
        RECT 75.380 215.900 79.330 216.050 ;
        RECT 70.130 215.450 70.730 215.900 ;
        RECT 78.730 215.450 79.330 215.900 ;
        RECT 70.130 215.300 74.080 215.450 ;
        RECT 75.380 215.300 79.330 215.450 ;
        RECT 70.130 214.850 70.730 215.300 ;
        RECT 78.730 214.850 79.330 215.300 ;
        RECT 70.130 214.700 74.080 214.850 ;
        RECT 75.380 214.700 79.330 214.850 ;
        RECT 70.130 214.250 70.730 214.700 ;
        RECT 78.730 214.250 79.330 214.700 ;
        RECT 70.130 214.100 74.080 214.250 ;
        RECT 75.380 214.100 79.330 214.250 ;
        RECT 70.130 213.650 70.730 214.100 ;
        RECT 78.730 213.650 79.330 214.100 ;
        RECT 70.130 213.500 74.080 213.650 ;
        RECT 75.380 213.500 79.330 213.650 ;
        RECT 70.130 213.050 70.730 213.500 ;
        RECT 78.730 213.050 79.330 213.500 ;
        RECT 70.130 212.900 74.080 213.050 ;
        RECT 75.380 212.900 79.330 213.050 ;
        RECT 70.130 212.450 70.730 212.900 ;
        RECT 78.730 212.450 79.330 212.900 ;
        RECT 70.130 212.300 74.080 212.450 ;
        RECT 75.380 212.300 79.330 212.450 ;
        RECT 70.130 211.850 70.730 212.300 ;
        RECT 78.730 211.850 79.330 212.300 ;
        RECT 70.130 211.700 74.080 211.850 ;
        RECT 75.380 211.700 79.330 211.850 ;
        RECT 70.130 211.250 70.730 211.700 ;
        RECT 78.730 211.250 79.330 211.700 ;
        RECT 70.130 211.100 74.080 211.250 ;
        RECT 75.380 211.100 79.330 211.250 ;
        RECT 70.130 210.650 70.730 211.100 ;
        RECT 78.730 210.650 79.330 211.100 ;
        RECT 70.130 210.450 74.080 210.650 ;
        RECT 75.380 210.450 79.330 210.650 ;
        RECT 79.780 210.450 79.930 218.000 ;
        RECT 80.380 210.450 80.530 218.000 ;
        RECT 80.980 210.450 81.130 218.000 ;
        RECT 81.580 210.450 81.730 218.000 ;
        RECT 82.180 210.450 82.330 218.000 ;
        RECT 82.780 215.150 82.930 218.000 ;
        RECT 83.530 215.600 85.930 218.800 ;
        RECT 89.280 218.650 90.730 218.950 ;
        RECT 86.530 218.450 90.730 218.650 ;
        RECT 98.730 218.950 110.730 219.800 ;
        RECT 98.730 218.900 109.130 218.950 ;
        RECT 98.730 218.650 100.180 218.900 ;
        RECT 100.330 218.800 109.130 218.900 ;
        RECT 98.730 218.450 102.930 218.650 ;
        RECT 86.530 218.300 94.080 218.450 ;
        RECT 95.430 218.300 102.930 218.450 ;
        RECT 86.530 218.000 90.730 218.300 ;
        RECT 86.530 215.150 86.680 218.000 ;
        RECT 87.130 210.450 87.280 218.000 ;
        RECT 87.730 210.450 87.880 218.000 ;
        RECT 88.330 210.450 88.480 218.000 ;
        RECT 88.930 210.450 89.080 218.000 ;
        RECT 89.530 210.450 89.680 218.000 ;
        RECT 90.130 217.850 90.730 218.000 ;
        RECT 98.730 218.000 102.930 218.300 ;
        RECT 98.730 217.850 99.330 218.000 ;
        RECT 90.130 217.700 94.080 217.850 ;
        RECT 95.380 217.700 99.330 217.850 ;
        RECT 90.130 217.250 90.730 217.700 ;
        RECT 98.730 217.250 99.330 217.700 ;
        RECT 90.130 217.100 94.080 217.250 ;
        RECT 95.380 217.100 99.330 217.250 ;
        RECT 90.130 216.650 90.730 217.100 ;
        RECT 98.730 216.650 99.330 217.100 ;
        RECT 90.130 216.500 94.080 216.650 ;
        RECT 95.380 216.500 99.330 216.650 ;
        RECT 90.130 216.050 90.730 216.500 ;
        RECT 98.730 216.050 99.330 216.500 ;
        RECT 90.130 215.900 94.080 216.050 ;
        RECT 95.380 215.900 99.330 216.050 ;
        RECT 90.130 215.450 90.730 215.900 ;
        RECT 98.730 215.450 99.330 215.900 ;
        RECT 90.130 215.300 94.080 215.450 ;
        RECT 95.380 215.300 99.330 215.450 ;
        RECT 90.130 214.850 90.730 215.300 ;
        RECT 98.730 214.850 99.330 215.300 ;
        RECT 90.130 214.700 94.080 214.850 ;
        RECT 95.380 214.700 99.330 214.850 ;
        RECT 90.130 214.250 90.730 214.700 ;
        RECT 98.730 214.250 99.330 214.700 ;
        RECT 90.130 214.100 94.080 214.250 ;
        RECT 95.380 214.100 99.330 214.250 ;
        RECT 90.130 213.650 90.730 214.100 ;
        RECT 98.730 213.650 99.330 214.100 ;
        RECT 90.130 213.500 94.080 213.650 ;
        RECT 95.380 213.500 99.330 213.650 ;
        RECT 90.130 213.050 90.730 213.500 ;
        RECT 98.730 213.050 99.330 213.500 ;
        RECT 90.130 212.900 94.080 213.050 ;
        RECT 95.380 212.900 99.330 213.050 ;
        RECT 90.130 212.450 90.730 212.900 ;
        RECT 98.730 212.450 99.330 212.900 ;
        RECT 90.130 212.300 94.080 212.450 ;
        RECT 95.380 212.300 99.330 212.450 ;
        RECT 90.130 211.850 90.730 212.300 ;
        RECT 98.730 211.850 99.330 212.300 ;
        RECT 90.130 211.700 94.080 211.850 ;
        RECT 95.380 211.700 99.330 211.850 ;
        RECT 90.130 211.250 90.730 211.700 ;
        RECT 98.730 211.250 99.330 211.700 ;
        RECT 90.130 211.100 94.080 211.250 ;
        RECT 95.380 211.100 99.330 211.250 ;
        RECT 90.130 210.650 90.730 211.100 ;
        RECT 98.730 210.650 99.330 211.100 ;
        RECT 90.130 210.450 94.080 210.650 ;
        RECT 95.380 210.450 99.330 210.650 ;
        RECT 99.780 210.450 99.930 218.000 ;
        RECT 100.380 210.450 100.530 218.000 ;
        RECT 100.980 210.450 101.130 218.000 ;
        RECT 101.580 210.450 101.730 218.000 ;
        RECT 102.180 210.450 102.330 218.000 ;
        RECT 102.780 215.150 102.930 218.000 ;
        RECT 103.530 215.600 105.930 218.800 ;
        RECT 109.280 218.650 110.730 218.950 ;
        RECT 106.530 218.450 110.730 218.650 ;
        RECT 118.730 218.900 124.730 219.800 ;
        RECT 118.730 218.650 120.180 218.900 ;
        RECT 120.330 218.800 124.730 218.900 ;
        RECT 118.730 218.450 122.930 218.650 ;
        RECT 106.530 218.300 114.080 218.450 ;
        RECT 115.430 218.300 122.930 218.450 ;
        RECT 106.530 218.000 110.730 218.300 ;
        RECT 106.530 215.150 106.680 218.000 ;
        RECT 107.130 210.450 107.280 218.000 ;
        RECT 107.730 210.450 107.880 218.000 ;
        RECT 108.330 210.450 108.480 218.000 ;
        RECT 108.930 210.450 109.080 218.000 ;
        RECT 109.530 210.450 109.680 218.000 ;
        RECT 110.130 217.850 110.730 218.000 ;
        RECT 118.730 218.000 122.930 218.300 ;
        RECT 118.730 217.850 119.330 218.000 ;
        RECT 110.130 217.700 114.080 217.850 ;
        RECT 115.380 217.700 119.330 217.850 ;
        RECT 110.130 217.250 110.730 217.700 ;
        RECT 118.730 217.250 119.330 217.700 ;
        RECT 110.130 217.100 114.080 217.250 ;
        RECT 115.380 217.100 119.330 217.250 ;
        RECT 110.130 216.650 110.730 217.100 ;
        RECT 118.730 216.650 119.330 217.100 ;
        RECT 110.130 216.500 114.080 216.650 ;
        RECT 115.380 216.500 119.330 216.650 ;
        RECT 110.130 216.050 110.730 216.500 ;
        RECT 118.730 216.050 119.330 216.500 ;
        RECT 110.130 215.900 114.080 216.050 ;
        RECT 115.380 215.900 119.330 216.050 ;
        RECT 110.130 215.450 110.730 215.900 ;
        RECT 118.730 215.450 119.330 215.900 ;
        RECT 110.130 215.300 114.080 215.450 ;
        RECT 115.380 215.300 119.330 215.450 ;
        RECT 110.130 214.850 110.730 215.300 ;
        RECT 118.730 214.850 119.330 215.300 ;
        RECT 110.130 214.700 114.080 214.850 ;
        RECT 115.380 214.700 119.330 214.850 ;
        RECT 110.130 214.250 110.730 214.700 ;
        RECT 118.730 214.250 119.330 214.700 ;
        RECT 110.130 214.100 114.080 214.250 ;
        RECT 115.380 214.100 119.330 214.250 ;
        RECT 110.130 213.650 110.730 214.100 ;
        RECT 118.730 213.650 119.330 214.100 ;
        RECT 110.130 213.500 114.080 213.650 ;
        RECT 115.380 213.500 119.330 213.650 ;
        RECT 110.130 213.050 110.730 213.500 ;
        RECT 118.730 213.050 119.330 213.500 ;
        RECT 110.130 212.900 114.080 213.050 ;
        RECT 115.380 212.900 119.330 213.050 ;
        RECT 110.130 212.450 110.730 212.900 ;
        RECT 118.730 212.450 119.330 212.900 ;
        RECT 110.130 212.300 114.080 212.450 ;
        RECT 115.380 212.300 119.330 212.450 ;
        RECT 110.130 211.850 110.730 212.300 ;
        RECT 118.730 211.850 119.330 212.300 ;
        RECT 110.130 211.700 114.080 211.850 ;
        RECT 115.380 211.700 119.330 211.850 ;
        RECT 110.130 211.250 110.730 211.700 ;
        RECT 118.730 211.250 119.330 211.700 ;
        RECT 110.130 211.100 114.080 211.250 ;
        RECT 115.380 211.100 119.330 211.250 ;
        RECT 110.130 210.650 110.730 211.100 ;
        RECT 118.730 210.650 119.330 211.100 ;
        RECT 110.130 210.450 114.080 210.650 ;
        RECT 115.380 210.450 119.330 210.650 ;
        RECT 119.780 210.450 119.930 218.000 ;
        RECT 120.380 210.450 120.530 218.000 ;
        RECT 120.980 210.450 121.130 218.000 ;
        RECT 121.580 210.450 121.730 218.000 ;
        RECT 122.180 210.450 122.330 218.000 ;
        RECT 122.780 215.150 122.930 218.000 ;
        RECT 123.530 217.765 124.730 218.800 ;
        RECT 123.530 216.490 127.140 217.765 ;
        RECT 123.530 215.600 124.730 216.490 ;
        RECT 2.315 204.455 4.315 206.750 ;
        RECT 2.315 204.450 4.180 204.455 ;
        RECT 4.730 202.670 5.930 204.400 ;
        RECT 2.315 201.395 5.930 202.670 ;
        RECT 4.730 201.200 5.930 201.395 ;
        RECT 6.530 202.000 6.680 204.900 ;
        RECT 7.130 202.000 7.280 209.550 ;
        RECT 7.730 202.000 7.880 209.550 ;
        RECT 8.330 202.000 8.480 209.550 ;
        RECT 8.930 202.000 9.080 209.550 ;
        RECT 9.530 202.000 9.680 209.550 ;
        RECT 10.130 209.350 14.080 209.550 ;
        RECT 15.380 209.350 19.330 209.550 ;
        RECT 10.130 208.900 10.730 209.350 ;
        RECT 18.730 208.900 19.330 209.350 ;
        RECT 10.130 208.750 14.080 208.900 ;
        RECT 15.380 208.750 19.330 208.900 ;
        RECT 10.130 208.300 10.730 208.750 ;
        RECT 18.730 208.300 19.330 208.750 ;
        RECT 10.130 208.150 14.080 208.300 ;
        RECT 15.380 208.150 19.330 208.300 ;
        RECT 10.130 207.700 10.730 208.150 ;
        RECT 18.730 207.700 19.330 208.150 ;
        RECT 10.130 207.550 14.080 207.700 ;
        RECT 15.380 207.550 19.330 207.700 ;
        RECT 10.130 207.100 10.730 207.550 ;
        RECT 18.730 207.100 19.330 207.550 ;
        RECT 10.130 206.950 14.080 207.100 ;
        RECT 15.380 206.950 19.330 207.100 ;
        RECT 10.130 206.500 10.730 206.950 ;
        RECT 18.730 206.500 19.330 206.950 ;
        RECT 10.130 206.350 14.080 206.500 ;
        RECT 15.380 206.350 19.330 206.500 ;
        RECT 10.130 205.900 10.730 206.350 ;
        RECT 18.730 205.900 19.330 206.350 ;
        RECT 10.130 205.750 14.080 205.900 ;
        RECT 15.380 205.750 19.330 205.900 ;
        RECT 10.130 205.300 10.730 205.750 ;
        RECT 18.730 205.300 19.330 205.750 ;
        RECT 10.130 205.150 14.080 205.300 ;
        RECT 15.380 205.150 19.330 205.300 ;
        RECT 10.130 204.700 10.730 205.150 ;
        RECT 18.730 204.700 19.330 205.150 ;
        RECT 10.130 204.550 14.080 204.700 ;
        RECT 15.380 204.550 19.330 204.700 ;
        RECT 10.130 204.100 10.730 204.550 ;
        RECT 18.730 204.100 19.330 204.550 ;
        RECT 10.130 203.950 14.080 204.100 ;
        RECT 15.380 203.950 19.330 204.100 ;
        RECT 10.130 203.500 10.730 203.950 ;
        RECT 18.730 203.500 19.330 203.950 ;
        RECT 10.130 203.350 14.080 203.500 ;
        RECT 15.380 203.350 19.330 203.500 ;
        RECT 10.130 202.900 10.730 203.350 ;
        RECT 18.730 202.900 19.330 203.350 ;
        RECT 10.130 202.750 14.080 202.900 ;
        RECT 15.380 202.750 19.330 202.900 ;
        RECT 10.130 202.300 10.730 202.750 ;
        RECT 18.730 202.300 19.330 202.750 ;
        RECT 10.130 202.150 14.080 202.300 ;
        RECT 15.380 202.150 19.330 202.300 ;
        RECT 10.130 202.000 10.730 202.150 ;
        RECT 6.530 201.700 10.730 202.000 ;
        RECT 18.730 202.000 19.330 202.150 ;
        RECT 19.780 202.000 19.930 209.550 ;
        RECT 20.380 202.000 20.530 209.550 ;
        RECT 20.980 202.000 21.130 209.550 ;
        RECT 21.580 202.000 21.730 209.550 ;
        RECT 22.180 202.000 22.330 209.550 ;
        RECT 22.780 202.000 22.930 204.900 ;
        RECT 18.730 201.700 22.930 202.000 ;
        RECT 6.530 201.550 14.080 201.700 ;
        RECT 15.380 201.550 22.930 201.700 ;
        RECT 6.530 201.350 10.730 201.550 ;
        RECT 4.730 201.050 9.130 201.200 ;
        RECT 9.280 201.050 10.730 201.350 ;
        RECT 4.730 200.150 10.730 201.050 ;
        RECT 18.730 201.350 22.930 201.550 ;
        RECT 18.730 201.050 20.180 201.350 ;
        RECT 23.530 201.200 25.930 204.400 ;
        RECT 26.530 202.000 26.680 204.900 ;
        RECT 27.130 202.000 27.280 209.550 ;
        RECT 27.730 202.000 27.880 209.550 ;
        RECT 28.330 202.000 28.480 209.550 ;
        RECT 28.930 202.000 29.080 209.550 ;
        RECT 29.530 202.000 29.680 209.550 ;
        RECT 30.130 209.350 34.080 209.550 ;
        RECT 35.380 209.350 39.330 209.550 ;
        RECT 30.130 208.900 30.730 209.350 ;
        RECT 38.730 208.900 39.330 209.350 ;
        RECT 30.130 208.750 34.080 208.900 ;
        RECT 35.380 208.750 39.330 208.900 ;
        RECT 30.130 208.300 30.730 208.750 ;
        RECT 38.730 208.300 39.330 208.750 ;
        RECT 30.130 208.150 34.080 208.300 ;
        RECT 35.380 208.150 39.330 208.300 ;
        RECT 30.130 207.700 30.730 208.150 ;
        RECT 38.730 207.700 39.330 208.150 ;
        RECT 30.130 207.550 34.080 207.700 ;
        RECT 35.380 207.550 39.330 207.700 ;
        RECT 30.130 207.100 30.730 207.550 ;
        RECT 38.730 207.100 39.330 207.550 ;
        RECT 30.130 206.950 34.080 207.100 ;
        RECT 35.380 206.950 39.330 207.100 ;
        RECT 30.130 206.500 30.730 206.950 ;
        RECT 38.730 206.500 39.330 206.950 ;
        RECT 30.130 206.350 34.080 206.500 ;
        RECT 35.380 206.350 39.330 206.500 ;
        RECT 30.130 205.900 30.730 206.350 ;
        RECT 38.730 205.900 39.330 206.350 ;
        RECT 30.130 205.750 34.080 205.900 ;
        RECT 35.380 205.750 39.330 205.900 ;
        RECT 30.130 205.300 30.730 205.750 ;
        RECT 38.730 205.300 39.330 205.750 ;
        RECT 30.130 205.150 34.080 205.300 ;
        RECT 35.380 205.150 39.330 205.300 ;
        RECT 30.130 204.700 30.730 205.150 ;
        RECT 38.730 204.700 39.330 205.150 ;
        RECT 30.130 204.550 34.080 204.700 ;
        RECT 35.380 204.550 39.330 204.700 ;
        RECT 30.130 204.100 30.730 204.550 ;
        RECT 38.730 204.100 39.330 204.550 ;
        RECT 30.130 203.950 34.080 204.100 ;
        RECT 35.380 203.950 39.330 204.100 ;
        RECT 30.130 203.500 30.730 203.950 ;
        RECT 38.730 203.500 39.330 203.950 ;
        RECT 30.130 203.350 34.080 203.500 ;
        RECT 35.380 203.350 39.330 203.500 ;
        RECT 30.130 202.900 30.730 203.350 ;
        RECT 38.730 202.900 39.330 203.350 ;
        RECT 30.130 202.750 34.080 202.900 ;
        RECT 35.380 202.750 39.330 202.900 ;
        RECT 30.130 202.300 30.730 202.750 ;
        RECT 38.730 202.300 39.330 202.750 ;
        RECT 30.130 202.150 34.080 202.300 ;
        RECT 35.380 202.150 39.330 202.300 ;
        RECT 30.130 202.000 30.730 202.150 ;
        RECT 26.530 201.700 30.730 202.000 ;
        RECT 38.730 202.000 39.330 202.150 ;
        RECT 39.780 202.000 39.930 209.550 ;
        RECT 40.380 202.000 40.530 209.550 ;
        RECT 40.980 202.000 41.130 209.550 ;
        RECT 41.580 202.000 41.730 209.550 ;
        RECT 42.180 202.000 42.330 209.550 ;
        RECT 42.780 202.000 42.930 204.900 ;
        RECT 38.730 201.700 42.930 202.000 ;
        RECT 26.530 201.550 34.080 201.700 ;
        RECT 35.380 201.550 42.930 201.700 ;
        RECT 26.530 201.350 30.730 201.550 ;
        RECT 20.330 201.050 29.130 201.200 ;
        RECT 29.280 201.050 30.730 201.350 ;
        RECT 18.730 200.150 30.730 201.050 ;
        RECT 38.730 201.350 42.930 201.550 ;
        RECT 38.730 201.050 40.180 201.350 ;
        RECT 43.530 201.200 45.930 204.400 ;
        RECT 46.530 202.000 46.680 204.900 ;
        RECT 47.130 202.000 47.280 209.550 ;
        RECT 47.730 202.000 47.880 209.550 ;
        RECT 48.330 202.000 48.480 209.550 ;
        RECT 48.930 202.000 49.080 209.550 ;
        RECT 49.530 202.000 49.680 209.550 ;
        RECT 50.130 209.350 54.080 209.550 ;
        RECT 55.380 209.350 59.330 209.550 ;
        RECT 50.130 208.900 50.730 209.350 ;
        RECT 58.730 208.900 59.330 209.350 ;
        RECT 50.130 208.750 54.080 208.900 ;
        RECT 55.380 208.750 59.330 208.900 ;
        RECT 50.130 208.300 50.730 208.750 ;
        RECT 58.730 208.300 59.330 208.750 ;
        RECT 50.130 208.150 54.080 208.300 ;
        RECT 55.380 208.150 59.330 208.300 ;
        RECT 50.130 207.700 50.730 208.150 ;
        RECT 58.730 207.700 59.330 208.150 ;
        RECT 50.130 207.550 54.080 207.700 ;
        RECT 55.380 207.550 59.330 207.700 ;
        RECT 50.130 207.100 50.730 207.550 ;
        RECT 58.730 207.100 59.330 207.550 ;
        RECT 50.130 206.950 54.080 207.100 ;
        RECT 55.380 206.950 59.330 207.100 ;
        RECT 50.130 206.500 50.730 206.950 ;
        RECT 58.730 206.500 59.330 206.950 ;
        RECT 50.130 206.350 54.080 206.500 ;
        RECT 55.380 206.350 59.330 206.500 ;
        RECT 50.130 205.900 50.730 206.350 ;
        RECT 58.730 205.900 59.330 206.350 ;
        RECT 50.130 205.750 54.080 205.900 ;
        RECT 55.380 205.750 59.330 205.900 ;
        RECT 50.130 205.300 50.730 205.750 ;
        RECT 58.730 205.300 59.330 205.750 ;
        RECT 50.130 205.150 54.080 205.300 ;
        RECT 55.380 205.150 59.330 205.300 ;
        RECT 50.130 204.700 50.730 205.150 ;
        RECT 58.730 204.700 59.330 205.150 ;
        RECT 50.130 204.550 54.080 204.700 ;
        RECT 55.380 204.550 59.330 204.700 ;
        RECT 50.130 204.100 50.730 204.550 ;
        RECT 58.730 204.100 59.330 204.550 ;
        RECT 50.130 203.950 54.080 204.100 ;
        RECT 55.380 203.950 59.330 204.100 ;
        RECT 50.130 203.500 50.730 203.950 ;
        RECT 58.730 203.500 59.330 203.950 ;
        RECT 50.130 203.350 54.080 203.500 ;
        RECT 55.380 203.350 59.330 203.500 ;
        RECT 50.130 202.900 50.730 203.350 ;
        RECT 58.730 202.900 59.330 203.350 ;
        RECT 50.130 202.750 54.080 202.900 ;
        RECT 55.380 202.750 59.330 202.900 ;
        RECT 50.130 202.300 50.730 202.750 ;
        RECT 58.730 202.300 59.330 202.750 ;
        RECT 50.130 202.150 54.080 202.300 ;
        RECT 55.380 202.150 59.330 202.300 ;
        RECT 50.130 202.000 50.730 202.150 ;
        RECT 46.530 201.700 50.730 202.000 ;
        RECT 58.730 202.000 59.330 202.150 ;
        RECT 59.780 202.000 59.930 209.550 ;
        RECT 60.380 202.000 60.530 209.550 ;
        RECT 60.980 202.000 61.130 209.550 ;
        RECT 61.580 202.000 61.730 209.550 ;
        RECT 62.180 202.000 62.330 209.550 ;
        RECT 62.780 202.000 62.930 204.900 ;
        RECT 58.730 201.700 62.930 202.000 ;
        RECT 46.530 201.550 54.080 201.700 ;
        RECT 55.380 201.550 62.930 201.700 ;
        RECT 46.530 201.350 50.730 201.550 ;
        RECT 40.330 201.050 49.130 201.200 ;
        RECT 49.280 201.050 50.730 201.350 ;
        RECT 38.730 200.150 50.730 201.050 ;
        RECT 58.730 201.350 62.930 201.550 ;
        RECT 58.730 201.050 60.180 201.350 ;
        RECT 63.530 201.200 65.930 204.400 ;
        RECT 66.530 202.000 66.680 204.900 ;
        RECT 67.130 202.000 67.280 209.550 ;
        RECT 67.730 202.000 67.880 209.550 ;
        RECT 68.330 202.000 68.480 209.550 ;
        RECT 68.930 202.000 69.080 209.550 ;
        RECT 69.530 202.000 69.680 209.550 ;
        RECT 70.130 209.350 74.080 209.550 ;
        RECT 75.380 209.350 79.330 209.550 ;
        RECT 70.130 208.900 70.730 209.350 ;
        RECT 78.730 208.900 79.330 209.350 ;
        RECT 70.130 208.750 74.080 208.900 ;
        RECT 75.380 208.750 79.330 208.900 ;
        RECT 70.130 208.300 70.730 208.750 ;
        RECT 78.730 208.300 79.330 208.750 ;
        RECT 70.130 208.150 74.080 208.300 ;
        RECT 75.380 208.150 79.330 208.300 ;
        RECT 70.130 207.700 70.730 208.150 ;
        RECT 78.730 207.700 79.330 208.150 ;
        RECT 70.130 207.550 74.080 207.700 ;
        RECT 75.380 207.550 79.330 207.700 ;
        RECT 70.130 207.100 70.730 207.550 ;
        RECT 78.730 207.100 79.330 207.550 ;
        RECT 70.130 206.950 74.080 207.100 ;
        RECT 75.380 206.950 79.330 207.100 ;
        RECT 70.130 206.500 70.730 206.950 ;
        RECT 78.730 206.500 79.330 206.950 ;
        RECT 70.130 206.350 74.080 206.500 ;
        RECT 75.380 206.350 79.330 206.500 ;
        RECT 70.130 205.900 70.730 206.350 ;
        RECT 78.730 205.900 79.330 206.350 ;
        RECT 70.130 205.750 74.080 205.900 ;
        RECT 75.380 205.750 79.330 205.900 ;
        RECT 70.130 205.300 70.730 205.750 ;
        RECT 78.730 205.300 79.330 205.750 ;
        RECT 70.130 205.150 74.080 205.300 ;
        RECT 75.380 205.150 79.330 205.300 ;
        RECT 70.130 204.700 70.730 205.150 ;
        RECT 78.730 204.700 79.330 205.150 ;
        RECT 70.130 204.550 74.080 204.700 ;
        RECT 75.380 204.550 79.330 204.700 ;
        RECT 70.130 204.100 70.730 204.550 ;
        RECT 78.730 204.100 79.330 204.550 ;
        RECT 70.130 203.950 74.080 204.100 ;
        RECT 75.380 203.950 79.330 204.100 ;
        RECT 70.130 203.500 70.730 203.950 ;
        RECT 78.730 203.500 79.330 203.950 ;
        RECT 70.130 203.350 74.080 203.500 ;
        RECT 75.380 203.350 79.330 203.500 ;
        RECT 70.130 202.900 70.730 203.350 ;
        RECT 78.730 202.900 79.330 203.350 ;
        RECT 70.130 202.750 74.080 202.900 ;
        RECT 75.380 202.750 79.330 202.900 ;
        RECT 70.130 202.300 70.730 202.750 ;
        RECT 78.730 202.300 79.330 202.750 ;
        RECT 70.130 202.150 74.080 202.300 ;
        RECT 75.380 202.150 79.330 202.300 ;
        RECT 70.130 202.000 70.730 202.150 ;
        RECT 66.530 201.700 70.730 202.000 ;
        RECT 78.730 202.000 79.330 202.150 ;
        RECT 79.780 202.000 79.930 209.550 ;
        RECT 80.380 202.000 80.530 209.550 ;
        RECT 80.980 202.000 81.130 209.550 ;
        RECT 81.580 202.000 81.730 209.550 ;
        RECT 82.180 202.000 82.330 209.550 ;
        RECT 82.780 202.000 82.930 204.900 ;
        RECT 78.730 201.700 82.930 202.000 ;
        RECT 66.530 201.550 74.080 201.700 ;
        RECT 75.380 201.550 82.930 201.700 ;
        RECT 66.530 201.350 70.730 201.550 ;
        RECT 60.330 201.050 69.130 201.200 ;
        RECT 69.280 201.050 70.730 201.350 ;
        RECT 58.730 200.150 70.730 201.050 ;
        RECT 78.730 201.350 82.930 201.550 ;
        RECT 78.730 201.050 80.180 201.350 ;
        RECT 83.530 201.200 85.930 204.400 ;
        RECT 86.530 202.000 86.680 204.900 ;
        RECT 87.130 202.000 87.280 209.550 ;
        RECT 87.730 202.000 87.880 209.550 ;
        RECT 88.330 202.000 88.480 209.550 ;
        RECT 88.930 202.000 89.080 209.550 ;
        RECT 89.530 202.000 89.680 209.550 ;
        RECT 90.130 209.350 94.080 209.550 ;
        RECT 95.380 209.350 99.330 209.550 ;
        RECT 90.130 208.900 90.730 209.350 ;
        RECT 98.730 208.900 99.330 209.350 ;
        RECT 90.130 208.750 94.080 208.900 ;
        RECT 95.380 208.750 99.330 208.900 ;
        RECT 90.130 208.300 90.730 208.750 ;
        RECT 98.730 208.300 99.330 208.750 ;
        RECT 90.130 208.150 94.080 208.300 ;
        RECT 95.380 208.150 99.330 208.300 ;
        RECT 90.130 207.700 90.730 208.150 ;
        RECT 98.730 207.700 99.330 208.150 ;
        RECT 90.130 207.550 94.080 207.700 ;
        RECT 95.380 207.550 99.330 207.700 ;
        RECT 90.130 207.100 90.730 207.550 ;
        RECT 98.730 207.100 99.330 207.550 ;
        RECT 90.130 206.950 94.080 207.100 ;
        RECT 95.380 206.950 99.330 207.100 ;
        RECT 90.130 206.500 90.730 206.950 ;
        RECT 98.730 206.500 99.330 206.950 ;
        RECT 90.130 206.350 94.080 206.500 ;
        RECT 95.380 206.350 99.330 206.500 ;
        RECT 90.130 205.900 90.730 206.350 ;
        RECT 98.730 205.900 99.330 206.350 ;
        RECT 90.130 205.750 94.080 205.900 ;
        RECT 95.380 205.750 99.330 205.900 ;
        RECT 90.130 205.300 90.730 205.750 ;
        RECT 98.730 205.300 99.330 205.750 ;
        RECT 90.130 205.150 94.080 205.300 ;
        RECT 95.380 205.150 99.330 205.300 ;
        RECT 90.130 204.700 90.730 205.150 ;
        RECT 98.730 204.700 99.330 205.150 ;
        RECT 90.130 204.550 94.080 204.700 ;
        RECT 95.380 204.550 99.330 204.700 ;
        RECT 90.130 204.100 90.730 204.550 ;
        RECT 98.730 204.100 99.330 204.550 ;
        RECT 90.130 203.950 94.080 204.100 ;
        RECT 95.380 203.950 99.330 204.100 ;
        RECT 90.130 203.500 90.730 203.950 ;
        RECT 98.730 203.500 99.330 203.950 ;
        RECT 90.130 203.350 94.080 203.500 ;
        RECT 95.380 203.350 99.330 203.500 ;
        RECT 90.130 202.900 90.730 203.350 ;
        RECT 98.730 202.900 99.330 203.350 ;
        RECT 90.130 202.750 94.080 202.900 ;
        RECT 95.380 202.750 99.330 202.900 ;
        RECT 90.130 202.300 90.730 202.750 ;
        RECT 98.730 202.300 99.330 202.750 ;
        RECT 90.130 202.150 94.080 202.300 ;
        RECT 95.380 202.150 99.330 202.300 ;
        RECT 90.130 202.000 90.730 202.150 ;
        RECT 86.530 201.700 90.730 202.000 ;
        RECT 98.730 202.000 99.330 202.150 ;
        RECT 99.780 202.000 99.930 209.550 ;
        RECT 100.380 202.000 100.530 209.550 ;
        RECT 100.980 202.000 101.130 209.550 ;
        RECT 101.580 202.000 101.730 209.550 ;
        RECT 102.180 202.000 102.330 209.550 ;
        RECT 102.780 202.000 102.930 204.900 ;
        RECT 98.730 201.700 102.930 202.000 ;
        RECT 86.530 201.550 94.080 201.700 ;
        RECT 95.380 201.550 102.930 201.700 ;
        RECT 86.530 201.350 90.730 201.550 ;
        RECT 80.330 201.050 89.130 201.200 ;
        RECT 89.280 201.050 90.730 201.350 ;
        RECT 78.730 200.150 90.730 201.050 ;
        RECT 98.730 201.350 102.930 201.550 ;
        RECT 98.730 201.050 100.180 201.350 ;
        RECT 103.530 201.200 105.930 204.400 ;
        RECT 106.530 202.000 106.680 204.900 ;
        RECT 107.130 202.000 107.280 209.550 ;
        RECT 107.730 202.000 107.880 209.550 ;
        RECT 108.330 202.000 108.480 209.550 ;
        RECT 108.930 202.000 109.080 209.550 ;
        RECT 109.530 202.000 109.680 209.550 ;
        RECT 110.130 209.350 114.080 209.550 ;
        RECT 115.380 209.350 119.330 209.550 ;
        RECT 110.130 208.900 110.730 209.350 ;
        RECT 118.730 208.900 119.330 209.350 ;
        RECT 110.130 208.750 114.080 208.900 ;
        RECT 115.380 208.750 119.330 208.900 ;
        RECT 110.130 208.300 110.730 208.750 ;
        RECT 118.730 208.300 119.330 208.750 ;
        RECT 110.130 208.150 114.080 208.300 ;
        RECT 115.380 208.150 119.330 208.300 ;
        RECT 110.130 207.700 110.730 208.150 ;
        RECT 118.730 207.700 119.330 208.150 ;
        RECT 110.130 207.550 114.080 207.700 ;
        RECT 115.380 207.550 119.330 207.700 ;
        RECT 110.130 207.100 110.730 207.550 ;
        RECT 118.730 207.100 119.330 207.550 ;
        RECT 110.130 206.950 114.080 207.100 ;
        RECT 115.380 206.950 119.330 207.100 ;
        RECT 110.130 206.500 110.730 206.950 ;
        RECT 118.730 206.500 119.330 206.950 ;
        RECT 110.130 206.350 114.080 206.500 ;
        RECT 115.380 206.350 119.330 206.500 ;
        RECT 110.130 205.900 110.730 206.350 ;
        RECT 118.730 205.900 119.330 206.350 ;
        RECT 110.130 205.750 114.080 205.900 ;
        RECT 115.380 205.750 119.330 205.900 ;
        RECT 110.130 205.300 110.730 205.750 ;
        RECT 118.730 205.300 119.330 205.750 ;
        RECT 110.130 205.150 114.080 205.300 ;
        RECT 115.380 205.150 119.330 205.300 ;
        RECT 110.130 204.700 110.730 205.150 ;
        RECT 118.730 204.700 119.330 205.150 ;
        RECT 110.130 204.550 114.080 204.700 ;
        RECT 115.380 204.550 119.330 204.700 ;
        RECT 110.130 204.100 110.730 204.550 ;
        RECT 118.730 204.100 119.330 204.550 ;
        RECT 110.130 203.950 114.080 204.100 ;
        RECT 115.380 203.950 119.330 204.100 ;
        RECT 110.130 203.500 110.730 203.950 ;
        RECT 118.730 203.500 119.330 203.950 ;
        RECT 110.130 203.350 114.080 203.500 ;
        RECT 115.380 203.350 119.330 203.500 ;
        RECT 110.130 202.900 110.730 203.350 ;
        RECT 118.730 202.900 119.330 203.350 ;
        RECT 110.130 202.750 114.080 202.900 ;
        RECT 115.380 202.750 119.330 202.900 ;
        RECT 110.130 202.300 110.730 202.750 ;
        RECT 118.730 202.300 119.330 202.750 ;
        RECT 110.130 202.150 114.080 202.300 ;
        RECT 115.380 202.150 119.330 202.300 ;
        RECT 110.130 202.000 110.730 202.150 ;
        RECT 106.530 201.700 110.730 202.000 ;
        RECT 118.730 202.000 119.330 202.150 ;
        RECT 119.780 202.000 119.930 209.550 ;
        RECT 120.380 202.000 120.530 209.550 ;
        RECT 120.980 202.000 121.130 209.550 ;
        RECT 121.580 202.000 121.730 209.550 ;
        RECT 122.180 202.000 122.330 209.550 ;
        RECT 122.780 202.000 122.930 204.900 ;
        RECT 118.730 201.700 122.930 202.000 ;
        RECT 106.530 201.550 114.080 201.700 ;
        RECT 115.380 201.550 122.930 201.700 ;
        RECT 106.530 201.350 110.730 201.550 ;
        RECT 100.330 201.050 109.130 201.200 ;
        RECT 109.280 201.050 110.730 201.350 ;
        RECT 98.730 200.150 110.730 201.050 ;
        RECT 118.730 201.350 122.930 201.550 ;
        RECT 123.530 202.185 124.730 204.400 ;
        RECT 118.730 201.050 120.180 201.350 ;
        RECT 123.530 201.200 127.140 202.185 ;
        RECT 120.330 201.050 127.140 201.200 ;
        RECT 118.730 200.910 127.140 201.050 ;
        RECT 118.730 200.150 124.730 200.910 ;
        RECT 4.730 200.000 9.130 200.150 ;
        RECT 20.330 200.000 29.130 200.150 ;
        RECT 40.330 200.000 49.130 200.150 ;
        RECT 60.330 200.000 69.130 200.150 ;
        RECT 80.330 200.000 89.130 200.150 ;
        RECT 100.330 200.000 109.130 200.150 ;
        RECT 120.330 200.000 124.730 200.150 ;
        RECT 42.635 176.510 47.035 176.660 ;
        RECT 58.235 176.510 67.035 176.660 ;
        RECT 78.235 176.510 87.035 176.660 ;
        RECT 98.235 176.510 107.035 176.660 ;
        RECT 4.720 175.695 6.190 175.865 ;
        RECT 7.100 175.695 7.560 175.700 ;
        RECT 2.315 175.215 23.605 175.695 ;
        RECT 42.635 175.610 48.635 176.510 ;
        RECT 58.235 176.460 68.635 176.510 ;
        RECT 78.235 176.460 88.635 176.510 ;
        RECT 98.235 176.460 108.635 176.510 ;
        RECT 118.235 176.460 122.635 176.660 ;
        RECT 42.635 175.460 47.035 175.610 ;
        RECT 4.720 174.615 6.190 175.215 ;
        RECT 7.960 174.410 9.830 174.770 ;
        RECT 42.635 172.260 43.835 175.460 ;
        RECT 47.185 175.310 48.635 175.610 ;
        RECT 44.435 175.110 48.635 175.310 ;
        RECT 56.635 175.610 68.635 176.460 ;
        RECT 56.635 175.560 67.035 175.610 ;
        RECT 56.635 175.310 58.085 175.560 ;
        RECT 58.235 175.460 67.035 175.560 ;
        RECT 56.635 175.110 60.835 175.310 ;
        RECT 44.435 174.960 51.985 175.110 ;
        RECT 53.335 174.960 60.835 175.110 ;
        RECT 44.435 174.660 48.635 174.960 ;
        RECT 44.435 171.810 44.585 174.660 ;
        RECT 2.315 169.775 24.065 170.255 ;
        RECT 45.035 167.110 45.185 174.660 ;
        RECT 45.635 167.110 45.785 174.660 ;
        RECT 46.235 167.110 46.385 174.660 ;
        RECT 46.835 167.110 46.985 174.660 ;
        RECT 47.435 167.110 47.585 174.660 ;
        RECT 48.035 174.510 48.635 174.660 ;
        RECT 56.635 174.660 60.835 174.960 ;
        RECT 56.635 174.510 57.235 174.660 ;
        RECT 48.035 174.360 51.985 174.510 ;
        RECT 53.285 174.360 57.235 174.510 ;
        RECT 48.035 173.910 48.635 174.360 ;
        RECT 56.635 173.910 57.235 174.360 ;
        RECT 48.035 173.760 51.985 173.910 ;
        RECT 53.285 173.760 57.235 173.910 ;
        RECT 48.035 173.310 48.635 173.760 ;
        RECT 56.635 173.310 57.235 173.760 ;
        RECT 48.035 173.160 51.985 173.310 ;
        RECT 53.285 173.160 57.235 173.310 ;
        RECT 48.035 172.710 48.635 173.160 ;
        RECT 56.635 172.710 57.235 173.160 ;
        RECT 48.035 172.560 51.985 172.710 ;
        RECT 53.285 172.560 57.235 172.710 ;
        RECT 48.035 172.110 48.635 172.560 ;
        RECT 56.635 172.110 57.235 172.560 ;
        RECT 48.035 171.960 51.985 172.110 ;
        RECT 53.285 171.960 57.235 172.110 ;
        RECT 48.035 171.510 48.635 171.960 ;
        RECT 56.635 171.510 57.235 171.960 ;
        RECT 48.035 171.360 51.985 171.510 ;
        RECT 53.285 171.360 57.235 171.510 ;
        RECT 48.035 170.910 48.635 171.360 ;
        RECT 56.635 170.910 57.235 171.360 ;
        RECT 48.035 170.760 51.985 170.910 ;
        RECT 53.285 170.760 57.235 170.910 ;
        RECT 48.035 170.310 48.635 170.760 ;
        RECT 56.635 170.310 57.235 170.760 ;
        RECT 48.035 170.160 51.985 170.310 ;
        RECT 53.285 170.160 57.235 170.310 ;
        RECT 48.035 169.710 48.635 170.160 ;
        RECT 56.635 169.710 57.235 170.160 ;
        RECT 48.035 169.560 51.985 169.710 ;
        RECT 53.285 169.560 57.235 169.710 ;
        RECT 48.035 169.110 48.635 169.560 ;
        RECT 56.635 169.110 57.235 169.560 ;
        RECT 48.035 168.960 51.985 169.110 ;
        RECT 53.285 168.960 57.235 169.110 ;
        RECT 48.035 168.510 48.635 168.960 ;
        RECT 56.635 168.510 57.235 168.960 ;
        RECT 48.035 168.360 51.985 168.510 ;
        RECT 53.285 168.360 57.235 168.510 ;
        RECT 48.035 167.910 48.635 168.360 ;
        RECT 56.635 167.910 57.235 168.360 ;
        RECT 48.035 167.760 51.985 167.910 ;
        RECT 53.285 167.760 57.235 167.910 ;
        RECT 48.035 167.310 48.635 167.760 ;
        RECT 56.635 167.310 57.235 167.760 ;
        RECT 48.035 167.110 51.985 167.310 ;
        RECT 53.285 167.110 57.235 167.310 ;
        RECT 57.685 167.110 57.835 174.660 ;
        RECT 58.285 167.110 58.435 174.660 ;
        RECT 58.885 167.110 59.035 174.660 ;
        RECT 59.485 167.110 59.635 174.660 ;
        RECT 60.085 167.110 60.235 174.660 ;
        RECT 60.685 171.810 60.835 174.660 ;
        RECT 61.435 172.260 63.835 175.460 ;
        RECT 67.185 175.310 68.635 175.610 ;
        RECT 64.435 175.110 68.635 175.310 ;
        RECT 76.635 175.610 88.635 176.460 ;
        RECT 76.635 175.560 87.035 175.610 ;
        RECT 76.635 175.310 78.085 175.560 ;
        RECT 78.235 175.460 87.035 175.560 ;
        RECT 76.635 175.110 80.835 175.310 ;
        RECT 64.435 174.960 71.985 175.110 ;
        RECT 73.335 174.960 80.835 175.110 ;
        RECT 64.435 174.660 68.635 174.960 ;
        RECT 64.435 171.810 64.585 174.660 ;
        RECT 65.035 167.110 65.185 174.660 ;
        RECT 65.635 167.110 65.785 174.660 ;
        RECT 66.235 167.110 66.385 174.660 ;
        RECT 66.835 167.110 66.985 174.660 ;
        RECT 67.435 167.110 67.585 174.660 ;
        RECT 68.035 174.510 68.635 174.660 ;
        RECT 76.635 174.660 80.835 174.960 ;
        RECT 76.635 174.510 77.235 174.660 ;
        RECT 68.035 174.360 71.985 174.510 ;
        RECT 73.285 174.360 77.235 174.510 ;
        RECT 68.035 173.910 68.635 174.360 ;
        RECT 76.635 173.910 77.235 174.360 ;
        RECT 68.035 173.760 71.985 173.910 ;
        RECT 73.285 173.760 77.235 173.910 ;
        RECT 68.035 173.310 68.635 173.760 ;
        RECT 76.635 173.310 77.235 173.760 ;
        RECT 68.035 173.160 71.985 173.310 ;
        RECT 73.285 173.160 77.235 173.310 ;
        RECT 68.035 172.710 68.635 173.160 ;
        RECT 76.635 172.710 77.235 173.160 ;
        RECT 68.035 172.560 71.985 172.710 ;
        RECT 73.285 172.560 77.235 172.710 ;
        RECT 68.035 172.110 68.635 172.560 ;
        RECT 76.635 172.110 77.235 172.560 ;
        RECT 68.035 171.960 71.985 172.110 ;
        RECT 73.285 171.960 77.235 172.110 ;
        RECT 68.035 171.510 68.635 171.960 ;
        RECT 76.635 171.510 77.235 171.960 ;
        RECT 68.035 171.360 71.985 171.510 ;
        RECT 73.285 171.360 77.235 171.510 ;
        RECT 68.035 170.910 68.635 171.360 ;
        RECT 76.635 170.910 77.235 171.360 ;
        RECT 68.035 170.760 71.985 170.910 ;
        RECT 73.285 170.760 77.235 170.910 ;
        RECT 68.035 170.310 68.635 170.760 ;
        RECT 76.635 170.310 77.235 170.760 ;
        RECT 68.035 170.160 71.985 170.310 ;
        RECT 73.285 170.160 77.235 170.310 ;
        RECT 68.035 169.710 68.635 170.160 ;
        RECT 76.635 169.710 77.235 170.160 ;
        RECT 68.035 169.560 71.985 169.710 ;
        RECT 73.285 169.560 77.235 169.710 ;
        RECT 68.035 169.110 68.635 169.560 ;
        RECT 76.635 169.110 77.235 169.560 ;
        RECT 68.035 168.960 71.985 169.110 ;
        RECT 73.285 168.960 77.235 169.110 ;
        RECT 68.035 168.510 68.635 168.960 ;
        RECT 76.635 168.510 77.235 168.960 ;
        RECT 68.035 168.360 71.985 168.510 ;
        RECT 73.285 168.360 77.235 168.510 ;
        RECT 68.035 167.910 68.635 168.360 ;
        RECT 76.635 167.910 77.235 168.360 ;
        RECT 68.035 167.760 71.985 167.910 ;
        RECT 73.285 167.760 77.235 167.910 ;
        RECT 68.035 167.310 68.635 167.760 ;
        RECT 76.635 167.310 77.235 167.760 ;
        RECT 68.035 167.110 71.985 167.310 ;
        RECT 73.285 167.110 77.235 167.310 ;
        RECT 77.685 167.110 77.835 174.660 ;
        RECT 78.285 167.110 78.435 174.660 ;
        RECT 78.885 167.110 79.035 174.660 ;
        RECT 79.485 167.110 79.635 174.660 ;
        RECT 80.085 167.110 80.235 174.660 ;
        RECT 80.685 171.810 80.835 174.660 ;
        RECT 81.435 172.260 83.835 175.460 ;
        RECT 87.185 175.310 88.635 175.610 ;
        RECT 84.435 175.110 88.635 175.310 ;
        RECT 96.635 175.610 108.635 176.460 ;
        RECT 96.635 175.560 107.035 175.610 ;
        RECT 96.635 175.310 98.085 175.560 ;
        RECT 98.235 175.460 107.035 175.560 ;
        RECT 96.635 175.110 100.835 175.310 ;
        RECT 84.435 174.960 91.985 175.110 ;
        RECT 93.335 174.960 100.835 175.110 ;
        RECT 84.435 174.660 88.635 174.960 ;
        RECT 84.435 171.810 84.585 174.660 ;
        RECT 85.035 167.110 85.185 174.660 ;
        RECT 85.635 167.110 85.785 174.660 ;
        RECT 86.235 167.110 86.385 174.660 ;
        RECT 86.835 167.110 86.985 174.660 ;
        RECT 87.435 167.110 87.585 174.660 ;
        RECT 88.035 174.510 88.635 174.660 ;
        RECT 96.635 174.660 100.835 174.960 ;
        RECT 96.635 174.510 97.235 174.660 ;
        RECT 88.035 174.360 91.985 174.510 ;
        RECT 93.285 174.360 97.235 174.510 ;
        RECT 88.035 173.910 88.635 174.360 ;
        RECT 96.635 173.910 97.235 174.360 ;
        RECT 88.035 173.760 91.985 173.910 ;
        RECT 93.285 173.760 97.235 173.910 ;
        RECT 88.035 173.310 88.635 173.760 ;
        RECT 96.635 173.310 97.235 173.760 ;
        RECT 88.035 173.160 91.985 173.310 ;
        RECT 93.285 173.160 97.235 173.310 ;
        RECT 88.035 172.710 88.635 173.160 ;
        RECT 96.635 172.710 97.235 173.160 ;
        RECT 88.035 172.560 91.985 172.710 ;
        RECT 93.285 172.560 97.235 172.710 ;
        RECT 88.035 172.110 88.635 172.560 ;
        RECT 96.635 172.110 97.235 172.560 ;
        RECT 88.035 171.960 91.985 172.110 ;
        RECT 93.285 171.960 97.235 172.110 ;
        RECT 88.035 171.510 88.635 171.960 ;
        RECT 96.635 171.510 97.235 171.960 ;
        RECT 88.035 171.360 91.985 171.510 ;
        RECT 93.285 171.360 97.235 171.510 ;
        RECT 88.035 170.910 88.635 171.360 ;
        RECT 96.635 170.910 97.235 171.360 ;
        RECT 88.035 170.760 91.985 170.910 ;
        RECT 93.285 170.760 97.235 170.910 ;
        RECT 88.035 170.310 88.635 170.760 ;
        RECT 96.635 170.310 97.235 170.760 ;
        RECT 88.035 170.160 91.985 170.310 ;
        RECT 93.285 170.160 97.235 170.310 ;
        RECT 88.035 169.710 88.635 170.160 ;
        RECT 96.635 169.710 97.235 170.160 ;
        RECT 88.035 169.560 91.985 169.710 ;
        RECT 93.285 169.560 97.235 169.710 ;
        RECT 88.035 169.110 88.635 169.560 ;
        RECT 96.635 169.110 97.235 169.560 ;
        RECT 88.035 168.960 91.985 169.110 ;
        RECT 93.285 168.960 97.235 169.110 ;
        RECT 88.035 168.510 88.635 168.960 ;
        RECT 96.635 168.510 97.235 168.960 ;
        RECT 88.035 168.360 91.985 168.510 ;
        RECT 93.285 168.360 97.235 168.510 ;
        RECT 88.035 167.910 88.635 168.360 ;
        RECT 96.635 167.910 97.235 168.360 ;
        RECT 88.035 167.760 91.985 167.910 ;
        RECT 93.285 167.760 97.235 167.910 ;
        RECT 88.035 167.310 88.635 167.760 ;
        RECT 96.635 167.310 97.235 167.760 ;
        RECT 88.035 167.110 91.985 167.310 ;
        RECT 93.285 167.110 97.235 167.310 ;
        RECT 97.685 167.110 97.835 174.660 ;
        RECT 98.285 167.110 98.435 174.660 ;
        RECT 98.885 167.110 99.035 174.660 ;
        RECT 99.485 167.110 99.635 174.660 ;
        RECT 100.085 167.110 100.235 174.660 ;
        RECT 100.685 171.810 100.835 174.660 ;
        RECT 101.435 172.260 103.835 175.460 ;
        RECT 107.185 175.310 108.635 175.610 ;
        RECT 104.435 175.110 108.635 175.310 ;
        RECT 116.635 175.560 122.635 176.460 ;
        RECT 116.635 175.310 118.085 175.560 ;
        RECT 118.235 175.460 122.635 175.560 ;
        RECT 116.635 175.110 120.835 175.310 ;
        RECT 104.435 174.960 111.985 175.110 ;
        RECT 113.335 174.960 120.835 175.110 ;
        RECT 104.435 174.660 108.635 174.960 ;
        RECT 104.435 171.810 104.585 174.660 ;
        RECT 105.035 167.110 105.185 174.660 ;
        RECT 105.635 167.110 105.785 174.660 ;
        RECT 106.235 167.110 106.385 174.660 ;
        RECT 106.835 167.110 106.985 174.660 ;
        RECT 107.435 167.110 107.585 174.660 ;
        RECT 108.035 174.510 108.635 174.660 ;
        RECT 116.635 174.660 120.835 174.960 ;
        RECT 116.635 174.510 117.235 174.660 ;
        RECT 108.035 174.360 111.985 174.510 ;
        RECT 113.285 174.360 117.235 174.510 ;
        RECT 108.035 173.910 108.635 174.360 ;
        RECT 116.635 173.910 117.235 174.360 ;
        RECT 108.035 173.760 111.985 173.910 ;
        RECT 113.285 173.760 117.235 173.910 ;
        RECT 108.035 173.310 108.635 173.760 ;
        RECT 116.635 173.310 117.235 173.760 ;
        RECT 108.035 173.160 111.985 173.310 ;
        RECT 113.285 173.160 117.235 173.310 ;
        RECT 108.035 172.710 108.635 173.160 ;
        RECT 116.635 172.710 117.235 173.160 ;
        RECT 108.035 172.560 111.985 172.710 ;
        RECT 113.285 172.560 117.235 172.710 ;
        RECT 108.035 172.110 108.635 172.560 ;
        RECT 116.635 172.110 117.235 172.560 ;
        RECT 108.035 171.960 111.985 172.110 ;
        RECT 113.285 171.960 117.235 172.110 ;
        RECT 108.035 171.510 108.635 171.960 ;
        RECT 116.635 171.510 117.235 171.960 ;
        RECT 108.035 171.360 111.985 171.510 ;
        RECT 113.285 171.360 117.235 171.510 ;
        RECT 108.035 170.910 108.635 171.360 ;
        RECT 116.635 170.910 117.235 171.360 ;
        RECT 108.035 170.760 111.985 170.910 ;
        RECT 113.285 170.760 117.235 170.910 ;
        RECT 108.035 170.310 108.635 170.760 ;
        RECT 116.635 170.310 117.235 170.760 ;
        RECT 108.035 170.160 111.985 170.310 ;
        RECT 113.285 170.160 117.235 170.310 ;
        RECT 108.035 169.710 108.635 170.160 ;
        RECT 116.635 169.710 117.235 170.160 ;
        RECT 108.035 169.560 111.985 169.710 ;
        RECT 113.285 169.560 117.235 169.710 ;
        RECT 108.035 169.110 108.635 169.560 ;
        RECT 116.635 169.110 117.235 169.560 ;
        RECT 108.035 168.960 111.985 169.110 ;
        RECT 113.285 168.960 117.235 169.110 ;
        RECT 108.035 168.510 108.635 168.960 ;
        RECT 116.635 168.510 117.235 168.960 ;
        RECT 108.035 168.360 111.985 168.510 ;
        RECT 113.285 168.360 117.235 168.510 ;
        RECT 108.035 167.910 108.635 168.360 ;
        RECT 116.635 167.910 117.235 168.360 ;
        RECT 108.035 167.760 111.985 167.910 ;
        RECT 113.285 167.760 117.235 167.910 ;
        RECT 108.035 167.310 108.635 167.760 ;
        RECT 116.635 167.310 117.235 167.760 ;
        RECT 108.035 167.110 111.985 167.310 ;
        RECT 113.285 167.110 117.235 167.310 ;
        RECT 117.685 167.110 117.835 174.660 ;
        RECT 118.285 167.110 118.435 174.660 ;
        RECT 118.885 167.110 119.035 174.660 ;
        RECT 119.485 167.110 119.635 174.660 ;
        RECT 120.085 167.110 120.235 174.660 ;
        RECT 120.685 171.810 120.835 174.660 ;
        RECT 121.435 174.990 122.635 175.460 ;
        RECT 121.435 173.715 127.140 174.990 ;
        RECT 121.435 172.260 122.635 173.715 ;
        RECT 125.140 169.915 127.140 172.210 ;
        RECT 125.140 169.910 127.005 169.915 ;
        RECT 4.720 164.815 6.190 165.555 ;
        RECT 2.315 164.335 23.605 164.815 ;
        RECT 4.720 164.175 6.190 164.335 ;
        RECT 42.635 157.860 43.835 161.060 ;
        RECT 44.435 158.660 44.585 161.560 ;
        RECT 45.035 158.660 45.185 166.210 ;
        RECT 45.635 158.660 45.785 166.210 ;
        RECT 46.235 158.660 46.385 166.210 ;
        RECT 46.835 158.660 46.985 166.210 ;
        RECT 47.435 158.660 47.585 166.210 ;
        RECT 48.035 166.010 51.985 166.210 ;
        RECT 53.285 166.010 57.235 166.210 ;
        RECT 48.035 165.560 48.635 166.010 ;
        RECT 56.635 165.560 57.235 166.010 ;
        RECT 48.035 165.410 51.985 165.560 ;
        RECT 53.285 165.410 57.235 165.560 ;
        RECT 48.035 164.960 48.635 165.410 ;
        RECT 56.635 164.960 57.235 165.410 ;
        RECT 48.035 164.810 51.985 164.960 ;
        RECT 53.285 164.810 57.235 164.960 ;
        RECT 48.035 164.360 48.635 164.810 ;
        RECT 56.635 164.360 57.235 164.810 ;
        RECT 48.035 164.210 51.985 164.360 ;
        RECT 53.285 164.210 57.235 164.360 ;
        RECT 48.035 163.760 48.635 164.210 ;
        RECT 56.635 163.760 57.235 164.210 ;
        RECT 48.035 163.610 51.985 163.760 ;
        RECT 53.285 163.610 57.235 163.760 ;
        RECT 48.035 163.160 48.635 163.610 ;
        RECT 56.635 163.160 57.235 163.610 ;
        RECT 48.035 163.010 51.985 163.160 ;
        RECT 53.285 163.010 57.235 163.160 ;
        RECT 48.035 162.560 48.635 163.010 ;
        RECT 56.635 162.560 57.235 163.010 ;
        RECT 48.035 162.410 51.985 162.560 ;
        RECT 53.285 162.410 57.235 162.560 ;
        RECT 48.035 161.960 48.635 162.410 ;
        RECT 56.635 161.960 57.235 162.410 ;
        RECT 48.035 161.810 51.985 161.960 ;
        RECT 53.285 161.810 57.235 161.960 ;
        RECT 48.035 161.360 48.635 161.810 ;
        RECT 56.635 161.360 57.235 161.810 ;
        RECT 48.035 161.210 51.985 161.360 ;
        RECT 53.285 161.210 57.235 161.360 ;
        RECT 48.035 160.760 48.635 161.210 ;
        RECT 56.635 160.760 57.235 161.210 ;
        RECT 48.035 160.610 51.985 160.760 ;
        RECT 53.285 160.610 57.235 160.760 ;
        RECT 48.035 160.160 48.635 160.610 ;
        RECT 56.635 160.160 57.235 160.610 ;
        RECT 48.035 160.010 51.985 160.160 ;
        RECT 53.285 160.010 57.235 160.160 ;
        RECT 48.035 159.560 48.635 160.010 ;
        RECT 56.635 159.560 57.235 160.010 ;
        RECT 48.035 159.410 51.985 159.560 ;
        RECT 53.285 159.410 57.235 159.560 ;
        RECT 48.035 158.960 48.635 159.410 ;
        RECT 56.635 158.960 57.235 159.410 ;
        RECT 48.035 158.810 51.985 158.960 ;
        RECT 53.285 158.810 57.235 158.960 ;
        RECT 48.035 158.660 48.635 158.810 ;
        RECT 44.435 158.360 48.635 158.660 ;
        RECT 56.635 158.660 57.235 158.810 ;
        RECT 57.685 158.660 57.835 166.210 ;
        RECT 58.285 158.660 58.435 166.210 ;
        RECT 58.885 158.660 59.035 166.210 ;
        RECT 59.485 158.660 59.635 166.210 ;
        RECT 60.085 158.660 60.235 166.210 ;
        RECT 60.685 158.660 60.835 161.560 ;
        RECT 56.635 158.360 60.835 158.660 ;
        RECT 44.435 158.210 51.985 158.360 ;
        RECT 53.285 158.210 60.835 158.360 ;
        RECT 44.435 158.010 48.635 158.210 ;
        RECT 42.635 157.710 47.035 157.860 ;
        RECT 47.185 157.710 48.635 158.010 ;
        RECT 42.635 156.810 48.635 157.710 ;
        RECT 56.635 158.010 60.835 158.210 ;
        RECT 56.635 157.710 58.085 158.010 ;
        RECT 61.435 157.860 63.835 161.060 ;
        RECT 64.435 158.660 64.585 161.560 ;
        RECT 65.035 158.660 65.185 166.210 ;
        RECT 65.635 158.660 65.785 166.210 ;
        RECT 66.235 158.660 66.385 166.210 ;
        RECT 66.835 158.660 66.985 166.210 ;
        RECT 67.435 158.660 67.585 166.210 ;
        RECT 68.035 166.010 71.985 166.210 ;
        RECT 73.285 166.010 77.235 166.210 ;
        RECT 68.035 165.560 68.635 166.010 ;
        RECT 76.635 165.560 77.235 166.010 ;
        RECT 68.035 165.410 71.985 165.560 ;
        RECT 73.285 165.410 77.235 165.560 ;
        RECT 68.035 164.960 68.635 165.410 ;
        RECT 76.635 164.960 77.235 165.410 ;
        RECT 68.035 164.810 71.985 164.960 ;
        RECT 73.285 164.810 77.235 164.960 ;
        RECT 68.035 164.360 68.635 164.810 ;
        RECT 76.635 164.360 77.235 164.810 ;
        RECT 68.035 164.210 71.985 164.360 ;
        RECT 73.285 164.210 77.235 164.360 ;
        RECT 68.035 163.760 68.635 164.210 ;
        RECT 76.635 163.760 77.235 164.210 ;
        RECT 68.035 163.610 71.985 163.760 ;
        RECT 73.285 163.610 77.235 163.760 ;
        RECT 68.035 163.160 68.635 163.610 ;
        RECT 76.635 163.160 77.235 163.610 ;
        RECT 68.035 163.010 71.985 163.160 ;
        RECT 73.285 163.010 77.235 163.160 ;
        RECT 68.035 162.560 68.635 163.010 ;
        RECT 76.635 162.560 77.235 163.010 ;
        RECT 68.035 162.410 71.985 162.560 ;
        RECT 73.285 162.410 77.235 162.560 ;
        RECT 68.035 161.960 68.635 162.410 ;
        RECT 76.635 161.960 77.235 162.410 ;
        RECT 68.035 161.810 71.985 161.960 ;
        RECT 73.285 161.810 77.235 161.960 ;
        RECT 68.035 161.360 68.635 161.810 ;
        RECT 76.635 161.360 77.235 161.810 ;
        RECT 68.035 161.210 71.985 161.360 ;
        RECT 73.285 161.210 77.235 161.360 ;
        RECT 68.035 160.760 68.635 161.210 ;
        RECT 76.635 160.760 77.235 161.210 ;
        RECT 68.035 160.610 71.985 160.760 ;
        RECT 73.285 160.610 77.235 160.760 ;
        RECT 68.035 160.160 68.635 160.610 ;
        RECT 76.635 160.160 77.235 160.610 ;
        RECT 68.035 160.010 71.985 160.160 ;
        RECT 73.285 160.010 77.235 160.160 ;
        RECT 68.035 159.560 68.635 160.010 ;
        RECT 76.635 159.560 77.235 160.010 ;
        RECT 68.035 159.410 71.985 159.560 ;
        RECT 73.285 159.410 77.235 159.560 ;
        RECT 68.035 158.960 68.635 159.410 ;
        RECT 76.635 158.960 77.235 159.410 ;
        RECT 68.035 158.810 71.985 158.960 ;
        RECT 73.285 158.810 77.235 158.960 ;
        RECT 68.035 158.660 68.635 158.810 ;
        RECT 64.435 158.360 68.635 158.660 ;
        RECT 76.635 158.660 77.235 158.810 ;
        RECT 77.685 158.660 77.835 166.210 ;
        RECT 78.285 158.660 78.435 166.210 ;
        RECT 78.885 158.660 79.035 166.210 ;
        RECT 79.485 158.660 79.635 166.210 ;
        RECT 80.085 158.660 80.235 166.210 ;
        RECT 80.685 158.660 80.835 161.560 ;
        RECT 76.635 158.360 80.835 158.660 ;
        RECT 64.435 158.210 71.985 158.360 ;
        RECT 73.285 158.210 80.835 158.360 ;
        RECT 64.435 158.010 68.635 158.210 ;
        RECT 58.235 157.710 67.035 157.860 ;
        RECT 67.185 157.710 68.635 158.010 ;
        RECT 56.635 156.810 68.635 157.710 ;
        RECT 76.635 158.010 80.835 158.210 ;
        RECT 76.635 157.710 78.085 158.010 ;
        RECT 81.435 157.860 83.835 161.060 ;
        RECT 84.435 158.660 84.585 161.560 ;
        RECT 85.035 158.660 85.185 166.210 ;
        RECT 85.635 158.660 85.785 166.210 ;
        RECT 86.235 158.660 86.385 166.210 ;
        RECT 86.835 158.660 86.985 166.210 ;
        RECT 87.435 158.660 87.585 166.210 ;
        RECT 88.035 166.010 91.985 166.210 ;
        RECT 93.285 166.010 97.235 166.210 ;
        RECT 88.035 165.560 88.635 166.010 ;
        RECT 96.635 165.560 97.235 166.010 ;
        RECT 88.035 165.410 91.985 165.560 ;
        RECT 93.285 165.410 97.235 165.560 ;
        RECT 88.035 164.960 88.635 165.410 ;
        RECT 96.635 164.960 97.235 165.410 ;
        RECT 88.035 164.810 91.985 164.960 ;
        RECT 93.285 164.810 97.235 164.960 ;
        RECT 88.035 164.360 88.635 164.810 ;
        RECT 96.635 164.360 97.235 164.810 ;
        RECT 88.035 164.210 91.985 164.360 ;
        RECT 93.285 164.210 97.235 164.360 ;
        RECT 88.035 163.760 88.635 164.210 ;
        RECT 96.635 163.760 97.235 164.210 ;
        RECT 88.035 163.610 91.985 163.760 ;
        RECT 93.285 163.610 97.235 163.760 ;
        RECT 88.035 163.160 88.635 163.610 ;
        RECT 96.635 163.160 97.235 163.610 ;
        RECT 88.035 163.010 91.985 163.160 ;
        RECT 93.285 163.010 97.235 163.160 ;
        RECT 88.035 162.560 88.635 163.010 ;
        RECT 96.635 162.560 97.235 163.010 ;
        RECT 88.035 162.410 91.985 162.560 ;
        RECT 93.285 162.410 97.235 162.560 ;
        RECT 88.035 161.960 88.635 162.410 ;
        RECT 96.635 161.960 97.235 162.410 ;
        RECT 88.035 161.810 91.985 161.960 ;
        RECT 93.285 161.810 97.235 161.960 ;
        RECT 88.035 161.360 88.635 161.810 ;
        RECT 96.635 161.360 97.235 161.810 ;
        RECT 88.035 161.210 91.985 161.360 ;
        RECT 93.285 161.210 97.235 161.360 ;
        RECT 88.035 160.760 88.635 161.210 ;
        RECT 96.635 160.760 97.235 161.210 ;
        RECT 88.035 160.610 91.985 160.760 ;
        RECT 93.285 160.610 97.235 160.760 ;
        RECT 88.035 160.160 88.635 160.610 ;
        RECT 96.635 160.160 97.235 160.610 ;
        RECT 88.035 160.010 91.985 160.160 ;
        RECT 93.285 160.010 97.235 160.160 ;
        RECT 88.035 159.560 88.635 160.010 ;
        RECT 96.635 159.560 97.235 160.010 ;
        RECT 88.035 159.410 91.985 159.560 ;
        RECT 93.285 159.410 97.235 159.560 ;
        RECT 88.035 158.960 88.635 159.410 ;
        RECT 96.635 158.960 97.235 159.410 ;
        RECT 88.035 158.810 91.985 158.960 ;
        RECT 93.285 158.810 97.235 158.960 ;
        RECT 88.035 158.660 88.635 158.810 ;
        RECT 84.435 158.360 88.635 158.660 ;
        RECT 96.635 158.660 97.235 158.810 ;
        RECT 97.685 158.660 97.835 166.210 ;
        RECT 98.285 158.660 98.435 166.210 ;
        RECT 98.885 158.660 99.035 166.210 ;
        RECT 99.485 158.660 99.635 166.210 ;
        RECT 100.085 158.660 100.235 166.210 ;
        RECT 100.685 158.660 100.835 161.560 ;
        RECT 96.635 158.360 100.835 158.660 ;
        RECT 84.435 158.210 91.985 158.360 ;
        RECT 93.285 158.210 100.835 158.360 ;
        RECT 84.435 158.010 88.635 158.210 ;
        RECT 78.235 157.710 87.035 157.860 ;
        RECT 87.185 157.710 88.635 158.010 ;
        RECT 76.635 156.810 88.635 157.710 ;
        RECT 96.635 158.010 100.835 158.210 ;
        RECT 96.635 157.710 98.085 158.010 ;
        RECT 101.435 157.860 103.835 161.060 ;
        RECT 104.435 158.660 104.585 161.560 ;
        RECT 105.035 158.660 105.185 166.210 ;
        RECT 105.635 158.660 105.785 166.210 ;
        RECT 106.235 158.660 106.385 166.210 ;
        RECT 106.835 158.660 106.985 166.210 ;
        RECT 107.435 158.660 107.585 166.210 ;
        RECT 108.035 166.010 111.985 166.210 ;
        RECT 113.285 166.010 117.235 166.210 ;
        RECT 108.035 165.560 108.635 166.010 ;
        RECT 116.635 165.560 117.235 166.010 ;
        RECT 108.035 165.410 111.985 165.560 ;
        RECT 113.285 165.410 117.235 165.560 ;
        RECT 108.035 164.960 108.635 165.410 ;
        RECT 116.635 164.960 117.235 165.410 ;
        RECT 108.035 164.810 111.985 164.960 ;
        RECT 113.285 164.810 117.235 164.960 ;
        RECT 108.035 164.360 108.635 164.810 ;
        RECT 116.635 164.360 117.235 164.810 ;
        RECT 108.035 164.210 111.985 164.360 ;
        RECT 113.285 164.210 117.235 164.360 ;
        RECT 108.035 163.760 108.635 164.210 ;
        RECT 116.635 163.760 117.235 164.210 ;
        RECT 108.035 163.610 111.985 163.760 ;
        RECT 113.285 163.610 117.235 163.760 ;
        RECT 108.035 163.160 108.635 163.610 ;
        RECT 116.635 163.160 117.235 163.610 ;
        RECT 108.035 163.010 111.985 163.160 ;
        RECT 113.285 163.010 117.235 163.160 ;
        RECT 108.035 162.560 108.635 163.010 ;
        RECT 116.635 162.560 117.235 163.010 ;
        RECT 108.035 162.410 111.985 162.560 ;
        RECT 113.285 162.410 117.235 162.560 ;
        RECT 108.035 161.960 108.635 162.410 ;
        RECT 116.635 161.960 117.235 162.410 ;
        RECT 108.035 161.810 111.985 161.960 ;
        RECT 113.285 161.810 117.235 161.960 ;
        RECT 108.035 161.360 108.635 161.810 ;
        RECT 116.635 161.360 117.235 161.810 ;
        RECT 108.035 161.210 111.985 161.360 ;
        RECT 113.285 161.210 117.235 161.360 ;
        RECT 108.035 160.760 108.635 161.210 ;
        RECT 116.635 160.760 117.235 161.210 ;
        RECT 108.035 160.610 111.985 160.760 ;
        RECT 113.285 160.610 117.235 160.760 ;
        RECT 108.035 160.160 108.635 160.610 ;
        RECT 116.635 160.160 117.235 160.610 ;
        RECT 108.035 160.010 111.985 160.160 ;
        RECT 113.285 160.010 117.235 160.160 ;
        RECT 108.035 159.560 108.635 160.010 ;
        RECT 116.635 159.560 117.235 160.010 ;
        RECT 108.035 159.410 111.985 159.560 ;
        RECT 113.285 159.410 117.235 159.560 ;
        RECT 108.035 158.960 108.635 159.410 ;
        RECT 116.635 158.960 117.235 159.410 ;
        RECT 108.035 158.810 111.985 158.960 ;
        RECT 113.285 158.810 117.235 158.960 ;
        RECT 108.035 158.660 108.635 158.810 ;
        RECT 104.435 158.360 108.635 158.660 ;
        RECT 116.635 158.660 117.235 158.810 ;
        RECT 117.685 158.660 117.835 166.210 ;
        RECT 118.285 158.660 118.435 166.210 ;
        RECT 118.885 158.660 119.035 166.210 ;
        RECT 119.485 158.660 119.635 166.210 ;
        RECT 120.085 158.660 120.235 166.210 ;
        RECT 120.685 158.660 120.835 161.560 ;
        RECT 125.140 161.115 127.140 163.410 ;
        RECT 125.140 161.110 127.005 161.115 ;
        RECT 116.635 158.360 120.835 158.660 ;
        RECT 104.435 158.210 111.985 158.360 ;
        RECT 113.285 158.210 120.835 158.360 ;
        RECT 104.435 158.010 108.635 158.210 ;
        RECT 98.235 157.710 107.035 157.860 ;
        RECT 107.185 157.710 108.635 158.010 ;
        RECT 96.635 156.810 108.635 157.710 ;
        RECT 116.635 158.010 120.835 158.210 ;
        RECT 121.435 159.715 122.635 161.060 ;
        RECT 121.435 158.440 127.135 159.715 ;
        RECT 116.635 157.710 118.085 158.010 ;
        RECT 121.435 157.860 122.635 158.440 ;
        RECT 118.235 157.710 122.635 157.860 ;
        RECT 116.635 156.810 122.635 157.710 ;
        RECT 42.635 156.660 47.035 156.810 ;
        RECT 58.235 156.660 67.035 156.810 ;
        RECT 78.235 156.660 87.035 156.810 ;
        RECT 98.235 156.660 107.035 156.810 ;
        RECT 118.235 156.660 122.635 156.810 ;
        RECT 2.315 140.365 127.140 141.800 ;
        RECT 2.315 140.360 9.125 140.365 ;
        RECT 11.565 140.360 127.140 140.365 ;
        RECT 4.730 139.850 9.130 140.000 ;
        RECT 20.330 139.850 29.130 140.000 ;
        RECT 40.330 139.850 49.130 140.000 ;
        RECT 60.330 139.850 69.130 140.000 ;
        RECT 80.330 139.850 89.130 140.000 ;
        RECT 100.330 139.850 109.130 140.000 ;
        RECT 4.730 138.950 10.730 139.850 ;
        RECT 20.330 139.800 30.730 139.850 ;
        RECT 40.330 139.800 50.730 139.850 ;
        RECT 60.330 139.800 70.730 139.850 ;
        RECT 80.330 139.800 90.730 139.850 ;
        RECT 100.330 139.800 110.730 139.850 ;
        RECT 120.330 139.800 124.730 140.000 ;
        RECT 4.730 138.800 9.130 138.950 ;
        RECT 4.730 137.725 5.930 138.800 ;
        RECT 9.280 138.650 10.730 138.950 ;
        RECT 2.315 136.450 5.930 137.725 ;
        RECT 4.730 135.600 5.930 136.450 ;
        RECT 6.530 138.450 10.730 138.650 ;
        RECT 18.730 138.950 30.730 139.800 ;
        RECT 18.730 138.900 29.130 138.950 ;
        RECT 18.730 138.650 20.180 138.900 ;
        RECT 20.330 138.800 29.130 138.900 ;
        RECT 18.730 138.450 22.930 138.650 ;
        RECT 6.530 138.300 14.080 138.450 ;
        RECT 15.430 138.300 22.930 138.450 ;
        RECT 6.530 138.000 10.730 138.300 ;
        RECT 2.315 133.255 4.315 135.555 ;
        RECT 6.530 135.150 6.680 138.000 ;
        RECT 7.130 130.450 7.280 138.000 ;
        RECT 7.730 130.450 7.880 138.000 ;
        RECT 8.330 130.450 8.480 138.000 ;
        RECT 8.930 130.450 9.080 138.000 ;
        RECT 9.530 130.450 9.680 138.000 ;
        RECT 10.130 137.850 10.730 138.000 ;
        RECT 18.730 138.000 22.930 138.300 ;
        RECT 18.730 137.850 19.330 138.000 ;
        RECT 10.130 137.700 14.080 137.850 ;
        RECT 15.380 137.700 19.330 137.850 ;
        RECT 10.130 137.250 10.730 137.700 ;
        RECT 18.730 137.250 19.330 137.700 ;
        RECT 10.130 137.100 14.080 137.250 ;
        RECT 15.380 137.100 19.330 137.250 ;
        RECT 10.130 136.650 10.730 137.100 ;
        RECT 18.730 136.650 19.330 137.100 ;
        RECT 10.130 136.500 14.080 136.650 ;
        RECT 15.380 136.500 19.330 136.650 ;
        RECT 10.130 136.050 10.730 136.500 ;
        RECT 18.730 136.050 19.330 136.500 ;
        RECT 10.130 135.900 14.080 136.050 ;
        RECT 15.380 135.900 19.330 136.050 ;
        RECT 10.130 135.450 10.730 135.900 ;
        RECT 18.730 135.450 19.330 135.900 ;
        RECT 10.130 135.300 14.080 135.450 ;
        RECT 15.380 135.300 19.330 135.450 ;
        RECT 10.130 134.850 10.730 135.300 ;
        RECT 18.730 134.850 19.330 135.300 ;
        RECT 10.130 134.700 14.080 134.850 ;
        RECT 15.380 134.700 19.330 134.850 ;
        RECT 10.130 134.250 10.730 134.700 ;
        RECT 18.730 134.250 19.330 134.700 ;
        RECT 10.130 134.100 14.080 134.250 ;
        RECT 15.380 134.100 19.330 134.250 ;
        RECT 10.130 133.650 10.730 134.100 ;
        RECT 18.730 133.650 19.330 134.100 ;
        RECT 10.130 133.500 14.080 133.650 ;
        RECT 15.380 133.500 19.330 133.650 ;
        RECT 10.130 133.050 10.730 133.500 ;
        RECT 18.730 133.050 19.330 133.500 ;
        RECT 10.130 132.900 14.080 133.050 ;
        RECT 15.380 132.900 19.330 133.050 ;
        RECT 10.130 132.450 10.730 132.900 ;
        RECT 18.730 132.450 19.330 132.900 ;
        RECT 10.130 132.300 14.080 132.450 ;
        RECT 15.380 132.300 19.330 132.450 ;
        RECT 10.130 131.850 10.730 132.300 ;
        RECT 18.730 131.850 19.330 132.300 ;
        RECT 10.130 131.700 14.080 131.850 ;
        RECT 15.380 131.700 19.330 131.850 ;
        RECT 10.130 131.250 10.730 131.700 ;
        RECT 18.730 131.250 19.330 131.700 ;
        RECT 10.130 131.100 14.080 131.250 ;
        RECT 15.380 131.100 19.330 131.250 ;
        RECT 10.130 130.650 10.730 131.100 ;
        RECT 18.730 130.650 19.330 131.100 ;
        RECT 10.130 130.450 14.080 130.650 ;
        RECT 15.380 130.450 19.330 130.650 ;
        RECT 19.780 130.450 19.930 138.000 ;
        RECT 20.380 130.450 20.530 138.000 ;
        RECT 20.980 130.450 21.130 138.000 ;
        RECT 21.580 130.450 21.730 138.000 ;
        RECT 22.180 130.450 22.330 138.000 ;
        RECT 22.780 135.150 22.930 138.000 ;
        RECT 23.530 135.600 25.930 138.800 ;
        RECT 29.280 138.650 30.730 138.950 ;
        RECT 26.530 138.450 30.730 138.650 ;
        RECT 38.730 138.950 50.730 139.800 ;
        RECT 38.730 138.900 49.130 138.950 ;
        RECT 38.730 138.650 40.180 138.900 ;
        RECT 40.330 138.800 49.130 138.900 ;
        RECT 38.730 138.450 42.930 138.650 ;
        RECT 26.530 138.300 34.080 138.450 ;
        RECT 35.430 138.300 42.930 138.450 ;
        RECT 26.530 138.000 30.730 138.300 ;
        RECT 26.530 135.150 26.680 138.000 ;
        RECT 27.130 130.450 27.280 138.000 ;
        RECT 27.730 130.450 27.880 138.000 ;
        RECT 28.330 130.450 28.480 138.000 ;
        RECT 28.930 130.450 29.080 138.000 ;
        RECT 29.530 130.450 29.680 138.000 ;
        RECT 30.130 137.850 30.730 138.000 ;
        RECT 38.730 138.000 42.930 138.300 ;
        RECT 38.730 137.850 39.330 138.000 ;
        RECT 30.130 137.700 34.080 137.850 ;
        RECT 35.380 137.700 39.330 137.850 ;
        RECT 30.130 137.250 30.730 137.700 ;
        RECT 38.730 137.250 39.330 137.700 ;
        RECT 30.130 137.100 34.080 137.250 ;
        RECT 35.380 137.100 39.330 137.250 ;
        RECT 30.130 136.650 30.730 137.100 ;
        RECT 38.730 136.650 39.330 137.100 ;
        RECT 30.130 136.500 34.080 136.650 ;
        RECT 35.380 136.500 39.330 136.650 ;
        RECT 30.130 136.050 30.730 136.500 ;
        RECT 38.730 136.050 39.330 136.500 ;
        RECT 30.130 135.900 34.080 136.050 ;
        RECT 35.380 135.900 39.330 136.050 ;
        RECT 30.130 135.450 30.730 135.900 ;
        RECT 38.730 135.450 39.330 135.900 ;
        RECT 30.130 135.300 34.080 135.450 ;
        RECT 35.380 135.300 39.330 135.450 ;
        RECT 30.130 134.850 30.730 135.300 ;
        RECT 38.730 134.850 39.330 135.300 ;
        RECT 30.130 134.700 34.080 134.850 ;
        RECT 35.380 134.700 39.330 134.850 ;
        RECT 30.130 134.250 30.730 134.700 ;
        RECT 38.730 134.250 39.330 134.700 ;
        RECT 30.130 134.100 34.080 134.250 ;
        RECT 35.380 134.100 39.330 134.250 ;
        RECT 30.130 133.650 30.730 134.100 ;
        RECT 38.730 133.650 39.330 134.100 ;
        RECT 30.130 133.500 34.080 133.650 ;
        RECT 35.380 133.500 39.330 133.650 ;
        RECT 30.130 133.050 30.730 133.500 ;
        RECT 38.730 133.050 39.330 133.500 ;
        RECT 30.130 132.900 34.080 133.050 ;
        RECT 35.380 132.900 39.330 133.050 ;
        RECT 30.130 132.450 30.730 132.900 ;
        RECT 38.730 132.450 39.330 132.900 ;
        RECT 30.130 132.300 34.080 132.450 ;
        RECT 35.380 132.300 39.330 132.450 ;
        RECT 30.130 131.850 30.730 132.300 ;
        RECT 38.730 131.850 39.330 132.300 ;
        RECT 30.130 131.700 34.080 131.850 ;
        RECT 35.380 131.700 39.330 131.850 ;
        RECT 30.130 131.250 30.730 131.700 ;
        RECT 38.730 131.250 39.330 131.700 ;
        RECT 30.130 131.100 34.080 131.250 ;
        RECT 35.380 131.100 39.330 131.250 ;
        RECT 30.130 130.650 30.730 131.100 ;
        RECT 38.730 130.650 39.330 131.100 ;
        RECT 30.130 130.450 34.080 130.650 ;
        RECT 35.380 130.450 39.330 130.650 ;
        RECT 39.780 130.450 39.930 138.000 ;
        RECT 40.380 130.450 40.530 138.000 ;
        RECT 40.980 130.450 41.130 138.000 ;
        RECT 41.580 130.450 41.730 138.000 ;
        RECT 42.180 130.450 42.330 138.000 ;
        RECT 42.780 135.150 42.930 138.000 ;
        RECT 43.530 135.600 45.930 138.800 ;
        RECT 49.280 138.650 50.730 138.950 ;
        RECT 46.530 138.450 50.730 138.650 ;
        RECT 58.730 138.950 70.730 139.800 ;
        RECT 58.730 138.900 69.130 138.950 ;
        RECT 58.730 138.650 60.180 138.900 ;
        RECT 60.330 138.800 69.130 138.900 ;
        RECT 58.730 138.450 62.930 138.650 ;
        RECT 46.530 138.300 54.080 138.450 ;
        RECT 55.430 138.300 62.930 138.450 ;
        RECT 46.530 138.000 50.730 138.300 ;
        RECT 46.530 135.150 46.680 138.000 ;
        RECT 47.130 130.450 47.280 138.000 ;
        RECT 47.730 130.450 47.880 138.000 ;
        RECT 48.330 130.450 48.480 138.000 ;
        RECT 48.930 130.450 49.080 138.000 ;
        RECT 49.530 130.450 49.680 138.000 ;
        RECT 50.130 137.850 50.730 138.000 ;
        RECT 58.730 138.000 62.930 138.300 ;
        RECT 58.730 137.850 59.330 138.000 ;
        RECT 50.130 137.700 54.080 137.850 ;
        RECT 55.380 137.700 59.330 137.850 ;
        RECT 50.130 137.250 50.730 137.700 ;
        RECT 58.730 137.250 59.330 137.700 ;
        RECT 50.130 137.100 54.080 137.250 ;
        RECT 55.380 137.100 59.330 137.250 ;
        RECT 50.130 136.650 50.730 137.100 ;
        RECT 58.730 136.650 59.330 137.100 ;
        RECT 50.130 136.500 54.080 136.650 ;
        RECT 55.380 136.500 59.330 136.650 ;
        RECT 50.130 136.050 50.730 136.500 ;
        RECT 58.730 136.050 59.330 136.500 ;
        RECT 50.130 135.900 54.080 136.050 ;
        RECT 55.380 135.900 59.330 136.050 ;
        RECT 50.130 135.450 50.730 135.900 ;
        RECT 58.730 135.450 59.330 135.900 ;
        RECT 50.130 135.300 54.080 135.450 ;
        RECT 55.380 135.300 59.330 135.450 ;
        RECT 50.130 134.850 50.730 135.300 ;
        RECT 58.730 134.850 59.330 135.300 ;
        RECT 50.130 134.700 54.080 134.850 ;
        RECT 55.380 134.700 59.330 134.850 ;
        RECT 50.130 134.250 50.730 134.700 ;
        RECT 58.730 134.250 59.330 134.700 ;
        RECT 50.130 134.100 54.080 134.250 ;
        RECT 55.380 134.100 59.330 134.250 ;
        RECT 50.130 133.650 50.730 134.100 ;
        RECT 58.730 133.650 59.330 134.100 ;
        RECT 50.130 133.500 54.080 133.650 ;
        RECT 55.380 133.500 59.330 133.650 ;
        RECT 50.130 133.050 50.730 133.500 ;
        RECT 58.730 133.050 59.330 133.500 ;
        RECT 50.130 132.900 54.080 133.050 ;
        RECT 55.380 132.900 59.330 133.050 ;
        RECT 50.130 132.450 50.730 132.900 ;
        RECT 58.730 132.450 59.330 132.900 ;
        RECT 50.130 132.300 54.080 132.450 ;
        RECT 55.380 132.300 59.330 132.450 ;
        RECT 50.130 131.850 50.730 132.300 ;
        RECT 58.730 131.850 59.330 132.300 ;
        RECT 50.130 131.700 54.080 131.850 ;
        RECT 55.380 131.700 59.330 131.850 ;
        RECT 50.130 131.250 50.730 131.700 ;
        RECT 58.730 131.250 59.330 131.700 ;
        RECT 50.130 131.100 54.080 131.250 ;
        RECT 55.380 131.100 59.330 131.250 ;
        RECT 50.130 130.650 50.730 131.100 ;
        RECT 58.730 130.650 59.330 131.100 ;
        RECT 50.130 130.450 54.080 130.650 ;
        RECT 55.380 130.450 59.330 130.650 ;
        RECT 59.780 130.450 59.930 138.000 ;
        RECT 60.380 130.450 60.530 138.000 ;
        RECT 60.980 130.450 61.130 138.000 ;
        RECT 61.580 130.450 61.730 138.000 ;
        RECT 62.180 130.450 62.330 138.000 ;
        RECT 62.780 135.150 62.930 138.000 ;
        RECT 63.530 135.600 65.930 138.800 ;
        RECT 69.280 138.650 70.730 138.950 ;
        RECT 66.530 138.450 70.730 138.650 ;
        RECT 78.730 138.950 90.730 139.800 ;
        RECT 78.730 138.900 89.130 138.950 ;
        RECT 78.730 138.650 80.180 138.900 ;
        RECT 80.330 138.800 89.130 138.900 ;
        RECT 78.730 138.450 82.930 138.650 ;
        RECT 66.530 138.300 74.080 138.450 ;
        RECT 75.430 138.300 82.930 138.450 ;
        RECT 66.530 138.000 70.730 138.300 ;
        RECT 66.530 135.150 66.680 138.000 ;
        RECT 67.130 130.450 67.280 138.000 ;
        RECT 67.730 130.450 67.880 138.000 ;
        RECT 68.330 130.450 68.480 138.000 ;
        RECT 68.930 130.450 69.080 138.000 ;
        RECT 69.530 130.450 69.680 138.000 ;
        RECT 70.130 137.850 70.730 138.000 ;
        RECT 78.730 138.000 82.930 138.300 ;
        RECT 78.730 137.850 79.330 138.000 ;
        RECT 70.130 137.700 74.080 137.850 ;
        RECT 75.380 137.700 79.330 137.850 ;
        RECT 70.130 137.250 70.730 137.700 ;
        RECT 78.730 137.250 79.330 137.700 ;
        RECT 70.130 137.100 74.080 137.250 ;
        RECT 75.380 137.100 79.330 137.250 ;
        RECT 70.130 136.650 70.730 137.100 ;
        RECT 78.730 136.650 79.330 137.100 ;
        RECT 70.130 136.500 74.080 136.650 ;
        RECT 75.380 136.500 79.330 136.650 ;
        RECT 70.130 136.050 70.730 136.500 ;
        RECT 78.730 136.050 79.330 136.500 ;
        RECT 70.130 135.900 74.080 136.050 ;
        RECT 75.380 135.900 79.330 136.050 ;
        RECT 70.130 135.450 70.730 135.900 ;
        RECT 78.730 135.450 79.330 135.900 ;
        RECT 70.130 135.300 74.080 135.450 ;
        RECT 75.380 135.300 79.330 135.450 ;
        RECT 70.130 134.850 70.730 135.300 ;
        RECT 78.730 134.850 79.330 135.300 ;
        RECT 70.130 134.700 74.080 134.850 ;
        RECT 75.380 134.700 79.330 134.850 ;
        RECT 70.130 134.250 70.730 134.700 ;
        RECT 78.730 134.250 79.330 134.700 ;
        RECT 70.130 134.100 74.080 134.250 ;
        RECT 75.380 134.100 79.330 134.250 ;
        RECT 70.130 133.650 70.730 134.100 ;
        RECT 78.730 133.650 79.330 134.100 ;
        RECT 70.130 133.500 74.080 133.650 ;
        RECT 75.380 133.500 79.330 133.650 ;
        RECT 70.130 133.050 70.730 133.500 ;
        RECT 78.730 133.050 79.330 133.500 ;
        RECT 70.130 132.900 74.080 133.050 ;
        RECT 75.380 132.900 79.330 133.050 ;
        RECT 70.130 132.450 70.730 132.900 ;
        RECT 78.730 132.450 79.330 132.900 ;
        RECT 70.130 132.300 74.080 132.450 ;
        RECT 75.380 132.300 79.330 132.450 ;
        RECT 70.130 131.850 70.730 132.300 ;
        RECT 78.730 131.850 79.330 132.300 ;
        RECT 70.130 131.700 74.080 131.850 ;
        RECT 75.380 131.700 79.330 131.850 ;
        RECT 70.130 131.250 70.730 131.700 ;
        RECT 78.730 131.250 79.330 131.700 ;
        RECT 70.130 131.100 74.080 131.250 ;
        RECT 75.380 131.100 79.330 131.250 ;
        RECT 70.130 130.650 70.730 131.100 ;
        RECT 78.730 130.650 79.330 131.100 ;
        RECT 70.130 130.450 74.080 130.650 ;
        RECT 75.380 130.450 79.330 130.650 ;
        RECT 79.780 130.450 79.930 138.000 ;
        RECT 80.380 130.450 80.530 138.000 ;
        RECT 80.980 130.450 81.130 138.000 ;
        RECT 81.580 130.450 81.730 138.000 ;
        RECT 82.180 130.450 82.330 138.000 ;
        RECT 82.780 135.150 82.930 138.000 ;
        RECT 83.530 135.600 85.930 138.800 ;
        RECT 89.280 138.650 90.730 138.950 ;
        RECT 86.530 138.450 90.730 138.650 ;
        RECT 98.730 138.950 110.730 139.800 ;
        RECT 98.730 138.900 109.130 138.950 ;
        RECT 98.730 138.650 100.180 138.900 ;
        RECT 100.330 138.800 109.130 138.900 ;
        RECT 98.730 138.450 102.930 138.650 ;
        RECT 86.530 138.300 94.080 138.450 ;
        RECT 95.430 138.300 102.930 138.450 ;
        RECT 86.530 138.000 90.730 138.300 ;
        RECT 86.530 135.150 86.680 138.000 ;
        RECT 87.130 130.450 87.280 138.000 ;
        RECT 87.730 130.450 87.880 138.000 ;
        RECT 88.330 130.450 88.480 138.000 ;
        RECT 88.930 130.450 89.080 138.000 ;
        RECT 89.530 130.450 89.680 138.000 ;
        RECT 90.130 137.850 90.730 138.000 ;
        RECT 98.730 138.000 102.930 138.300 ;
        RECT 98.730 137.850 99.330 138.000 ;
        RECT 90.130 137.700 94.080 137.850 ;
        RECT 95.380 137.700 99.330 137.850 ;
        RECT 90.130 137.250 90.730 137.700 ;
        RECT 98.730 137.250 99.330 137.700 ;
        RECT 90.130 137.100 94.080 137.250 ;
        RECT 95.380 137.100 99.330 137.250 ;
        RECT 90.130 136.650 90.730 137.100 ;
        RECT 98.730 136.650 99.330 137.100 ;
        RECT 90.130 136.500 94.080 136.650 ;
        RECT 95.380 136.500 99.330 136.650 ;
        RECT 90.130 136.050 90.730 136.500 ;
        RECT 98.730 136.050 99.330 136.500 ;
        RECT 90.130 135.900 94.080 136.050 ;
        RECT 95.380 135.900 99.330 136.050 ;
        RECT 90.130 135.450 90.730 135.900 ;
        RECT 98.730 135.450 99.330 135.900 ;
        RECT 90.130 135.300 94.080 135.450 ;
        RECT 95.380 135.300 99.330 135.450 ;
        RECT 90.130 134.850 90.730 135.300 ;
        RECT 98.730 134.850 99.330 135.300 ;
        RECT 90.130 134.700 94.080 134.850 ;
        RECT 95.380 134.700 99.330 134.850 ;
        RECT 90.130 134.250 90.730 134.700 ;
        RECT 98.730 134.250 99.330 134.700 ;
        RECT 90.130 134.100 94.080 134.250 ;
        RECT 95.380 134.100 99.330 134.250 ;
        RECT 90.130 133.650 90.730 134.100 ;
        RECT 98.730 133.650 99.330 134.100 ;
        RECT 90.130 133.500 94.080 133.650 ;
        RECT 95.380 133.500 99.330 133.650 ;
        RECT 90.130 133.050 90.730 133.500 ;
        RECT 98.730 133.050 99.330 133.500 ;
        RECT 90.130 132.900 94.080 133.050 ;
        RECT 95.380 132.900 99.330 133.050 ;
        RECT 90.130 132.450 90.730 132.900 ;
        RECT 98.730 132.450 99.330 132.900 ;
        RECT 90.130 132.300 94.080 132.450 ;
        RECT 95.380 132.300 99.330 132.450 ;
        RECT 90.130 131.850 90.730 132.300 ;
        RECT 98.730 131.850 99.330 132.300 ;
        RECT 90.130 131.700 94.080 131.850 ;
        RECT 95.380 131.700 99.330 131.850 ;
        RECT 90.130 131.250 90.730 131.700 ;
        RECT 98.730 131.250 99.330 131.700 ;
        RECT 90.130 131.100 94.080 131.250 ;
        RECT 95.380 131.100 99.330 131.250 ;
        RECT 90.130 130.650 90.730 131.100 ;
        RECT 98.730 130.650 99.330 131.100 ;
        RECT 90.130 130.450 94.080 130.650 ;
        RECT 95.380 130.450 99.330 130.650 ;
        RECT 99.780 130.450 99.930 138.000 ;
        RECT 100.380 130.450 100.530 138.000 ;
        RECT 100.980 130.450 101.130 138.000 ;
        RECT 101.580 130.450 101.730 138.000 ;
        RECT 102.180 130.450 102.330 138.000 ;
        RECT 102.780 135.150 102.930 138.000 ;
        RECT 103.530 135.600 105.930 138.800 ;
        RECT 109.280 138.650 110.730 138.950 ;
        RECT 106.530 138.450 110.730 138.650 ;
        RECT 118.730 138.900 124.730 139.800 ;
        RECT 118.730 138.650 120.180 138.900 ;
        RECT 120.330 138.800 124.730 138.900 ;
        RECT 118.730 138.450 122.930 138.650 ;
        RECT 106.530 138.300 114.080 138.450 ;
        RECT 115.430 138.300 122.930 138.450 ;
        RECT 106.530 138.000 110.730 138.300 ;
        RECT 106.530 135.150 106.680 138.000 ;
        RECT 107.130 130.450 107.280 138.000 ;
        RECT 107.730 130.450 107.880 138.000 ;
        RECT 108.330 130.450 108.480 138.000 ;
        RECT 108.930 130.450 109.080 138.000 ;
        RECT 109.530 130.450 109.680 138.000 ;
        RECT 110.130 137.850 110.730 138.000 ;
        RECT 118.730 138.000 122.930 138.300 ;
        RECT 118.730 137.850 119.330 138.000 ;
        RECT 110.130 137.700 114.080 137.850 ;
        RECT 115.380 137.700 119.330 137.850 ;
        RECT 110.130 137.250 110.730 137.700 ;
        RECT 118.730 137.250 119.330 137.700 ;
        RECT 110.130 137.100 114.080 137.250 ;
        RECT 115.380 137.100 119.330 137.250 ;
        RECT 110.130 136.650 110.730 137.100 ;
        RECT 118.730 136.650 119.330 137.100 ;
        RECT 110.130 136.500 114.080 136.650 ;
        RECT 115.380 136.500 119.330 136.650 ;
        RECT 110.130 136.050 110.730 136.500 ;
        RECT 118.730 136.050 119.330 136.500 ;
        RECT 110.130 135.900 114.080 136.050 ;
        RECT 115.380 135.900 119.330 136.050 ;
        RECT 110.130 135.450 110.730 135.900 ;
        RECT 118.730 135.450 119.330 135.900 ;
        RECT 110.130 135.300 114.080 135.450 ;
        RECT 115.380 135.300 119.330 135.450 ;
        RECT 110.130 134.850 110.730 135.300 ;
        RECT 118.730 134.850 119.330 135.300 ;
        RECT 110.130 134.700 114.080 134.850 ;
        RECT 115.380 134.700 119.330 134.850 ;
        RECT 110.130 134.250 110.730 134.700 ;
        RECT 118.730 134.250 119.330 134.700 ;
        RECT 110.130 134.100 114.080 134.250 ;
        RECT 115.380 134.100 119.330 134.250 ;
        RECT 110.130 133.650 110.730 134.100 ;
        RECT 118.730 133.650 119.330 134.100 ;
        RECT 110.130 133.500 114.080 133.650 ;
        RECT 115.380 133.500 119.330 133.650 ;
        RECT 110.130 133.050 110.730 133.500 ;
        RECT 118.730 133.050 119.330 133.500 ;
        RECT 110.130 132.900 114.080 133.050 ;
        RECT 115.380 132.900 119.330 133.050 ;
        RECT 110.130 132.450 110.730 132.900 ;
        RECT 118.730 132.450 119.330 132.900 ;
        RECT 110.130 132.300 114.080 132.450 ;
        RECT 115.380 132.300 119.330 132.450 ;
        RECT 110.130 131.850 110.730 132.300 ;
        RECT 118.730 131.850 119.330 132.300 ;
        RECT 110.130 131.700 114.080 131.850 ;
        RECT 115.380 131.700 119.330 131.850 ;
        RECT 110.130 131.250 110.730 131.700 ;
        RECT 118.730 131.250 119.330 131.700 ;
        RECT 110.130 131.100 114.080 131.250 ;
        RECT 115.380 131.100 119.330 131.250 ;
        RECT 110.130 130.650 110.730 131.100 ;
        RECT 118.730 130.650 119.330 131.100 ;
        RECT 110.130 130.450 114.080 130.650 ;
        RECT 115.380 130.450 119.330 130.650 ;
        RECT 119.780 130.450 119.930 138.000 ;
        RECT 120.380 130.450 120.530 138.000 ;
        RECT 120.980 130.450 121.130 138.000 ;
        RECT 121.580 130.450 121.730 138.000 ;
        RECT 122.180 130.450 122.330 138.000 ;
        RECT 122.780 135.150 122.930 138.000 ;
        RECT 123.530 137.725 124.730 138.800 ;
        RECT 123.530 136.450 127.140 137.725 ;
        RECT 123.530 135.600 124.730 136.450 ;
        RECT 2.315 124.425 4.315 126.750 ;
        RECT 2.315 124.420 4.310 124.425 ;
        RECT 4.720 123.405 5.930 124.400 ;
        RECT 4.730 123.165 5.930 123.405 ;
        RECT 2.315 121.890 5.930 123.165 ;
        RECT 4.730 121.200 5.930 121.890 ;
        RECT 6.530 122.000 6.680 124.900 ;
        RECT 7.130 122.000 7.280 129.550 ;
        RECT 7.730 122.000 7.880 129.550 ;
        RECT 8.330 122.000 8.480 129.550 ;
        RECT 8.930 122.000 9.080 129.550 ;
        RECT 9.530 122.000 9.680 129.550 ;
        RECT 10.130 129.350 14.080 129.550 ;
        RECT 15.380 129.350 19.330 129.550 ;
        RECT 10.130 128.900 10.730 129.350 ;
        RECT 18.730 128.900 19.330 129.350 ;
        RECT 10.130 128.750 14.080 128.900 ;
        RECT 15.380 128.750 19.330 128.900 ;
        RECT 10.130 128.300 10.730 128.750 ;
        RECT 18.730 128.300 19.330 128.750 ;
        RECT 10.130 128.150 14.080 128.300 ;
        RECT 15.380 128.150 19.330 128.300 ;
        RECT 10.130 127.700 10.730 128.150 ;
        RECT 18.730 127.700 19.330 128.150 ;
        RECT 10.130 127.550 14.080 127.700 ;
        RECT 15.380 127.550 19.330 127.700 ;
        RECT 10.130 127.100 10.730 127.550 ;
        RECT 18.730 127.100 19.330 127.550 ;
        RECT 10.130 126.950 14.080 127.100 ;
        RECT 15.380 126.950 19.330 127.100 ;
        RECT 10.130 126.500 10.730 126.950 ;
        RECT 18.730 126.500 19.330 126.950 ;
        RECT 10.130 126.350 14.080 126.500 ;
        RECT 15.380 126.350 19.330 126.500 ;
        RECT 10.130 125.900 10.730 126.350 ;
        RECT 18.730 125.900 19.330 126.350 ;
        RECT 10.130 125.750 14.080 125.900 ;
        RECT 15.380 125.750 19.330 125.900 ;
        RECT 10.130 125.300 10.730 125.750 ;
        RECT 18.730 125.300 19.330 125.750 ;
        RECT 10.130 125.150 14.080 125.300 ;
        RECT 15.380 125.150 19.330 125.300 ;
        RECT 10.130 124.700 10.730 125.150 ;
        RECT 18.730 124.700 19.330 125.150 ;
        RECT 10.130 124.550 14.080 124.700 ;
        RECT 15.380 124.550 19.330 124.700 ;
        RECT 10.130 124.100 10.730 124.550 ;
        RECT 18.730 124.100 19.330 124.550 ;
        RECT 10.130 123.950 14.080 124.100 ;
        RECT 15.380 123.950 19.330 124.100 ;
        RECT 10.130 123.500 10.730 123.950 ;
        RECT 18.730 123.500 19.330 123.950 ;
        RECT 10.130 123.350 14.080 123.500 ;
        RECT 15.380 123.350 19.330 123.500 ;
        RECT 10.130 122.900 10.730 123.350 ;
        RECT 18.730 122.900 19.330 123.350 ;
        RECT 10.130 122.750 14.080 122.900 ;
        RECT 15.380 122.750 19.330 122.900 ;
        RECT 10.130 122.300 10.730 122.750 ;
        RECT 18.730 122.300 19.330 122.750 ;
        RECT 10.130 122.150 14.080 122.300 ;
        RECT 15.380 122.150 19.330 122.300 ;
        RECT 10.130 122.000 10.730 122.150 ;
        RECT 6.530 121.700 10.730 122.000 ;
        RECT 18.730 122.000 19.330 122.150 ;
        RECT 19.780 122.000 19.930 129.550 ;
        RECT 20.380 122.000 20.530 129.550 ;
        RECT 20.980 122.000 21.130 129.550 ;
        RECT 21.580 122.000 21.730 129.550 ;
        RECT 22.180 122.000 22.330 129.550 ;
        RECT 22.780 122.000 22.930 124.900 ;
        RECT 18.730 121.700 22.930 122.000 ;
        RECT 6.530 121.550 14.080 121.700 ;
        RECT 15.380 121.550 22.930 121.700 ;
        RECT 6.530 121.350 10.730 121.550 ;
        RECT 4.730 121.050 9.130 121.200 ;
        RECT 9.280 121.050 10.730 121.350 ;
        RECT 4.730 120.150 10.730 121.050 ;
        RECT 18.730 121.350 22.930 121.550 ;
        RECT 18.730 121.050 20.180 121.350 ;
        RECT 23.530 121.200 25.930 124.400 ;
        RECT 26.530 122.000 26.680 124.900 ;
        RECT 27.130 122.000 27.280 129.550 ;
        RECT 27.730 122.000 27.880 129.550 ;
        RECT 28.330 122.000 28.480 129.550 ;
        RECT 28.930 122.000 29.080 129.550 ;
        RECT 29.530 122.000 29.680 129.550 ;
        RECT 30.130 129.350 34.080 129.550 ;
        RECT 35.380 129.350 39.330 129.550 ;
        RECT 30.130 128.900 30.730 129.350 ;
        RECT 38.730 128.900 39.330 129.350 ;
        RECT 30.130 128.750 34.080 128.900 ;
        RECT 35.380 128.750 39.330 128.900 ;
        RECT 30.130 128.300 30.730 128.750 ;
        RECT 38.730 128.300 39.330 128.750 ;
        RECT 30.130 128.150 34.080 128.300 ;
        RECT 35.380 128.150 39.330 128.300 ;
        RECT 30.130 127.700 30.730 128.150 ;
        RECT 38.730 127.700 39.330 128.150 ;
        RECT 30.130 127.550 34.080 127.700 ;
        RECT 35.380 127.550 39.330 127.700 ;
        RECT 30.130 127.100 30.730 127.550 ;
        RECT 38.730 127.100 39.330 127.550 ;
        RECT 30.130 126.950 34.080 127.100 ;
        RECT 35.380 126.950 39.330 127.100 ;
        RECT 30.130 126.500 30.730 126.950 ;
        RECT 38.730 126.500 39.330 126.950 ;
        RECT 30.130 126.350 34.080 126.500 ;
        RECT 35.380 126.350 39.330 126.500 ;
        RECT 30.130 125.900 30.730 126.350 ;
        RECT 38.730 125.900 39.330 126.350 ;
        RECT 30.130 125.750 34.080 125.900 ;
        RECT 35.380 125.750 39.330 125.900 ;
        RECT 30.130 125.300 30.730 125.750 ;
        RECT 38.730 125.300 39.330 125.750 ;
        RECT 30.130 125.150 34.080 125.300 ;
        RECT 35.380 125.150 39.330 125.300 ;
        RECT 30.130 124.700 30.730 125.150 ;
        RECT 38.730 124.700 39.330 125.150 ;
        RECT 30.130 124.550 34.080 124.700 ;
        RECT 35.380 124.550 39.330 124.700 ;
        RECT 30.130 124.100 30.730 124.550 ;
        RECT 38.730 124.100 39.330 124.550 ;
        RECT 30.130 123.950 34.080 124.100 ;
        RECT 35.380 123.950 39.330 124.100 ;
        RECT 30.130 123.500 30.730 123.950 ;
        RECT 38.730 123.500 39.330 123.950 ;
        RECT 30.130 123.350 34.080 123.500 ;
        RECT 35.380 123.350 39.330 123.500 ;
        RECT 30.130 122.900 30.730 123.350 ;
        RECT 38.730 122.900 39.330 123.350 ;
        RECT 30.130 122.750 34.080 122.900 ;
        RECT 35.380 122.750 39.330 122.900 ;
        RECT 30.130 122.300 30.730 122.750 ;
        RECT 38.730 122.300 39.330 122.750 ;
        RECT 30.130 122.150 34.080 122.300 ;
        RECT 35.380 122.150 39.330 122.300 ;
        RECT 30.130 122.000 30.730 122.150 ;
        RECT 26.530 121.700 30.730 122.000 ;
        RECT 38.730 122.000 39.330 122.150 ;
        RECT 39.780 122.000 39.930 129.550 ;
        RECT 40.380 122.000 40.530 129.550 ;
        RECT 40.980 122.000 41.130 129.550 ;
        RECT 41.580 122.000 41.730 129.550 ;
        RECT 42.180 122.000 42.330 129.550 ;
        RECT 42.780 122.000 42.930 124.900 ;
        RECT 38.730 121.700 42.930 122.000 ;
        RECT 26.530 121.550 34.080 121.700 ;
        RECT 35.380 121.550 42.930 121.700 ;
        RECT 26.530 121.350 30.730 121.550 ;
        RECT 20.330 121.050 29.130 121.200 ;
        RECT 29.280 121.050 30.730 121.350 ;
        RECT 18.730 120.150 30.730 121.050 ;
        RECT 38.730 121.350 42.930 121.550 ;
        RECT 38.730 121.050 40.180 121.350 ;
        RECT 43.530 121.200 45.930 124.400 ;
        RECT 46.530 122.000 46.680 124.900 ;
        RECT 47.130 122.000 47.280 129.550 ;
        RECT 47.730 122.000 47.880 129.550 ;
        RECT 48.330 122.000 48.480 129.550 ;
        RECT 48.930 122.000 49.080 129.550 ;
        RECT 49.530 122.000 49.680 129.550 ;
        RECT 50.130 129.350 54.080 129.550 ;
        RECT 55.380 129.350 59.330 129.550 ;
        RECT 50.130 128.900 50.730 129.350 ;
        RECT 58.730 128.900 59.330 129.350 ;
        RECT 50.130 128.750 54.080 128.900 ;
        RECT 55.380 128.750 59.330 128.900 ;
        RECT 50.130 128.300 50.730 128.750 ;
        RECT 58.730 128.300 59.330 128.750 ;
        RECT 50.130 128.150 54.080 128.300 ;
        RECT 55.380 128.150 59.330 128.300 ;
        RECT 50.130 127.700 50.730 128.150 ;
        RECT 58.730 127.700 59.330 128.150 ;
        RECT 50.130 127.550 54.080 127.700 ;
        RECT 55.380 127.550 59.330 127.700 ;
        RECT 50.130 127.100 50.730 127.550 ;
        RECT 58.730 127.100 59.330 127.550 ;
        RECT 50.130 126.950 54.080 127.100 ;
        RECT 55.380 126.950 59.330 127.100 ;
        RECT 50.130 126.500 50.730 126.950 ;
        RECT 58.730 126.500 59.330 126.950 ;
        RECT 50.130 126.350 54.080 126.500 ;
        RECT 55.380 126.350 59.330 126.500 ;
        RECT 50.130 125.900 50.730 126.350 ;
        RECT 58.730 125.900 59.330 126.350 ;
        RECT 50.130 125.750 54.080 125.900 ;
        RECT 55.380 125.750 59.330 125.900 ;
        RECT 50.130 125.300 50.730 125.750 ;
        RECT 58.730 125.300 59.330 125.750 ;
        RECT 50.130 125.150 54.080 125.300 ;
        RECT 55.380 125.150 59.330 125.300 ;
        RECT 50.130 124.700 50.730 125.150 ;
        RECT 58.730 124.700 59.330 125.150 ;
        RECT 50.130 124.550 54.080 124.700 ;
        RECT 55.380 124.550 59.330 124.700 ;
        RECT 50.130 124.100 50.730 124.550 ;
        RECT 58.730 124.100 59.330 124.550 ;
        RECT 50.130 123.950 54.080 124.100 ;
        RECT 55.380 123.950 59.330 124.100 ;
        RECT 50.130 123.500 50.730 123.950 ;
        RECT 58.730 123.500 59.330 123.950 ;
        RECT 50.130 123.350 54.080 123.500 ;
        RECT 55.380 123.350 59.330 123.500 ;
        RECT 50.130 122.900 50.730 123.350 ;
        RECT 58.730 122.900 59.330 123.350 ;
        RECT 50.130 122.750 54.080 122.900 ;
        RECT 55.380 122.750 59.330 122.900 ;
        RECT 50.130 122.300 50.730 122.750 ;
        RECT 58.730 122.300 59.330 122.750 ;
        RECT 50.130 122.150 54.080 122.300 ;
        RECT 55.380 122.150 59.330 122.300 ;
        RECT 50.130 122.000 50.730 122.150 ;
        RECT 46.530 121.700 50.730 122.000 ;
        RECT 58.730 122.000 59.330 122.150 ;
        RECT 59.780 122.000 59.930 129.550 ;
        RECT 60.380 122.000 60.530 129.550 ;
        RECT 60.980 122.000 61.130 129.550 ;
        RECT 61.580 122.000 61.730 129.550 ;
        RECT 62.180 122.000 62.330 129.550 ;
        RECT 62.780 122.000 62.930 124.900 ;
        RECT 58.730 121.700 62.930 122.000 ;
        RECT 46.530 121.550 54.080 121.700 ;
        RECT 55.380 121.550 62.930 121.700 ;
        RECT 46.530 121.350 50.730 121.550 ;
        RECT 40.330 121.050 49.130 121.200 ;
        RECT 49.280 121.050 50.730 121.350 ;
        RECT 38.730 120.150 50.730 121.050 ;
        RECT 58.730 121.350 62.930 121.550 ;
        RECT 58.730 121.050 60.180 121.350 ;
        RECT 63.530 121.200 65.930 124.400 ;
        RECT 66.530 122.000 66.680 124.900 ;
        RECT 67.130 122.000 67.280 129.550 ;
        RECT 67.730 122.000 67.880 129.550 ;
        RECT 68.330 122.000 68.480 129.550 ;
        RECT 68.930 122.000 69.080 129.550 ;
        RECT 69.530 122.000 69.680 129.550 ;
        RECT 70.130 129.350 74.080 129.550 ;
        RECT 75.380 129.350 79.330 129.550 ;
        RECT 70.130 128.900 70.730 129.350 ;
        RECT 78.730 128.900 79.330 129.350 ;
        RECT 70.130 128.750 74.080 128.900 ;
        RECT 75.380 128.750 79.330 128.900 ;
        RECT 70.130 128.300 70.730 128.750 ;
        RECT 78.730 128.300 79.330 128.750 ;
        RECT 70.130 128.150 74.080 128.300 ;
        RECT 75.380 128.150 79.330 128.300 ;
        RECT 70.130 127.700 70.730 128.150 ;
        RECT 78.730 127.700 79.330 128.150 ;
        RECT 70.130 127.550 74.080 127.700 ;
        RECT 75.380 127.550 79.330 127.700 ;
        RECT 70.130 127.100 70.730 127.550 ;
        RECT 78.730 127.100 79.330 127.550 ;
        RECT 70.130 126.950 74.080 127.100 ;
        RECT 75.380 126.950 79.330 127.100 ;
        RECT 70.130 126.500 70.730 126.950 ;
        RECT 78.730 126.500 79.330 126.950 ;
        RECT 70.130 126.350 74.080 126.500 ;
        RECT 75.380 126.350 79.330 126.500 ;
        RECT 70.130 125.900 70.730 126.350 ;
        RECT 78.730 125.900 79.330 126.350 ;
        RECT 70.130 125.750 74.080 125.900 ;
        RECT 75.380 125.750 79.330 125.900 ;
        RECT 70.130 125.300 70.730 125.750 ;
        RECT 78.730 125.300 79.330 125.750 ;
        RECT 70.130 125.150 74.080 125.300 ;
        RECT 75.380 125.150 79.330 125.300 ;
        RECT 70.130 124.700 70.730 125.150 ;
        RECT 78.730 124.700 79.330 125.150 ;
        RECT 70.130 124.550 74.080 124.700 ;
        RECT 75.380 124.550 79.330 124.700 ;
        RECT 70.130 124.100 70.730 124.550 ;
        RECT 78.730 124.100 79.330 124.550 ;
        RECT 70.130 123.950 74.080 124.100 ;
        RECT 75.380 123.950 79.330 124.100 ;
        RECT 70.130 123.500 70.730 123.950 ;
        RECT 78.730 123.500 79.330 123.950 ;
        RECT 70.130 123.350 74.080 123.500 ;
        RECT 75.380 123.350 79.330 123.500 ;
        RECT 70.130 122.900 70.730 123.350 ;
        RECT 78.730 122.900 79.330 123.350 ;
        RECT 70.130 122.750 74.080 122.900 ;
        RECT 75.380 122.750 79.330 122.900 ;
        RECT 70.130 122.300 70.730 122.750 ;
        RECT 78.730 122.300 79.330 122.750 ;
        RECT 70.130 122.150 74.080 122.300 ;
        RECT 75.380 122.150 79.330 122.300 ;
        RECT 70.130 122.000 70.730 122.150 ;
        RECT 66.530 121.700 70.730 122.000 ;
        RECT 78.730 122.000 79.330 122.150 ;
        RECT 79.780 122.000 79.930 129.550 ;
        RECT 80.380 122.000 80.530 129.550 ;
        RECT 80.980 122.000 81.130 129.550 ;
        RECT 81.580 122.000 81.730 129.550 ;
        RECT 82.180 122.000 82.330 129.550 ;
        RECT 82.780 122.000 82.930 124.900 ;
        RECT 78.730 121.700 82.930 122.000 ;
        RECT 66.530 121.550 74.080 121.700 ;
        RECT 75.380 121.550 82.930 121.700 ;
        RECT 66.530 121.350 70.730 121.550 ;
        RECT 60.330 121.050 69.130 121.200 ;
        RECT 69.280 121.050 70.730 121.350 ;
        RECT 58.730 120.150 70.730 121.050 ;
        RECT 78.730 121.350 82.930 121.550 ;
        RECT 78.730 121.050 80.180 121.350 ;
        RECT 83.530 121.200 85.930 124.400 ;
        RECT 86.530 122.000 86.680 124.900 ;
        RECT 87.130 122.000 87.280 129.550 ;
        RECT 87.730 122.000 87.880 129.550 ;
        RECT 88.330 122.000 88.480 129.550 ;
        RECT 88.930 122.000 89.080 129.550 ;
        RECT 89.530 122.000 89.680 129.550 ;
        RECT 90.130 129.350 94.080 129.550 ;
        RECT 95.380 129.350 99.330 129.550 ;
        RECT 90.130 128.900 90.730 129.350 ;
        RECT 98.730 128.900 99.330 129.350 ;
        RECT 90.130 128.750 94.080 128.900 ;
        RECT 95.380 128.750 99.330 128.900 ;
        RECT 90.130 128.300 90.730 128.750 ;
        RECT 98.730 128.300 99.330 128.750 ;
        RECT 90.130 128.150 94.080 128.300 ;
        RECT 95.380 128.150 99.330 128.300 ;
        RECT 90.130 127.700 90.730 128.150 ;
        RECT 98.730 127.700 99.330 128.150 ;
        RECT 90.130 127.550 94.080 127.700 ;
        RECT 95.380 127.550 99.330 127.700 ;
        RECT 90.130 127.100 90.730 127.550 ;
        RECT 98.730 127.100 99.330 127.550 ;
        RECT 90.130 126.950 94.080 127.100 ;
        RECT 95.380 126.950 99.330 127.100 ;
        RECT 90.130 126.500 90.730 126.950 ;
        RECT 98.730 126.500 99.330 126.950 ;
        RECT 90.130 126.350 94.080 126.500 ;
        RECT 95.380 126.350 99.330 126.500 ;
        RECT 90.130 125.900 90.730 126.350 ;
        RECT 98.730 125.900 99.330 126.350 ;
        RECT 90.130 125.750 94.080 125.900 ;
        RECT 95.380 125.750 99.330 125.900 ;
        RECT 90.130 125.300 90.730 125.750 ;
        RECT 98.730 125.300 99.330 125.750 ;
        RECT 90.130 125.150 94.080 125.300 ;
        RECT 95.380 125.150 99.330 125.300 ;
        RECT 90.130 124.700 90.730 125.150 ;
        RECT 98.730 124.700 99.330 125.150 ;
        RECT 90.130 124.550 94.080 124.700 ;
        RECT 95.380 124.550 99.330 124.700 ;
        RECT 90.130 124.100 90.730 124.550 ;
        RECT 98.730 124.100 99.330 124.550 ;
        RECT 90.130 123.950 94.080 124.100 ;
        RECT 95.380 123.950 99.330 124.100 ;
        RECT 90.130 123.500 90.730 123.950 ;
        RECT 98.730 123.500 99.330 123.950 ;
        RECT 90.130 123.350 94.080 123.500 ;
        RECT 95.380 123.350 99.330 123.500 ;
        RECT 90.130 122.900 90.730 123.350 ;
        RECT 98.730 122.900 99.330 123.350 ;
        RECT 90.130 122.750 94.080 122.900 ;
        RECT 95.380 122.750 99.330 122.900 ;
        RECT 90.130 122.300 90.730 122.750 ;
        RECT 98.730 122.300 99.330 122.750 ;
        RECT 90.130 122.150 94.080 122.300 ;
        RECT 95.380 122.150 99.330 122.300 ;
        RECT 90.130 122.000 90.730 122.150 ;
        RECT 86.530 121.700 90.730 122.000 ;
        RECT 98.730 122.000 99.330 122.150 ;
        RECT 99.780 122.000 99.930 129.550 ;
        RECT 100.380 122.000 100.530 129.550 ;
        RECT 100.980 122.000 101.130 129.550 ;
        RECT 101.580 122.000 101.730 129.550 ;
        RECT 102.180 122.000 102.330 129.550 ;
        RECT 102.780 122.000 102.930 124.900 ;
        RECT 98.730 121.700 102.930 122.000 ;
        RECT 86.530 121.550 94.080 121.700 ;
        RECT 95.380 121.550 102.930 121.700 ;
        RECT 86.530 121.350 90.730 121.550 ;
        RECT 80.330 121.050 89.130 121.200 ;
        RECT 89.280 121.050 90.730 121.350 ;
        RECT 78.730 120.150 90.730 121.050 ;
        RECT 98.730 121.350 102.930 121.550 ;
        RECT 98.730 121.050 100.180 121.350 ;
        RECT 103.530 121.200 105.930 124.400 ;
        RECT 106.530 122.000 106.680 124.900 ;
        RECT 107.130 122.000 107.280 129.550 ;
        RECT 107.730 122.000 107.880 129.550 ;
        RECT 108.330 122.000 108.480 129.550 ;
        RECT 108.930 122.000 109.080 129.550 ;
        RECT 109.530 122.000 109.680 129.550 ;
        RECT 110.130 129.350 114.080 129.550 ;
        RECT 115.380 129.350 119.330 129.550 ;
        RECT 110.130 128.900 110.730 129.350 ;
        RECT 118.730 128.900 119.330 129.350 ;
        RECT 110.130 128.750 114.080 128.900 ;
        RECT 115.380 128.750 119.330 128.900 ;
        RECT 110.130 128.300 110.730 128.750 ;
        RECT 118.730 128.300 119.330 128.750 ;
        RECT 110.130 128.150 114.080 128.300 ;
        RECT 115.380 128.150 119.330 128.300 ;
        RECT 110.130 127.700 110.730 128.150 ;
        RECT 118.730 127.700 119.330 128.150 ;
        RECT 110.130 127.550 114.080 127.700 ;
        RECT 115.380 127.550 119.330 127.700 ;
        RECT 110.130 127.100 110.730 127.550 ;
        RECT 118.730 127.100 119.330 127.550 ;
        RECT 110.130 126.950 114.080 127.100 ;
        RECT 115.380 126.950 119.330 127.100 ;
        RECT 110.130 126.500 110.730 126.950 ;
        RECT 118.730 126.500 119.330 126.950 ;
        RECT 110.130 126.350 114.080 126.500 ;
        RECT 115.380 126.350 119.330 126.500 ;
        RECT 110.130 125.900 110.730 126.350 ;
        RECT 118.730 125.900 119.330 126.350 ;
        RECT 110.130 125.750 114.080 125.900 ;
        RECT 115.380 125.750 119.330 125.900 ;
        RECT 110.130 125.300 110.730 125.750 ;
        RECT 118.730 125.300 119.330 125.750 ;
        RECT 110.130 125.150 114.080 125.300 ;
        RECT 115.380 125.150 119.330 125.300 ;
        RECT 110.130 124.700 110.730 125.150 ;
        RECT 118.730 124.700 119.330 125.150 ;
        RECT 110.130 124.550 114.080 124.700 ;
        RECT 115.380 124.550 119.330 124.700 ;
        RECT 110.130 124.100 110.730 124.550 ;
        RECT 118.730 124.100 119.330 124.550 ;
        RECT 110.130 123.950 114.080 124.100 ;
        RECT 115.380 123.950 119.330 124.100 ;
        RECT 110.130 123.500 110.730 123.950 ;
        RECT 118.730 123.500 119.330 123.950 ;
        RECT 110.130 123.350 114.080 123.500 ;
        RECT 115.380 123.350 119.330 123.500 ;
        RECT 110.130 122.900 110.730 123.350 ;
        RECT 118.730 122.900 119.330 123.350 ;
        RECT 110.130 122.750 114.080 122.900 ;
        RECT 115.380 122.750 119.330 122.900 ;
        RECT 110.130 122.300 110.730 122.750 ;
        RECT 118.730 122.300 119.330 122.750 ;
        RECT 110.130 122.150 114.080 122.300 ;
        RECT 115.380 122.150 119.330 122.300 ;
        RECT 110.130 122.000 110.730 122.150 ;
        RECT 106.530 121.700 110.730 122.000 ;
        RECT 118.730 122.000 119.330 122.150 ;
        RECT 119.780 122.000 119.930 129.550 ;
        RECT 120.380 122.000 120.530 129.550 ;
        RECT 120.980 122.000 121.130 129.550 ;
        RECT 121.580 122.000 121.730 129.550 ;
        RECT 122.180 122.000 122.330 129.550 ;
        RECT 122.780 122.000 122.930 124.900 ;
        RECT 118.730 121.700 122.930 122.000 ;
        RECT 106.530 121.550 114.080 121.700 ;
        RECT 115.380 121.550 122.930 121.700 ;
        RECT 106.530 121.350 110.730 121.550 ;
        RECT 100.330 121.050 109.130 121.200 ;
        RECT 109.280 121.050 110.730 121.350 ;
        RECT 98.730 120.150 110.730 121.050 ;
        RECT 118.730 121.350 122.930 121.550 ;
        RECT 123.530 122.920 124.730 124.400 ;
        RECT 123.530 121.645 127.140 122.920 ;
        RECT 118.730 121.050 120.180 121.350 ;
        RECT 123.530 121.200 124.730 121.645 ;
        RECT 120.330 121.050 124.730 121.200 ;
        RECT 118.730 120.150 124.730 121.050 ;
        RECT 4.730 119.850 9.130 120.150 ;
        RECT 20.330 119.850 29.130 120.150 ;
        RECT 40.330 119.850 49.130 120.150 ;
        RECT 60.330 119.850 69.130 120.150 ;
        RECT 80.330 119.850 89.130 120.150 ;
        RECT 100.330 119.850 109.130 120.150 ;
        RECT 4.730 118.950 10.730 119.850 ;
        RECT 20.330 119.800 30.730 119.850 ;
        RECT 40.330 119.800 50.730 119.850 ;
        RECT 60.330 119.800 70.730 119.850 ;
        RECT 80.330 119.800 90.730 119.850 ;
        RECT 100.330 119.800 110.730 119.850 ;
        RECT 120.330 119.800 124.730 120.150 ;
        RECT 4.730 118.800 9.130 118.950 ;
        RECT 4.730 118.145 5.930 118.800 ;
        RECT 9.280 118.650 10.730 118.950 ;
        RECT 2.315 116.870 5.930 118.145 ;
        RECT 4.730 115.600 5.930 116.870 ;
        RECT 6.530 118.450 10.730 118.650 ;
        RECT 18.730 118.950 30.730 119.800 ;
        RECT 18.730 118.900 29.130 118.950 ;
        RECT 18.730 118.650 20.180 118.900 ;
        RECT 20.330 118.800 29.130 118.900 ;
        RECT 18.730 118.450 22.930 118.650 ;
        RECT 6.530 118.300 14.080 118.450 ;
        RECT 15.430 118.300 22.930 118.450 ;
        RECT 6.530 118.000 10.730 118.300 ;
        RECT 2.315 113.250 4.315 115.545 ;
        RECT 6.530 115.150 6.680 118.000 ;
        RECT 7.130 110.450 7.280 118.000 ;
        RECT 7.730 110.450 7.880 118.000 ;
        RECT 8.330 110.450 8.480 118.000 ;
        RECT 8.930 110.450 9.080 118.000 ;
        RECT 9.530 110.450 9.680 118.000 ;
        RECT 10.130 117.850 10.730 118.000 ;
        RECT 18.730 118.000 22.930 118.300 ;
        RECT 18.730 117.850 19.330 118.000 ;
        RECT 10.130 117.700 14.080 117.850 ;
        RECT 15.380 117.700 19.330 117.850 ;
        RECT 10.130 117.250 10.730 117.700 ;
        RECT 18.730 117.250 19.330 117.700 ;
        RECT 10.130 117.100 14.080 117.250 ;
        RECT 15.380 117.100 19.330 117.250 ;
        RECT 10.130 116.650 10.730 117.100 ;
        RECT 18.730 116.650 19.330 117.100 ;
        RECT 10.130 116.500 14.080 116.650 ;
        RECT 15.380 116.500 19.330 116.650 ;
        RECT 10.130 116.050 10.730 116.500 ;
        RECT 18.730 116.050 19.330 116.500 ;
        RECT 10.130 115.900 14.080 116.050 ;
        RECT 15.380 115.900 19.330 116.050 ;
        RECT 10.130 115.450 10.730 115.900 ;
        RECT 18.730 115.450 19.330 115.900 ;
        RECT 10.130 115.300 14.080 115.450 ;
        RECT 15.380 115.300 19.330 115.450 ;
        RECT 10.130 114.850 10.730 115.300 ;
        RECT 18.730 114.850 19.330 115.300 ;
        RECT 10.130 114.700 14.080 114.850 ;
        RECT 15.380 114.700 19.330 114.850 ;
        RECT 10.130 114.250 10.730 114.700 ;
        RECT 18.730 114.250 19.330 114.700 ;
        RECT 10.130 114.100 14.080 114.250 ;
        RECT 15.380 114.100 19.330 114.250 ;
        RECT 10.130 113.650 10.730 114.100 ;
        RECT 18.730 113.650 19.330 114.100 ;
        RECT 10.130 113.500 14.080 113.650 ;
        RECT 15.380 113.500 19.330 113.650 ;
        RECT 10.130 113.050 10.730 113.500 ;
        RECT 18.730 113.050 19.330 113.500 ;
        RECT 10.130 112.900 14.080 113.050 ;
        RECT 15.380 112.900 19.330 113.050 ;
        RECT 10.130 112.450 10.730 112.900 ;
        RECT 18.730 112.450 19.330 112.900 ;
        RECT 10.130 112.300 14.080 112.450 ;
        RECT 15.380 112.300 19.330 112.450 ;
        RECT 10.130 111.850 10.730 112.300 ;
        RECT 18.730 111.850 19.330 112.300 ;
        RECT 10.130 111.700 14.080 111.850 ;
        RECT 15.380 111.700 19.330 111.850 ;
        RECT 10.130 111.250 10.730 111.700 ;
        RECT 18.730 111.250 19.330 111.700 ;
        RECT 10.130 111.100 14.080 111.250 ;
        RECT 15.380 111.100 19.330 111.250 ;
        RECT 10.130 110.650 10.730 111.100 ;
        RECT 18.730 110.650 19.330 111.100 ;
        RECT 10.130 110.450 14.080 110.650 ;
        RECT 15.380 110.450 19.330 110.650 ;
        RECT 19.780 110.450 19.930 118.000 ;
        RECT 20.380 110.450 20.530 118.000 ;
        RECT 20.980 110.450 21.130 118.000 ;
        RECT 21.580 110.450 21.730 118.000 ;
        RECT 22.180 110.450 22.330 118.000 ;
        RECT 22.780 115.150 22.930 118.000 ;
        RECT 23.530 115.600 25.930 118.800 ;
        RECT 29.280 118.650 30.730 118.950 ;
        RECT 26.530 118.450 30.730 118.650 ;
        RECT 38.730 118.950 50.730 119.800 ;
        RECT 38.730 118.900 49.130 118.950 ;
        RECT 38.730 118.650 40.180 118.900 ;
        RECT 40.330 118.800 49.130 118.900 ;
        RECT 38.730 118.450 42.930 118.650 ;
        RECT 26.530 118.300 34.080 118.450 ;
        RECT 35.430 118.300 42.930 118.450 ;
        RECT 26.530 118.000 30.730 118.300 ;
        RECT 26.530 115.150 26.680 118.000 ;
        RECT 27.130 110.450 27.280 118.000 ;
        RECT 27.730 110.450 27.880 118.000 ;
        RECT 28.330 110.450 28.480 118.000 ;
        RECT 28.930 110.450 29.080 118.000 ;
        RECT 29.530 110.450 29.680 118.000 ;
        RECT 30.130 117.850 30.730 118.000 ;
        RECT 38.730 118.000 42.930 118.300 ;
        RECT 38.730 117.850 39.330 118.000 ;
        RECT 30.130 117.700 34.080 117.850 ;
        RECT 35.380 117.700 39.330 117.850 ;
        RECT 30.130 117.250 30.730 117.700 ;
        RECT 38.730 117.250 39.330 117.700 ;
        RECT 30.130 117.100 34.080 117.250 ;
        RECT 35.380 117.100 39.330 117.250 ;
        RECT 30.130 116.650 30.730 117.100 ;
        RECT 38.730 116.650 39.330 117.100 ;
        RECT 30.130 116.500 34.080 116.650 ;
        RECT 35.380 116.500 39.330 116.650 ;
        RECT 30.130 116.050 30.730 116.500 ;
        RECT 38.730 116.050 39.330 116.500 ;
        RECT 30.130 115.900 34.080 116.050 ;
        RECT 35.380 115.900 39.330 116.050 ;
        RECT 30.130 115.450 30.730 115.900 ;
        RECT 38.730 115.450 39.330 115.900 ;
        RECT 30.130 115.300 34.080 115.450 ;
        RECT 35.380 115.300 39.330 115.450 ;
        RECT 30.130 114.850 30.730 115.300 ;
        RECT 38.730 114.850 39.330 115.300 ;
        RECT 30.130 114.700 34.080 114.850 ;
        RECT 35.380 114.700 39.330 114.850 ;
        RECT 30.130 114.250 30.730 114.700 ;
        RECT 38.730 114.250 39.330 114.700 ;
        RECT 30.130 114.100 34.080 114.250 ;
        RECT 35.380 114.100 39.330 114.250 ;
        RECT 30.130 113.650 30.730 114.100 ;
        RECT 38.730 113.650 39.330 114.100 ;
        RECT 30.130 113.500 34.080 113.650 ;
        RECT 35.380 113.500 39.330 113.650 ;
        RECT 30.130 113.050 30.730 113.500 ;
        RECT 38.730 113.050 39.330 113.500 ;
        RECT 30.130 112.900 34.080 113.050 ;
        RECT 35.380 112.900 39.330 113.050 ;
        RECT 30.130 112.450 30.730 112.900 ;
        RECT 38.730 112.450 39.330 112.900 ;
        RECT 30.130 112.300 34.080 112.450 ;
        RECT 35.380 112.300 39.330 112.450 ;
        RECT 30.130 111.850 30.730 112.300 ;
        RECT 38.730 111.850 39.330 112.300 ;
        RECT 30.130 111.700 34.080 111.850 ;
        RECT 35.380 111.700 39.330 111.850 ;
        RECT 30.130 111.250 30.730 111.700 ;
        RECT 38.730 111.250 39.330 111.700 ;
        RECT 30.130 111.100 34.080 111.250 ;
        RECT 35.380 111.100 39.330 111.250 ;
        RECT 30.130 110.650 30.730 111.100 ;
        RECT 38.730 110.650 39.330 111.100 ;
        RECT 30.130 110.450 34.080 110.650 ;
        RECT 35.380 110.450 39.330 110.650 ;
        RECT 39.780 110.450 39.930 118.000 ;
        RECT 40.380 110.450 40.530 118.000 ;
        RECT 40.980 110.450 41.130 118.000 ;
        RECT 41.580 110.450 41.730 118.000 ;
        RECT 42.180 110.450 42.330 118.000 ;
        RECT 42.780 115.150 42.930 118.000 ;
        RECT 43.530 115.600 45.930 118.800 ;
        RECT 49.280 118.650 50.730 118.950 ;
        RECT 46.530 118.450 50.730 118.650 ;
        RECT 58.730 118.950 70.730 119.800 ;
        RECT 58.730 118.900 69.130 118.950 ;
        RECT 58.730 118.650 60.180 118.900 ;
        RECT 60.330 118.800 69.130 118.900 ;
        RECT 58.730 118.450 62.930 118.650 ;
        RECT 46.530 118.300 54.080 118.450 ;
        RECT 55.430 118.300 62.930 118.450 ;
        RECT 46.530 118.000 50.730 118.300 ;
        RECT 46.530 115.150 46.680 118.000 ;
        RECT 47.130 110.450 47.280 118.000 ;
        RECT 47.730 110.450 47.880 118.000 ;
        RECT 48.330 110.450 48.480 118.000 ;
        RECT 48.930 110.450 49.080 118.000 ;
        RECT 49.530 110.450 49.680 118.000 ;
        RECT 50.130 117.850 50.730 118.000 ;
        RECT 58.730 118.000 62.930 118.300 ;
        RECT 58.730 117.850 59.330 118.000 ;
        RECT 50.130 117.700 54.080 117.850 ;
        RECT 55.380 117.700 59.330 117.850 ;
        RECT 50.130 117.250 50.730 117.700 ;
        RECT 58.730 117.250 59.330 117.700 ;
        RECT 50.130 117.100 54.080 117.250 ;
        RECT 55.380 117.100 59.330 117.250 ;
        RECT 50.130 116.650 50.730 117.100 ;
        RECT 58.730 116.650 59.330 117.100 ;
        RECT 50.130 116.500 54.080 116.650 ;
        RECT 55.380 116.500 59.330 116.650 ;
        RECT 50.130 116.050 50.730 116.500 ;
        RECT 58.730 116.050 59.330 116.500 ;
        RECT 50.130 115.900 54.080 116.050 ;
        RECT 55.380 115.900 59.330 116.050 ;
        RECT 50.130 115.450 50.730 115.900 ;
        RECT 58.730 115.450 59.330 115.900 ;
        RECT 50.130 115.300 54.080 115.450 ;
        RECT 55.380 115.300 59.330 115.450 ;
        RECT 50.130 114.850 50.730 115.300 ;
        RECT 58.730 114.850 59.330 115.300 ;
        RECT 50.130 114.700 54.080 114.850 ;
        RECT 55.380 114.700 59.330 114.850 ;
        RECT 50.130 114.250 50.730 114.700 ;
        RECT 58.730 114.250 59.330 114.700 ;
        RECT 50.130 114.100 54.080 114.250 ;
        RECT 55.380 114.100 59.330 114.250 ;
        RECT 50.130 113.650 50.730 114.100 ;
        RECT 58.730 113.650 59.330 114.100 ;
        RECT 50.130 113.500 54.080 113.650 ;
        RECT 55.380 113.500 59.330 113.650 ;
        RECT 50.130 113.050 50.730 113.500 ;
        RECT 58.730 113.050 59.330 113.500 ;
        RECT 50.130 112.900 54.080 113.050 ;
        RECT 55.380 112.900 59.330 113.050 ;
        RECT 50.130 112.450 50.730 112.900 ;
        RECT 58.730 112.450 59.330 112.900 ;
        RECT 50.130 112.300 54.080 112.450 ;
        RECT 55.380 112.300 59.330 112.450 ;
        RECT 50.130 111.850 50.730 112.300 ;
        RECT 58.730 111.850 59.330 112.300 ;
        RECT 50.130 111.700 54.080 111.850 ;
        RECT 55.380 111.700 59.330 111.850 ;
        RECT 50.130 111.250 50.730 111.700 ;
        RECT 58.730 111.250 59.330 111.700 ;
        RECT 50.130 111.100 54.080 111.250 ;
        RECT 55.380 111.100 59.330 111.250 ;
        RECT 50.130 110.650 50.730 111.100 ;
        RECT 58.730 110.650 59.330 111.100 ;
        RECT 50.130 110.450 54.080 110.650 ;
        RECT 55.380 110.450 59.330 110.650 ;
        RECT 59.780 110.450 59.930 118.000 ;
        RECT 60.380 110.450 60.530 118.000 ;
        RECT 60.980 110.450 61.130 118.000 ;
        RECT 61.580 110.450 61.730 118.000 ;
        RECT 62.180 110.450 62.330 118.000 ;
        RECT 62.780 115.150 62.930 118.000 ;
        RECT 63.530 115.600 65.930 118.800 ;
        RECT 69.280 118.650 70.730 118.950 ;
        RECT 66.530 118.450 70.730 118.650 ;
        RECT 78.730 118.950 90.730 119.800 ;
        RECT 78.730 118.900 89.130 118.950 ;
        RECT 78.730 118.650 80.180 118.900 ;
        RECT 80.330 118.800 89.130 118.900 ;
        RECT 78.730 118.450 82.930 118.650 ;
        RECT 66.530 118.300 74.080 118.450 ;
        RECT 75.430 118.300 82.930 118.450 ;
        RECT 66.530 118.000 70.730 118.300 ;
        RECT 66.530 115.150 66.680 118.000 ;
        RECT 67.130 110.450 67.280 118.000 ;
        RECT 67.730 110.450 67.880 118.000 ;
        RECT 68.330 110.450 68.480 118.000 ;
        RECT 68.930 110.450 69.080 118.000 ;
        RECT 69.530 110.450 69.680 118.000 ;
        RECT 70.130 117.850 70.730 118.000 ;
        RECT 78.730 118.000 82.930 118.300 ;
        RECT 78.730 117.850 79.330 118.000 ;
        RECT 70.130 117.700 74.080 117.850 ;
        RECT 75.380 117.700 79.330 117.850 ;
        RECT 70.130 117.250 70.730 117.700 ;
        RECT 78.730 117.250 79.330 117.700 ;
        RECT 70.130 117.100 74.080 117.250 ;
        RECT 75.380 117.100 79.330 117.250 ;
        RECT 70.130 116.650 70.730 117.100 ;
        RECT 78.730 116.650 79.330 117.100 ;
        RECT 70.130 116.500 74.080 116.650 ;
        RECT 75.380 116.500 79.330 116.650 ;
        RECT 70.130 116.050 70.730 116.500 ;
        RECT 78.730 116.050 79.330 116.500 ;
        RECT 70.130 115.900 74.080 116.050 ;
        RECT 75.380 115.900 79.330 116.050 ;
        RECT 70.130 115.450 70.730 115.900 ;
        RECT 78.730 115.450 79.330 115.900 ;
        RECT 70.130 115.300 74.080 115.450 ;
        RECT 75.380 115.300 79.330 115.450 ;
        RECT 70.130 114.850 70.730 115.300 ;
        RECT 78.730 114.850 79.330 115.300 ;
        RECT 70.130 114.700 74.080 114.850 ;
        RECT 75.380 114.700 79.330 114.850 ;
        RECT 70.130 114.250 70.730 114.700 ;
        RECT 78.730 114.250 79.330 114.700 ;
        RECT 70.130 114.100 74.080 114.250 ;
        RECT 75.380 114.100 79.330 114.250 ;
        RECT 70.130 113.650 70.730 114.100 ;
        RECT 78.730 113.650 79.330 114.100 ;
        RECT 70.130 113.500 74.080 113.650 ;
        RECT 75.380 113.500 79.330 113.650 ;
        RECT 70.130 113.050 70.730 113.500 ;
        RECT 78.730 113.050 79.330 113.500 ;
        RECT 70.130 112.900 74.080 113.050 ;
        RECT 75.380 112.900 79.330 113.050 ;
        RECT 70.130 112.450 70.730 112.900 ;
        RECT 78.730 112.450 79.330 112.900 ;
        RECT 70.130 112.300 74.080 112.450 ;
        RECT 75.380 112.300 79.330 112.450 ;
        RECT 70.130 111.850 70.730 112.300 ;
        RECT 78.730 111.850 79.330 112.300 ;
        RECT 70.130 111.700 74.080 111.850 ;
        RECT 75.380 111.700 79.330 111.850 ;
        RECT 70.130 111.250 70.730 111.700 ;
        RECT 78.730 111.250 79.330 111.700 ;
        RECT 70.130 111.100 74.080 111.250 ;
        RECT 75.380 111.100 79.330 111.250 ;
        RECT 70.130 110.650 70.730 111.100 ;
        RECT 78.730 110.650 79.330 111.100 ;
        RECT 70.130 110.450 74.080 110.650 ;
        RECT 75.380 110.450 79.330 110.650 ;
        RECT 79.780 110.450 79.930 118.000 ;
        RECT 80.380 110.450 80.530 118.000 ;
        RECT 80.980 110.450 81.130 118.000 ;
        RECT 81.580 110.450 81.730 118.000 ;
        RECT 82.180 110.450 82.330 118.000 ;
        RECT 82.780 115.150 82.930 118.000 ;
        RECT 83.530 115.600 85.930 118.800 ;
        RECT 89.280 118.650 90.730 118.950 ;
        RECT 86.530 118.450 90.730 118.650 ;
        RECT 98.730 118.950 110.730 119.800 ;
        RECT 98.730 118.900 109.130 118.950 ;
        RECT 98.730 118.650 100.180 118.900 ;
        RECT 100.330 118.800 109.130 118.900 ;
        RECT 98.730 118.450 102.930 118.650 ;
        RECT 86.530 118.300 94.080 118.450 ;
        RECT 95.430 118.300 102.930 118.450 ;
        RECT 86.530 118.000 90.730 118.300 ;
        RECT 86.530 115.150 86.680 118.000 ;
        RECT 87.130 110.450 87.280 118.000 ;
        RECT 87.730 110.450 87.880 118.000 ;
        RECT 88.330 110.450 88.480 118.000 ;
        RECT 88.930 110.450 89.080 118.000 ;
        RECT 89.530 110.450 89.680 118.000 ;
        RECT 90.130 117.850 90.730 118.000 ;
        RECT 98.730 118.000 102.930 118.300 ;
        RECT 98.730 117.850 99.330 118.000 ;
        RECT 90.130 117.700 94.080 117.850 ;
        RECT 95.380 117.700 99.330 117.850 ;
        RECT 90.130 117.250 90.730 117.700 ;
        RECT 98.730 117.250 99.330 117.700 ;
        RECT 90.130 117.100 94.080 117.250 ;
        RECT 95.380 117.100 99.330 117.250 ;
        RECT 90.130 116.650 90.730 117.100 ;
        RECT 98.730 116.650 99.330 117.100 ;
        RECT 90.130 116.500 94.080 116.650 ;
        RECT 95.380 116.500 99.330 116.650 ;
        RECT 90.130 116.050 90.730 116.500 ;
        RECT 98.730 116.050 99.330 116.500 ;
        RECT 90.130 115.900 94.080 116.050 ;
        RECT 95.380 115.900 99.330 116.050 ;
        RECT 90.130 115.450 90.730 115.900 ;
        RECT 98.730 115.450 99.330 115.900 ;
        RECT 90.130 115.300 94.080 115.450 ;
        RECT 95.380 115.300 99.330 115.450 ;
        RECT 90.130 114.850 90.730 115.300 ;
        RECT 98.730 114.850 99.330 115.300 ;
        RECT 90.130 114.700 94.080 114.850 ;
        RECT 95.380 114.700 99.330 114.850 ;
        RECT 90.130 114.250 90.730 114.700 ;
        RECT 98.730 114.250 99.330 114.700 ;
        RECT 90.130 114.100 94.080 114.250 ;
        RECT 95.380 114.100 99.330 114.250 ;
        RECT 90.130 113.650 90.730 114.100 ;
        RECT 98.730 113.650 99.330 114.100 ;
        RECT 90.130 113.500 94.080 113.650 ;
        RECT 95.380 113.500 99.330 113.650 ;
        RECT 90.130 113.050 90.730 113.500 ;
        RECT 98.730 113.050 99.330 113.500 ;
        RECT 90.130 112.900 94.080 113.050 ;
        RECT 95.380 112.900 99.330 113.050 ;
        RECT 90.130 112.450 90.730 112.900 ;
        RECT 98.730 112.450 99.330 112.900 ;
        RECT 90.130 112.300 94.080 112.450 ;
        RECT 95.380 112.300 99.330 112.450 ;
        RECT 90.130 111.850 90.730 112.300 ;
        RECT 98.730 111.850 99.330 112.300 ;
        RECT 90.130 111.700 94.080 111.850 ;
        RECT 95.380 111.700 99.330 111.850 ;
        RECT 90.130 111.250 90.730 111.700 ;
        RECT 98.730 111.250 99.330 111.700 ;
        RECT 90.130 111.100 94.080 111.250 ;
        RECT 95.380 111.100 99.330 111.250 ;
        RECT 90.130 110.650 90.730 111.100 ;
        RECT 98.730 110.650 99.330 111.100 ;
        RECT 90.130 110.450 94.080 110.650 ;
        RECT 95.380 110.450 99.330 110.650 ;
        RECT 99.780 110.450 99.930 118.000 ;
        RECT 100.380 110.450 100.530 118.000 ;
        RECT 100.980 110.450 101.130 118.000 ;
        RECT 101.580 110.450 101.730 118.000 ;
        RECT 102.180 110.450 102.330 118.000 ;
        RECT 102.780 115.150 102.930 118.000 ;
        RECT 103.530 115.600 105.930 118.800 ;
        RECT 109.280 118.650 110.730 118.950 ;
        RECT 106.530 118.450 110.730 118.650 ;
        RECT 118.730 118.900 124.730 119.800 ;
        RECT 118.730 118.650 120.180 118.900 ;
        RECT 120.330 118.800 124.730 118.900 ;
        RECT 118.730 118.450 122.930 118.650 ;
        RECT 106.530 118.300 114.080 118.450 ;
        RECT 115.430 118.300 122.930 118.450 ;
        RECT 106.530 118.000 110.730 118.300 ;
        RECT 106.530 115.150 106.680 118.000 ;
        RECT 107.130 110.450 107.280 118.000 ;
        RECT 107.730 110.450 107.880 118.000 ;
        RECT 108.330 110.450 108.480 118.000 ;
        RECT 108.930 110.450 109.080 118.000 ;
        RECT 109.530 110.450 109.680 118.000 ;
        RECT 110.130 117.850 110.730 118.000 ;
        RECT 118.730 118.000 122.930 118.300 ;
        RECT 118.730 117.850 119.330 118.000 ;
        RECT 110.130 117.700 114.080 117.850 ;
        RECT 115.380 117.700 119.330 117.850 ;
        RECT 110.130 117.250 110.730 117.700 ;
        RECT 118.730 117.250 119.330 117.700 ;
        RECT 110.130 117.100 114.080 117.250 ;
        RECT 115.380 117.100 119.330 117.250 ;
        RECT 110.130 116.650 110.730 117.100 ;
        RECT 118.730 116.650 119.330 117.100 ;
        RECT 110.130 116.500 114.080 116.650 ;
        RECT 115.380 116.500 119.330 116.650 ;
        RECT 110.130 116.050 110.730 116.500 ;
        RECT 118.730 116.050 119.330 116.500 ;
        RECT 110.130 115.900 114.080 116.050 ;
        RECT 115.380 115.900 119.330 116.050 ;
        RECT 110.130 115.450 110.730 115.900 ;
        RECT 118.730 115.450 119.330 115.900 ;
        RECT 110.130 115.300 114.080 115.450 ;
        RECT 115.380 115.300 119.330 115.450 ;
        RECT 110.130 114.850 110.730 115.300 ;
        RECT 118.730 114.850 119.330 115.300 ;
        RECT 110.130 114.700 114.080 114.850 ;
        RECT 115.380 114.700 119.330 114.850 ;
        RECT 110.130 114.250 110.730 114.700 ;
        RECT 118.730 114.250 119.330 114.700 ;
        RECT 110.130 114.100 114.080 114.250 ;
        RECT 115.380 114.100 119.330 114.250 ;
        RECT 110.130 113.650 110.730 114.100 ;
        RECT 118.730 113.650 119.330 114.100 ;
        RECT 110.130 113.500 114.080 113.650 ;
        RECT 115.380 113.500 119.330 113.650 ;
        RECT 110.130 113.050 110.730 113.500 ;
        RECT 118.730 113.050 119.330 113.500 ;
        RECT 110.130 112.900 114.080 113.050 ;
        RECT 115.380 112.900 119.330 113.050 ;
        RECT 110.130 112.450 110.730 112.900 ;
        RECT 118.730 112.450 119.330 112.900 ;
        RECT 110.130 112.300 114.080 112.450 ;
        RECT 115.380 112.300 119.330 112.450 ;
        RECT 110.130 111.850 110.730 112.300 ;
        RECT 118.730 111.850 119.330 112.300 ;
        RECT 110.130 111.700 114.080 111.850 ;
        RECT 115.380 111.700 119.330 111.850 ;
        RECT 110.130 111.250 110.730 111.700 ;
        RECT 118.730 111.250 119.330 111.700 ;
        RECT 110.130 111.100 114.080 111.250 ;
        RECT 115.380 111.100 119.330 111.250 ;
        RECT 110.130 110.650 110.730 111.100 ;
        RECT 118.730 110.650 119.330 111.100 ;
        RECT 110.130 110.450 114.080 110.650 ;
        RECT 115.380 110.450 119.330 110.650 ;
        RECT 119.780 110.450 119.930 118.000 ;
        RECT 120.380 110.450 120.530 118.000 ;
        RECT 120.980 110.450 121.130 118.000 ;
        RECT 121.580 110.450 121.730 118.000 ;
        RECT 122.180 110.450 122.330 118.000 ;
        RECT 122.780 115.150 122.930 118.000 ;
        RECT 123.530 117.335 124.730 118.800 ;
        RECT 123.530 116.060 127.135 117.335 ;
        RECT 123.530 115.600 124.730 116.060 ;
        RECT 2.315 104.450 4.315 106.745 ;
        RECT 4.730 103.255 5.930 104.400 ;
        RECT 2.315 101.980 5.930 103.255 ;
        RECT 4.730 101.200 5.930 101.980 ;
        RECT 6.530 102.000 6.680 104.900 ;
        RECT 7.130 102.000 7.280 109.550 ;
        RECT 7.730 102.000 7.880 109.550 ;
        RECT 8.330 102.000 8.480 109.550 ;
        RECT 8.930 102.000 9.080 109.550 ;
        RECT 9.530 102.000 9.680 109.550 ;
        RECT 10.130 109.350 14.080 109.550 ;
        RECT 15.380 109.350 19.330 109.550 ;
        RECT 10.130 108.900 10.730 109.350 ;
        RECT 18.730 108.900 19.330 109.350 ;
        RECT 10.130 108.750 14.080 108.900 ;
        RECT 15.380 108.750 19.330 108.900 ;
        RECT 10.130 108.300 10.730 108.750 ;
        RECT 18.730 108.300 19.330 108.750 ;
        RECT 10.130 108.150 14.080 108.300 ;
        RECT 15.380 108.150 19.330 108.300 ;
        RECT 10.130 107.700 10.730 108.150 ;
        RECT 18.730 107.700 19.330 108.150 ;
        RECT 10.130 107.550 14.080 107.700 ;
        RECT 15.380 107.550 19.330 107.700 ;
        RECT 10.130 107.100 10.730 107.550 ;
        RECT 18.730 107.100 19.330 107.550 ;
        RECT 10.130 106.950 14.080 107.100 ;
        RECT 15.380 106.950 19.330 107.100 ;
        RECT 10.130 106.500 10.730 106.950 ;
        RECT 18.730 106.500 19.330 106.950 ;
        RECT 10.130 106.350 14.080 106.500 ;
        RECT 15.380 106.350 19.330 106.500 ;
        RECT 10.130 105.900 10.730 106.350 ;
        RECT 18.730 105.900 19.330 106.350 ;
        RECT 10.130 105.750 14.080 105.900 ;
        RECT 15.380 105.750 19.330 105.900 ;
        RECT 10.130 105.300 10.730 105.750 ;
        RECT 18.730 105.300 19.330 105.750 ;
        RECT 10.130 105.150 14.080 105.300 ;
        RECT 15.380 105.150 19.330 105.300 ;
        RECT 10.130 104.700 10.730 105.150 ;
        RECT 18.730 104.700 19.330 105.150 ;
        RECT 10.130 104.550 14.080 104.700 ;
        RECT 15.380 104.550 19.330 104.700 ;
        RECT 10.130 104.100 10.730 104.550 ;
        RECT 18.730 104.100 19.330 104.550 ;
        RECT 10.130 103.950 14.080 104.100 ;
        RECT 15.380 103.950 19.330 104.100 ;
        RECT 10.130 103.500 10.730 103.950 ;
        RECT 18.730 103.500 19.330 103.950 ;
        RECT 10.130 103.350 14.080 103.500 ;
        RECT 15.380 103.350 19.330 103.500 ;
        RECT 10.130 102.900 10.730 103.350 ;
        RECT 18.730 102.900 19.330 103.350 ;
        RECT 10.130 102.750 14.080 102.900 ;
        RECT 15.380 102.750 19.330 102.900 ;
        RECT 10.130 102.300 10.730 102.750 ;
        RECT 18.730 102.300 19.330 102.750 ;
        RECT 10.130 102.150 14.080 102.300 ;
        RECT 15.380 102.150 19.330 102.300 ;
        RECT 10.130 102.000 10.730 102.150 ;
        RECT 6.530 101.700 10.730 102.000 ;
        RECT 18.730 102.000 19.330 102.150 ;
        RECT 19.780 102.000 19.930 109.550 ;
        RECT 20.380 102.000 20.530 109.550 ;
        RECT 20.980 102.000 21.130 109.550 ;
        RECT 21.580 102.000 21.730 109.550 ;
        RECT 22.180 102.000 22.330 109.550 ;
        RECT 22.780 102.000 22.930 104.900 ;
        RECT 18.730 101.700 22.930 102.000 ;
        RECT 6.530 101.550 14.080 101.700 ;
        RECT 15.380 101.550 22.930 101.700 ;
        RECT 6.530 101.350 10.730 101.550 ;
        RECT 4.730 101.050 9.130 101.200 ;
        RECT 9.280 101.050 10.730 101.350 ;
        RECT 4.730 100.150 10.730 101.050 ;
        RECT 18.730 101.350 22.930 101.550 ;
        RECT 18.730 101.050 20.180 101.350 ;
        RECT 23.530 101.200 25.930 104.400 ;
        RECT 26.530 102.000 26.680 104.900 ;
        RECT 27.130 102.000 27.280 109.550 ;
        RECT 27.730 102.000 27.880 109.550 ;
        RECT 28.330 102.000 28.480 109.550 ;
        RECT 28.930 102.000 29.080 109.550 ;
        RECT 29.530 102.000 29.680 109.550 ;
        RECT 30.130 109.350 34.080 109.550 ;
        RECT 35.380 109.350 39.330 109.550 ;
        RECT 30.130 108.900 30.730 109.350 ;
        RECT 38.730 108.900 39.330 109.350 ;
        RECT 30.130 108.750 34.080 108.900 ;
        RECT 35.380 108.750 39.330 108.900 ;
        RECT 30.130 108.300 30.730 108.750 ;
        RECT 38.730 108.300 39.330 108.750 ;
        RECT 30.130 108.150 34.080 108.300 ;
        RECT 35.380 108.150 39.330 108.300 ;
        RECT 30.130 107.700 30.730 108.150 ;
        RECT 38.730 107.700 39.330 108.150 ;
        RECT 30.130 107.550 34.080 107.700 ;
        RECT 35.380 107.550 39.330 107.700 ;
        RECT 30.130 107.100 30.730 107.550 ;
        RECT 38.730 107.100 39.330 107.550 ;
        RECT 30.130 106.950 34.080 107.100 ;
        RECT 35.380 106.950 39.330 107.100 ;
        RECT 30.130 106.500 30.730 106.950 ;
        RECT 38.730 106.500 39.330 106.950 ;
        RECT 30.130 106.350 34.080 106.500 ;
        RECT 35.380 106.350 39.330 106.500 ;
        RECT 30.130 105.900 30.730 106.350 ;
        RECT 38.730 105.900 39.330 106.350 ;
        RECT 30.130 105.750 34.080 105.900 ;
        RECT 35.380 105.750 39.330 105.900 ;
        RECT 30.130 105.300 30.730 105.750 ;
        RECT 38.730 105.300 39.330 105.750 ;
        RECT 30.130 105.150 34.080 105.300 ;
        RECT 35.380 105.150 39.330 105.300 ;
        RECT 30.130 104.700 30.730 105.150 ;
        RECT 38.730 104.700 39.330 105.150 ;
        RECT 30.130 104.550 34.080 104.700 ;
        RECT 35.380 104.550 39.330 104.700 ;
        RECT 30.130 104.100 30.730 104.550 ;
        RECT 38.730 104.100 39.330 104.550 ;
        RECT 30.130 103.950 34.080 104.100 ;
        RECT 35.380 103.950 39.330 104.100 ;
        RECT 30.130 103.500 30.730 103.950 ;
        RECT 38.730 103.500 39.330 103.950 ;
        RECT 30.130 103.350 34.080 103.500 ;
        RECT 35.380 103.350 39.330 103.500 ;
        RECT 30.130 102.900 30.730 103.350 ;
        RECT 38.730 102.900 39.330 103.350 ;
        RECT 30.130 102.750 34.080 102.900 ;
        RECT 35.380 102.750 39.330 102.900 ;
        RECT 30.130 102.300 30.730 102.750 ;
        RECT 38.730 102.300 39.330 102.750 ;
        RECT 30.130 102.150 34.080 102.300 ;
        RECT 35.380 102.150 39.330 102.300 ;
        RECT 30.130 102.000 30.730 102.150 ;
        RECT 26.530 101.700 30.730 102.000 ;
        RECT 38.730 102.000 39.330 102.150 ;
        RECT 39.780 102.000 39.930 109.550 ;
        RECT 40.380 102.000 40.530 109.550 ;
        RECT 40.980 102.000 41.130 109.550 ;
        RECT 41.580 102.000 41.730 109.550 ;
        RECT 42.180 102.000 42.330 109.550 ;
        RECT 42.780 102.000 42.930 104.900 ;
        RECT 38.730 101.700 42.930 102.000 ;
        RECT 26.530 101.550 34.080 101.700 ;
        RECT 35.380 101.550 42.930 101.700 ;
        RECT 26.530 101.350 30.730 101.550 ;
        RECT 20.330 101.050 29.130 101.200 ;
        RECT 29.280 101.050 30.730 101.350 ;
        RECT 18.730 100.150 30.730 101.050 ;
        RECT 38.730 101.350 42.930 101.550 ;
        RECT 38.730 101.050 40.180 101.350 ;
        RECT 43.530 101.200 45.930 104.400 ;
        RECT 46.530 102.000 46.680 104.900 ;
        RECT 47.130 102.000 47.280 109.550 ;
        RECT 47.730 102.000 47.880 109.550 ;
        RECT 48.330 102.000 48.480 109.550 ;
        RECT 48.930 102.000 49.080 109.550 ;
        RECT 49.530 102.000 49.680 109.550 ;
        RECT 50.130 109.350 54.080 109.550 ;
        RECT 55.380 109.350 59.330 109.550 ;
        RECT 50.130 108.900 50.730 109.350 ;
        RECT 58.730 108.900 59.330 109.350 ;
        RECT 50.130 108.750 54.080 108.900 ;
        RECT 55.380 108.750 59.330 108.900 ;
        RECT 50.130 108.300 50.730 108.750 ;
        RECT 58.730 108.300 59.330 108.750 ;
        RECT 50.130 108.150 54.080 108.300 ;
        RECT 55.380 108.150 59.330 108.300 ;
        RECT 50.130 107.700 50.730 108.150 ;
        RECT 58.730 107.700 59.330 108.150 ;
        RECT 50.130 107.550 54.080 107.700 ;
        RECT 55.380 107.550 59.330 107.700 ;
        RECT 50.130 107.100 50.730 107.550 ;
        RECT 58.730 107.100 59.330 107.550 ;
        RECT 50.130 106.950 54.080 107.100 ;
        RECT 55.380 106.950 59.330 107.100 ;
        RECT 50.130 106.500 50.730 106.950 ;
        RECT 58.730 106.500 59.330 106.950 ;
        RECT 50.130 106.350 54.080 106.500 ;
        RECT 55.380 106.350 59.330 106.500 ;
        RECT 50.130 105.900 50.730 106.350 ;
        RECT 58.730 105.900 59.330 106.350 ;
        RECT 50.130 105.750 54.080 105.900 ;
        RECT 55.380 105.750 59.330 105.900 ;
        RECT 50.130 105.300 50.730 105.750 ;
        RECT 58.730 105.300 59.330 105.750 ;
        RECT 50.130 105.150 54.080 105.300 ;
        RECT 55.380 105.150 59.330 105.300 ;
        RECT 50.130 104.700 50.730 105.150 ;
        RECT 58.730 104.700 59.330 105.150 ;
        RECT 50.130 104.550 54.080 104.700 ;
        RECT 55.380 104.550 59.330 104.700 ;
        RECT 50.130 104.100 50.730 104.550 ;
        RECT 58.730 104.100 59.330 104.550 ;
        RECT 50.130 103.950 54.080 104.100 ;
        RECT 55.380 103.950 59.330 104.100 ;
        RECT 50.130 103.500 50.730 103.950 ;
        RECT 58.730 103.500 59.330 103.950 ;
        RECT 50.130 103.350 54.080 103.500 ;
        RECT 55.380 103.350 59.330 103.500 ;
        RECT 50.130 102.900 50.730 103.350 ;
        RECT 58.730 102.900 59.330 103.350 ;
        RECT 50.130 102.750 54.080 102.900 ;
        RECT 55.380 102.750 59.330 102.900 ;
        RECT 50.130 102.300 50.730 102.750 ;
        RECT 58.730 102.300 59.330 102.750 ;
        RECT 50.130 102.150 54.080 102.300 ;
        RECT 55.380 102.150 59.330 102.300 ;
        RECT 50.130 102.000 50.730 102.150 ;
        RECT 46.530 101.700 50.730 102.000 ;
        RECT 58.730 102.000 59.330 102.150 ;
        RECT 59.780 102.000 59.930 109.550 ;
        RECT 60.380 102.000 60.530 109.550 ;
        RECT 60.980 102.000 61.130 109.550 ;
        RECT 61.580 102.000 61.730 109.550 ;
        RECT 62.180 102.000 62.330 109.550 ;
        RECT 62.780 102.000 62.930 104.900 ;
        RECT 58.730 101.700 62.930 102.000 ;
        RECT 46.530 101.550 54.080 101.700 ;
        RECT 55.380 101.550 62.930 101.700 ;
        RECT 46.530 101.350 50.730 101.550 ;
        RECT 40.330 101.050 49.130 101.200 ;
        RECT 49.280 101.050 50.730 101.350 ;
        RECT 38.730 100.150 50.730 101.050 ;
        RECT 58.730 101.350 62.930 101.550 ;
        RECT 58.730 101.050 60.180 101.350 ;
        RECT 63.530 101.200 65.930 104.400 ;
        RECT 66.530 102.000 66.680 104.900 ;
        RECT 67.130 102.000 67.280 109.550 ;
        RECT 67.730 102.000 67.880 109.550 ;
        RECT 68.330 102.000 68.480 109.550 ;
        RECT 68.930 102.000 69.080 109.550 ;
        RECT 69.530 102.000 69.680 109.550 ;
        RECT 70.130 109.350 74.080 109.550 ;
        RECT 75.380 109.350 79.330 109.550 ;
        RECT 70.130 108.900 70.730 109.350 ;
        RECT 78.730 108.900 79.330 109.350 ;
        RECT 70.130 108.750 74.080 108.900 ;
        RECT 75.380 108.750 79.330 108.900 ;
        RECT 70.130 108.300 70.730 108.750 ;
        RECT 78.730 108.300 79.330 108.750 ;
        RECT 70.130 108.150 74.080 108.300 ;
        RECT 75.380 108.150 79.330 108.300 ;
        RECT 70.130 107.700 70.730 108.150 ;
        RECT 78.730 107.700 79.330 108.150 ;
        RECT 70.130 107.550 74.080 107.700 ;
        RECT 75.380 107.550 79.330 107.700 ;
        RECT 70.130 107.100 70.730 107.550 ;
        RECT 78.730 107.100 79.330 107.550 ;
        RECT 70.130 106.950 74.080 107.100 ;
        RECT 75.380 106.950 79.330 107.100 ;
        RECT 70.130 106.500 70.730 106.950 ;
        RECT 78.730 106.500 79.330 106.950 ;
        RECT 70.130 106.350 74.080 106.500 ;
        RECT 75.380 106.350 79.330 106.500 ;
        RECT 70.130 105.900 70.730 106.350 ;
        RECT 78.730 105.900 79.330 106.350 ;
        RECT 70.130 105.750 74.080 105.900 ;
        RECT 75.380 105.750 79.330 105.900 ;
        RECT 70.130 105.300 70.730 105.750 ;
        RECT 78.730 105.300 79.330 105.750 ;
        RECT 70.130 105.150 74.080 105.300 ;
        RECT 75.380 105.150 79.330 105.300 ;
        RECT 70.130 104.700 70.730 105.150 ;
        RECT 78.730 104.700 79.330 105.150 ;
        RECT 70.130 104.550 74.080 104.700 ;
        RECT 75.380 104.550 79.330 104.700 ;
        RECT 70.130 104.100 70.730 104.550 ;
        RECT 78.730 104.100 79.330 104.550 ;
        RECT 70.130 103.950 74.080 104.100 ;
        RECT 75.380 103.950 79.330 104.100 ;
        RECT 70.130 103.500 70.730 103.950 ;
        RECT 78.730 103.500 79.330 103.950 ;
        RECT 70.130 103.350 74.080 103.500 ;
        RECT 75.380 103.350 79.330 103.500 ;
        RECT 70.130 102.900 70.730 103.350 ;
        RECT 78.730 102.900 79.330 103.350 ;
        RECT 70.130 102.750 74.080 102.900 ;
        RECT 75.380 102.750 79.330 102.900 ;
        RECT 70.130 102.300 70.730 102.750 ;
        RECT 78.730 102.300 79.330 102.750 ;
        RECT 70.130 102.150 74.080 102.300 ;
        RECT 75.380 102.150 79.330 102.300 ;
        RECT 70.130 102.000 70.730 102.150 ;
        RECT 66.530 101.700 70.730 102.000 ;
        RECT 78.730 102.000 79.330 102.150 ;
        RECT 79.780 102.000 79.930 109.550 ;
        RECT 80.380 102.000 80.530 109.550 ;
        RECT 80.980 102.000 81.130 109.550 ;
        RECT 81.580 102.000 81.730 109.550 ;
        RECT 82.180 102.000 82.330 109.550 ;
        RECT 82.780 102.000 82.930 104.900 ;
        RECT 78.730 101.700 82.930 102.000 ;
        RECT 66.530 101.550 74.080 101.700 ;
        RECT 75.380 101.550 82.930 101.700 ;
        RECT 66.530 101.350 70.730 101.550 ;
        RECT 60.330 101.050 69.130 101.200 ;
        RECT 69.280 101.050 70.730 101.350 ;
        RECT 58.730 100.150 70.730 101.050 ;
        RECT 78.730 101.350 82.930 101.550 ;
        RECT 78.730 101.050 80.180 101.350 ;
        RECT 83.530 101.200 85.930 104.400 ;
        RECT 86.530 102.000 86.680 104.900 ;
        RECT 87.130 102.000 87.280 109.550 ;
        RECT 87.730 102.000 87.880 109.550 ;
        RECT 88.330 102.000 88.480 109.550 ;
        RECT 88.930 102.000 89.080 109.550 ;
        RECT 89.530 102.000 89.680 109.550 ;
        RECT 90.130 109.350 94.080 109.550 ;
        RECT 95.380 109.350 99.330 109.550 ;
        RECT 90.130 108.900 90.730 109.350 ;
        RECT 98.730 108.900 99.330 109.350 ;
        RECT 90.130 108.750 94.080 108.900 ;
        RECT 95.380 108.750 99.330 108.900 ;
        RECT 90.130 108.300 90.730 108.750 ;
        RECT 98.730 108.300 99.330 108.750 ;
        RECT 90.130 108.150 94.080 108.300 ;
        RECT 95.380 108.150 99.330 108.300 ;
        RECT 90.130 107.700 90.730 108.150 ;
        RECT 98.730 107.700 99.330 108.150 ;
        RECT 90.130 107.550 94.080 107.700 ;
        RECT 95.380 107.550 99.330 107.700 ;
        RECT 90.130 107.100 90.730 107.550 ;
        RECT 98.730 107.100 99.330 107.550 ;
        RECT 90.130 106.950 94.080 107.100 ;
        RECT 95.380 106.950 99.330 107.100 ;
        RECT 90.130 106.500 90.730 106.950 ;
        RECT 98.730 106.500 99.330 106.950 ;
        RECT 90.130 106.350 94.080 106.500 ;
        RECT 95.380 106.350 99.330 106.500 ;
        RECT 90.130 105.900 90.730 106.350 ;
        RECT 98.730 105.900 99.330 106.350 ;
        RECT 90.130 105.750 94.080 105.900 ;
        RECT 95.380 105.750 99.330 105.900 ;
        RECT 90.130 105.300 90.730 105.750 ;
        RECT 98.730 105.300 99.330 105.750 ;
        RECT 90.130 105.150 94.080 105.300 ;
        RECT 95.380 105.150 99.330 105.300 ;
        RECT 90.130 104.700 90.730 105.150 ;
        RECT 98.730 104.700 99.330 105.150 ;
        RECT 90.130 104.550 94.080 104.700 ;
        RECT 95.380 104.550 99.330 104.700 ;
        RECT 90.130 104.100 90.730 104.550 ;
        RECT 98.730 104.100 99.330 104.550 ;
        RECT 90.130 103.950 94.080 104.100 ;
        RECT 95.380 103.950 99.330 104.100 ;
        RECT 90.130 103.500 90.730 103.950 ;
        RECT 98.730 103.500 99.330 103.950 ;
        RECT 90.130 103.350 94.080 103.500 ;
        RECT 95.380 103.350 99.330 103.500 ;
        RECT 90.130 102.900 90.730 103.350 ;
        RECT 98.730 102.900 99.330 103.350 ;
        RECT 90.130 102.750 94.080 102.900 ;
        RECT 95.380 102.750 99.330 102.900 ;
        RECT 90.130 102.300 90.730 102.750 ;
        RECT 98.730 102.300 99.330 102.750 ;
        RECT 90.130 102.150 94.080 102.300 ;
        RECT 95.380 102.150 99.330 102.300 ;
        RECT 90.130 102.000 90.730 102.150 ;
        RECT 86.530 101.700 90.730 102.000 ;
        RECT 98.730 102.000 99.330 102.150 ;
        RECT 99.780 102.000 99.930 109.550 ;
        RECT 100.380 102.000 100.530 109.550 ;
        RECT 100.980 102.000 101.130 109.550 ;
        RECT 101.580 102.000 101.730 109.550 ;
        RECT 102.180 102.000 102.330 109.550 ;
        RECT 102.780 102.000 102.930 104.900 ;
        RECT 98.730 101.700 102.930 102.000 ;
        RECT 86.530 101.550 94.080 101.700 ;
        RECT 95.380 101.550 102.930 101.700 ;
        RECT 86.530 101.350 90.730 101.550 ;
        RECT 80.330 101.050 89.130 101.200 ;
        RECT 89.280 101.050 90.730 101.350 ;
        RECT 78.730 100.150 90.730 101.050 ;
        RECT 98.730 101.350 102.930 101.550 ;
        RECT 98.730 101.050 100.180 101.350 ;
        RECT 103.530 101.200 105.930 104.400 ;
        RECT 106.530 102.000 106.680 104.900 ;
        RECT 107.130 102.000 107.280 109.550 ;
        RECT 107.730 102.000 107.880 109.550 ;
        RECT 108.330 102.000 108.480 109.550 ;
        RECT 108.930 102.000 109.080 109.550 ;
        RECT 109.530 102.000 109.680 109.550 ;
        RECT 110.130 109.350 114.080 109.550 ;
        RECT 115.380 109.350 119.330 109.550 ;
        RECT 110.130 108.900 110.730 109.350 ;
        RECT 118.730 108.900 119.330 109.350 ;
        RECT 110.130 108.750 114.080 108.900 ;
        RECT 115.380 108.750 119.330 108.900 ;
        RECT 110.130 108.300 110.730 108.750 ;
        RECT 118.730 108.300 119.330 108.750 ;
        RECT 110.130 108.150 114.080 108.300 ;
        RECT 115.380 108.150 119.330 108.300 ;
        RECT 110.130 107.700 110.730 108.150 ;
        RECT 118.730 107.700 119.330 108.150 ;
        RECT 110.130 107.550 114.080 107.700 ;
        RECT 115.380 107.550 119.330 107.700 ;
        RECT 110.130 107.100 110.730 107.550 ;
        RECT 118.730 107.100 119.330 107.550 ;
        RECT 110.130 106.950 114.080 107.100 ;
        RECT 115.380 106.950 119.330 107.100 ;
        RECT 110.130 106.500 110.730 106.950 ;
        RECT 118.730 106.500 119.330 106.950 ;
        RECT 110.130 106.350 114.080 106.500 ;
        RECT 115.380 106.350 119.330 106.500 ;
        RECT 110.130 105.900 110.730 106.350 ;
        RECT 118.730 105.900 119.330 106.350 ;
        RECT 110.130 105.750 114.080 105.900 ;
        RECT 115.380 105.750 119.330 105.900 ;
        RECT 110.130 105.300 110.730 105.750 ;
        RECT 118.730 105.300 119.330 105.750 ;
        RECT 110.130 105.150 114.080 105.300 ;
        RECT 115.380 105.150 119.330 105.300 ;
        RECT 110.130 104.700 110.730 105.150 ;
        RECT 118.730 104.700 119.330 105.150 ;
        RECT 110.130 104.550 114.080 104.700 ;
        RECT 115.380 104.550 119.330 104.700 ;
        RECT 110.130 104.100 110.730 104.550 ;
        RECT 118.730 104.100 119.330 104.550 ;
        RECT 110.130 103.950 114.080 104.100 ;
        RECT 115.380 103.950 119.330 104.100 ;
        RECT 110.130 103.500 110.730 103.950 ;
        RECT 118.730 103.500 119.330 103.950 ;
        RECT 110.130 103.350 114.080 103.500 ;
        RECT 115.380 103.350 119.330 103.500 ;
        RECT 110.130 102.900 110.730 103.350 ;
        RECT 118.730 102.900 119.330 103.350 ;
        RECT 110.130 102.750 114.080 102.900 ;
        RECT 115.380 102.750 119.330 102.900 ;
        RECT 110.130 102.300 110.730 102.750 ;
        RECT 118.730 102.300 119.330 102.750 ;
        RECT 110.130 102.150 114.080 102.300 ;
        RECT 115.380 102.150 119.330 102.300 ;
        RECT 110.130 102.000 110.730 102.150 ;
        RECT 106.530 101.700 110.730 102.000 ;
        RECT 118.730 102.000 119.330 102.150 ;
        RECT 119.780 102.000 119.930 109.550 ;
        RECT 120.380 102.000 120.530 109.550 ;
        RECT 120.980 102.000 121.130 109.550 ;
        RECT 121.580 102.000 121.730 109.550 ;
        RECT 122.180 102.000 122.330 109.550 ;
        RECT 122.780 102.000 122.930 104.900 ;
        RECT 118.730 101.700 122.930 102.000 ;
        RECT 106.530 101.550 114.080 101.700 ;
        RECT 115.380 101.550 122.930 101.700 ;
        RECT 106.530 101.350 110.730 101.550 ;
        RECT 100.330 101.050 109.130 101.200 ;
        RECT 109.280 101.050 110.730 101.350 ;
        RECT 98.730 100.150 110.730 101.050 ;
        RECT 118.730 101.350 122.930 101.550 ;
        RECT 123.530 103.120 124.730 104.400 ;
        RECT 123.530 101.845 127.140 103.120 ;
        RECT 118.730 101.050 120.180 101.350 ;
        RECT 123.530 101.200 124.730 101.845 ;
        RECT 120.330 101.050 124.730 101.200 ;
        RECT 118.730 100.150 124.730 101.050 ;
        RECT 4.730 99.850 9.130 100.150 ;
        RECT 20.330 99.850 29.130 100.150 ;
        RECT 40.330 99.850 49.130 100.150 ;
        RECT 60.330 99.850 69.130 100.150 ;
        RECT 80.330 99.850 89.130 100.150 ;
        RECT 100.330 99.850 109.130 100.150 ;
        RECT 4.730 98.950 10.730 99.850 ;
        RECT 20.330 99.800 30.730 99.850 ;
        RECT 40.330 99.800 50.730 99.850 ;
        RECT 60.330 99.800 70.730 99.850 ;
        RECT 80.330 99.800 90.730 99.850 ;
        RECT 100.330 99.800 110.730 99.850 ;
        RECT 120.330 99.800 124.730 100.150 ;
        RECT 4.730 98.800 9.130 98.950 ;
        RECT 4.730 97.845 5.930 98.800 ;
        RECT 9.280 98.650 10.730 98.950 ;
        RECT 2.315 96.570 5.930 97.845 ;
        RECT 4.730 95.600 5.930 96.570 ;
        RECT 6.530 98.450 10.730 98.650 ;
        RECT 18.730 98.950 30.730 99.800 ;
        RECT 18.730 98.900 29.130 98.950 ;
        RECT 18.730 98.650 20.180 98.900 ;
        RECT 20.330 98.800 29.130 98.900 ;
        RECT 18.730 98.450 22.930 98.650 ;
        RECT 6.530 98.300 14.080 98.450 ;
        RECT 15.430 98.300 22.930 98.450 ;
        RECT 6.530 98.000 10.730 98.300 ;
        RECT 2.315 93.250 4.315 95.545 ;
        RECT 6.530 95.150 6.680 98.000 ;
        RECT 7.130 90.450 7.280 98.000 ;
        RECT 7.730 90.450 7.880 98.000 ;
        RECT 8.330 90.450 8.480 98.000 ;
        RECT 8.930 90.450 9.080 98.000 ;
        RECT 9.530 90.450 9.680 98.000 ;
        RECT 10.130 97.850 10.730 98.000 ;
        RECT 18.730 98.000 22.930 98.300 ;
        RECT 18.730 97.850 19.330 98.000 ;
        RECT 10.130 97.700 14.080 97.850 ;
        RECT 15.380 97.700 19.330 97.850 ;
        RECT 10.130 97.250 10.730 97.700 ;
        RECT 18.730 97.250 19.330 97.700 ;
        RECT 10.130 97.100 14.080 97.250 ;
        RECT 15.380 97.100 19.330 97.250 ;
        RECT 10.130 96.650 10.730 97.100 ;
        RECT 18.730 96.650 19.330 97.100 ;
        RECT 10.130 96.500 14.080 96.650 ;
        RECT 15.380 96.500 19.330 96.650 ;
        RECT 10.130 96.050 10.730 96.500 ;
        RECT 18.730 96.050 19.330 96.500 ;
        RECT 10.130 95.900 14.080 96.050 ;
        RECT 15.380 95.900 19.330 96.050 ;
        RECT 10.130 95.450 10.730 95.900 ;
        RECT 18.730 95.450 19.330 95.900 ;
        RECT 10.130 95.300 14.080 95.450 ;
        RECT 15.380 95.300 19.330 95.450 ;
        RECT 10.130 94.850 10.730 95.300 ;
        RECT 18.730 94.850 19.330 95.300 ;
        RECT 10.130 94.700 14.080 94.850 ;
        RECT 15.380 94.700 19.330 94.850 ;
        RECT 10.130 94.250 10.730 94.700 ;
        RECT 18.730 94.250 19.330 94.700 ;
        RECT 10.130 94.100 14.080 94.250 ;
        RECT 15.380 94.100 19.330 94.250 ;
        RECT 10.130 93.650 10.730 94.100 ;
        RECT 18.730 93.650 19.330 94.100 ;
        RECT 10.130 93.500 14.080 93.650 ;
        RECT 15.380 93.500 19.330 93.650 ;
        RECT 10.130 93.050 10.730 93.500 ;
        RECT 18.730 93.050 19.330 93.500 ;
        RECT 10.130 92.900 14.080 93.050 ;
        RECT 15.380 92.900 19.330 93.050 ;
        RECT 10.130 92.450 10.730 92.900 ;
        RECT 18.730 92.450 19.330 92.900 ;
        RECT 10.130 92.300 14.080 92.450 ;
        RECT 15.380 92.300 19.330 92.450 ;
        RECT 10.130 91.850 10.730 92.300 ;
        RECT 18.730 91.850 19.330 92.300 ;
        RECT 10.130 91.700 14.080 91.850 ;
        RECT 15.380 91.700 19.330 91.850 ;
        RECT 10.130 91.250 10.730 91.700 ;
        RECT 18.730 91.250 19.330 91.700 ;
        RECT 10.130 91.100 14.080 91.250 ;
        RECT 15.380 91.100 19.330 91.250 ;
        RECT 10.130 90.650 10.730 91.100 ;
        RECT 18.730 90.650 19.330 91.100 ;
        RECT 10.130 90.450 14.080 90.650 ;
        RECT 15.380 90.450 19.330 90.650 ;
        RECT 19.780 90.450 19.930 98.000 ;
        RECT 20.380 90.450 20.530 98.000 ;
        RECT 20.980 90.450 21.130 98.000 ;
        RECT 21.580 90.450 21.730 98.000 ;
        RECT 22.180 90.450 22.330 98.000 ;
        RECT 22.780 95.150 22.930 98.000 ;
        RECT 23.530 95.600 25.930 98.800 ;
        RECT 29.280 98.650 30.730 98.950 ;
        RECT 26.530 98.450 30.730 98.650 ;
        RECT 38.730 98.950 50.730 99.800 ;
        RECT 38.730 98.900 49.130 98.950 ;
        RECT 38.730 98.650 40.180 98.900 ;
        RECT 40.330 98.800 49.130 98.900 ;
        RECT 38.730 98.450 42.930 98.650 ;
        RECT 26.530 98.300 34.080 98.450 ;
        RECT 35.430 98.300 42.930 98.450 ;
        RECT 26.530 98.000 30.730 98.300 ;
        RECT 26.530 95.150 26.680 98.000 ;
        RECT 27.130 90.450 27.280 98.000 ;
        RECT 27.730 90.450 27.880 98.000 ;
        RECT 28.330 90.450 28.480 98.000 ;
        RECT 28.930 90.450 29.080 98.000 ;
        RECT 29.530 90.450 29.680 98.000 ;
        RECT 30.130 97.850 30.730 98.000 ;
        RECT 38.730 98.000 42.930 98.300 ;
        RECT 38.730 97.850 39.330 98.000 ;
        RECT 30.130 97.700 34.080 97.850 ;
        RECT 35.380 97.700 39.330 97.850 ;
        RECT 30.130 97.250 30.730 97.700 ;
        RECT 38.730 97.250 39.330 97.700 ;
        RECT 30.130 97.100 34.080 97.250 ;
        RECT 35.380 97.100 39.330 97.250 ;
        RECT 30.130 96.650 30.730 97.100 ;
        RECT 38.730 96.650 39.330 97.100 ;
        RECT 30.130 96.500 34.080 96.650 ;
        RECT 35.380 96.500 39.330 96.650 ;
        RECT 30.130 96.050 30.730 96.500 ;
        RECT 38.730 96.050 39.330 96.500 ;
        RECT 30.130 95.900 34.080 96.050 ;
        RECT 35.380 95.900 39.330 96.050 ;
        RECT 30.130 95.450 30.730 95.900 ;
        RECT 38.730 95.450 39.330 95.900 ;
        RECT 30.130 95.300 34.080 95.450 ;
        RECT 35.380 95.300 39.330 95.450 ;
        RECT 30.130 94.850 30.730 95.300 ;
        RECT 38.730 94.850 39.330 95.300 ;
        RECT 30.130 94.700 34.080 94.850 ;
        RECT 35.380 94.700 39.330 94.850 ;
        RECT 30.130 94.250 30.730 94.700 ;
        RECT 38.730 94.250 39.330 94.700 ;
        RECT 30.130 94.100 34.080 94.250 ;
        RECT 35.380 94.100 39.330 94.250 ;
        RECT 30.130 93.650 30.730 94.100 ;
        RECT 38.730 93.650 39.330 94.100 ;
        RECT 30.130 93.500 34.080 93.650 ;
        RECT 35.380 93.500 39.330 93.650 ;
        RECT 30.130 93.050 30.730 93.500 ;
        RECT 38.730 93.050 39.330 93.500 ;
        RECT 30.130 92.900 34.080 93.050 ;
        RECT 35.380 92.900 39.330 93.050 ;
        RECT 30.130 92.450 30.730 92.900 ;
        RECT 38.730 92.450 39.330 92.900 ;
        RECT 30.130 92.300 34.080 92.450 ;
        RECT 35.380 92.300 39.330 92.450 ;
        RECT 30.130 91.850 30.730 92.300 ;
        RECT 38.730 91.850 39.330 92.300 ;
        RECT 30.130 91.700 34.080 91.850 ;
        RECT 35.380 91.700 39.330 91.850 ;
        RECT 30.130 91.250 30.730 91.700 ;
        RECT 38.730 91.250 39.330 91.700 ;
        RECT 30.130 91.100 34.080 91.250 ;
        RECT 35.380 91.100 39.330 91.250 ;
        RECT 30.130 90.650 30.730 91.100 ;
        RECT 38.730 90.650 39.330 91.100 ;
        RECT 30.130 90.450 34.080 90.650 ;
        RECT 35.380 90.450 39.330 90.650 ;
        RECT 39.780 90.450 39.930 98.000 ;
        RECT 40.380 90.450 40.530 98.000 ;
        RECT 40.980 90.450 41.130 98.000 ;
        RECT 41.580 90.450 41.730 98.000 ;
        RECT 42.180 90.450 42.330 98.000 ;
        RECT 42.780 95.150 42.930 98.000 ;
        RECT 43.530 95.600 45.930 98.800 ;
        RECT 49.280 98.650 50.730 98.950 ;
        RECT 46.530 98.450 50.730 98.650 ;
        RECT 58.730 98.950 70.730 99.800 ;
        RECT 58.730 98.900 69.130 98.950 ;
        RECT 58.730 98.650 60.180 98.900 ;
        RECT 60.330 98.800 69.130 98.900 ;
        RECT 58.730 98.450 62.930 98.650 ;
        RECT 46.530 98.300 54.080 98.450 ;
        RECT 55.430 98.300 62.930 98.450 ;
        RECT 46.530 98.000 50.730 98.300 ;
        RECT 46.530 95.150 46.680 98.000 ;
        RECT 47.130 90.450 47.280 98.000 ;
        RECT 47.730 90.450 47.880 98.000 ;
        RECT 48.330 90.450 48.480 98.000 ;
        RECT 48.930 90.450 49.080 98.000 ;
        RECT 49.530 90.450 49.680 98.000 ;
        RECT 50.130 97.850 50.730 98.000 ;
        RECT 58.730 98.000 62.930 98.300 ;
        RECT 58.730 97.850 59.330 98.000 ;
        RECT 50.130 97.700 54.080 97.850 ;
        RECT 55.380 97.700 59.330 97.850 ;
        RECT 50.130 97.250 50.730 97.700 ;
        RECT 58.730 97.250 59.330 97.700 ;
        RECT 50.130 97.100 54.080 97.250 ;
        RECT 55.380 97.100 59.330 97.250 ;
        RECT 50.130 96.650 50.730 97.100 ;
        RECT 58.730 96.650 59.330 97.100 ;
        RECT 50.130 96.500 54.080 96.650 ;
        RECT 55.380 96.500 59.330 96.650 ;
        RECT 50.130 96.050 50.730 96.500 ;
        RECT 58.730 96.050 59.330 96.500 ;
        RECT 50.130 95.900 54.080 96.050 ;
        RECT 55.380 95.900 59.330 96.050 ;
        RECT 50.130 95.450 50.730 95.900 ;
        RECT 58.730 95.450 59.330 95.900 ;
        RECT 50.130 95.300 54.080 95.450 ;
        RECT 55.380 95.300 59.330 95.450 ;
        RECT 50.130 94.850 50.730 95.300 ;
        RECT 58.730 94.850 59.330 95.300 ;
        RECT 50.130 94.700 54.080 94.850 ;
        RECT 55.380 94.700 59.330 94.850 ;
        RECT 50.130 94.250 50.730 94.700 ;
        RECT 58.730 94.250 59.330 94.700 ;
        RECT 50.130 94.100 54.080 94.250 ;
        RECT 55.380 94.100 59.330 94.250 ;
        RECT 50.130 93.650 50.730 94.100 ;
        RECT 58.730 93.650 59.330 94.100 ;
        RECT 50.130 93.500 54.080 93.650 ;
        RECT 55.380 93.500 59.330 93.650 ;
        RECT 50.130 93.050 50.730 93.500 ;
        RECT 58.730 93.050 59.330 93.500 ;
        RECT 50.130 92.900 54.080 93.050 ;
        RECT 55.380 92.900 59.330 93.050 ;
        RECT 50.130 92.450 50.730 92.900 ;
        RECT 58.730 92.450 59.330 92.900 ;
        RECT 50.130 92.300 54.080 92.450 ;
        RECT 55.380 92.300 59.330 92.450 ;
        RECT 50.130 91.850 50.730 92.300 ;
        RECT 58.730 91.850 59.330 92.300 ;
        RECT 50.130 91.700 54.080 91.850 ;
        RECT 55.380 91.700 59.330 91.850 ;
        RECT 50.130 91.250 50.730 91.700 ;
        RECT 58.730 91.250 59.330 91.700 ;
        RECT 50.130 91.100 54.080 91.250 ;
        RECT 55.380 91.100 59.330 91.250 ;
        RECT 50.130 90.650 50.730 91.100 ;
        RECT 58.730 90.650 59.330 91.100 ;
        RECT 50.130 90.450 54.080 90.650 ;
        RECT 55.380 90.450 59.330 90.650 ;
        RECT 59.780 90.450 59.930 98.000 ;
        RECT 60.380 90.450 60.530 98.000 ;
        RECT 60.980 90.450 61.130 98.000 ;
        RECT 61.580 90.450 61.730 98.000 ;
        RECT 62.180 90.450 62.330 98.000 ;
        RECT 62.780 95.150 62.930 98.000 ;
        RECT 63.530 95.600 65.930 98.800 ;
        RECT 69.280 98.650 70.730 98.950 ;
        RECT 66.530 98.450 70.730 98.650 ;
        RECT 78.730 98.950 90.730 99.800 ;
        RECT 78.730 98.900 89.130 98.950 ;
        RECT 78.730 98.650 80.180 98.900 ;
        RECT 80.330 98.800 89.130 98.900 ;
        RECT 78.730 98.450 82.930 98.650 ;
        RECT 66.530 98.300 74.080 98.450 ;
        RECT 75.430 98.300 82.930 98.450 ;
        RECT 66.530 98.000 70.730 98.300 ;
        RECT 66.530 95.150 66.680 98.000 ;
        RECT 67.130 90.450 67.280 98.000 ;
        RECT 67.730 90.450 67.880 98.000 ;
        RECT 68.330 90.450 68.480 98.000 ;
        RECT 68.930 90.450 69.080 98.000 ;
        RECT 69.530 90.450 69.680 98.000 ;
        RECT 70.130 97.850 70.730 98.000 ;
        RECT 78.730 98.000 82.930 98.300 ;
        RECT 78.730 97.850 79.330 98.000 ;
        RECT 70.130 97.700 74.080 97.850 ;
        RECT 75.380 97.700 79.330 97.850 ;
        RECT 70.130 97.250 70.730 97.700 ;
        RECT 78.730 97.250 79.330 97.700 ;
        RECT 70.130 97.100 74.080 97.250 ;
        RECT 75.380 97.100 79.330 97.250 ;
        RECT 70.130 96.650 70.730 97.100 ;
        RECT 78.730 96.650 79.330 97.100 ;
        RECT 70.130 96.500 74.080 96.650 ;
        RECT 75.380 96.500 79.330 96.650 ;
        RECT 70.130 96.050 70.730 96.500 ;
        RECT 78.730 96.050 79.330 96.500 ;
        RECT 70.130 95.900 74.080 96.050 ;
        RECT 75.380 95.900 79.330 96.050 ;
        RECT 70.130 95.450 70.730 95.900 ;
        RECT 78.730 95.450 79.330 95.900 ;
        RECT 70.130 95.300 74.080 95.450 ;
        RECT 75.380 95.300 79.330 95.450 ;
        RECT 70.130 94.850 70.730 95.300 ;
        RECT 78.730 94.850 79.330 95.300 ;
        RECT 70.130 94.700 74.080 94.850 ;
        RECT 75.380 94.700 79.330 94.850 ;
        RECT 70.130 94.250 70.730 94.700 ;
        RECT 78.730 94.250 79.330 94.700 ;
        RECT 70.130 94.100 74.080 94.250 ;
        RECT 75.380 94.100 79.330 94.250 ;
        RECT 70.130 93.650 70.730 94.100 ;
        RECT 78.730 93.650 79.330 94.100 ;
        RECT 70.130 93.500 74.080 93.650 ;
        RECT 75.380 93.500 79.330 93.650 ;
        RECT 70.130 93.050 70.730 93.500 ;
        RECT 78.730 93.050 79.330 93.500 ;
        RECT 70.130 92.900 74.080 93.050 ;
        RECT 75.380 92.900 79.330 93.050 ;
        RECT 70.130 92.450 70.730 92.900 ;
        RECT 78.730 92.450 79.330 92.900 ;
        RECT 70.130 92.300 74.080 92.450 ;
        RECT 75.380 92.300 79.330 92.450 ;
        RECT 70.130 91.850 70.730 92.300 ;
        RECT 78.730 91.850 79.330 92.300 ;
        RECT 70.130 91.700 74.080 91.850 ;
        RECT 75.380 91.700 79.330 91.850 ;
        RECT 70.130 91.250 70.730 91.700 ;
        RECT 78.730 91.250 79.330 91.700 ;
        RECT 70.130 91.100 74.080 91.250 ;
        RECT 75.380 91.100 79.330 91.250 ;
        RECT 70.130 90.650 70.730 91.100 ;
        RECT 78.730 90.650 79.330 91.100 ;
        RECT 70.130 90.450 74.080 90.650 ;
        RECT 75.380 90.450 79.330 90.650 ;
        RECT 79.780 90.450 79.930 98.000 ;
        RECT 80.380 90.450 80.530 98.000 ;
        RECT 80.980 90.450 81.130 98.000 ;
        RECT 81.580 90.450 81.730 98.000 ;
        RECT 82.180 90.450 82.330 98.000 ;
        RECT 82.780 95.150 82.930 98.000 ;
        RECT 83.530 95.600 85.930 98.800 ;
        RECT 89.280 98.650 90.730 98.950 ;
        RECT 86.530 98.450 90.730 98.650 ;
        RECT 98.730 98.950 110.730 99.800 ;
        RECT 98.730 98.900 109.130 98.950 ;
        RECT 98.730 98.650 100.180 98.900 ;
        RECT 100.330 98.800 109.130 98.900 ;
        RECT 98.730 98.450 102.930 98.650 ;
        RECT 86.530 98.300 94.080 98.450 ;
        RECT 95.430 98.300 102.930 98.450 ;
        RECT 86.530 98.000 90.730 98.300 ;
        RECT 86.530 95.150 86.680 98.000 ;
        RECT 87.130 90.450 87.280 98.000 ;
        RECT 87.730 90.450 87.880 98.000 ;
        RECT 88.330 90.450 88.480 98.000 ;
        RECT 88.930 90.450 89.080 98.000 ;
        RECT 89.530 90.450 89.680 98.000 ;
        RECT 90.130 97.850 90.730 98.000 ;
        RECT 98.730 98.000 102.930 98.300 ;
        RECT 98.730 97.850 99.330 98.000 ;
        RECT 90.130 97.700 94.080 97.850 ;
        RECT 95.380 97.700 99.330 97.850 ;
        RECT 90.130 97.250 90.730 97.700 ;
        RECT 98.730 97.250 99.330 97.700 ;
        RECT 90.130 97.100 94.080 97.250 ;
        RECT 95.380 97.100 99.330 97.250 ;
        RECT 90.130 96.650 90.730 97.100 ;
        RECT 98.730 96.650 99.330 97.100 ;
        RECT 90.130 96.500 94.080 96.650 ;
        RECT 95.380 96.500 99.330 96.650 ;
        RECT 90.130 96.050 90.730 96.500 ;
        RECT 98.730 96.050 99.330 96.500 ;
        RECT 90.130 95.900 94.080 96.050 ;
        RECT 95.380 95.900 99.330 96.050 ;
        RECT 90.130 95.450 90.730 95.900 ;
        RECT 98.730 95.450 99.330 95.900 ;
        RECT 90.130 95.300 94.080 95.450 ;
        RECT 95.380 95.300 99.330 95.450 ;
        RECT 90.130 94.850 90.730 95.300 ;
        RECT 98.730 94.850 99.330 95.300 ;
        RECT 90.130 94.700 94.080 94.850 ;
        RECT 95.380 94.700 99.330 94.850 ;
        RECT 90.130 94.250 90.730 94.700 ;
        RECT 98.730 94.250 99.330 94.700 ;
        RECT 90.130 94.100 94.080 94.250 ;
        RECT 95.380 94.100 99.330 94.250 ;
        RECT 90.130 93.650 90.730 94.100 ;
        RECT 98.730 93.650 99.330 94.100 ;
        RECT 90.130 93.500 94.080 93.650 ;
        RECT 95.380 93.500 99.330 93.650 ;
        RECT 90.130 93.050 90.730 93.500 ;
        RECT 98.730 93.050 99.330 93.500 ;
        RECT 90.130 92.900 94.080 93.050 ;
        RECT 95.380 92.900 99.330 93.050 ;
        RECT 90.130 92.450 90.730 92.900 ;
        RECT 98.730 92.450 99.330 92.900 ;
        RECT 90.130 92.300 94.080 92.450 ;
        RECT 95.380 92.300 99.330 92.450 ;
        RECT 90.130 91.850 90.730 92.300 ;
        RECT 98.730 91.850 99.330 92.300 ;
        RECT 90.130 91.700 94.080 91.850 ;
        RECT 95.380 91.700 99.330 91.850 ;
        RECT 90.130 91.250 90.730 91.700 ;
        RECT 98.730 91.250 99.330 91.700 ;
        RECT 90.130 91.100 94.080 91.250 ;
        RECT 95.380 91.100 99.330 91.250 ;
        RECT 90.130 90.650 90.730 91.100 ;
        RECT 98.730 90.650 99.330 91.100 ;
        RECT 90.130 90.450 94.080 90.650 ;
        RECT 95.380 90.450 99.330 90.650 ;
        RECT 99.780 90.450 99.930 98.000 ;
        RECT 100.380 90.450 100.530 98.000 ;
        RECT 100.980 90.450 101.130 98.000 ;
        RECT 101.580 90.450 101.730 98.000 ;
        RECT 102.180 90.450 102.330 98.000 ;
        RECT 102.780 95.150 102.930 98.000 ;
        RECT 103.530 95.600 105.930 98.800 ;
        RECT 109.280 98.650 110.730 98.950 ;
        RECT 106.530 98.450 110.730 98.650 ;
        RECT 118.730 98.900 124.730 99.800 ;
        RECT 118.730 98.650 120.180 98.900 ;
        RECT 120.330 98.800 124.730 98.900 ;
        RECT 118.730 98.450 122.930 98.650 ;
        RECT 106.530 98.300 114.080 98.450 ;
        RECT 115.430 98.300 122.930 98.450 ;
        RECT 106.530 98.000 110.730 98.300 ;
        RECT 106.530 95.150 106.680 98.000 ;
        RECT 107.130 90.450 107.280 98.000 ;
        RECT 107.730 90.450 107.880 98.000 ;
        RECT 108.330 90.450 108.480 98.000 ;
        RECT 108.930 90.450 109.080 98.000 ;
        RECT 109.530 90.450 109.680 98.000 ;
        RECT 110.130 97.850 110.730 98.000 ;
        RECT 118.730 98.000 122.930 98.300 ;
        RECT 118.730 97.850 119.330 98.000 ;
        RECT 110.130 97.700 114.080 97.850 ;
        RECT 115.380 97.700 119.330 97.850 ;
        RECT 110.130 97.250 110.730 97.700 ;
        RECT 118.730 97.250 119.330 97.700 ;
        RECT 110.130 97.100 114.080 97.250 ;
        RECT 115.380 97.100 119.330 97.250 ;
        RECT 110.130 96.650 110.730 97.100 ;
        RECT 118.730 96.650 119.330 97.100 ;
        RECT 110.130 96.500 114.080 96.650 ;
        RECT 115.380 96.500 119.330 96.650 ;
        RECT 110.130 96.050 110.730 96.500 ;
        RECT 118.730 96.050 119.330 96.500 ;
        RECT 110.130 95.900 114.080 96.050 ;
        RECT 115.380 95.900 119.330 96.050 ;
        RECT 110.130 95.450 110.730 95.900 ;
        RECT 118.730 95.450 119.330 95.900 ;
        RECT 110.130 95.300 114.080 95.450 ;
        RECT 115.380 95.300 119.330 95.450 ;
        RECT 110.130 94.850 110.730 95.300 ;
        RECT 118.730 94.850 119.330 95.300 ;
        RECT 110.130 94.700 114.080 94.850 ;
        RECT 115.380 94.700 119.330 94.850 ;
        RECT 110.130 94.250 110.730 94.700 ;
        RECT 118.730 94.250 119.330 94.700 ;
        RECT 110.130 94.100 114.080 94.250 ;
        RECT 115.380 94.100 119.330 94.250 ;
        RECT 110.130 93.650 110.730 94.100 ;
        RECT 118.730 93.650 119.330 94.100 ;
        RECT 110.130 93.500 114.080 93.650 ;
        RECT 115.380 93.500 119.330 93.650 ;
        RECT 110.130 93.050 110.730 93.500 ;
        RECT 118.730 93.050 119.330 93.500 ;
        RECT 110.130 92.900 114.080 93.050 ;
        RECT 115.380 92.900 119.330 93.050 ;
        RECT 110.130 92.450 110.730 92.900 ;
        RECT 118.730 92.450 119.330 92.900 ;
        RECT 110.130 92.300 114.080 92.450 ;
        RECT 115.380 92.300 119.330 92.450 ;
        RECT 110.130 91.850 110.730 92.300 ;
        RECT 118.730 91.850 119.330 92.300 ;
        RECT 110.130 91.700 114.080 91.850 ;
        RECT 115.380 91.700 119.330 91.850 ;
        RECT 110.130 91.250 110.730 91.700 ;
        RECT 118.730 91.250 119.330 91.700 ;
        RECT 110.130 91.100 114.080 91.250 ;
        RECT 115.380 91.100 119.330 91.250 ;
        RECT 110.130 90.650 110.730 91.100 ;
        RECT 118.730 90.650 119.330 91.100 ;
        RECT 110.130 90.450 114.080 90.650 ;
        RECT 115.380 90.450 119.330 90.650 ;
        RECT 119.780 90.450 119.930 98.000 ;
        RECT 120.380 90.450 120.530 98.000 ;
        RECT 120.980 90.450 121.130 98.000 ;
        RECT 121.580 90.450 121.730 98.000 ;
        RECT 122.180 90.450 122.330 98.000 ;
        RECT 122.780 95.150 122.930 98.000 ;
        RECT 123.530 97.245 124.730 98.800 ;
        RECT 123.530 95.970 127.140 97.245 ;
        RECT 123.530 95.600 124.730 95.970 ;
        RECT 2.315 84.455 4.315 86.750 ;
        RECT 4.730 83.470 5.930 84.400 ;
        RECT 2.315 82.195 5.930 83.470 ;
        RECT 4.730 81.200 5.930 82.195 ;
        RECT 6.530 82.000 6.680 84.900 ;
        RECT 7.130 82.000 7.280 89.550 ;
        RECT 7.730 82.000 7.880 89.550 ;
        RECT 8.330 82.000 8.480 89.550 ;
        RECT 8.930 82.000 9.080 89.550 ;
        RECT 9.530 82.000 9.680 89.550 ;
        RECT 10.130 89.350 14.080 89.550 ;
        RECT 15.380 89.350 19.330 89.550 ;
        RECT 10.130 88.900 10.730 89.350 ;
        RECT 18.730 88.900 19.330 89.350 ;
        RECT 10.130 88.750 14.080 88.900 ;
        RECT 15.380 88.750 19.330 88.900 ;
        RECT 10.130 88.300 10.730 88.750 ;
        RECT 18.730 88.300 19.330 88.750 ;
        RECT 10.130 88.150 14.080 88.300 ;
        RECT 15.380 88.150 19.330 88.300 ;
        RECT 10.130 87.700 10.730 88.150 ;
        RECT 18.730 87.700 19.330 88.150 ;
        RECT 10.130 87.550 14.080 87.700 ;
        RECT 15.380 87.550 19.330 87.700 ;
        RECT 10.130 87.100 10.730 87.550 ;
        RECT 18.730 87.100 19.330 87.550 ;
        RECT 10.130 86.950 14.080 87.100 ;
        RECT 15.380 86.950 19.330 87.100 ;
        RECT 10.130 86.500 10.730 86.950 ;
        RECT 18.730 86.500 19.330 86.950 ;
        RECT 10.130 86.350 14.080 86.500 ;
        RECT 15.380 86.350 19.330 86.500 ;
        RECT 10.130 85.900 10.730 86.350 ;
        RECT 18.730 85.900 19.330 86.350 ;
        RECT 10.130 85.750 14.080 85.900 ;
        RECT 15.380 85.750 19.330 85.900 ;
        RECT 10.130 85.300 10.730 85.750 ;
        RECT 18.730 85.300 19.330 85.750 ;
        RECT 10.130 85.150 14.080 85.300 ;
        RECT 15.380 85.150 19.330 85.300 ;
        RECT 10.130 84.700 10.730 85.150 ;
        RECT 18.730 84.700 19.330 85.150 ;
        RECT 10.130 84.550 14.080 84.700 ;
        RECT 15.380 84.550 19.330 84.700 ;
        RECT 10.130 84.100 10.730 84.550 ;
        RECT 18.730 84.100 19.330 84.550 ;
        RECT 10.130 83.950 14.080 84.100 ;
        RECT 15.380 83.950 19.330 84.100 ;
        RECT 10.130 83.500 10.730 83.950 ;
        RECT 18.730 83.500 19.330 83.950 ;
        RECT 10.130 83.350 14.080 83.500 ;
        RECT 15.380 83.350 19.330 83.500 ;
        RECT 10.130 82.900 10.730 83.350 ;
        RECT 18.730 82.900 19.330 83.350 ;
        RECT 10.130 82.750 14.080 82.900 ;
        RECT 15.380 82.750 19.330 82.900 ;
        RECT 10.130 82.300 10.730 82.750 ;
        RECT 18.730 82.300 19.330 82.750 ;
        RECT 10.130 82.150 14.080 82.300 ;
        RECT 15.380 82.150 19.330 82.300 ;
        RECT 10.130 82.000 10.730 82.150 ;
        RECT 6.530 81.700 10.730 82.000 ;
        RECT 18.730 82.000 19.330 82.150 ;
        RECT 19.780 82.000 19.930 89.550 ;
        RECT 20.380 82.000 20.530 89.550 ;
        RECT 20.980 82.000 21.130 89.550 ;
        RECT 21.580 82.000 21.730 89.550 ;
        RECT 22.180 82.000 22.330 89.550 ;
        RECT 22.780 82.000 22.930 84.900 ;
        RECT 18.730 81.700 22.930 82.000 ;
        RECT 6.530 81.550 14.080 81.700 ;
        RECT 15.380 81.550 22.930 81.700 ;
        RECT 6.530 81.350 10.730 81.550 ;
        RECT 4.730 81.050 9.130 81.200 ;
        RECT 9.280 81.050 10.730 81.350 ;
        RECT 4.730 80.150 10.730 81.050 ;
        RECT 18.730 81.350 22.930 81.550 ;
        RECT 18.730 81.050 20.180 81.350 ;
        RECT 23.530 81.200 25.930 84.400 ;
        RECT 26.530 82.000 26.680 84.900 ;
        RECT 27.130 82.000 27.280 89.550 ;
        RECT 27.730 82.000 27.880 89.550 ;
        RECT 28.330 82.000 28.480 89.550 ;
        RECT 28.930 82.000 29.080 89.550 ;
        RECT 29.530 82.000 29.680 89.550 ;
        RECT 30.130 89.350 34.080 89.550 ;
        RECT 35.380 89.350 39.330 89.550 ;
        RECT 30.130 88.900 30.730 89.350 ;
        RECT 38.730 88.900 39.330 89.350 ;
        RECT 30.130 88.750 34.080 88.900 ;
        RECT 35.380 88.750 39.330 88.900 ;
        RECT 30.130 88.300 30.730 88.750 ;
        RECT 38.730 88.300 39.330 88.750 ;
        RECT 30.130 88.150 34.080 88.300 ;
        RECT 35.380 88.150 39.330 88.300 ;
        RECT 30.130 87.700 30.730 88.150 ;
        RECT 38.730 87.700 39.330 88.150 ;
        RECT 30.130 87.550 34.080 87.700 ;
        RECT 35.380 87.550 39.330 87.700 ;
        RECT 30.130 87.100 30.730 87.550 ;
        RECT 38.730 87.100 39.330 87.550 ;
        RECT 30.130 86.950 34.080 87.100 ;
        RECT 35.380 86.950 39.330 87.100 ;
        RECT 30.130 86.500 30.730 86.950 ;
        RECT 38.730 86.500 39.330 86.950 ;
        RECT 30.130 86.350 34.080 86.500 ;
        RECT 35.380 86.350 39.330 86.500 ;
        RECT 30.130 85.900 30.730 86.350 ;
        RECT 38.730 85.900 39.330 86.350 ;
        RECT 30.130 85.750 34.080 85.900 ;
        RECT 35.380 85.750 39.330 85.900 ;
        RECT 30.130 85.300 30.730 85.750 ;
        RECT 38.730 85.300 39.330 85.750 ;
        RECT 30.130 85.150 34.080 85.300 ;
        RECT 35.380 85.150 39.330 85.300 ;
        RECT 30.130 84.700 30.730 85.150 ;
        RECT 38.730 84.700 39.330 85.150 ;
        RECT 30.130 84.550 34.080 84.700 ;
        RECT 35.380 84.550 39.330 84.700 ;
        RECT 30.130 84.100 30.730 84.550 ;
        RECT 38.730 84.100 39.330 84.550 ;
        RECT 30.130 83.950 34.080 84.100 ;
        RECT 35.380 83.950 39.330 84.100 ;
        RECT 30.130 83.500 30.730 83.950 ;
        RECT 38.730 83.500 39.330 83.950 ;
        RECT 30.130 83.350 34.080 83.500 ;
        RECT 35.380 83.350 39.330 83.500 ;
        RECT 30.130 82.900 30.730 83.350 ;
        RECT 38.730 82.900 39.330 83.350 ;
        RECT 30.130 82.750 34.080 82.900 ;
        RECT 35.380 82.750 39.330 82.900 ;
        RECT 30.130 82.300 30.730 82.750 ;
        RECT 38.730 82.300 39.330 82.750 ;
        RECT 30.130 82.150 34.080 82.300 ;
        RECT 35.380 82.150 39.330 82.300 ;
        RECT 30.130 82.000 30.730 82.150 ;
        RECT 26.530 81.700 30.730 82.000 ;
        RECT 38.730 82.000 39.330 82.150 ;
        RECT 39.780 82.000 39.930 89.550 ;
        RECT 40.380 82.000 40.530 89.550 ;
        RECT 40.980 82.000 41.130 89.550 ;
        RECT 41.580 82.000 41.730 89.550 ;
        RECT 42.180 82.000 42.330 89.550 ;
        RECT 42.780 82.000 42.930 84.900 ;
        RECT 38.730 81.700 42.930 82.000 ;
        RECT 26.530 81.550 34.080 81.700 ;
        RECT 35.380 81.550 42.930 81.700 ;
        RECT 26.530 81.350 30.730 81.550 ;
        RECT 20.330 81.050 29.130 81.200 ;
        RECT 29.280 81.050 30.730 81.350 ;
        RECT 18.730 80.150 30.730 81.050 ;
        RECT 38.730 81.350 42.930 81.550 ;
        RECT 38.730 81.050 40.180 81.350 ;
        RECT 43.530 81.200 45.930 84.400 ;
        RECT 46.530 82.000 46.680 84.900 ;
        RECT 47.130 82.000 47.280 89.550 ;
        RECT 47.730 82.000 47.880 89.550 ;
        RECT 48.330 82.000 48.480 89.550 ;
        RECT 48.930 82.000 49.080 89.550 ;
        RECT 49.530 82.000 49.680 89.550 ;
        RECT 50.130 89.350 54.080 89.550 ;
        RECT 55.380 89.350 59.330 89.550 ;
        RECT 50.130 88.900 50.730 89.350 ;
        RECT 58.730 88.900 59.330 89.350 ;
        RECT 50.130 88.750 54.080 88.900 ;
        RECT 55.380 88.750 59.330 88.900 ;
        RECT 50.130 88.300 50.730 88.750 ;
        RECT 58.730 88.300 59.330 88.750 ;
        RECT 50.130 88.150 54.080 88.300 ;
        RECT 55.380 88.150 59.330 88.300 ;
        RECT 50.130 87.700 50.730 88.150 ;
        RECT 58.730 87.700 59.330 88.150 ;
        RECT 50.130 87.550 54.080 87.700 ;
        RECT 55.380 87.550 59.330 87.700 ;
        RECT 50.130 87.100 50.730 87.550 ;
        RECT 58.730 87.100 59.330 87.550 ;
        RECT 50.130 86.950 54.080 87.100 ;
        RECT 55.380 86.950 59.330 87.100 ;
        RECT 50.130 86.500 50.730 86.950 ;
        RECT 58.730 86.500 59.330 86.950 ;
        RECT 50.130 86.350 54.080 86.500 ;
        RECT 55.380 86.350 59.330 86.500 ;
        RECT 50.130 85.900 50.730 86.350 ;
        RECT 58.730 85.900 59.330 86.350 ;
        RECT 50.130 85.750 54.080 85.900 ;
        RECT 55.380 85.750 59.330 85.900 ;
        RECT 50.130 85.300 50.730 85.750 ;
        RECT 58.730 85.300 59.330 85.750 ;
        RECT 50.130 85.150 54.080 85.300 ;
        RECT 55.380 85.150 59.330 85.300 ;
        RECT 50.130 84.700 50.730 85.150 ;
        RECT 58.730 84.700 59.330 85.150 ;
        RECT 50.130 84.550 54.080 84.700 ;
        RECT 55.380 84.550 59.330 84.700 ;
        RECT 50.130 84.100 50.730 84.550 ;
        RECT 58.730 84.100 59.330 84.550 ;
        RECT 50.130 83.950 54.080 84.100 ;
        RECT 55.380 83.950 59.330 84.100 ;
        RECT 50.130 83.500 50.730 83.950 ;
        RECT 58.730 83.500 59.330 83.950 ;
        RECT 50.130 83.350 54.080 83.500 ;
        RECT 55.380 83.350 59.330 83.500 ;
        RECT 50.130 82.900 50.730 83.350 ;
        RECT 58.730 82.900 59.330 83.350 ;
        RECT 50.130 82.750 54.080 82.900 ;
        RECT 55.380 82.750 59.330 82.900 ;
        RECT 50.130 82.300 50.730 82.750 ;
        RECT 58.730 82.300 59.330 82.750 ;
        RECT 50.130 82.150 54.080 82.300 ;
        RECT 55.380 82.150 59.330 82.300 ;
        RECT 50.130 82.000 50.730 82.150 ;
        RECT 46.530 81.700 50.730 82.000 ;
        RECT 58.730 82.000 59.330 82.150 ;
        RECT 59.780 82.000 59.930 89.550 ;
        RECT 60.380 82.000 60.530 89.550 ;
        RECT 60.980 82.000 61.130 89.550 ;
        RECT 61.580 82.000 61.730 89.550 ;
        RECT 62.180 82.000 62.330 89.550 ;
        RECT 62.780 82.000 62.930 84.900 ;
        RECT 58.730 81.700 62.930 82.000 ;
        RECT 46.530 81.550 54.080 81.700 ;
        RECT 55.380 81.550 62.930 81.700 ;
        RECT 46.530 81.350 50.730 81.550 ;
        RECT 40.330 81.050 49.130 81.200 ;
        RECT 49.280 81.050 50.730 81.350 ;
        RECT 38.730 80.150 50.730 81.050 ;
        RECT 58.730 81.350 62.930 81.550 ;
        RECT 58.730 81.050 60.180 81.350 ;
        RECT 63.530 81.200 65.930 84.400 ;
        RECT 66.530 82.000 66.680 84.900 ;
        RECT 67.130 82.000 67.280 89.550 ;
        RECT 67.730 82.000 67.880 89.550 ;
        RECT 68.330 82.000 68.480 89.550 ;
        RECT 68.930 82.000 69.080 89.550 ;
        RECT 69.530 82.000 69.680 89.550 ;
        RECT 70.130 89.350 74.080 89.550 ;
        RECT 75.380 89.350 79.330 89.550 ;
        RECT 70.130 88.900 70.730 89.350 ;
        RECT 78.730 88.900 79.330 89.350 ;
        RECT 70.130 88.750 74.080 88.900 ;
        RECT 75.380 88.750 79.330 88.900 ;
        RECT 70.130 88.300 70.730 88.750 ;
        RECT 78.730 88.300 79.330 88.750 ;
        RECT 70.130 88.150 74.080 88.300 ;
        RECT 75.380 88.150 79.330 88.300 ;
        RECT 70.130 87.700 70.730 88.150 ;
        RECT 78.730 87.700 79.330 88.150 ;
        RECT 70.130 87.550 74.080 87.700 ;
        RECT 75.380 87.550 79.330 87.700 ;
        RECT 70.130 87.100 70.730 87.550 ;
        RECT 78.730 87.100 79.330 87.550 ;
        RECT 70.130 86.950 74.080 87.100 ;
        RECT 75.380 86.950 79.330 87.100 ;
        RECT 70.130 86.500 70.730 86.950 ;
        RECT 78.730 86.500 79.330 86.950 ;
        RECT 70.130 86.350 74.080 86.500 ;
        RECT 75.380 86.350 79.330 86.500 ;
        RECT 70.130 85.900 70.730 86.350 ;
        RECT 78.730 85.900 79.330 86.350 ;
        RECT 70.130 85.750 74.080 85.900 ;
        RECT 75.380 85.750 79.330 85.900 ;
        RECT 70.130 85.300 70.730 85.750 ;
        RECT 78.730 85.300 79.330 85.750 ;
        RECT 70.130 85.150 74.080 85.300 ;
        RECT 75.380 85.150 79.330 85.300 ;
        RECT 70.130 84.700 70.730 85.150 ;
        RECT 78.730 84.700 79.330 85.150 ;
        RECT 70.130 84.550 74.080 84.700 ;
        RECT 75.380 84.550 79.330 84.700 ;
        RECT 70.130 84.100 70.730 84.550 ;
        RECT 78.730 84.100 79.330 84.550 ;
        RECT 70.130 83.950 74.080 84.100 ;
        RECT 75.380 83.950 79.330 84.100 ;
        RECT 70.130 83.500 70.730 83.950 ;
        RECT 78.730 83.500 79.330 83.950 ;
        RECT 70.130 83.350 74.080 83.500 ;
        RECT 75.380 83.350 79.330 83.500 ;
        RECT 70.130 82.900 70.730 83.350 ;
        RECT 78.730 82.900 79.330 83.350 ;
        RECT 70.130 82.750 74.080 82.900 ;
        RECT 75.380 82.750 79.330 82.900 ;
        RECT 70.130 82.300 70.730 82.750 ;
        RECT 78.730 82.300 79.330 82.750 ;
        RECT 70.130 82.150 74.080 82.300 ;
        RECT 75.380 82.150 79.330 82.300 ;
        RECT 70.130 82.000 70.730 82.150 ;
        RECT 66.530 81.700 70.730 82.000 ;
        RECT 78.730 82.000 79.330 82.150 ;
        RECT 79.780 82.000 79.930 89.550 ;
        RECT 80.380 82.000 80.530 89.550 ;
        RECT 80.980 82.000 81.130 89.550 ;
        RECT 81.580 82.000 81.730 89.550 ;
        RECT 82.180 82.000 82.330 89.550 ;
        RECT 82.780 82.000 82.930 84.900 ;
        RECT 78.730 81.700 82.930 82.000 ;
        RECT 66.530 81.550 74.080 81.700 ;
        RECT 75.380 81.550 82.930 81.700 ;
        RECT 66.530 81.350 70.730 81.550 ;
        RECT 60.330 81.050 69.130 81.200 ;
        RECT 69.280 81.050 70.730 81.350 ;
        RECT 58.730 80.150 70.730 81.050 ;
        RECT 78.730 81.350 82.930 81.550 ;
        RECT 78.730 81.050 80.180 81.350 ;
        RECT 83.530 81.200 85.930 84.400 ;
        RECT 86.530 82.000 86.680 84.900 ;
        RECT 87.130 82.000 87.280 89.550 ;
        RECT 87.730 82.000 87.880 89.550 ;
        RECT 88.330 82.000 88.480 89.550 ;
        RECT 88.930 82.000 89.080 89.550 ;
        RECT 89.530 82.000 89.680 89.550 ;
        RECT 90.130 89.350 94.080 89.550 ;
        RECT 95.380 89.350 99.330 89.550 ;
        RECT 90.130 88.900 90.730 89.350 ;
        RECT 98.730 88.900 99.330 89.350 ;
        RECT 90.130 88.750 94.080 88.900 ;
        RECT 95.380 88.750 99.330 88.900 ;
        RECT 90.130 88.300 90.730 88.750 ;
        RECT 98.730 88.300 99.330 88.750 ;
        RECT 90.130 88.150 94.080 88.300 ;
        RECT 95.380 88.150 99.330 88.300 ;
        RECT 90.130 87.700 90.730 88.150 ;
        RECT 98.730 87.700 99.330 88.150 ;
        RECT 90.130 87.550 94.080 87.700 ;
        RECT 95.380 87.550 99.330 87.700 ;
        RECT 90.130 87.100 90.730 87.550 ;
        RECT 98.730 87.100 99.330 87.550 ;
        RECT 90.130 86.950 94.080 87.100 ;
        RECT 95.380 86.950 99.330 87.100 ;
        RECT 90.130 86.500 90.730 86.950 ;
        RECT 98.730 86.500 99.330 86.950 ;
        RECT 90.130 86.350 94.080 86.500 ;
        RECT 95.380 86.350 99.330 86.500 ;
        RECT 90.130 85.900 90.730 86.350 ;
        RECT 98.730 85.900 99.330 86.350 ;
        RECT 90.130 85.750 94.080 85.900 ;
        RECT 95.380 85.750 99.330 85.900 ;
        RECT 90.130 85.300 90.730 85.750 ;
        RECT 98.730 85.300 99.330 85.750 ;
        RECT 90.130 85.150 94.080 85.300 ;
        RECT 95.380 85.150 99.330 85.300 ;
        RECT 90.130 84.700 90.730 85.150 ;
        RECT 98.730 84.700 99.330 85.150 ;
        RECT 90.130 84.550 94.080 84.700 ;
        RECT 95.380 84.550 99.330 84.700 ;
        RECT 90.130 84.100 90.730 84.550 ;
        RECT 98.730 84.100 99.330 84.550 ;
        RECT 90.130 83.950 94.080 84.100 ;
        RECT 95.380 83.950 99.330 84.100 ;
        RECT 90.130 83.500 90.730 83.950 ;
        RECT 98.730 83.500 99.330 83.950 ;
        RECT 90.130 83.350 94.080 83.500 ;
        RECT 95.380 83.350 99.330 83.500 ;
        RECT 90.130 82.900 90.730 83.350 ;
        RECT 98.730 82.900 99.330 83.350 ;
        RECT 90.130 82.750 94.080 82.900 ;
        RECT 95.380 82.750 99.330 82.900 ;
        RECT 90.130 82.300 90.730 82.750 ;
        RECT 98.730 82.300 99.330 82.750 ;
        RECT 90.130 82.150 94.080 82.300 ;
        RECT 95.380 82.150 99.330 82.300 ;
        RECT 90.130 82.000 90.730 82.150 ;
        RECT 86.530 81.700 90.730 82.000 ;
        RECT 98.730 82.000 99.330 82.150 ;
        RECT 99.780 82.000 99.930 89.550 ;
        RECT 100.380 82.000 100.530 89.550 ;
        RECT 100.980 82.000 101.130 89.550 ;
        RECT 101.580 82.000 101.730 89.550 ;
        RECT 102.180 82.000 102.330 89.550 ;
        RECT 102.780 82.000 102.930 84.900 ;
        RECT 98.730 81.700 102.930 82.000 ;
        RECT 86.530 81.550 94.080 81.700 ;
        RECT 95.380 81.550 102.930 81.700 ;
        RECT 86.530 81.350 90.730 81.550 ;
        RECT 80.330 81.050 89.130 81.200 ;
        RECT 89.280 81.050 90.730 81.350 ;
        RECT 78.730 80.150 90.730 81.050 ;
        RECT 98.730 81.350 102.930 81.550 ;
        RECT 98.730 81.050 100.180 81.350 ;
        RECT 103.530 81.200 105.930 84.400 ;
        RECT 106.530 82.000 106.680 84.900 ;
        RECT 107.130 82.000 107.280 89.550 ;
        RECT 107.730 82.000 107.880 89.550 ;
        RECT 108.330 82.000 108.480 89.550 ;
        RECT 108.930 82.000 109.080 89.550 ;
        RECT 109.530 82.000 109.680 89.550 ;
        RECT 110.130 89.350 114.080 89.550 ;
        RECT 115.380 89.350 119.330 89.550 ;
        RECT 110.130 88.900 110.730 89.350 ;
        RECT 118.730 88.900 119.330 89.350 ;
        RECT 110.130 88.750 114.080 88.900 ;
        RECT 115.380 88.750 119.330 88.900 ;
        RECT 110.130 88.300 110.730 88.750 ;
        RECT 118.730 88.300 119.330 88.750 ;
        RECT 110.130 88.150 114.080 88.300 ;
        RECT 115.380 88.150 119.330 88.300 ;
        RECT 110.130 87.700 110.730 88.150 ;
        RECT 118.730 87.700 119.330 88.150 ;
        RECT 110.130 87.550 114.080 87.700 ;
        RECT 115.380 87.550 119.330 87.700 ;
        RECT 110.130 87.100 110.730 87.550 ;
        RECT 118.730 87.100 119.330 87.550 ;
        RECT 110.130 86.950 114.080 87.100 ;
        RECT 115.380 86.950 119.330 87.100 ;
        RECT 110.130 86.500 110.730 86.950 ;
        RECT 118.730 86.500 119.330 86.950 ;
        RECT 110.130 86.350 114.080 86.500 ;
        RECT 115.380 86.350 119.330 86.500 ;
        RECT 110.130 85.900 110.730 86.350 ;
        RECT 118.730 85.900 119.330 86.350 ;
        RECT 110.130 85.750 114.080 85.900 ;
        RECT 115.380 85.750 119.330 85.900 ;
        RECT 110.130 85.300 110.730 85.750 ;
        RECT 118.730 85.300 119.330 85.750 ;
        RECT 110.130 85.150 114.080 85.300 ;
        RECT 115.380 85.150 119.330 85.300 ;
        RECT 110.130 84.700 110.730 85.150 ;
        RECT 118.730 84.700 119.330 85.150 ;
        RECT 110.130 84.550 114.080 84.700 ;
        RECT 115.380 84.550 119.330 84.700 ;
        RECT 110.130 84.100 110.730 84.550 ;
        RECT 118.730 84.100 119.330 84.550 ;
        RECT 110.130 83.950 114.080 84.100 ;
        RECT 115.380 83.950 119.330 84.100 ;
        RECT 110.130 83.500 110.730 83.950 ;
        RECT 118.730 83.500 119.330 83.950 ;
        RECT 110.130 83.350 114.080 83.500 ;
        RECT 115.380 83.350 119.330 83.500 ;
        RECT 110.130 82.900 110.730 83.350 ;
        RECT 118.730 82.900 119.330 83.350 ;
        RECT 110.130 82.750 114.080 82.900 ;
        RECT 115.380 82.750 119.330 82.900 ;
        RECT 110.130 82.300 110.730 82.750 ;
        RECT 118.730 82.300 119.330 82.750 ;
        RECT 110.130 82.150 114.080 82.300 ;
        RECT 115.380 82.150 119.330 82.300 ;
        RECT 110.130 82.000 110.730 82.150 ;
        RECT 106.530 81.700 110.730 82.000 ;
        RECT 118.730 82.000 119.330 82.150 ;
        RECT 119.780 82.000 119.930 89.550 ;
        RECT 120.380 82.000 120.530 89.550 ;
        RECT 120.980 82.000 121.130 89.550 ;
        RECT 121.580 82.000 121.730 89.550 ;
        RECT 122.180 82.000 122.330 89.550 ;
        RECT 122.780 82.000 122.930 84.900 ;
        RECT 118.730 81.700 122.930 82.000 ;
        RECT 106.530 81.550 114.080 81.700 ;
        RECT 115.380 81.550 122.930 81.700 ;
        RECT 106.530 81.350 110.730 81.550 ;
        RECT 100.330 81.050 109.130 81.200 ;
        RECT 109.280 81.050 110.730 81.350 ;
        RECT 98.730 80.150 110.730 81.050 ;
        RECT 118.730 81.350 122.930 81.550 ;
        RECT 123.530 83.040 124.730 84.400 ;
        RECT 123.530 81.765 127.135 83.040 ;
        RECT 118.730 81.050 120.180 81.350 ;
        RECT 123.530 81.200 124.730 81.765 ;
        RECT 120.330 81.050 124.730 81.200 ;
        RECT 118.730 80.150 124.730 81.050 ;
        RECT 4.730 79.850 9.130 80.150 ;
        RECT 20.330 79.850 29.130 80.150 ;
        RECT 40.330 79.850 49.130 80.150 ;
        RECT 60.330 79.850 69.130 80.150 ;
        RECT 80.330 79.850 89.130 80.150 ;
        RECT 100.330 79.850 109.130 80.150 ;
        RECT 4.730 78.950 10.730 79.850 ;
        RECT 20.330 79.800 30.730 79.850 ;
        RECT 40.330 79.800 50.730 79.850 ;
        RECT 60.330 79.800 70.730 79.850 ;
        RECT 80.330 79.800 90.730 79.850 ;
        RECT 100.330 79.800 110.730 79.850 ;
        RECT 120.330 79.800 124.730 80.150 ;
        RECT 4.730 78.800 9.130 78.950 ;
        RECT 4.730 77.965 5.930 78.800 ;
        RECT 9.280 78.650 10.730 78.950 ;
        RECT 2.315 76.690 5.930 77.965 ;
        RECT 4.730 75.600 5.930 76.690 ;
        RECT 6.530 78.450 10.730 78.650 ;
        RECT 18.730 78.950 30.730 79.800 ;
        RECT 18.730 78.900 29.130 78.950 ;
        RECT 18.730 78.650 20.180 78.900 ;
        RECT 20.330 78.800 29.130 78.900 ;
        RECT 18.730 78.450 22.930 78.650 ;
        RECT 6.530 78.300 14.080 78.450 ;
        RECT 15.430 78.300 22.930 78.450 ;
        RECT 6.530 78.000 10.730 78.300 ;
        RECT 2.315 73.250 4.315 75.545 ;
        RECT 6.530 75.150 6.680 78.000 ;
        RECT 7.130 70.450 7.280 78.000 ;
        RECT 7.730 70.450 7.880 78.000 ;
        RECT 8.330 70.450 8.480 78.000 ;
        RECT 8.930 70.450 9.080 78.000 ;
        RECT 9.530 70.450 9.680 78.000 ;
        RECT 10.130 77.850 10.730 78.000 ;
        RECT 18.730 78.000 22.930 78.300 ;
        RECT 18.730 77.850 19.330 78.000 ;
        RECT 10.130 77.700 14.080 77.850 ;
        RECT 15.380 77.700 19.330 77.850 ;
        RECT 10.130 77.250 10.730 77.700 ;
        RECT 18.730 77.250 19.330 77.700 ;
        RECT 10.130 77.100 14.080 77.250 ;
        RECT 15.380 77.100 19.330 77.250 ;
        RECT 10.130 76.650 10.730 77.100 ;
        RECT 18.730 76.650 19.330 77.100 ;
        RECT 10.130 76.500 14.080 76.650 ;
        RECT 15.380 76.500 19.330 76.650 ;
        RECT 10.130 76.050 10.730 76.500 ;
        RECT 18.730 76.050 19.330 76.500 ;
        RECT 10.130 75.900 14.080 76.050 ;
        RECT 15.380 75.900 19.330 76.050 ;
        RECT 10.130 75.450 10.730 75.900 ;
        RECT 18.730 75.450 19.330 75.900 ;
        RECT 10.130 75.300 14.080 75.450 ;
        RECT 15.380 75.300 19.330 75.450 ;
        RECT 10.130 74.850 10.730 75.300 ;
        RECT 18.730 74.850 19.330 75.300 ;
        RECT 10.130 74.700 14.080 74.850 ;
        RECT 15.380 74.700 19.330 74.850 ;
        RECT 10.130 74.250 10.730 74.700 ;
        RECT 18.730 74.250 19.330 74.700 ;
        RECT 10.130 74.100 14.080 74.250 ;
        RECT 15.380 74.100 19.330 74.250 ;
        RECT 10.130 73.650 10.730 74.100 ;
        RECT 18.730 73.650 19.330 74.100 ;
        RECT 10.130 73.500 14.080 73.650 ;
        RECT 15.380 73.500 19.330 73.650 ;
        RECT 10.130 73.050 10.730 73.500 ;
        RECT 18.730 73.050 19.330 73.500 ;
        RECT 10.130 72.900 14.080 73.050 ;
        RECT 15.380 72.900 19.330 73.050 ;
        RECT 10.130 72.450 10.730 72.900 ;
        RECT 18.730 72.450 19.330 72.900 ;
        RECT 10.130 72.300 14.080 72.450 ;
        RECT 15.380 72.300 19.330 72.450 ;
        RECT 10.130 71.850 10.730 72.300 ;
        RECT 18.730 71.850 19.330 72.300 ;
        RECT 10.130 71.700 14.080 71.850 ;
        RECT 15.380 71.700 19.330 71.850 ;
        RECT 10.130 71.250 10.730 71.700 ;
        RECT 18.730 71.250 19.330 71.700 ;
        RECT 10.130 71.100 14.080 71.250 ;
        RECT 15.380 71.100 19.330 71.250 ;
        RECT 10.130 70.650 10.730 71.100 ;
        RECT 18.730 70.650 19.330 71.100 ;
        RECT 10.130 70.450 14.080 70.650 ;
        RECT 15.380 70.450 19.330 70.650 ;
        RECT 19.780 70.450 19.930 78.000 ;
        RECT 20.380 70.450 20.530 78.000 ;
        RECT 20.980 70.450 21.130 78.000 ;
        RECT 21.580 70.450 21.730 78.000 ;
        RECT 22.180 70.450 22.330 78.000 ;
        RECT 22.780 75.150 22.930 78.000 ;
        RECT 23.530 75.600 25.930 78.800 ;
        RECT 29.280 78.650 30.730 78.950 ;
        RECT 26.530 78.450 30.730 78.650 ;
        RECT 38.730 78.950 50.730 79.800 ;
        RECT 38.730 78.900 49.130 78.950 ;
        RECT 38.730 78.650 40.180 78.900 ;
        RECT 40.330 78.800 49.130 78.900 ;
        RECT 38.730 78.450 42.930 78.650 ;
        RECT 26.530 78.300 34.080 78.450 ;
        RECT 35.430 78.300 42.930 78.450 ;
        RECT 26.530 78.000 30.730 78.300 ;
        RECT 26.530 75.150 26.680 78.000 ;
        RECT 27.130 70.450 27.280 78.000 ;
        RECT 27.730 70.450 27.880 78.000 ;
        RECT 28.330 70.450 28.480 78.000 ;
        RECT 28.930 70.450 29.080 78.000 ;
        RECT 29.530 70.450 29.680 78.000 ;
        RECT 30.130 77.850 30.730 78.000 ;
        RECT 38.730 78.000 42.930 78.300 ;
        RECT 38.730 77.850 39.330 78.000 ;
        RECT 30.130 77.700 34.080 77.850 ;
        RECT 35.380 77.700 39.330 77.850 ;
        RECT 30.130 77.250 30.730 77.700 ;
        RECT 38.730 77.250 39.330 77.700 ;
        RECT 30.130 77.100 34.080 77.250 ;
        RECT 35.380 77.100 39.330 77.250 ;
        RECT 30.130 76.650 30.730 77.100 ;
        RECT 38.730 76.650 39.330 77.100 ;
        RECT 30.130 76.500 34.080 76.650 ;
        RECT 35.380 76.500 39.330 76.650 ;
        RECT 30.130 76.050 30.730 76.500 ;
        RECT 38.730 76.050 39.330 76.500 ;
        RECT 30.130 75.900 34.080 76.050 ;
        RECT 35.380 75.900 39.330 76.050 ;
        RECT 30.130 75.450 30.730 75.900 ;
        RECT 38.730 75.450 39.330 75.900 ;
        RECT 30.130 75.300 34.080 75.450 ;
        RECT 35.380 75.300 39.330 75.450 ;
        RECT 30.130 74.850 30.730 75.300 ;
        RECT 38.730 74.850 39.330 75.300 ;
        RECT 30.130 74.700 34.080 74.850 ;
        RECT 35.380 74.700 39.330 74.850 ;
        RECT 30.130 74.250 30.730 74.700 ;
        RECT 38.730 74.250 39.330 74.700 ;
        RECT 30.130 74.100 34.080 74.250 ;
        RECT 35.380 74.100 39.330 74.250 ;
        RECT 30.130 73.650 30.730 74.100 ;
        RECT 38.730 73.650 39.330 74.100 ;
        RECT 30.130 73.500 34.080 73.650 ;
        RECT 35.380 73.500 39.330 73.650 ;
        RECT 30.130 73.050 30.730 73.500 ;
        RECT 38.730 73.050 39.330 73.500 ;
        RECT 30.130 72.900 34.080 73.050 ;
        RECT 35.380 72.900 39.330 73.050 ;
        RECT 30.130 72.450 30.730 72.900 ;
        RECT 38.730 72.450 39.330 72.900 ;
        RECT 30.130 72.300 34.080 72.450 ;
        RECT 35.380 72.300 39.330 72.450 ;
        RECT 30.130 71.850 30.730 72.300 ;
        RECT 38.730 71.850 39.330 72.300 ;
        RECT 30.130 71.700 34.080 71.850 ;
        RECT 35.380 71.700 39.330 71.850 ;
        RECT 30.130 71.250 30.730 71.700 ;
        RECT 38.730 71.250 39.330 71.700 ;
        RECT 30.130 71.100 34.080 71.250 ;
        RECT 35.380 71.100 39.330 71.250 ;
        RECT 30.130 70.650 30.730 71.100 ;
        RECT 38.730 70.650 39.330 71.100 ;
        RECT 30.130 70.450 34.080 70.650 ;
        RECT 35.380 70.450 39.330 70.650 ;
        RECT 39.780 70.450 39.930 78.000 ;
        RECT 40.380 70.450 40.530 78.000 ;
        RECT 40.980 70.450 41.130 78.000 ;
        RECT 41.580 70.450 41.730 78.000 ;
        RECT 42.180 70.450 42.330 78.000 ;
        RECT 42.780 75.150 42.930 78.000 ;
        RECT 43.530 75.600 45.930 78.800 ;
        RECT 49.280 78.650 50.730 78.950 ;
        RECT 46.530 78.450 50.730 78.650 ;
        RECT 58.730 78.950 70.730 79.800 ;
        RECT 58.730 78.900 69.130 78.950 ;
        RECT 58.730 78.650 60.180 78.900 ;
        RECT 60.330 78.800 69.130 78.900 ;
        RECT 58.730 78.450 62.930 78.650 ;
        RECT 46.530 78.300 54.080 78.450 ;
        RECT 55.430 78.300 62.930 78.450 ;
        RECT 46.530 78.000 50.730 78.300 ;
        RECT 46.530 75.150 46.680 78.000 ;
        RECT 47.130 70.450 47.280 78.000 ;
        RECT 47.730 70.450 47.880 78.000 ;
        RECT 48.330 70.450 48.480 78.000 ;
        RECT 48.930 70.450 49.080 78.000 ;
        RECT 49.530 70.450 49.680 78.000 ;
        RECT 50.130 77.850 50.730 78.000 ;
        RECT 58.730 78.000 62.930 78.300 ;
        RECT 58.730 77.850 59.330 78.000 ;
        RECT 50.130 77.700 54.080 77.850 ;
        RECT 55.380 77.700 59.330 77.850 ;
        RECT 50.130 77.250 50.730 77.700 ;
        RECT 58.730 77.250 59.330 77.700 ;
        RECT 50.130 77.100 54.080 77.250 ;
        RECT 55.380 77.100 59.330 77.250 ;
        RECT 50.130 76.650 50.730 77.100 ;
        RECT 58.730 76.650 59.330 77.100 ;
        RECT 50.130 76.500 54.080 76.650 ;
        RECT 55.380 76.500 59.330 76.650 ;
        RECT 50.130 76.050 50.730 76.500 ;
        RECT 58.730 76.050 59.330 76.500 ;
        RECT 50.130 75.900 54.080 76.050 ;
        RECT 55.380 75.900 59.330 76.050 ;
        RECT 50.130 75.450 50.730 75.900 ;
        RECT 58.730 75.450 59.330 75.900 ;
        RECT 50.130 75.300 54.080 75.450 ;
        RECT 55.380 75.300 59.330 75.450 ;
        RECT 50.130 74.850 50.730 75.300 ;
        RECT 58.730 74.850 59.330 75.300 ;
        RECT 50.130 74.700 54.080 74.850 ;
        RECT 55.380 74.700 59.330 74.850 ;
        RECT 50.130 74.250 50.730 74.700 ;
        RECT 58.730 74.250 59.330 74.700 ;
        RECT 50.130 74.100 54.080 74.250 ;
        RECT 55.380 74.100 59.330 74.250 ;
        RECT 50.130 73.650 50.730 74.100 ;
        RECT 58.730 73.650 59.330 74.100 ;
        RECT 50.130 73.500 54.080 73.650 ;
        RECT 55.380 73.500 59.330 73.650 ;
        RECT 50.130 73.050 50.730 73.500 ;
        RECT 58.730 73.050 59.330 73.500 ;
        RECT 50.130 72.900 54.080 73.050 ;
        RECT 55.380 72.900 59.330 73.050 ;
        RECT 50.130 72.450 50.730 72.900 ;
        RECT 58.730 72.450 59.330 72.900 ;
        RECT 50.130 72.300 54.080 72.450 ;
        RECT 55.380 72.300 59.330 72.450 ;
        RECT 50.130 71.850 50.730 72.300 ;
        RECT 58.730 71.850 59.330 72.300 ;
        RECT 50.130 71.700 54.080 71.850 ;
        RECT 55.380 71.700 59.330 71.850 ;
        RECT 50.130 71.250 50.730 71.700 ;
        RECT 58.730 71.250 59.330 71.700 ;
        RECT 50.130 71.100 54.080 71.250 ;
        RECT 55.380 71.100 59.330 71.250 ;
        RECT 50.130 70.650 50.730 71.100 ;
        RECT 58.730 70.650 59.330 71.100 ;
        RECT 50.130 70.450 54.080 70.650 ;
        RECT 55.380 70.450 59.330 70.650 ;
        RECT 59.780 70.450 59.930 78.000 ;
        RECT 60.380 70.450 60.530 78.000 ;
        RECT 60.980 70.450 61.130 78.000 ;
        RECT 61.580 70.450 61.730 78.000 ;
        RECT 62.180 70.450 62.330 78.000 ;
        RECT 62.780 75.150 62.930 78.000 ;
        RECT 63.530 75.600 65.930 78.800 ;
        RECT 69.280 78.650 70.730 78.950 ;
        RECT 66.530 78.450 70.730 78.650 ;
        RECT 78.730 78.950 90.730 79.800 ;
        RECT 78.730 78.900 89.130 78.950 ;
        RECT 78.730 78.650 80.180 78.900 ;
        RECT 80.330 78.800 89.130 78.900 ;
        RECT 78.730 78.450 82.930 78.650 ;
        RECT 66.530 78.300 74.080 78.450 ;
        RECT 75.430 78.300 82.930 78.450 ;
        RECT 66.530 78.000 70.730 78.300 ;
        RECT 66.530 75.150 66.680 78.000 ;
        RECT 67.130 70.450 67.280 78.000 ;
        RECT 67.730 70.450 67.880 78.000 ;
        RECT 68.330 70.450 68.480 78.000 ;
        RECT 68.930 70.450 69.080 78.000 ;
        RECT 69.530 70.450 69.680 78.000 ;
        RECT 70.130 77.850 70.730 78.000 ;
        RECT 78.730 78.000 82.930 78.300 ;
        RECT 78.730 77.850 79.330 78.000 ;
        RECT 70.130 77.700 74.080 77.850 ;
        RECT 75.380 77.700 79.330 77.850 ;
        RECT 70.130 77.250 70.730 77.700 ;
        RECT 78.730 77.250 79.330 77.700 ;
        RECT 70.130 77.100 74.080 77.250 ;
        RECT 75.380 77.100 79.330 77.250 ;
        RECT 70.130 76.650 70.730 77.100 ;
        RECT 78.730 76.650 79.330 77.100 ;
        RECT 70.130 76.500 74.080 76.650 ;
        RECT 75.380 76.500 79.330 76.650 ;
        RECT 70.130 76.050 70.730 76.500 ;
        RECT 78.730 76.050 79.330 76.500 ;
        RECT 70.130 75.900 74.080 76.050 ;
        RECT 75.380 75.900 79.330 76.050 ;
        RECT 70.130 75.450 70.730 75.900 ;
        RECT 78.730 75.450 79.330 75.900 ;
        RECT 70.130 75.300 74.080 75.450 ;
        RECT 75.380 75.300 79.330 75.450 ;
        RECT 70.130 74.850 70.730 75.300 ;
        RECT 78.730 74.850 79.330 75.300 ;
        RECT 70.130 74.700 74.080 74.850 ;
        RECT 75.380 74.700 79.330 74.850 ;
        RECT 70.130 74.250 70.730 74.700 ;
        RECT 78.730 74.250 79.330 74.700 ;
        RECT 70.130 74.100 74.080 74.250 ;
        RECT 75.380 74.100 79.330 74.250 ;
        RECT 70.130 73.650 70.730 74.100 ;
        RECT 78.730 73.650 79.330 74.100 ;
        RECT 70.130 73.500 74.080 73.650 ;
        RECT 75.380 73.500 79.330 73.650 ;
        RECT 70.130 73.050 70.730 73.500 ;
        RECT 78.730 73.050 79.330 73.500 ;
        RECT 70.130 72.900 74.080 73.050 ;
        RECT 75.380 72.900 79.330 73.050 ;
        RECT 70.130 72.450 70.730 72.900 ;
        RECT 78.730 72.450 79.330 72.900 ;
        RECT 70.130 72.300 74.080 72.450 ;
        RECT 75.380 72.300 79.330 72.450 ;
        RECT 70.130 71.850 70.730 72.300 ;
        RECT 78.730 71.850 79.330 72.300 ;
        RECT 70.130 71.700 74.080 71.850 ;
        RECT 75.380 71.700 79.330 71.850 ;
        RECT 70.130 71.250 70.730 71.700 ;
        RECT 78.730 71.250 79.330 71.700 ;
        RECT 70.130 71.100 74.080 71.250 ;
        RECT 75.380 71.100 79.330 71.250 ;
        RECT 70.130 70.650 70.730 71.100 ;
        RECT 78.730 70.650 79.330 71.100 ;
        RECT 70.130 70.450 74.080 70.650 ;
        RECT 75.380 70.450 79.330 70.650 ;
        RECT 79.780 70.450 79.930 78.000 ;
        RECT 80.380 70.450 80.530 78.000 ;
        RECT 80.980 70.450 81.130 78.000 ;
        RECT 81.580 70.450 81.730 78.000 ;
        RECT 82.180 70.450 82.330 78.000 ;
        RECT 82.780 75.150 82.930 78.000 ;
        RECT 83.530 75.600 85.930 78.800 ;
        RECT 89.280 78.650 90.730 78.950 ;
        RECT 86.530 78.450 90.730 78.650 ;
        RECT 98.730 78.950 110.730 79.800 ;
        RECT 98.730 78.900 109.130 78.950 ;
        RECT 98.730 78.650 100.180 78.900 ;
        RECT 100.330 78.800 109.130 78.900 ;
        RECT 98.730 78.450 102.930 78.650 ;
        RECT 86.530 78.300 94.080 78.450 ;
        RECT 95.430 78.300 102.930 78.450 ;
        RECT 86.530 78.000 90.730 78.300 ;
        RECT 86.530 75.150 86.680 78.000 ;
        RECT 87.130 70.450 87.280 78.000 ;
        RECT 87.730 70.450 87.880 78.000 ;
        RECT 88.330 70.450 88.480 78.000 ;
        RECT 88.930 70.450 89.080 78.000 ;
        RECT 89.530 70.450 89.680 78.000 ;
        RECT 90.130 77.850 90.730 78.000 ;
        RECT 98.730 78.000 102.930 78.300 ;
        RECT 98.730 77.850 99.330 78.000 ;
        RECT 90.130 77.700 94.080 77.850 ;
        RECT 95.380 77.700 99.330 77.850 ;
        RECT 90.130 77.250 90.730 77.700 ;
        RECT 98.730 77.250 99.330 77.700 ;
        RECT 90.130 77.100 94.080 77.250 ;
        RECT 95.380 77.100 99.330 77.250 ;
        RECT 90.130 76.650 90.730 77.100 ;
        RECT 98.730 76.650 99.330 77.100 ;
        RECT 90.130 76.500 94.080 76.650 ;
        RECT 95.380 76.500 99.330 76.650 ;
        RECT 90.130 76.050 90.730 76.500 ;
        RECT 98.730 76.050 99.330 76.500 ;
        RECT 90.130 75.900 94.080 76.050 ;
        RECT 95.380 75.900 99.330 76.050 ;
        RECT 90.130 75.450 90.730 75.900 ;
        RECT 98.730 75.450 99.330 75.900 ;
        RECT 90.130 75.300 94.080 75.450 ;
        RECT 95.380 75.300 99.330 75.450 ;
        RECT 90.130 74.850 90.730 75.300 ;
        RECT 98.730 74.850 99.330 75.300 ;
        RECT 90.130 74.700 94.080 74.850 ;
        RECT 95.380 74.700 99.330 74.850 ;
        RECT 90.130 74.250 90.730 74.700 ;
        RECT 98.730 74.250 99.330 74.700 ;
        RECT 90.130 74.100 94.080 74.250 ;
        RECT 95.380 74.100 99.330 74.250 ;
        RECT 90.130 73.650 90.730 74.100 ;
        RECT 98.730 73.650 99.330 74.100 ;
        RECT 90.130 73.500 94.080 73.650 ;
        RECT 95.380 73.500 99.330 73.650 ;
        RECT 90.130 73.050 90.730 73.500 ;
        RECT 98.730 73.050 99.330 73.500 ;
        RECT 90.130 72.900 94.080 73.050 ;
        RECT 95.380 72.900 99.330 73.050 ;
        RECT 90.130 72.450 90.730 72.900 ;
        RECT 98.730 72.450 99.330 72.900 ;
        RECT 90.130 72.300 94.080 72.450 ;
        RECT 95.380 72.300 99.330 72.450 ;
        RECT 90.130 71.850 90.730 72.300 ;
        RECT 98.730 71.850 99.330 72.300 ;
        RECT 90.130 71.700 94.080 71.850 ;
        RECT 95.380 71.700 99.330 71.850 ;
        RECT 90.130 71.250 90.730 71.700 ;
        RECT 98.730 71.250 99.330 71.700 ;
        RECT 90.130 71.100 94.080 71.250 ;
        RECT 95.380 71.100 99.330 71.250 ;
        RECT 90.130 70.650 90.730 71.100 ;
        RECT 98.730 70.650 99.330 71.100 ;
        RECT 90.130 70.450 94.080 70.650 ;
        RECT 95.380 70.450 99.330 70.650 ;
        RECT 99.780 70.450 99.930 78.000 ;
        RECT 100.380 70.450 100.530 78.000 ;
        RECT 100.980 70.450 101.130 78.000 ;
        RECT 101.580 70.450 101.730 78.000 ;
        RECT 102.180 70.450 102.330 78.000 ;
        RECT 102.780 75.150 102.930 78.000 ;
        RECT 103.530 75.600 105.930 78.800 ;
        RECT 109.280 78.650 110.730 78.950 ;
        RECT 106.530 78.450 110.730 78.650 ;
        RECT 118.730 78.900 124.730 79.800 ;
        RECT 118.730 78.650 120.180 78.900 ;
        RECT 120.330 78.800 124.730 78.900 ;
        RECT 118.730 78.450 122.930 78.650 ;
        RECT 106.530 78.300 114.080 78.450 ;
        RECT 115.430 78.300 122.930 78.450 ;
        RECT 106.530 78.000 110.730 78.300 ;
        RECT 106.530 75.150 106.680 78.000 ;
        RECT 107.130 70.450 107.280 78.000 ;
        RECT 107.730 70.450 107.880 78.000 ;
        RECT 108.330 70.450 108.480 78.000 ;
        RECT 108.930 70.450 109.080 78.000 ;
        RECT 109.530 70.450 109.680 78.000 ;
        RECT 110.130 77.850 110.730 78.000 ;
        RECT 118.730 78.000 122.930 78.300 ;
        RECT 118.730 77.850 119.330 78.000 ;
        RECT 110.130 77.700 114.080 77.850 ;
        RECT 115.380 77.700 119.330 77.850 ;
        RECT 110.130 77.250 110.730 77.700 ;
        RECT 118.730 77.250 119.330 77.700 ;
        RECT 110.130 77.100 114.080 77.250 ;
        RECT 115.380 77.100 119.330 77.250 ;
        RECT 110.130 76.650 110.730 77.100 ;
        RECT 118.730 76.650 119.330 77.100 ;
        RECT 110.130 76.500 114.080 76.650 ;
        RECT 115.380 76.500 119.330 76.650 ;
        RECT 110.130 76.050 110.730 76.500 ;
        RECT 118.730 76.050 119.330 76.500 ;
        RECT 110.130 75.900 114.080 76.050 ;
        RECT 115.380 75.900 119.330 76.050 ;
        RECT 110.130 75.450 110.730 75.900 ;
        RECT 118.730 75.450 119.330 75.900 ;
        RECT 110.130 75.300 114.080 75.450 ;
        RECT 115.380 75.300 119.330 75.450 ;
        RECT 110.130 74.850 110.730 75.300 ;
        RECT 118.730 74.850 119.330 75.300 ;
        RECT 110.130 74.700 114.080 74.850 ;
        RECT 115.380 74.700 119.330 74.850 ;
        RECT 110.130 74.250 110.730 74.700 ;
        RECT 118.730 74.250 119.330 74.700 ;
        RECT 110.130 74.100 114.080 74.250 ;
        RECT 115.380 74.100 119.330 74.250 ;
        RECT 110.130 73.650 110.730 74.100 ;
        RECT 118.730 73.650 119.330 74.100 ;
        RECT 110.130 73.500 114.080 73.650 ;
        RECT 115.380 73.500 119.330 73.650 ;
        RECT 110.130 73.050 110.730 73.500 ;
        RECT 118.730 73.050 119.330 73.500 ;
        RECT 110.130 72.900 114.080 73.050 ;
        RECT 115.380 72.900 119.330 73.050 ;
        RECT 110.130 72.450 110.730 72.900 ;
        RECT 118.730 72.450 119.330 72.900 ;
        RECT 110.130 72.300 114.080 72.450 ;
        RECT 115.380 72.300 119.330 72.450 ;
        RECT 110.130 71.850 110.730 72.300 ;
        RECT 118.730 71.850 119.330 72.300 ;
        RECT 110.130 71.700 114.080 71.850 ;
        RECT 115.380 71.700 119.330 71.850 ;
        RECT 110.130 71.250 110.730 71.700 ;
        RECT 118.730 71.250 119.330 71.700 ;
        RECT 110.130 71.100 114.080 71.250 ;
        RECT 115.380 71.100 119.330 71.250 ;
        RECT 110.130 70.650 110.730 71.100 ;
        RECT 118.730 70.650 119.330 71.100 ;
        RECT 110.130 70.450 114.080 70.650 ;
        RECT 115.380 70.450 119.330 70.650 ;
        RECT 119.780 70.450 119.930 78.000 ;
        RECT 120.380 70.450 120.530 78.000 ;
        RECT 120.980 70.450 121.130 78.000 ;
        RECT 121.580 70.450 121.730 78.000 ;
        RECT 122.180 70.450 122.330 78.000 ;
        RECT 122.780 75.150 122.930 78.000 ;
        RECT 123.530 77.185 124.730 78.800 ;
        RECT 123.530 75.910 127.135 77.185 ;
        RECT 123.530 75.600 124.730 75.910 ;
        RECT 2.315 64.450 4.315 66.745 ;
        RECT 4.730 63.635 5.930 64.400 ;
        RECT 2.315 62.360 5.930 63.635 ;
        RECT 4.730 61.200 5.930 62.360 ;
        RECT 6.530 62.000 6.680 64.900 ;
        RECT 7.130 62.000 7.280 69.550 ;
        RECT 7.730 62.000 7.880 69.550 ;
        RECT 8.330 62.000 8.480 69.550 ;
        RECT 8.930 62.000 9.080 69.550 ;
        RECT 9.530 62.000 9.680 69.550 ;
        RECT 10.130 69.350 14.080 69.550 ;
        RECT 15.380 69.350 19.330 69.550 ;
        RECT 10.130 68.900 10.730 69.350 ;
        RECT 18.730 68.900 19.330 69.350 ;
        RECT 10.130 68.750 14.080 68.900 ;
        RECT 15.380 68.750 19.330 68.900 ;
        RECT 10.130 68.300 10.730 68.750 ;
        RECT 18.730 68.300 19.330 68.750 ;
        RECT 10.130 68.150 14.080 68.300 ;
        RECT 15.380 68.150 19.330 68.300 ;
        RECT 10.130 67.700 10.730 68.150 ;
        RECT 18.730 67.700 19.330 68.150 ;
        RECT 10.130 67.550 14.080 67.700 ;
        RECT 15.380 67.550 19.330 67.700 ;
        RECT 10.130 67.100 10.730 67.550 ;
        RECT 18.730 67.100 19.330 67.550 ;
        RECT 10.130 66.950 14.080 67.100 ;
        RECT 15.380 66.950 19.330 67.100 ;
        RECT 10.130 66.500 10.730 66.950 ;
        RECT 18.730 66.500 19.330 66.950 ;
        RECT 10.130 66.350 14.080 66.500 ;
        RECT 15.380 66.350 19.330 66.500 ;
        RECT 10.130 65.900 10.730 66.350 ;
        RECT 18.730 65.900 19.330 66.350 ;
        RECT 10.130 65.750 14.080 65.900 ;
        RECT 15.380 65.750 19.330 65.900 ;
        RECT 10.130 65.300 10.730 65.750 ;
        RECT 18.730 65.300 19.330 65.750 ;
        RECT 10.130 65.150 14.080 65.300 ;
        RECT 15.380 65.150 19.330 65.300 ;
        RECT 10.130 64.700 10.730 65.150 ;
        RECT 18.730 64.700 19.330 65.150 ;
        RECT 10.130 64.550 14.080 64.700 ;
        RECT 15.380 64.550 19.330 64.700 ;
        RECT 10.130 64.100 10.730 64.550 ;
        RECT 18.730 64.100 19.330 64.550 ;
        RECT 10.130 63.950 14.080 64.100 ;
        RECT 15.380 63.950 19.330 64.100 ;
        RECT 10.130 63.500 10.730 63.950 ;
        RECT 18.730 63.500 19.330 63.950 ;
        RECT 10.130 63.350 14.080 63.500 ;
        RECT 15.380 63.350 19.330 63.500 ;
        RECT 10.130 62.900 10.730 63.350 ;
        RECT 18.730 62.900 19.330 63.350 ;
        RECT 10.130 62.750 14.080 62.900 ;
        RECT 15.380 62.750 19.330 62.900 ;
        RECT 10.130 62.300 10.730 62.750 ;
        RECT 18.730 62.300 19.330 62.750 ;
        RECT 10.130 62.150 14.080 62.300 ;
        RECT 15.380 62.150 19.330 62.300 ;
        RECT 10.130 62.000 10.730 62.150 ;
        RECT 6.530 61.700 10.730 62.000 ;
        RECT 18.730 62.000 19.330 62.150 ;
        RECT 19.780 62.000 19.930 69.550 ;
        RECT 20.380 62.000 20.530 69.550 ;
        RECT 20.980 62.000 21.130 69.550 ;
        RECT 21.580 62.000 21.730 69.550 ;
        RECT 22.180 62.000 22.330 69.550 ;
        RECT 22.780 62.000 22.930 64.900 ;
        RECT 18.730 61.700 22.930 62.000 ;
        RECT 6.530 61.550 14.080 61.700 ;
        RECT 15.380 61.550 22.930 61.700 ;
        RECT 6.530 61.350 10.730 61.550 ;
        RECT 4.730 61.050 9.130 61.200 ;
        RECT 9.280 61.050 10.730 61.350 ;
        RECT 4.730 60.150 10.730 61.050 ;
        RECT 18.730 61.350 22.930 61.550 ;
        RECT 18.730 61.050 20.180 61.350 ;
        RECT 23.530 61.200 25.930 64.400 ;
        RECT 26.530 62.000 26.680 64.900 ;
        RECT 27.130 62.000 27.280 69.550 ;
        RECT 27.730 62.000 27.880 69.550 ;
        RECT 28.330 62.000 28.480 69.550 ;
        RECT 28.930 62.000 29.080 69.550 ;
        RECT 29.530 62.000 29.680 69.550 ;
        RECT 30.130 69.350 34.080 69.550 ;
        RECT 35.380 69.350 39.330 69.550 ;
        RECT 30.130 68.900 30.730 69.350 ;
        RECT 38.730 68.900 39.330 69.350 ;
        RECT 30.130 68.750 34.080 68.900 ;
        RECT 35.380 68.750 39.330 68.900 ;
        RECT 30.130 68.300 30.730 68.750 ;
        RECT 38.730 68.300 39.330 68.750 ;
        RECT 30.130 68.150 34.080 68.300 ;
        RECT 35.380 68.150 39.330 68.300 ;
        RECT 30.130 67.700 30.730 68.150 ;
        RECT 38.730 67.700 39.330 68.150 ;
        RECT 30.130 67.550 34.080 67.700 ;
        RECT 35.380 67.550 39.330 67.700 ;
        RECT 30.130 67.100 30.730 67.550 ;
        RECT 38.730 67.100 39.330 67.550 ;
        RECT 30.130 66.950 34.080 67.100 ;
        RECT 35.380 66.950 39.330 67.100 ;
        RECT 30.130 66.500 30.730 66.950 ;
        RECT 38.730 66.500 39.330 66.950 ;
        RECT 30.130 66.350 34.080 66.500 ;
        RECT 35.380 66.350 39.330 66.500 ;
        RECT 30.130 65.900 30.730 66.350 ;
        RECT 38.730 65.900 39.330 66.350 ;
        RECT 30.130 65.750 34.080 65.900 ;
        RECT 35.380 65.750 39.330 65.900 ;
        RECT 30.130 65.300 30.730 65.750 ;
        RECT 38.730 65.300 39.330 65.750 ;
        RECT 30.130 65.150 34.080 65.300 ;
        RECT 35.380 65.150 39.330 65.300 ;
        RECT 30.130 64.700 30.730 65.150 ;
        RECT 38.730 64.700 39.330 65.150 ;
        RECT 30.130 64.550 34.080 64.700 ;
        RECT 35.380 64.550 39.330 64.700 ;
        RECT 30.130 64.100 30.730 64.550 ;
        RECT 38.730 64.100 39.330 64.550 ;
        RECT 30.130 63.950 34.080 64.100 ;
        RECT 35.380 63.950 39.330 64.100 ;
        RECT 30.130 63.500 30.730 63.950 ;
        RECT 38.730 63.500 39.330 63.950 ;
        RECT 30.130 63.350 34.080 63.500 ;
        RECT 35.380 63.350 39.330 63.500 ;
        RECT 30.130 62.900 30.730 63.350 ;
        RECT 38.730 62.900 39.330 63.350 ;
        RECT 30.130 62.750 34.080 62.900 ;
        RECT 35.380 62.750 39.330 62.900 ;
        RECT 30.130 62.300 30.730 62.750 ;
        RECT 38.730 62.300 39.330 62.750 ;
        RECT 30.130 62.150 34.080 62.300 ;
        RECT 35.380 62.150 39.330 62.300 ;
        RECT 30.130 62.000 30.730 62.150 ;
        RECT 26.530 61.700 30.730 62.000 ;
        RECT 38.730 62.000 39.330 62.150 ;
        RECT 39.780 62.000 39.930 69.550 ;
        RECT 40.380 62.000 40.530 69.550 ;
        RECT 40.980 62.000 41.130 69.550 ;
        RECT 41.580 62.000 41.730 69.550 ;
        RECT 42.180 62.000 42.330 69.550 ;
        RECT 42.780 62.000 42.930 64.900 ;
        RECT 38.730 61.700 42.930 62.000 ;
        RECT 26.530 61.550 34.080 61.700 ;
        RECT 35.380 61.550 42.930 61.700 ;
        RECT 26.530 61.350 30.730 61.550 ;
        RECT 20.330 61.050 29.130 61.200 ;
        RECT 29.280 61.050 30.730 61.350 ;
        RECT 18.730 60.150 30.730 61.050 ;
        RECT 38.730 61.350 42.930 61.550 ;
        RECT 38.730 61.050 40.180 61.350 ;
        RECT 43.530 61.200 45.930 64.400 ;
        RECT 46.530 62.000 46.680 64.900 ;
        RECT 47.130 62.000 47.280 69.550 ;
        RECT 47.730 62.000 47.880 69.550 ;
        RECT 48.330 62.000 48.480 69.550 ;
        RECT 48.930 62.000 49.080 69.550 ;
        RECT 49.530 62.000 49.680 69.550 ;
        RECT 50.130 69.350 54.080 69.550 ;
        RECT 55.380 69.350 59.330 69.550 ;
        RECT 50.130 68.900 50.730 69.350 ;
        RECT 58.730 68.900 59.330 69.350 ;
        RECT 50.130 68.750 54.080 68.900 ;
        RECT 55.380 68.750 59.330 68.900 ;
        RECT 50.130 68.300 50.730 68.750 ;
        RECT 58.730 68.300 59.330 68.750 ;
        RECT 50.130 68.150 54.080 68.300 ;
        RECT 55.380 68.150 59.330 68.300 ;
        RECT 50.130 67.700 50.730 68.150 ;
        RECT 58.730 67.700 59.330 68.150 ;
        RECT 50.130 67.550 54.080 67.700 ;
        RECT 55.380 67.550 59.330 67.700 ;
        RECT 50.130 67.100 50.730 67.550 ;
        RECT 58.730 67.100 59.330 67.550 ;
        RECT 50.130 66.950 54.080 67.100 ;
        RECT 55.380 66.950 59.330 67.100 ;
        RECT 50.130 66.500 50.730 66.950 ;
        RECT 58.730 66.500 59.330 66.950 ;
        RECT 50.130 66.350 54.080 66.500 ;
        RECT 55.380 66.350 59.330 66.500 ;
        RECT 50.130 65.900 50.730 66.350 ;
        RECT 58.730 65.900 59.330 66.350 ;
        RECT 50.130 65.750 54.080 65.900 ;
        RECT 55.380 65.750 59.330 65.900 ;
        RECT 50.130 65.300 50.730 65.750 ;
        RECT 58.730 65.300 59.330 65.750 ;
        RECT 50.130 65.150 54.080 65.300 ;
        RECT 55.380 65.150 59.330 65.300 ;
        RECT 50.130 64.700 50.730 65.150 ;
        RECT 58.730 64.700 59.330 65.150 ;
        RECT 50.130 64.550 54.080 64.700 ;
        RECT 55.380 64.550 59.330 64.700 ;
        RECT 50.130 64.100 50.730 64.550 ;
        RECT 58.730 64.100 59.330 64.550 ;
        RECT 50.130 63.950 54.080 64.100 ;
        RECT 55.380 63.950 59.330 64.100 ;
        RECT 50.130 63.500 50.730 63.950 ;
        RECT 58.730 63.500 59.330 63.950 ;
        RECT 50.130 63.350 54.080 63.500 ;
        RECT 55.380 63.350 59.330 63.500 ;
        RECT 50.130 62.900 50.730 63.350 ;
        RECT 58.730 62.900 59.330 63.350 ;
        RECT 50.130 62.750 54.080 62.900 ;
        RECT 55.380 62.750 59.330 62.900 ;
        RECT 50.130 62.300 50.730 62.750 ;
        RECT 58.730 62.300 59.330 62.750 ;
        RECT 50.130 62.150 54.080 62.300 ;
        RECT 55.380 62.150 59.330 62.300 ;
        RECT 50.130 62.000 50.730 62.150 ;
        RECT 46.530 61.700 50.730 62.000 ;
        RECT 58.730 62.000 59.330 62.150 ;
        RECT 59.780 62.000 59.930 69.550 ;
        RECT 60.380 62.000 60.530 69.550 ;
        RECT 60.980 62.000 61.130 69.550 ;
        RECT 61.580 62.000 61.730 69.550 ;
        RECT 62.180 62.000 62.330 69.550 ;
        RECT 62.780 62.000 62.930 64.900 ;
        RECT 58.730 61.700 62.930 62.000 ;
        RECT 46.530 61.550 54.080 61.700 ;
        RECT 55.380 61.550 62.930 61.700 ;
        RECT 46.530 61.350 50.730 61.550 ;
        RECT 40.330 61.050 49.130 61.200 ;
        RECT 49.280 61.050 50.730 61.350 ;
        RECT 38.730 60.150 50.730 61.050 ;
        RECT 58.730 61.350 62.930 61.550 ;
        RECT 58.730 61.050 60.180 61.350 ;
        RECT 63.530 61.200 65.930 64.400 ;
        RECT 66.530 62.000 66.680 64.900 ;
        RECT 67.130 62.000 67.280 69.550 ;
        RECT 67.730 62.000 67.880 69.550 ;
        RECT 68.330 62.000 68.480 69.550 ;
        RECT 68.930 62.000 69.080 69.550 ;
        RECT 69.530 62.000 69.680 69.550 ;
        RECT 70.130 69.350 74.080 69.550 ;
        RECT 75.380 69.350 79.330 69.550 ;
        RECT 70.130 68.900 70.730 69.350 ;
        RECT 78.730 68.900 79.330 69.350 ;
        RECT 70.130 68.750 74.080 68.900 ;
        RECT 75.380 68.750 79.330 68.900 ;
        RECT 70.130 68.300 70.730 68.750 ;
        RECT 78.730 68.300 79.330 68.750 ;
        RECT 70.130 68.150 74.080 68.300 ;
        RECT 75.380 68.150 79.330 68.300 ;
        RECT 70.130 67.700 70.730 68.150 ;
        RECT 78.730 67.700 79.330 68.150 ;
        RECT 70.130 67.550 74.080 67.700 ;
        RECT 75.380 67.550 79.330 67.700 ;
        RECT 70.130 67.100 70.730 67.550 ;
        RECT 78.730 67.100 79.330 67.550 ;
        RECT 70.130 66.950 74.080 67.100 ;
        RECT 75.380 66.950 79.330 67.100 ;
        RECT 70.130 66.500 70.730 66.950 ;
        RECT 78.730 66.500 79.330 66.950 ;
        RECT 70.130 66.350 74.080 66.500 ;
        RECT 75.380 66.350 79.330 66.500 ;
        RECT 70.130 65.900 70.730 66.350 ;
        RECT 78.730 65.900 79.330 66.350 ;
        RECT 70.130 65.750 74.080 65.900 ;
        RECT 75.380 65.750 79.330 65.900 ;
        RECT 70.130 65.300 70.730 65.750 ;
        RECT 78.730 65.300 79.330 65.750 ;
        RECT 70.130 65.150 74.080 65.300 ;
        RECT 75.380 65.150 79.330 65.300 ;
        RECT 70.130 64.700 70.730 65.150 ;
        RECT 78.730 64.700 79.330 65.150 ;
        RECT 70.130 64.550 74.080 64.700 ;
        RECT 75.380 64.550 79.330 64.700 ;
        RECT 70.130 64.100 70.730 64.550 ;
        RECT 78.730 64.100 79.330 64.550 ;
        RECT 70.130 63.950 74.080 64.100 ;
        RECT 75.380 63.950 79.330 64.100 ;
        RECT 70.130 63.500 70.730 63.950 ;
        RECT 78.730 63.500 79.330 63.950 ;
        RECT 70.130 63.350 74.080 63.500 ;
        RECT 75.380 63.350 79.330 63.500 ;
        RECT 70.130 62.900 70.730 63.350 ;
        RECT 78.730 62.900 79.330 63.350 ;
        RECT 70.130 62.750 74.080 62.900 ;
        RECT 75.380 62.750 79.330 62.900 ;
        RECT 70.130 62.300 70.730 62.750 ;
        RECT 78.730 62.300 79.330 62.750 ;
        RECT 70.130 62.150 74.080 62.300 ;
        RECT 75.380 62.150 79.330 62.300 ;
        RECT 70.130 62.000 70.730 62.150 ;
        RECT 66.530 61.700 70.730 62.000 ;
        RECT 78.730 62.000 79.330 62.150 ;
        RECT 79.780 62.000 79.930 69.550 ;
        RECT 80.380 62.000 80.530 69.550 ;
        RECT 80.980 62.000 81.130 69.550 ;
        RECT 81.580 62.000 81.730 69.550 ;
        RECT 82.180 62.000 82.330 69.550 ;
        RECT 82.780 62.000 82.930 64.900 ;
        RECT 78.730 61.700 82.930 62.000 ;
        RECT 66.530 61.550 74.080 61.700 ;
        RECT 75.380 61.550 82.930 61.700 ;
        RECT 66.530 61.350 70.730 61.550 ;
        RECT 60.330 61.050 69.130 61.200 ;
        RECT 69.280 61.050 70.730 61.350 ;
        RECT 58.730 60.150 70.730 61.050 ;
        RECT 78.730 61.350 82.930 61.550 ;
        RECT 78.730 61.050 80.180 61.350 ;
        RECT 83.530 61.200 85.930 64.400 ;
        RECT 86.530 62.000 86.680 64.900 ;
        RECT 87.130 62.000 87.280 69.550 ;
        RECT 87.730 62.000 87.880 69.550 ;
        RECT 88.330 62.000 88.480 69.550 ;
        RECT 88.930 62.000 89.080 69.550 ;
        RECT 89.530 62.000 89.680 69.550 ;
        RECT 90.130 69.350 94.080 69.550 ;
        RECT 95.380 69.350 99.330 69.550 ;
        RECT 90.130 68.900 90.730 69.350 ;
        RECT 98.730 68.900 99.330 69.350 ;
        RECT 90.130 68.750 94.080 68.900 ;
        RECT 95.380 68.750 99.330 68.900 ;
        RECT 90.130 68.300 90.730 68.750 ;
        RECT 98.730 68.300 99.330 68.750 ;
        RECT 90.130 68.150 94.080 68.300 ;
        RECT 95.380 68.150 99.330 68.300 ;
        RECT 90.130 67.700 90.730 68.150 ;
        RECT 98.730 67.700 99.330 68.150 ;
        RECT 90.130 67.550 94.080 67.700 ;
        RECT 95.380 67.550 99.330 67.700 ;
        RECT 90.130 67.100 90.730 67.550 ;
        RECT 98.730 67.100 99.330 67.550 ;
        RECT 90.130 66.950 94.080 67.100 ;
        RECT 95.380 66.950 99.330 67.100 ;
        RECT 90.130 66.500 90.730 66.950 ;
        RECT 98.730 66.500 99.330 66.950 ;
        RECT 90.130 66.350 94.080 66.500 ;
        RECT 95.380 66.350 99.330 66.500 ;
        RECT 90.130 65.900 90.730 66.350 ;
        RECT 98.730 65.900 99.330 66.350 ;
        RECT 90.130 65.750 94.080 65.900 ;
        RECT 95.380 65.750 99.330 65.900 ;
        RECT 90.130 65.300 90.730 65.750 ;
        RECT 98.730 65.300 99.330 65.750 ;
        RECT 90.130 65.150 94.080 65.300 ;
        RECT 95.380 65.150 99.330 65.300 ;
        RECT 90.130 64.700 90.730 65.150 ;
        RECT 98.730 64.700 99.330 65.150 ;
        RECT 90.130 64.550 94.080 64.700 ;
        RECT 95.380 64.550 99.330 64.700 ;
        RECT 90.130 64.100 90.730 64.550 ;
        RECT 98.730 64.100 99.330 64.550 ;
        RECT 90.130 63.950 94.080 64.100 ;
        RECT 95.380 63.950 99.330 64.100 ;
        RECT 90.130 63.500 90.730 63.950 ;
        RECT 98.730 63.500 99.330 63.950 ;
        RECT 90.130 63.350 94.080 63.500 ;
        RECT 95.380 63.350 99.330 63.500 ;
        RECT 90.130 62.900 90.730 63.350 ;
        RECT 98.730 62.900 99.330 63.350 ;
        RECT 90.130 62.750 94.080 62.900 ;
        RECT 95.380 62.750 99.330 62.900 ;
        RECT 90.130 62.300 90.730 62.750 ;
        RECT 98.730 62.300 99.330 62.750 ;
        RECT 90.130 62.150 94.080 62.300 ;
        RECT 95.380 62.150 99.330 62.300 ;
        RECT 90.130 62.000 90.730 62.150 ;
        RECT 86.530 61.700 90.730 62.000 ;
        RECT 98.730 62.000 99.330 62.150 ;
        RECT 99.780 62.000 99.930 69.550 ;
        RECT 100.380 62.000 100.530 69.550 ;
        RECT 100.980 62.000 101.130 69.550 ;
        RECT 101.580 62.000 101.730 69.550 ;
        RECT 102.180 62.000 102.330 69.550 ;
        RECT 102.780 62.000 102.930 64.900 ;
        RECT 98.730 61.700 102.930 62.000 ;
        RECT 86.530 61.550 94.080 61.700 ;
        RECT 95.380 61.550 102.930 61.700 ;
        RECT 86.530 61.350 90.730 61.550 ;
        RECT 80.330 61.050 89.130 61.200 ;
        RECT 89.280 61.050 90.730 61.350 ;
        RECT 78.730 60.150 90.730 61.050 ;
        RECT 98.730 61.350 102.930 61.550 ;
        RECT 98.730 61.050 100.180 61.350 ;
        RECT 103.530 61.200 105.930 64.400 ;
        RECT 106.530 62.000 106.680 64.900 ;
        RECT 107.130 62.000 107.280 69.550 ;
        RECT 107.730 62.000 107.880 69.550 ;
        RECT 108.330 62.000 108.480 69.550 ;
        RECT 108.930 62.000 109.080 69.550 ;
        RECT 109.530 62.000 109.680 69.550 ;
        RECT 110.130 69.350 114.080 69.550 ;
        RECT 115.380 69.350 119.330 69.550 ;
        RECT 110.130 68.900 110.730 69.350 ;
        RECT 118.730 68.900 119.330 69.350 ;
        RECT 110.130 68.750 114.080 68.900 ;
        RECT 115.380 68.750 119.330 68.900 ;
        RECT 110.130 68.300 110.730 68.750 ;
        RECT 118.730 68.300 119.330 68.750 ;
        RECT 110.130 68.150 114.080 68.300 ;
        RECT 115.380 68.150 119.330 68.300 ;
        RECT 110.130 67.700 110.730 68.150 ;
        RECT 118.730 67.700 119.330 68.150 ;
        RECT 110.130 67.550 114.080 67.700 ;
        RECT 115.380 67.550 119.330 67.700 ;
        RECT 110.130 67.100 110.730 67.550 ;
        RECT 118.730 67.100 119.330 67.550 ;
        RECT 110.130 66.950 114.080 67.100 ;
        RECT 115.380 66.950 119.330 67.100 ;
        RECT 110.130 66.500 110.730 66.950 ;
        RECT 118.730 66.500 119.330 66.950 ;
        RECT 110.130 66.350 114.080 66.500 ;
        RECT 115.380 66.350 119.330 66.500 ;
        RECT 110.130 65.900 110.730 66.350 ;
        RECT 118.730 65.900 119.330 66.350 ;
        RECT 110.130 65.750 114.080 65.900 ;
        RECT 115.380 65.750 119.330 65.900 ;
        RECT 110.130 65.300 110.730 65.750 ;
        RECT 118.730 65.300 119.330 65.750 ;
        RECT 110.130 65.150 114.080 65.300 ;
        RECT 115.380 65.150 119.330 65.300 ;
        RECT 110.130 64.700 110.730 65.150 ;
        RECT 118.730 64.700 119.330 65.150 ;
        RECT 110.130 64.550 114.080 64.700 ;
        RECT 115.380 64.550 119.330 64.700 ;
        RECT 110.130 64.100 110.730 64.550 ;
        RECT 118.730 64.100 119.330 64.550 ;
        RECT 110.130 63.950 114.080 64.100 ;
        RECT 115.380 63.950 119.330 64.100 ;
        RECT 110.130 63.500 110.730 63.950 ;
        RECT 118.730 63.500 119.330 63.950 ;
        RECT 110.130 63.350 114.080 63.500 ;
        RECT 115.380 63.350 119.330 63.500 ;
        RECT 110.130 62.900 110.730 63.350 ;
        RECT 118.730 62.900 119.330 63.350 ;
        RECT 110.130 62.750 114.080 62.900 ;
        RECT 115.380 62.750 119.330 62.900 ;
        RECT 110.130 62.300 110.730 62.750 ;
        RECT 118.730 62.300 119.330 62.750 ;
        RECT 110.130 62.150 114.080 62.300 ;
        RECT 115.380 62.150 119.330 62.300 ;
        RECT 110.130 62.000 110.730 62.150 ;
        RECT 106.530 61.700 110.730 62.000 ;
        RECT 118.730 62.000 119.330 62.150 ;
        RECT 119.780 62.000 119.930 69.550 ;
        RECT 120.380 62.000 120.530 69.550 ;
        RECT 120.980 62.000 121.130 69.550 ;
        RECT 121.580 62.000 121.730 69.550 ;
        RECT 122.180 62.000 122.330 69.550 ;
        RECT 122.780 62.000 122.930 64.900 ;
        RECT 118.730 61.700 122.930 62.000 ;
        RECT 106.530 61.550 114.080 61.700 ;
        RECT 115.380 61.550 122.930 61.700 ;
        RECT 106.530 61.350 110.730 61.550 ;
        RECT 100.330 61.050 109.130 61.200 ;
        RECT 109.280 61.050 110.730 61.350 ;
        RECT 98.730 60.150 110.730 61.050 ;
        RECT 118.730 61.350 122.930 61.550 ;
        RECT 123.530 63.380 124.730 64.400 ;
        RECT 123.530 62.105 127.135 63.380 ;
        RECT 118.730 61.050 120.180 61.350 ;
        RECT 123.530 61.200 124.730 62.105 ;
        RECT 120.330 61.050 124.730 61.200 ;
        RECT 118.730 60.150 124.730 61.050 ;
        RECT 4.730 59.850 9.130 60.150 ;
        RECT 20.330 59.850 29.130 60.150 ;
        RECT 40.330 59.850 49.130 60.150 ;
        RECT 60.330 59.850 69.130 60.150 ;
        RECT 80.330 59.850 89.130 60.150 ;
        RECT 100.330 59.850 109.130 60.150 ;
        RECT 4.730 58.950 10.730 59.850 ;
        RECT 20.330 59.800 30.730 59.850 ;
        RECT 40.330 59.800 50.730 59.850 ;
        RECT 60.330 59.800 70.730 59.850 ;
        RECT 80.330 59.800 90.730 59.850 ;
        RECT 100.330 59.800 110.730 59.850 ;
        RECT 120.330 59.800 124.730 60.150 ;
        RECT 4.730 58.800 9.130 58.950 ;
        RECT 4.730 57.555 5.930 58.800 ;
        RECT 9.280 58.650 10.730 58.950 ;
        RECT 2.315 56.280 5.930 57.555 ;
        RECT 4.730 55.600 5.930 56.280 ;
        RECT 6.530 58.450 10.730 58.650 ;
        RECT 18.730 58.950 30.730 59.800 ;
        RECT 18.730 58.900 29.130 58.950 ;
        RECT 18.730 58.650 20.180 58.900 ;
        RECT 20.330 58.800 29.130 58.900 ;
        RECT 18.730 58.450 22.930 58.650 ;
        RECT 6.530 58.300 14.080 58.450 ;
        RECT 15.430 58.300 22.930 58.450 ;
        RECT 6.530 58.000 10.730 58.300 ;
        RECT 2.315 53.250 4.315 55.545 ;
        RECT 6.530 55.150 6.680 58.000 ;
        RECT 7.130 50.450 7.280 58.000 ;
        RECT 7.730 50.450 7.880 58.000 ;
        RECT 8.330 50.450 8.480 58.000 ;
        RECT 8.930 50.450 9.080 58.000 ;
        RECT 9.530 50.450 9.680 58.000 ;
        RECT 10.130 57.850 10.730 58.000 ;
        RECT 18.730 58.000 22.930 58.300 ;
        RECT 18.730 57.850 19.330 58.000 ;
        RECT 10.130 57.700 14.080 57.850 ;
        RECT 15.380 57.700 19.330 57.850 ;
        RECT 10.130 57.250 10.730 57.700 ;
        RECT 18.730 57.250 19.330 57.700 ;
        RECT 10.130 57.100 14.080 57.250 ;
        RECT 15.380 57.100 19.330 57.250 ;
        RECT 10.130 56.650 10.730 57.100 ;
        RECT 18.730 56.650 19.330 57.100 ;
        RECT 10.130 56.500 14.080 56.650 ;
        RECT 15.380 56.500 19.330 56.650 ;
        RECT 10.130 56.050 10.730 56.500 ;
        RECT 18.730 56.050 19.330 56.500 ;
        RECT 10.130 55.900 14.080 56.050 ;
        RECT 15.380 55.900 19.330 56.050 ;
        RECT 10.130 55.450 10.730 55.900 ;
        RECT 18.730 55.450 19.330 55.900 ;
        RECT 10.130 55.300 14.080 55.450 ;
        RECT 15.380 55.300 19.330 55.450 ;
        RECT 10.130 54.850 10.730 55.300 ;
        RECT 18.730 54.850 19.330 55.300 ;
        RECT 10.130 54.700 14.080 54.850 ;
        RECT 15.380 54.700 19.330 54.850 ;
        RECT 10.130 54.250 10.730 54.700 ;
        RECT 18.730 54.250 19.330 54.700 ;
        RECT 10.130 54.100 14.080 54.250 ;
        RECT 15.380 54.100 19.330 54.250 ;
        RECT 10.130 53.650 10.730 54.100 ;
        RECT 18.730 53.650 19.330 54.100 ;
        RECT 10.130 53.500 14.080 53.650 ;
        RECT 15.380 53.500 19.330 53.650 ;
        RECT 10.130 53.050 10.730 53.500 ;
        RECT 18.730 53.050 19.330 53.500 ;
        RECT 10.130 52.900 14.080 53.050 ;
        RECT 15.380 52.900 19.330 53.050 ;
        RECT 10.130 52.450 10.730 52.900 ;
        RECT 18.730 52.450 19.330 52.900 ;
        RECT 10.130 52.300 14.080 52.450 ;
        RECT 15.380 52.300 19.330 52.450 ;
        RECT 10.130 51.850 10.730 52.300 ;
        RECT 18.730 51.850 19.330 52.300 ;
        RECT 10.130 51.700 14.080 51.850 ;
        RECT 15.380 51.700 19.330 51.850 ;
        RECT 10.130 51.250 10.730 51.700 ;
        RECT 18.730 51.250 19.330 51.700 ;
        RECT 10.130 51.100 14.080 51.250 ;
        RECT 15.380 51.100 19.330 51.250 ;
        RECT 10.130 50.650 10.730 51.100 ;
        RECT 18.730 50.650 19.330 51.100 ;
        RECT 10.130 50.450 14.080 50.650 ;
        RECT 15.380 50.450 19.330 50.650 ;
        RECT 19.780 50.450 19.930 58.000 ;
        RECT 20.380 50.450 20.530 58.000 ;
        RECT 20.980 50.450 21.130 58.000 ;
        RECT 21.580 50.450 21.730 58.000 ;
        RECT 22.180 50.450 22.330 58.000 ;
        RECT 22.780 55.150 22.930 58.000 ;
        RECT 23.530 55.600 25.930 58.800 ;
        RECT 29.280 58.650 30.730 58.950 ;
        RECT 26.530 58.450 30.730 58.650 ;
        RECT 38.730 58.950 50.730 59.800 ;
        RECT 38.730 58.900 49.130 58.950 ;
        RECT 38.730 58.650 40.180 58.900 ;
        RECT 40.330 58.800 49.130 58.900 ;
        RECT 38.730 58.450 42.930 58.650 ;
        RECT 26.530 58.300 34.080 58.450 ;
        RECT 35.430 58.300 42.930 58.450 ;
        RECT 26.530 58.000 30.730 58.300 ;
        RECT 26.530 55.150 26.680 58.000 ;
        RECT 27.130 50.450 27.280 58.000 ;
        RECT 27.730 50.450 27.880 58.000 ;
        RECT 28.330 50.450 28.480 58.000 ;
        RECT 28.930 50.450 29.080 58.000 ;
        RECT 29.530 50.450 29.680 58.000 ;
        RECT 30.130 57.850 30.730 58.000 ;
        RECT 38.730 58.000 42.930 58.300 ;
        RECT 38.730 57.850 39.330 58.000 ;
        RECT 30.130 57.700 34.080 57.850 ;
        RECT 35.380 57.700 39.330 57.850 ;
        RECT 30.130 57.250 30.730 57.700 ;
        RECT 38.730 57.250 39.330 57.700 ;
        RECT 30.130 57.100 34.080 57.250 ;
        RECT 35.380 57.100 39.330 57.250 ;
        RECT 30.130 56.650 30.730 57.100 ;
        RECT 38.730 56.650 39.330 57.100 ;
        RECT 30.130 56.500 34.080 56.650 ;
        RECT 35.380 56.500 39.330 56.650 ;
        RECT 30.130 56.050 30.730 56.500 ;
        RECT 38.730 56.050 39.330 56.500 ;
        RECT 30.130 55.900 34.080 56.050 ;
        RECT 35.380 55.900 39.330 56.050 ;
        RECT 30.130 55.450 30.730 55.900 ;
        RECT 38.730 55.450 39.330 55.900 ;
        RECT 30.130 55.300 34.080 55.450 ;
        RECT 35.380 55.300 39.330 55.450 ;
        RECT 30.130 54.850 30.730 55.300 ;
        RECT 38.730 54.850 39.330 55.300 ;
        RECT 30.130 54.700 34.080 54.850 ;
        RECT 35.380 54.700 39.330 54.850 ;
        RECT 30.130 54.250 30.730 54.700 ;
        RECT 38.730 54.250 39.330 54.700 ;
        RECT 30.130 54.100 34.080 54.250 ;
        RECT 35.380 54.100 39.330 54.250 ;
        RECT 30.130 53.650 30.730 54.100 ;
        RECT 38.730 53.650 39.330 54.100 ;
        RECT 30.130 53.500 34.080 53.650 ;
        RECT 35.380 53.500 39.330 53.650 ;
        RECT 30.130 53.050 30.730 53.500 ;
        RECT 38.730 53.050 39.330 53.500 ;
        RECT 30.130 52.900 34.080 53.050 ;
        RECT 35.380 52.900 39.330 53.050 ;
        RECT 30.130 52.450 30.730 52.900 ;
        RECT 38.730 52.450 39.330 52.900 ;
        RECT 30.130 52.300 34.080 52.450 ;
        RECT 35.380 52.300 39.330 52.450 ;
        RECT 30.130 51.850 30.730 52.300 ;
        RECT 38.730 51.850 39.330 52.300 ;
        RECT 30.130 51.700 34.080 51.850 ;
        RECT 35.380 51.700 39.330 51.850 ;
        RECT 30.130 51.250 30.730 51.700 ;
        RECT 38.730 51.250 39.330 51.700 ;
        RECT 30.130 51.100 34.080 51.250 ;
        RECT 35.380 51.100 39.330 51.250 ;
        RECT 30.130 50.650 30.730 51.100 ;
        RECT 38.730 50.650 39.330 51.100 ;
        RECT 30.130 50.450 34.080 50.650 ;
        RECT 35.380 50.450 39.330 50.650 ;
        RECT 39.780 50.450 39.930 58.000 ;
        RECT 40.380 50.450 40.530 58.000 ;
        RECT 40.980 50.450 41.130 58.000 ;
        RECT 41.580 50.450 41.730 58.000 ;
        RECT 42.180 50.450 42.330 58.000 ;
        RECT 42.780 55.150 42.930 58.000 ;
        RECT 43.530 55.600 45.930 58.800 ;
        RECT 49.280 58.650 50.730 58.950 ;
        RECT 46.530 58.450 50.730 58.650 ;
        RECT 58.730 58.950 70.730 59.800 ;
        RECT 58.730 58.900 69.130 58.950 ;
        RECT 58.730 58.650 60.180 58.900 ;
        RECT 60.330 58.800 69.130 58.900 ;
        RECT 58.730 58.450 62.930 58.650 ;
        RECT 46.530 58.300 54.080 58.450 ;
        RECT 55.430 58.300 62.930 58.450 ;
        RECT 46.530 58.000 50.730 58.300 ;
        RECT 46.530 55.150 46.680 58.000 ;
        RECT 47.130 50.450 47.280 58.000 ;
        RECT 47.730 50.450 47.880 58.000 ;
        RECT 48.330 50.450 48.480 58.000 ;
        RECT 48.930 50.450 49.080 58.000 ;
        RECT 49.530 50.450 49.680 58.000 ;
        RECT 50.130 57.850 50.730 58.000 ;
        RECT 58.730 58.000 62.930 58.300 ;
        RECT 58.730 57.850 59.330 58.000 ;
        RECT 50.130 57.700 54.080 57.850 ;
        RECT 55.380 57.700 59.330 57.850 ;
        RECT 50.130 57.250 50.730 57.700 ;
        RECT 58.730 57.250 59.330 57.700 ;
        RECT 50.130 57.100 54.080 57.250 ;
        RECT 55.380 57.100 59.330 57.250 ;
        RECT 50.130 56.650 50.730 57.100 ;
        RECT 58.730 56.650 59.330 57.100 ;
        RECT 50.130 56.500 54.080 56.650 ;
        RECT 55.380 56.500 59.330 56.650 ;
        RECT 50.130 56.050 50.730 56.500 ;
        RECT 58.730 56.050 59.330 56.500 ;
        RECT 50.130 55.900 54.080 56.050 ;
        RECT 55.380 55.900 59.330 56.050 ;
        RECT 50.130 55.450 50.730 55.900 ;
        RECT 58.730 55.450 59.330 55.900 ;
        RECT 50.130 55.300 54.080 55.450 ;
        RECT 55.380 55.300 59.330 55.450 ;
        RECT 50.130 54.850 50.730 55.300 ;
        RECT 58.730 54.850 59.330 55.300 ;
        RECT 50.130 54.700 54.080 54.850 ;
        RECT 55.380 54.700 59.330 54.850 ;
        RECT 50.130 54.250 50.730 54.700 ;
        RECT 58.730 54.250 59.330 54.700 ;
        RECT 50.130 54.100 54.080 54.250 ;
        RECT 55.380 54.100 59.330 54.250 ;
        RECT 50.130 53.650 50.730 54.100 ;
        RECT 58.730 53.650 59.330 54.100 ;
        RECT 50.130 53.500 54.080 53.650 ;
        RECT 55.380 53.500 59.330 53.650 ;
        RECT 50.130 53.050 50.730 53.500 ;
        RECT 58.730 53.050 59.330 53.500 ;
        RECT 50.130 52.900 54.080 53.050 ;
        RECT 55.380 52.900 59.330 53.050 ;
        RECT 50.130 52.450 50.730 52.900 ;
        RECT 58.730 52.450 59.330 52.900 ;
        RECT 50.130 52.300 54.080 52.450 ;
        RECT 55.380 52.300 59.330 52.450 ;
        RECT 50.130 51.850 50.730 52.300 ;
        RECT 58.730 51.850 59.330 52.300 ;
        RECT 50.130 51.700 54.080 51.850 ;
        RECT 55.380 51.700 59.330 51.850 ;
        RECT 50.130 51.250 50.730 51.700 ;
        RECT 58.730 51.250 59.330 51.700 ;
        RECT 50.130 51.100 54.080 51.250 ;
        RECT 55.380 51.100 59.330 51.250 ;
        RECT 50.130 50.650 50.730 51.100 ;
        RECT 58.730 50.650 59.330 51.100 ;
        RECT 50.130 50.450 54.080 50.650 ;
        RECT 55.380 50.450 59.330 50.650 ;
        RECT 59.780 50.450 59.930 58.000 ;
        RECT 60.380 50.450 60.530 58.000 ;
        RECT 60.980 50.450 61.130 58.000 ;
        RECT 61.580 50.450 61.730 58.000 ;
        RECT 62.180 50.450 62.330 58.000 ;
        RECT 62.780 55.150 62.930 58.000 ;
        RECT 63.530 55.600 65.930 58.800 ;
        RECT 69.280 58.650 70.730 58.950 ;
        RECT 66.530 58.450 70.730 58.650 ;
        RECT 78.730 58.950 90.730 59.800 ;
        RECT 78.730 58.900 89.130 58.950 ;
        RECT 78.730 58.650 80.180 58.900 ;
        RECT 80.330 58.800 89.130 58.900 ;
        RECT 78.730 58.450 82.930 58.650 ;
        RECT 66.530 58.300 74.080 58.450 ;
        RECT 75.430 58.300 82.930 58.450 ;
        RECT 66.530 58.000 70.730 58.300 ;
        RECT 66.530 55.150 66.680 58.000 ;
        RECT 67.130 50.450 67.280 58.000 ;
        RECT 67.730 50.450 67.880 58.000 ;
        RECT 68.330 50.450 68.480 58.000 ;
        RECT 68.930 50.450 69.080 58.000 ;
        RECT 69.530 50.450 69.680 58.000 ;
        RECT 70.130 57.850 70.730 58.000 ;
        RECT 78.730 58.000 82.930 58.300 ;
        RECT 78.730 57.850 79.330 58.000 ;
        RECT 70.130 57.700 74.080 57.850 ;
        RECT 75.380 57.700 79.330 57.850 ;
        RECT 70.130 57.250 70.730 57.700 ;
        RECT 78.730 57.250 79.330 57.700 ;
        RECT 70.130 57.100 74.080 57.250 ;
        RECT 75.380 57.100 79.330 57.250 ;
        RECT 70.130 56.650 70.730 57.100 ;
        RECT 78.730 56.650 79.330 57.100 ;
        RECT 70.130 56.500 74.080 56.650 ;
        RECT 75.380 56.500 79.330 56.650 ;
        RECT 70.130 56.050 70.730 56.500 ;
        RECT 78.730 56.050 79.330 56.500 ;
        RECT 70.130 55.900 74.080 56.050 ;
        RECT 75.380 55.900 79.330 56.050 ;
        RECT 70.130 55.450 70.730 55.900 ;
        RECT 78.730 55.450 79.330 55.900 ;
        RECT 70.130 55.300 74.080 55.450 ;
        RECT 75.380 55.300 79.330 55.450 ;
        RECT 70.130 54.850 70.730 55.300 ;
        RECT 78.730 54.850 79.330 55.300 ;
        RECT 70.130 54.700 74.080 54.850 ;
        RECT 75.380 54.700 79.330 54.850 ;
        RECT 70.130 54.250 70.730 54.700 ;
        RECT 78.730 54.250 79.330 54.700 ;
        RECT 70.130 54.100 74.080 54.250 ;
        RECT 75.380 54.100 79.330 54.250 ;
        RECT 70.130 53.650 70.730 54.100 ;
        RECT 78.730 53.650 79.330 54.100 ;
        RECT 70.130 53.500 74.080 53.650 ;
        RECT 75.380 53.500 79.330 53.650 ;
        RECT 70.130 53.050 70.730 53.500 ;
        RECT 78.730 53.050 79.330 53.500 ;
        RECT 70.130 52.900 74.080 53.050 ;
        RECT 75.380 52.900 79.330 53.050 ;
        RECT 70.130 52.450 70.730 52.900 ;
        RECT 78.730 52.450 79.330 52.900 ;
        RECT 70.130 52.300 74.080 52.450 ;
        RECT 75.380 52.300 79.330 52.450 ;
        RECT 70.130 51.850 70.730 52.300 ;
        RECT 78.730 51.850 79.330 52.300 ;
        RECT 70.130 51.700 74.080 51.850 ;
        RECT 75.380 51.700 79.330 51.850 ;
        RECT 70.130 51.250 70.730 51.700 ;
        RECT 78.730 51.250 79.330 51.700 ;
        RECT 70.130 51.100 74.080 51.250 ;
        RECT 75.380 51.100 79.330 51.250 ;
        RECT 70.130 50.650 70.730 51.100 ;
        RECT 78.730 50.650 79.330 51.100 ;
        RECT 70.130 50.450 74.080 50.650 ;
        RECT 75.380 50.450 79.330 50.650 ;
        RECT 79.780 50.450 79.930 58.000 ;
        RECT 80.380 50.450 80.530 58.000 ;
        RECT 80.980 50.450 81.130 58.000 ;
        RECT 81.580 50.450 81.730 58.000 ;
        RECT 82.180 50.450 82.330 58.000 ;
        RECT 82.780 55.150 82.930 58.000 ;
        RECT 83.530 55.600 85.930 58.800 ;
        RECT 89.280 58.650 90.730 58.950 ;
        RECT 86.530 58.450 90.730 58.650 ;
        RECT 98.730 58.950 110.730 59.800 ;
        RECT 98.730 58.900 109.130 58.950 ;
        RECT 98.730 58.650 100.180 58.900 ;
        RECT 100.330 58.800 109.130 58.900 ;
        RECT 98.730 58.450 102.930 58.650 ;
        RECT 86.530 58.300 94.080 58.450 ;
        RECT 95.430 58.300 102.930 58.450 ;
        RECT 86.530 58.000 90.730 58.300 ;
        RECT 86.530 55.150 86.680 58.000 ;
        RECT 87.130 50.450 87.280 58.000 ;
        RECT 87.730 50.450 87.880 58.000 ;
        RECT 88.330 50.450 88.480 58.000 ;
        RECT 88.930 50.450 89.080 58.000 ;
        RECT 89.530 50.450 89.680 58.000 ;
        RECT 90.130 57.850 90.730 58.000 ;
        RECT 98.730 58.000 102.930 58.300 ;
        RECT 98.730 57.850 99.330 58.000 ;
        RECT 90.130 57.700 94.080 57.850 ;
        RECT 95.380 57.700 99.330 57.850 ;
        RECT 90.130 57.250 90.730 57.700 ;
        RECT 98.730 57.250 99.330 57.700 ;
        RECT 90.130 57.100 94.080 57.250 ;
        RECT 95.380 57.100 99.330 57.250 ;
        RECT 90.130 56.650 90.730 57.100 ;
        RECT 98.730 56.650 99.330 57.100 ;
        RECT 90.130 56.500 94.080 56.650 ;
        RECT 95.380 56.500 99.330 56.650 ;
        RECT 90.130 56.050 90.730 56.500 ;
        RECT 98.730 56.050 99.330 56.500 ;
        RECT 90.130 55.900 94.080 56.050 ;
        RECT 95.380 55.900 99.330 56.050 ;
        RECT 90.130 55.450 90.730 55.900 ;
        RECT 98.730 55.450 99.330 55.900 ;
        RECT 90.130 55.300 94.080 55.450 ;
        RECT 95.380 55.300 99.330 55.450 ;
        RECT 90.130 54.850 90.730 55.300 ;
        RECT 98.730 54.850 99.330 55.300 ;
        RECT 90.130 54.700 94.080 54.850 ;
        RECT 95.380 54.700 99.330 54.850 ;
        RECT 90.130 54.250 90.730 54.700 ;
        RECT 98.730 54.250 99.330 54.700 ;
        RECT 90.130 54.100 94.080 54.250 ;
        RECT 95.380 54.100 99.330 54.250 ;
        RECT 90.130 53.650 90.730 54.100 ;
        RECT 98.730 53.650 99.330 54.100 ;
        RECT 90.130 53.500 94.080 53.650 ;
        RECT 95.380 53.500 99.330 53.650 ;
        RECT 90.130 53.050 90.730 53.500 ;
        RECT 98.730 53.050 99.330 53.500 ;
        RECT 90.130 52.900 94.080 53.050 ;
        RECT 95.380 52.900 99.330 53.050 ;
        RECT 90.130 52.450 90.730 52.900 ;
        RECT 98.730 52.450 99.330 52.900 ;
        RECT 90.130 52.300 94.080 52.450 ;
        RECT 95.380 52.300 99.330 52.450 ;
        RECT 90.130 51.850 90.730 52.300 ;
        RECT 98.730 51.850 99.330 52.300 ;
        RECT 90.130 51.700 94.080 51.850 ;
        RECT 95.380 51.700 99.330 51.850 ;
        RECT 90.130 51.250 90.730 51.700 ;
        RECT 98.730 51.250 99.330 51.700 ;
        RECT 90.130 51.100 94.080 51.250 ;
        RECT 95.380 51.100 99.330 51.250 ;
        RECT 90.130 50.650 90.730 51.100 ;
        RECT 98.730 50.650 99.330 51.100 ;
        RECT 90.130 50.450 94.080 50.650 ;
        RECT 95.380 50.450 99.330 50.650 ;
        RECT 99.780 50.450 99.930 58.000 ;
        RECT 100.380 50.450 100.530 58.000 ;
        RECT 100.980 50.450 101.130 58.000 ;
        RECT 101.580 50.450 101.730 58.000 ;
        RECT 102.180 50.450 102.330 58.000 ;
        RECT 102.780 55.150 102.930 58.000 ;
        RECT 103.530 55.600 105.930 58.800 ;
        RECT 109.280 58.650 110.730 58.950 ;
        RECT 106.530 58.450 110.730 58.650 ;
        RECT 118.730 58.900 124.730 59.800 ;
        RECT 118.730 58.650 120.180 58.900 ;
        RECT 120.330 58.800 124.730 58.900 ;
        RECT 118.730 58.450 122.930 58.650 ;
        RECT 106.530 58.300 114.080 58.450 ;
        RECT 115.430 58.300 122.930 58.450 ;
        RECT 106.530 58.000 110.730 58.300 ;
        RECT 106.530 55.150 106.680 58.000 ;
        RECT 107.130 50.450 107.280 58.000 ;
        RECT 107.730 50.450 107.880 58.000 ;
        RECT 108.330 50.450 108.480 58.000 ;
        RECT 108.930 50.450 109.080 58.000 ;
        RECT 109.530 50.450 109.680 58.000 ;
        RECT 110.130 57.850 110.730 58.000 ;
        RECT 118.730 58.000 122.930 58.300 ;
        RECT 118.730 57.850 119.330 58.000 ;
        RECT 110.130 57.700 114.080 57.850 ;
        RECT 115.380 57.700 119.330 57.850 ;
        RECT 110.130 57.250 110.730 57.700 ;
        RECT 118.730 57.250 119.330 57.700 ;
        RECT 110.130 57.100 114.080 57.250 ;
        RECT 115.380 57.100 119.330 57.250 ;
        RECT 110.130 56.650 110.730 57.100 ;
        RECT 118.730 56.650 119.330 57.100 ;
        RECT 110.130 56.500 114.080 56.650 ;
        RECT 115.380 56.500 119.330 56.650 ;
        RECT 110.130 56.050 110.730 56.500 ;
        RECT 118.730 56.050 119.330 56.500 ;
        RECT 110.130 55.900 114.080 56.050 ;
        RECT 115.380 55.900 119.330 56.050 ;
        RECT 110.130 55.450 110.730 55.900 ;
        RECT 118.730 55.450 119.330 55.900 ;
        RECT 110.130 55.300 114.080 55.450 ;
        RECT 115.380 55.300 119.330 55.450 ;
        RECT 110.130 54.850 110.730 55.300 ;
        RECT 118.730 54.850 119.330 55.300 ;
        RECT 110.130 54.700 114.080 54.850 ;
        RECT 115.380 54.700 119.330 54.850 ;
        RECT 110.130 54.250 110.730 54.700 ;
        RECT 118.730 54.250 119.330 54.700 ;
        RECT 110.130 54.100 114.080 54.250 ;
        RECT 115.380 54.100 119.330 54.250 ;
        RECT 110.130 53.650 110.730 54.100 ;
        RECT 118.730 53.650 119.330 54.100 ;
        RECT 110.130 53.500 114.080 53.650 ;
        RECT 115.380 53.500 119.330 53.650 ;
        RECT 110.130 53.050 110.730 53.500 ;
        RECT 118.730 53.050 119.330 53.500 ;
        RECT 110.130 52.900 114.080 53.050 ;
        RECT 115.380 52.900 119.330 53.050 ;
        RECT 110.130 52.450 110.730 52.900 ;
        RECT 118.730 52.450 119.330 52.900 ;
        RECT 110.130 52.300 114.080 52.450 ;
        RECT 115.380 52.300 119.330 52.450 ;
        RECT 110.130 51.850 110.730 52.300 ;
        RECT 118.730 51.850 119.330 52.300 ;
        RECT 110.130 51.700 114.080 51.850 ;
        RECT 115.380 51.700 119.330 51.850 ;
        RECT 110.130 51.250 110.730 51.700 ;
        RECT 118.730 51.250 119.330 51.700 ;
        RECT 110.130 51.100 114.080 51.250 ;
        RECT 115.380 51.100 119.330 51.250 ;
        RECT 110.130 50.650 110.730 51.100 ;
        RECT 118.730 50.650 119.330 51.100 ;
        RECT 110.130 50.450 114.080 50.650 ;
        RECT 115.380 50.450 119.330 50.650 ;
        RECT 119.780 50.450 119.930 58.000 ;
        RECT 120.380 50.450 120.530 58.000 ;
        RECT 120.980 50.450 121.130 58.000 ;
        RECT 121.580 50.450 121.730 58.000 ;
        RECT 122.180 50.450 122.330 58.000 ;
        RECT 122.780 55.150 122.930 58.000 ;
        RECT 123.530 57.310 124.730 58.800 ;
        RECT 123.530 56.035 127.135 57.310 ;
        RECT 123.530 55.600 124.730 56.035 ;
        RECT 2.315 44.450 4.315 46.745 ;
        RECT 4.730 43.230 5.930 44.400 ;
        RECT 2.315 41.955 5.930 43.230 ;
        RECT 4.730 41.200 5.930 41.955 ;
        RECT 6.530 42.000 6.680 44.900 ;
        RECT 7.130 42.000 7.280 49.550 ;
        RECT 7.730 42.000 7.880 49.550 ;
        RECT 8.330 42.000 8.480 49.550 ;
        RECT 8.930 42.000 9.080 49.550 ;
        RECT 9.530 42.000 9.680 49.550 ;
        RECT 10.130 49.350 14.080 49.550 ;
        RECT 15.380 49.350 19.330 49.550 ;
        RECT 10.130 48.900 10.730 49.350 ;
        RECT 18.730 48.900 19.330 49.350 ;
        RECT 10.130 48.750 14.080 48.900 ;
        RECT 15.380 48.750 19.330 48.900 ;
        RECT 10.130 48.300 10.730 48.750 ;
        RECT 18.730 48.300 19.330 48.750 ;
        RECT 10.130 48.150 14.080 48.300 ;
        RECT 15.380 48.150 19.330 48.300 ;
        RECT 10.130 47.700 10.730 48.150 ;
        RECT 18.730 47.700 19.330 48.150 ;
        RECT 10.130 47.550 14.080 47.700 ;
        RECT 15.380 47.550 19.330 47.700 ;
        RECT 10.130 47.100 10.730 47.550 ;
        RECT 18.730 47.100 19.330 47.550 ;
        RECT 10.130 46.950 14.080 47.100 ;
        RECT 15.380 46.950 19.330 47.100 ;
        RECT 10.130 46.500 10.730 46.950 ;
        RECT 18.730 46.500 19.330 46.950 ;
        RECT 10.130 46.350 14.080 46.500 ;
        RECT 15.380 46.350 19.330 46.500 ;
        RECT 10.130 45.900 10.730 46.350 ;
        RECT 18.730 45.900 19.330 46.350 ;
        RECT 10.130 45.750 14.080 45.900 ;
        RECT 15.380 45.750 19.330 45.900 ;
        RECT 10.130 45.300 10.730 45.750 ;
        RECT 18.730 45.300 19.330 45.750 ;
        RECT 10.130 45.150 14.080 45.300 ;
        RECT 15.380 45.150 19.330 45.300 ;
        RECT 10.130 44.700 10.730 45.150 ;
        RECT 18.730 44.700 19.330 45.150 ;
        RECT 10.130 44.550 14.080 44.700 ;
        RECT 15.380 44.550 19.330 44.700 ;
        RECT 10.130 44.100 10.730 44.550 ;
        RECT 18.730 44.100 19.330 44.550 ;
        RECT 10.130 43.950 14.080 44.100 ;
        RECT 15.380 43.950 19.330 44.100 ;
        RECT 10.130 43.500 10.730 43.950 ;
        RECT 18.730 43.500 19.330 43.950 ;
        RECT 10.130 43.350 14.080 43.500 ;
        RECT 15.380 43.350 19.330 43.500 ;
        RECT 10.130 42.900 10.730 43.350 ;
        RECT 18.730 42.900 19.330 43.350 ;
        RECT 10.130 42.750 14.080 42.900 ;
        RECT 15.380 42.750 19.330 42.900 ;
        RECT 10.130 42.300 10.730 42.750 ;
        RECT 18.730 42.300 19.330 42.750 ;
        RECT 10.130 42.150 14.080 42.300 ;
        RECT 15.380 42.150 19.330 42.300 ;
        RECT 10.130 42.000 10.730 42.150 ;
        RECT 6.530 41.700 10.730 42.000 ;
        RECT 18.730 42.000 19.330 42.150 ;
        RECT 19.780 42.000 19.930 49.550 ;
        RECT 20.380 42.000 20.530 49.550 ;
        RECT 20.980 42.000 21.130 49.550 ;
        RECT 21.580 42.000 21.730 49.550 ;
        RECT 22.180 42.000 22.330 49.550 ;
        RECT 22.780 42.000 22.930 44.900 ;
        RECT 18.730 41.700 22.930 42.000 ;
        RECT 6.530 41.550 14.080 41.700 ;
        RECT 15.380 41.550 22.930 41.700 ;
        RECT 6.530 41.350 10.730 41.550 ;
        RECT 4.730 41.050 9.130 41.200 ;
        RECT 9.280 41.050 10.730 41.350 ;
        RECT 4.730 40.150 10.730 41.050 ;
        RECT 18.730 41.350 22.930 41.550 ;
        RECT 18.730 41.050 20.180 41.350 ;
        RECT 23.530 41.200 25.930 44.400 ;
        RECT 26.530 42.000 26.680 44.900 ;
        RECT 27.130 42.000 27.280 49.550 ;
        RECT 27.730 42.000 27.880 49.550 ;
        RECT 28.330 42.000 28.480 49.550 ;
        RECT 28.930 42.000 29.080 49.550 ;
        RECT 29.530 42.000 29.680 49.550 ;
        RECT 30.130 49.350 34.080 49.550 ;
        RECT 35.380 49.350 39.330 49.550 ;
        RECT 30.130 48.900 30.730 49.350 ;
        RECT 38.730 48.900 39.330 49.350 ;
        RECT 30.130 48.750 34.080 48.900 ;
        RECT 35.380 48.750 39.330 48.900 ;
        RECT 30.130 48.300 30.730 48.750 ;
        RECT 38.730 48.300 39.330 48.750 ;
        RECT 30.130 48.150 34.080 48.300 ;
        RECT 35.380 48.150 39.330 48.300 ;
        RECT 30.130 47.700 30.730 48.150 ;
        RECT 38.730 47.700 39.330 48.150 ;
        RECT 30.130 47.550 34.080 47.700 ;
        RECT 35.380 47.550 39.330 47.700 ;
        RECT 30.130 47.100 30.730 47.550 ;
        RECT 38.730 47.100 39.330 47.550 ;
        RECT 30.130 46.950 34.080 47.100 ;
        RECT 35.380 46.950 39.330 47.100 ;
        RECT 30.130 46.500 30.730 46.950 ;
        RECT 38.730 46.500 39.330 46.950 ;
        RECT 30.130 46.350 34.080 46.500 ;
        RECT 35.380 46.350 39.330 46.500 ;
        RECT 30.130 45.900 30.730 46.350 ;
        RECT 38.730 45.900 39.330 46.350 ;
        RECT 30.130 45.750 34.080 45.900 ;
        RECT 35.380 45.750 39.330 45.900 ;
        RECT 30.130 45.300 30.730 45.750 ;
        RECT 38.730 45.300 39.330 45.750 ;
        RECT 30.130 45.150 34.080 45.300 ;
        RECT 35.380 45.150 39.330 45.300 ;
        RECT 30.130 44.700 30.730 45.150 ;
        RECT 38.730 44.700 39.330 45.150 ;
        RECT 30.130 44.550 34.080 44.700 ;
        RECT 35.380 44.550 39.330 44.700 ;
        RECT 30.130 44.100 30.730 44.550 ;
        RECT 38.730 44.100 39.330 44.550 ;
        RECT 30.130 43.950 34.080 44.100 ;
        RECT 35.380 43.950 39.330 44.100 ;
        RECT 30.130 43.500 30.730 43.950 ;
        RECT 38.730 43.500 39.330 43.950 ;
        RECT 30.130 43.350 34.080 43.500 ;
        RECT 35.380 43.350 39.330 43.500 ;
        RECT 30.130 42.900 30.730 43.350 ;
        RECT 38.730 42.900 39.330 43.350 ;
        RECT 30.130 42.750 34.080 42.900 ;
        RECT 35.380 42.750 39.330 42.900 ;
        RECT 30.130 42.300 30.730 42.750 ;
        RECT 38.730 42.300 39.330 42.750 ;
        RECT 30.130 42.150 34.080 42.300 ;
        RECT 35.380 42.150 39.330 42.300 ;
        RECT 30.130 42.000 30.730 42.150 ;
        RECT 26.530 41.700 30.730 42.000 ;
        RECT 38.730 42.000 39.330 42.150 ;
        RECT 39.780 42.000 39.930 49.550 ;
        RECT 40.380 42.000 40.530 49.550 ;
        RECT 40.980 42.000 41.130 49.550 ;
        RECT 41.580 42.000 41.730 49.550 ;
        RECT 42.180 42.000 42.330 49.550 ;
        RECT 42.780 42.000 42.930 44.900 ;
        RECT 38.730 41.700 42.930 42.000 ;
        RECT 26.530 41.550 34.080 41.700 ;
        RECT 35.380 41.550 42.930 41.700 ;
        RECT 26.530 41.350 30.730 41.550 ;
        RECT 20.330 41.050 29.130 41.200 ;
        RECT 29.280 41.050 30.730 41.350 ;
        RECT 18.730 40.150 30.730 41.050 ;
        RECT 38.730 41.350 42.930 41.550 ;
        RECT 38.730 41.050 40.180 41.350 ;
        RECT 43.530 41.200 45.930 44.400 ;
        RECT 46.530 42.000 46.680 44.900 ;
        RECT 47.130 42.000 47.280 49.550 ;
        RECT 47.730 42.000 47.880 49.550 ;
        RECT 48.330 42.000 48.480 49.550 ;
        RECT 48.930 42.000 49.080 49.550 ;
        RECT 49.530 42.000 49.680 49.550 ;
        RECT 50.130 49.350 54.080 49.550 ;
        RECT 55.380 49.350 59.330 49.550 ;
        RECT 50.130 48.900 50.730 49.350 ;
        RECT 58.730 48.900 59.330 49.350 ;
        RECT 50.130 48.750 54.080 48.900 ;
        RECT 55.380 48.750 59.330 48.900 ;
        RECT 50.130 48.300 50.730 48.750 ;
        RECT 58.730 48.300 59.330 48.750 ;
        RECT 50.130 48.150 54.080 48.300 ;
        RECT 55.380 48.150 59.330 48.300 ;
        RECT 50.130 47.700 50.730 48.150 ;
        RECT 58.730 47.700 59.330 48.150 ;
        RECT 50.130 47.550 54.080 47.700 ;
        RECT 55.380 47.550 59.330 47.700 ;
        RECT 50.130 47.100 50.730 47.550 ;
        RECT 58.730 47.100 59.330 47.550 ;
        RECT 50.130 46.950 54.080 47.100 ;
        RECT 55.380 46.950 59.330 47.100 ;
        RECT 50.130 46.500 50.730 46.950 ;
        RECT 58.730 46.500 59.330 46.950 ;
        RECT 50.130 46.350 54.080 46.500 ;
        RECT 55.380 46.350 59.330 46.500 ;
        RECT 50.130 45.900 50.730 46.350 ;
        RECT 58.730 45.900 59.330 46.350 ;
        RECT 50.130 45.750 54.080 45.900 ;
        RECT 55.380 45.750 59.330 45.900 ;
        RECT 50.130 45.300 50.730 45.750 ;
        RECT 58.730 45.300 59.330 45.750 ;
        RECT 50.130 45.150 54.080 45.300 ;
        RECT 55.380 45.150 59.330 45.300 ;
        RECT 50.130 44.700 50.730 45.150 ;
        RECT 58.730 44.700 59.330 45.150 ;
        RECT 50.130 44.550 54.080 44.700 ;
        RECT 55.380 44.550 59.330 44.700 ;
        RECT 50.130 44.100 50.730 44.550 ;
        RECT 58.730 44.100 59.330 44.550 ;
        RECT 50.130 43.950 54.080 44.100 ;
        RECT 55.380 43.950 59.330 44.100 ;
        RECT 50.130 43.500 50.730 43.950 ;
        RECT 58.730 43.500 59.330 43.950 ;
        RECT 50.130 43.350 54.080 43.500 ;
        RECT 55.380 43.350 59.330 43.500 ;
        RECT 50.130 42.900 50.730 43.350 ;
        RECT 58.730 42.900 59.330 43.350 ;
        RECT 50.130 42.750 54.080 42.900 ;
        RECT 55.380 42.750 59.330 42.900 ;
        RECT 50.130 42.300 50.730 42.750 ;
        RECT 58.730 42.300 59.330 42.750 ;
        RECT 50.130 42.150 54.080 42.300 ;
        RECT 55.380 42.150 59.330 42.300 ;
        RECT 50.130 42.000 50.730 42.150 ;
        RECT 46.530 41.700 50.730 42.000 ;
        RECT 58.730 42.000 59.330 42.150 ;
        RECT 59.780 42.000 59.930 49.550 ;
        RECT 60.380 42.000 60.530 49.550 ;
        RECT 60.980 42.000 61.130 49.550 ;
        RECT 61.580 42.000 61.730 49.550 ;
        RECT 62.180 42.000 62.330 49.550 ;
        RECT 62.780 42.000 62.930 44.900 ;
        RECT 58.730 41.700 62.930 42.000 ;
        RECT 46.530 41.550 54.080 41.700 ;
        RECT 55.380 41.550 62.930 41.700 ;
        RECT 46.530 41.350 50.730 41.550 ;
        RECT 40.330 41.050 49.130 41.200 ;
        RECT 49.280 41.050 50.730 41.350 ;
        RECT 38.730 40.150 50.730 41.050 ;
        RECT 58.730 41.350 62.930 41.550 ;
        RECT 58.730 41.050 60.180 41.350 ;
        RECT 63.530 41.200 65.930 44.400 ;
        RECT 66.530 42.000 66.680 44.900 ;
        RECT 67.130 42.000 67.280 49.550 ;
        RECT 67.730 42.000 67.880 49.550 ;
        RECT 68.330 42.000 68.480 49.550 ;
        RECT 68.930 42.000 69.080 49.550 ;
        RECT 69.530 42.000 69.680 49.550 ;
        RECT 70.130 49.350 74.080 49.550 ;
        RECT 75.380 49.350 79.330 49.550 ;
        RECT 70.130 48.900 70.730 49.350 ;
        RECT 78.730 48.900 79.330 49.350 ;
        RECT 70.130 48.750 74.080 48.900 ;
        RECT 75.380 48.750 79.330 48.900 ;
        RECT 70.130 48.300 70.730 48.750 ;
        RECT 78.730 48.300 79.330 48.750 ;
        RECT 70.130 48.150 74.080 48.300 ;
        RECT 75.380 48.150 79.330 48.300 ;
        RECT 70.130 47.700 70.730 48.150 ;
        RECT 78.730 47.700 79.330 48.150 ;
        RECT 70.130 47.550 74.080 47.700 ;
        RECT 75.380 47.550 79.330 47.700 ;
        RECT 70.130 47.100 70.730 47.550 ;
        RECT 78.730 47.100 79.330 47.550 ;
        RECT 70.130 46.950 74.080 47.100 ;
        RECT 75.380 46.950 79.330 47.100 ;
        RECT 70.130 46.500 70.730 46.950 ;
        RECT 78.730 46.500 79.330 46.950 ;
        RECT 70.130 46.350 74.080 46.500 ;
        RECT 75.380 46.350 79.330 46.500 ;
        RECT 70.130 45.900 70.730 46.350 ;
        RECT 78.730 45.900 79.330 46.350 ;
        RECT 70.130 45.750 74.080 45.900 ;
        RECT 75.380 45.750 79.330 45.900 ;
        RECT 70.130 45.300 70.730 45.750 ;
        RECT 78.730 45.300 79.330 45.750 ;
        RECT 70.130 45.150 74.080 45.300 ;
        RECT 75.380 45.150 79.330 45.300 ;
        RECT 70.130 44.700 70.730 45.150 ;
        RECT 78.730 44.700 79.330 45.150 ;
        RECT 70.130 44.550 74.080 44.700 ;
        RECT 75.380 44.550 79.330 44.700 ;
        RECT 70.130 44.100 70.730 44.550 ;
        RECT 78.730 44.100 79.330 44.550 ;
        RECT 70.130 43.950 74.080 44.100 ;
        RECT 75.380 43.950 79.330 44.100 ;
        RECT 70.130 43.500 70.730 43.950 ;
        RECT 78.730 43.500 79.330 43.950 ;
        RECT 70.130 43.350 74.080 43.500 ;
        RECT 75.380 43.350 79.330 43.500 ;
        RECT 70.130 42.900 70.730 43.350 ;
        RECT 78.730 42.900 79.330 43.350 ;
        RECT 70.130 42.750 74.080 42.900 ;
        RECT 75.380 42.750 79.330 42.900 ;
        RECT 70.130 42.300 70.730 42.750 ;
        RECT 78.730 42.300 79.330 42.750 ;
        RECT 70.130 42.150 74.080 42.300 ;
        RECT 75.380 42.150 79.330 42.300 ;
        RECT 70.130 42.000 70.730 42.150 ;
        RECT 66.530 41.700 70.730 42.000 ;
        RECT 78.730 42.000 79.330 42.150 ;
        RECT 79.780 42.000 79.930 49.550 ;
        RECT 80.380 42.000 80.530 49.550 ;
        RECT 80.980 42.000 81.130 49.550 ;
        RECT 81.580 42.000 81.730 49.550 ;
        RECT 82.180 42.000 82.330 49.550 ;
        RECT 82.780 42.000 82.930 44.900 ;
        RECT 78.730 41.700 82.930 42.000 ;
        RECT 66.530 41.550 74.080 41.700 ;
        RECT 75.380 41.550 82.930 41.700 ;
        RECT 66.530 41.350 70.730 41.550 ;
        RECT 60.330 41.050 69.130 41.200 ;
        RECT 69.280 41.050 70.730 41.350 ;
        RECT 58.730 40.150 70.730 41.050 ;
        RECT 78.730 41.350 82.930 41.550 ;
        RECT 78.730 41.050 80.180 41.350 ;
        RECT 83.530 41.200 85.930 44.400 ;
        RECT 86.530 42.000 86.680 44.900 ;
        RECT 87.130 42.000 87.280 49.550 ;
        RECT 87.730 42.000 87.880 49.550 ;
        RECT 88.330 42.000 88.480 49.550 ;
        RECT 88.930 42.000 89.080 49.550 ;
        RECT 89.530 42.000 89.680 49.550 ;
        RECT 90.130 49.350 94.080 49.550 ;
        RECT 95.380 49.350 99.330 49.550 ;
        RECT 90.130 48.900 90.730 49.350 ;
        RECT 98.730 48.900 99.330 49.350 ;
        RECT 90.130 48.750 94.080 48.900 ;
        RECT 95.380 48.750 99.330 48.900 ;
        RECT 90.130 48.300 90.730 48.750 ;
        RECT 98.730 48.300 99.330 48.750 ;
        RECT 90.130 48.150 94.080 48.300 ;
        RECT 95.380 48.150 99.330 48.300 ;
        RECT 90.130 47.700 90.730 48.150 ;
        RECT 98.730 47.700 99.330 48.150 ;
        RECT 90.130 47.550 94.080 47.700 ;
        RECT 95.380 47.550 99.330 47.700 ;
        RECT 90.130 47.100 90.730 47.550 ;
        RECT 98.730 47.100 99.330 47.550 ;
        RECT 90.130 46.950 94.080 47.100 ;
        RECT 95.380 46.950 99.330 47.100 ;
        RECT 90.130 46.500 90.730 46.950 ;
        RECT 98.730 46.500 99.330 46.950 ;
        RECT 90.130 46.350 94.080 46.500 ;
        RECT 95.380 46.350 99.330 46.500 ;
        RECT 90.130 45.900 90.730 46.350 ;
        RECT 98.730 45.900 99.330 46.350 ;
        RECT 90.130 45.750 94.080 45.900 ;
        RECT 95.380 45.750 99.330 45.900 ;
        RECT 90.130 45.300 90.730 45.750 ;
        RECT 98.730 45.300 99.330 45.750 ;
        RECT 90.130 45.150 94.080 45.300 ;
        RECT 95.380 45.150 99.330 45.300 ;
        RECT 90.130 44.700 90.730 45.150 ;
        RECT 98.730 44.700 99.330 45.150 ;
        RECT 90.130 44.550 94.080 44.700 ;
        RECT 95.380 44.550 99.330 44.700 ;
        RECT 90.130 44.100 90.730 44.550 ;
        RECT 98.730 44.100 99.330 44.550 ;
        RECT 90.130 43.950 94.080 44.100 ;
        RECT 95.380 43.950 99.330 44.100 ;
        RECT 90.130 43.500 90.730 43.950 ;
        RECT 98.730 43.500 99.330 43.950 ;
        RECT 90.130 43.350 94.080 43.500 ;
        RECT 95.380 43.350 99.330 43.500 ;
        RECT 90.130 42.900 90.730 43.350 ;
        RECT 98.730 42.900 99.330 43.350 ;
        RECT 90.130 42.750 94.080 42.900 ;
        RECT 95.380 42.750 99.330 42.900 ;
        RECT 90.130 42.300 90.730 42.750 ;
        RECT 98.730 42.300 99.330 42.750 ;
        RECT 90.130 42.150 94.080 42.300 ;
        RECT 95.380 42.150 99.330 42.300 ;
        RECT 90.130 42.000 90.730 42.150 ;
        RECT 86.530 41.700 90.730 42.000 ;
        RECT 98.730 42.000 99.330 42.150 ;
        RECT 99.780 42.000 99.930 49.550 ;
        RECT 100.380 42.000 100.530 49.550 ;
        RECT 100.980 42.000 101.130 49.550 ;
        RECT 101.580 42.000 101.730 49.550 ;
        RECT 102.180 42.000 102.330 49.550 ;
        RECT 102.780 42.000 102.930 44.900 ;
        RECT 98.730 41.700 102.930 42.000 ;
        RECT 86.530 41.550 94.080 41.700 ;
        RECT 95.380 41.550 102.930 41.700 ;
        RECT 86.530 41.350 90.730 41.550 ;
        RECT 80.330 41.050 89.130 41.200 ;
        RECT 89.280 41.050 90.730 41.350 ;
        RECT 78.730 40.150 90.730 41.050 ;
        RECT 98.730 41.350 102.930 41.550 ;
        RECT 98.730 41.050 100.180 41.350 ;
        RECT 103.530 41.200 105.930 44.400 ;
        RECT 106.530 42.000 106.680 44.900 ;
        RECT 107.130 42.000 107.280 49.550 ;
        RECT 107.730 42.000 107.880 49.550 ;
        RECT 108.330 42.000 108.480 49.550 ;
        RECT 108.930 42.000 109.080 49.550 ;
        RECT 109.530 42.000 109.680 49.550 ;
        RECT 110.130 49.350 114.080 49.550 ;
        RECT 115.380 49.350 119.330 49.550 ;
        RECT 110.130 48.900 110.730 49.350 ;
        RECT 118.730 48.900 119.330 49.350 ;
        RECT 110.130 48.750 114.080 48.900 ;
        RECT 115.380 48.750 119.330 48.900 ;
        RECT 110.130 48.300 110.730 48.750 ;
        RECT 118.730 48.300 119.330 48.750 ;
        RECT 110.130 48.150 114.080 48.300 ;
        RECT 115.380 48.150 119.330 48.300 ;
        RECT 110.130 47.700 110.730 48.150 ;
        RECT 118.730 47.700 119.330 48.150 ;
        RECT 110.130 47.550 114.080 47.700 ;
        RECT 115.380 47.550 119.330 47.700 ;
        RECT 110.130 47.100 110.730 47.550 ;
        RECT 118.730 47.100 119.330 47.550 ;
        RECT 110.130 46.950 114.080 47.100 ;
        RECT 115.380 46.950 119.330 47.100 ;
        RECT 110.130 46.500 110.730 46.950 ;
        RECT 118.730 46.500 119.330 46.950 ;
        RECT 110.130 46.350 114.080 46.500 ;
        RECT 115.380 46.350 119.330 46.500 ;
        RECT 110.130 45.900 110.730 46.350 ;
        RECT 118.730 45.900 119.330 46.350 ;
        RECT 110.130 45.750 114.080 45.900 ;
        RECT 115.380 45.750 119.330 45.900 ;
        RECT 110.130 45.300 110.730 45.750 ;
        RECT 118.730 45.300 119.330 45.750 ;
        RECT 110.130 45.150 114.080 45.300 ;
        RECT 115.380 45.150 119.330 45.300 ;
        RECT 110.130 44.700 110.730 45.150 ;
        RECT 118.730 44.700 119.330 45.150 ;
        RECT 110.130 44.550 114.080 44.700 ;
        RECT 115.380 44.550 119.330 44.700 ;
        RECT 110.130 44.100 110.730 44.550 ;
        RECT 118.730 44.100 119.330 44.550 ;
        RECT 110.130 43.950 114.080 44.100 ;
        RECT 115.380 43.950 119.330 44.100 ;
        RECT 110.130 43.500 110.730 43.950 ;
        RECT 118.730 43.500 119.330 43.950 ;
        RECT 110.130 43.350 114.080 43.500 ;
        RECT 115.380 43.350 119.330 43.500 ;
        RECT 110.130 42.900 110.730 43.350 ;
        RECT 118.730 42.900 119.330 43.350 ;
        RECT 110.130 42.750 114.080 42.900 ;
        RECT 115.380 42.750 119.330 42.900 ;
        RECT 110.130 42.300 110.730 42.750 ;
        RECT 118.730 42.300 119.330 42.750 ;
        RECT 110.130 42.150 114.080 42.300 ;
        RECT 115.380 42.150 119.330 42.300 ;
        RECT 110.130 42.000 110.730 42.150 ;
        RECT 106.530 41.700 110.730 42.000 ;
        RECT 118.730 42.000 119.330 42.150 ;
        RECT 119.780 42.000 119.930 49.550 ;
        RECT 120.380 42.000 120.530 49.550 ;
        RECT 120.980 42.000 121.130 49.550 ;
        RECT 121.580 42.000 121.730 49.550 ;
        RECT 122.180 42.000 122.330 49.550 ;
        RECT 122.780 42.000 122.930 44.900 ;
        RECT 118.730 41.700 122.930 42.000 ;
        RECT 106.530 41.550 114.080 41.700 ;
        RECT 115.380 41.550 122.930 41.700 ;
        RECT 106.530 41.350 110.730 41.550 ;
        RECT 100.330 41.050 109.130 41.200 ;
        RECT 109.280 41.050 110.730 41.350 ;
        RECT 98.730 40.150 110.730 41.050 ;
        RECT 118.730 41.350 122.930 41.550 ;
        RECT 123.530 43.095 124.730 44.400 ;
        RECT 123.530 41.820 127.140 43.095 ;
        RECT 118.730 41.050 120.180 41.350 ;
        RECT 123.530 41.200 124.730 41.820 ;
        RECT 120.330 41.050 124.730 41.200 ;
        RECT 118.730 40.150 124.730 41.050 ;
        RECT 4.730 39.850 9.130 40.150 ;
        RECT 20.330 39.850 29.130 40.150 ;
        RECT 40.330 39.850 49.130 40.150 ;
        RECT 60.330 39.850 69.130 40.150 ;
        RECT 80.330 39.850 89.130 40.150 ;
        RECT 100.330 39.850 109.130 40.150 ;
        RECT 4.730 38.950 10.730 39.850 ;
        RECT 20.330 39.800 30.730 39.850 ;
        RECT 40.330 39.800 50.730 39.850 ;
        RECT 60.330 39.800 70.730 39.850 ;
        RECT 80.330 39.800 90.730 39.850 ;
        RECT 100.330 39.800 110.730 39.850 ;
        RECT 120.330 39.800 124.730 40.150 ;
        RECT 4.730 38.800 9.130 38.950 ;
        RECT 4.730 37.620 5.930 38.800 ;
        RECT 9.280 38.650 10.730 38.950 ;
        RECT 2.315 36.345 5.930 37.620 ;
        RECT 4.730 35.600 5.930 36.345 ;
        RECT 6.530 38.450 10.730 38.650 ;
        RECT 18.730 38.950 30.730 39.800 ;
        RECT 18.730 38.900 29.130 38.950 ;
        RECT 18.730 38.650 20.180 38.900 ;
        RECT 20.330 38.800 29.130 38.900 ;
        RECT 18.730 38.450 22.930 38.650 ;
        RECT 6.530 38.300 14.080 38.450 ;
        RECT 15.430 38.300 22.930 38.450 ;
        RECT 6.530 38.000 10.730 38.300 ;
        RECT 2.315 33.255 4.315 35.550 ;
        RECT 6.530 35.150 6.680 38.000 ;
        RECT 7.130 30.450 7.280 38.000 ;
        RECT 7.730 30.450 7.880 38.000 ;
        RECT 8.330 30.450 8.480 38.000 ;
        RECT 8.930 30.450 9.080 38.000 ;
        RECT 9.530 30.450 9.680 38.000 ;
        RECT 10.130 37.850 10.730 38.000 ;
        RECT 18.730 38.000 22.930 38.300 ;
        RECT 18.730 37.850 19.330 38.000 ;
        RECT 10.130 37.700 14.080 37.850 ;
        RECT 15.380 37.700 19.330 37.850 ;
        RECT 10.130 37.250 10.730 37.700 ;
        RECT 18.730 37.250 19.330 37.700 ;
        RECT 10.130 37.100 14.080 37.250 ;
        RECT 15.380 37.100 19.330 37.250 ;
        RECT 10.130 36.650 10.730 37.100 ;
        RECT 18.730 36.650 19.330 37.100 ;
        RECT 10.130 36.500 14.080 36.650 ;
        RECT 15.380 36.500 19.330 36.650 ;
        RECT 10.130 36.050 10.730 36.500 ;
        RECT 18.730 36.050 19.330 36.500 ;
        RECT 10.130 35.900 14.080 36.050 ;
        RECT 15.380 35.900 19.330 36.050 ;
        RECT 10.130 35.450 10.730 35.900 ;
        RECT 18.730 35.450 19.330 35.900 ;
        RECT 10.130 35.300 14.080 35.450 ;
        RECT 15.380 35.300 19.330 35.450 ;
        RECT 10.130 34.850 10.730 35.300 ;
        RECT 18.730 34.850 19.330 35.300 ;
        RECT 10.130 34.700 14.080 34.850 ;
        RECT 15.380 34.700 19.330 34.850 ;
        RECT 10.130 34.250 10.730 34.700 ;
        RECT 18.730 34.250 19.330 34.700 ;
        RECT 10.130 34.100 14.080 34.250 ;
        RECT 15.380 34.100 19.330 34.250 ;
        RECT 10.130 33.650 10.730 34.100 ;
        RECT 18.730 33.650 19.330 34.100 ;
        RECT 10.130 33.500 14.080 33.650 ;
        RECT 15.380 33.500 19.330 33.650 ;
        RECT 10.130 33.050 10.730 33.500 ;
        RECT 18.730 33.050 19.330 33.500 ;
        RECT 10.130 32.900 14.080 33.050 ;
        RECT 15.380 32.900 19.330 33.050 ;
        RECT 10.130 32.450 10.730 32.900 ;
        RECT 18.730 32.450 19.330 32.900 ;
        RECT 10.130 32.300 14.080 32.450 ;
        RECT 15.380 32.300 19.330 32.450 ;
        RECT 10.130 31.850 10.730 32.300 ;
        RECT 18.730 31.850 19.330 32.300 ;
        RECT 10.130 31.700 14.080 31.850 ;
        RECT 15.380 31.700 19.330 31.850 ;
        RECT 10.130 31.250 10.730 31.700 ;
        RECT 18.730 31.250 19.330 31.700 ;
        RECT 10.130 31.100 14.080 31.250 ;
        RECT 15.380 31.100 19.330 31.250 ;
        RECT 10.130 30.650 10.730 31.100 ;
        RECT 18.730 30.650 19.330 31.100 ;
        RECT 10.130 30.450 14.080 30.650 ;
        RECT 15.380 30.450 19.330 30.650 ;
        RECT 19.780 30.450 19.930 38.000 ;
        RECT 20.380 30.450 20.530 38.000 ;
        RECT 20.980 30.450 21.130 38.000 ;
        RECT 21.580 30.450 21.730 38.000 ;
        RECT 22.180 30.450 22.330 38.000 ;
        RECT 22.780 35.150 22.930 38.000 ;
        RECT 23.530 35.600 25.930 38.800 ;
        RECT 29.280 38.650 30.730 38.950 ;
        RECT 26.530 38.450 30.730 38.650 ;
        RECT 38.730 38.950 50.730 39.800 ;
        RECT 38.730 38.900 49.130 38.950 ;
        RECT 38.730 38.650 40.180 38.900 ;
        RECT 40.330 38.800 49.130 38.900 ;
        RECT 38.730 38.450 42.930 38.650 ;
        RECT 26.530 38.300 34.080 38.450 ;
        RECT 35.430 38.300 42.930 38.450 ;
        RECT 26.530 38.000 30.730 38.300 ;
        RECT 26.530 35.150 26.680 38.000 ;
        RECT 27.130 30.450 27.280 38.000 ;
        RECT 27.730 30.450 27.880 38.000 ;
        RECT 28.330 30.450 28.480 38.000 ;
        RECT 28.930 30.450 29.080 38.000 ;
        RECT 29.530 30.450 29.680 38.000 ;
        RECT 30.130 37.850 30.730 38.000 ;
        RECT 38.730 38.000 42.930 38.300 ;
        RECT 38.730 37.850 39.330 38.000 ;
        RECT 30.130 37.700 34.080 37.850 ;
        RECT 35.380 37.700 39.330 37.850 ;
        RECT 30.130 37.250 30.730 37.700 ;
        RECT 38.730 37.250 39.330 37.700 ;
        RECT 30.130 37.100 34.080 37.250 ;
        RECT 35.380 37.100 39.330 37.250 ;
        RECT 30.130 36.650 30.730 37.100 ;
        RECT 38.730 36.650 39.330 37.100 ;
        RECT 30.130 36.500 34.080 36.650 ;
        RECT 35.380 36.500 39.330 36.650 ;
        RECT 30.130 36.050 30.730 36.500 ;
        RECT 38.730 36.050 39.330 36.500 ;
        RECT 30.130 35.900 34.080 36.050 ;
        RECT 35.380 35.900 39.330 36.050 ;
        RECT 30.130 35.450 30.730 35.900 ;
        RECT 38.730 35.450 39.330 35.900 ;
        RECT 30.130 35.300 34.080 35.450 ;
        RECT 35.380 35.300 39.330 35.450 ;
        RECT 30.130 34.850 30.730 35.300 ;
        RECT 38.730 34.850 39.330 35.300 ;
        RECT 30.130 34.700 34.080 34.850 ;
        RECT 35.380 34.700 39.330 34.850 ;
        RECT 30.130 34.250 30.730 34.700 ;
        RECT 38.730 34.250 39.330 34.700 ;
        RECT 30.130 34.100 34.080 34.250 ;
        RECT 35.380 34.100 39.330 34.250 ;
        RECT 30.130 33.650 30.730 34.100 ;
        RECT 38.730 33.650 39.330 34.100 ;
        RECT 30.130 33.500 34.080 33.650 ;
        RECT 35.380 33.500 39.330 33.650 ;
        RECT 30.130 33.050 30.730 33.500 ;
        RECT 38.730 33.050 39.330 33.500 ;
        RECT 30.130 32.900 34.080 33.050 ;
        RECT 35.380 32.900 39.330 33.050 ;
        RECT 30.130 32.450 30.730 32.900 ;
        RECT 38.730 32.450 39.330 32.900 ;
        RECT 30.130 32.300 34.080 32.450 ;
        RECT 35.380 32.300 39.330 32.450 ;
        RECT 30.130 31.850 30.730 32.300 ;
        RECT 38.730 31.850 39.330 32.300 ;
        RECT 30.130 31.700 34.080 31.850 ;
        RECT 35.380 31.700 39.330 31.850 ;
        RECT 30.130 31.250 30.730 31.700 ;
        RECT 38.730 31.250 39.330 31.700 ;
        RECT 30.130 31.100 34.080 31.250 ;
        RECT 35.380 31.100 39.330 31.250 ;
        RECT 30.130 30.650 30.730 31.100 ;
        RECT 38.730 30.650 39.330 31.100 ;
        RECT 30.130 30.450 34.080 30.650 ;
        RECT 35.380 30.450 39.330 30.650 ;
        RECT 39.780 30.450 39.930 38.000 ;
        RECT 40.380 30.450 40.530 38.000 ;
        RECT 40.980 30.450 41.130 38.000 ;
        RECT 41.580 30.450 41.730 38.000 ;
        RECT 42.180 30.450 42.330 38.000 ;
        RECT 42.780 35.150 42.930 38.000 ;
        RECT 43.530 35.600 45.930 38.800 ;
        RECT 49.280 38.650 50.730 38.950 ;
        RECT 46.530 38.450 50.730 38.650 ;
        RECT 58.730 38.950 70.730 39.800 ;
        RECT 58.730 38.900 69.130 38.950 ;
        RECT 58.730 38.650 60.180 38.900 ;
        RECT 60.330 38.800 69.130 38.900 ;
        RECT 58.730 38.450 62.930 38.650 ;
        RECT 46.530 38.300 54.080 38.450 ;
        RECT 55.430 38.300 62.930 38.450 ;
        RECT 46.530 38.000 50.730 38.300 ;
        RECT 46.530 35.150 46.680 38.000 ;
        RECT 47.130 30.450 47.280 38.000 ;
        RECT 47.730 30.450 47.880 38.000 ;
        RECT 48.330 30.450 48.480 38.000 ;
        RECT 48.930 30.450 49.080 38.000 ;
        RECT 49.530 30.450 49.680 38.000 ;
        RECT 50.130 37.850 50.730 38.000 ;
        RECT 58.730 38.000 62.930 38.300 ;
        RECT 58.730 37.850 59.330 38.000 ;
        RECT 50.130 37.700 54.080 37.850 ;
        RECT 55.380 37.700 59.330 37.850 ;
        RECT 50.130 37.250 50.730 37.700 ;
        RECT 58.730 37.250 59.330 37.700 ;
        RECT 50.130 37.100 54.080 37.250 ;
        RECT 55.380 37.100 59.330 37.250 ;
        RECT 50.130 36.650 50.730 37.100 ;
        RECT 58.730 36.650 59.330 37.100 ;
        RECT 50.130 36.500 54.080 36.650 ;
        RECT 55.380 36.500 59.330 36.650 ;
        RECT 50.130 36.050 50.730 36.500 ;
        RECT 58.730 36.050 59.330 36.500 ;
        RECT 50.130 35.900 54.080 36.050 ;
        RECT 55.380 35.900 59.330 36.050 ;
        RECT 50.130 35.450 50.730 35.900 ;
        RECT 58.730 35.450 59.330 35.900 ;
        RECT 50.130 35.300 54.080 35.450 ;
        RECT 55.380 35.300 59.330 35.450 ;
        RECT 50.130 34.850 50.730 35.300 ;
        RECT 58.730 34.850 59.330 35.300 ;
        RECT 50.130 34.700 54.080 34.850 ;
        RECT 55.380 34.700 59.330 34.850 ;
        RECT 50.130 34.250 50.730 34.700 ;
        RECT 58.730 34.250 59.330 34.700 ;
        RECT 50.130 34.100 54.080 34.250 ;
        RECT 55.380 34.100 59.330 34.250 ;
        RECT 50.130 33.650 50.730 34.100 ;
        RECT 58.730 33.650 59.330 34.100 ;
        RECT 50.130 33.500 54.080 33.650 ;
        RECT 55.380 33.500 59.330 33.650 ;
        RECT 50.130 33.050 50.730 33.500 ;
        RECT 58.730 33.050 59.330 33.500 ;
        RECT 50.130 32.900 54.080 33.050 ;
        RECT 55.380 32.900 59.330 33.050 ;
        RECT 50.130 32.450 50.730 32.900 ;
        RECT 58.730 32.450 59.330 32.900 ;
        RECT 50.130 32.300 54.080 32.450 ;
        RECT 55.380 32.300 59.330 32.450 ;
        RECT 50.130 31.850 50.730 32.300 ;
        RECT 58.730 31.850 59.330 32.300 ;
        RECT 50.130 31.700 54.080 31.850 ;
        RECT 55.380 31.700 59.330 31.850 ;
        RECT 50.130 31.250 50.730 31.700 ;
        RECT 58.730 31.250 59.330 31.700 ;
        RECT 50.130 31.100 54.080 31.250 ;
        RECT 55.380 31.100 59.330 31.250 ;
        RECT 50.130 30.650 50.730 31.100 ;
        RECT 58.730 30.650 59.330 31.100 ;
        RECT 50.130 30.450 54.080 30.650 ;
        RECT 55.380 30.450 59.330 30.650 ;
        RECT 59.780 30.450 59.930 38.000 ;
        RECT 60.380 30.450 60.530 38.000 ;
        RECT 60.980 30.450 61.130 38.000 ;
        RECT 61.580 30.450 61.730 38.000 ;
        RECT 62.180 30.450 62.330 38.000 ;
        RECT 62.780 35.150 62.930 38.000 ;
        RECT 63.530 35.600 65.930 38.800 ;
        RECT 69.280 38.650 70.730 38.950 ;
        RECT 66.530 38.450 70.730 38.650 ;
        RECT 78.730 38.950 90.730 39.800 ;
        RECT 78.730 38.900 89.130 38.950 ;
        RECT 78.730 38.650 80.180 38.900 ;
        RECT 80.330 38.800 89.130 38.900 ;
        RECT 78.730 38.450 82.930 38.650 ;
        RECT 66.530 38.300 74.080 38.450 ;
        RECT 75.430 38.300 82.930 38.450 ;
        RECT 66.530 38.000 70.730 38.300 ;
        RECT 66.530 35.150 66.680 38.000 ;
        RECT 67.130 30.450 67.280 38.000 ;
        RECT 67.730 30.450 67.880 38.000 ;
        RECT 68.330 30.450 68.480 38.000 ;
        RECT 68.930 30.450 69.080 38.000 ;
        RECT 69.530 30.450 69.680 38.000 ;
        RECT 70.130 37.850 70.730 38.000 ;
        RECT 78.730 38.000 82.930 38.300 ;
        RECT 78.730 37.850 79.330 38.000 ;
        RECT 70.130 37.700 74.080 37.850 ;
        RECT 75.380 37.700 79.330 37.850 ;
        RECT 70.130 37.250 70.730 37.700 ;
        RECT 78.730 37.250 79.330 37.700 ;
        RECT 70.130 37.100 74.080 37.250 ;
        RECT 75.380 37.100 79.330 37.250 ;
        RECT 70.130 36.650 70.730 37.100 ;
        RECT 78.730 36.650 79.330 37.100 ;
        RECT 70.130 36.500 74.080 36.650 ;
        RECT 75.380 36.500 79.330 36.650 ;
        RECT 70.130 36.050 70.730 36.500 ;
        RECT 78.730 36.050 79.330 36.500 ;
        RECT 70.130 35.900 74.080 36.050 ;
        RECT 75.380 35.900 79.330 36.050 ;
        RECT 70.130 35.450 70.730 35.900 ;
        RECT 78.730 35.450 79.330 35.900 ;
        RECT 70.130 35.300 74.080 35.450 ;
        RECT 75.380 35.300 79.330 35.450 ;
        RECT 70.130 34.850 70.730 35.300 ;
        RECT 78.730 34.850 79.330 35.300 ;
        RECT 70.130 34.700 74.080 34.850 ;
        RECT 75.380 34.700 79.330 34.850 ;
        RECT 70.130 34.250 70.730 34.700 ;
        RECT 78.730 34.250 79.330 34.700 ;
        RECT 70.130 34.100 74.080 34.250 ;
        RECT 75.380 34.100 79.330 34.250 ;
        RECT 70.130 33.650 70.730 34.100 ;
        RECT 78.730 33.650 79.330 34.100 ;
        RECT 70.130 33.500 74.080 33.650 ;
        RECT 75.380 33.500 79.330 33.650 ;
        RECT 70.130 33.050 70.730 33.500 ;
        RECT 78.730 33.050 79.330 33.500 ;
        RECT 70.130 32.900 74.080 33.050 ;
        RECT 75.380 32.900 79.330 33.050 ;
        RECT 70.130 32.450 70.730 32.900 ;
        RECT 78.730 32.450 79.330 32.900 ;
        RECT 70.130 32.300 74.080 32.450 ;
        RECT 75.380 32.300 79.330 32.450 ;
        RECT 70.130 31.850 70.730 32.300 ;
        RECT 78.730 31.850 79.330 32.300 ;
        RECT 70.130 31.700 74.080 31.850 ;
        RECT 75.380 31.700 79.330 31.850 ;
        RECT 70.130 31.250 70.730 31.700 ;
        RECT 78.730 31.250 79.330 31.700 ;
        RECT 70.130 31.100 74.080 31.250 ;
        RECT 75.380 31.100 79.330 31.250 ;
        RECT 70.130 30.650 70.730 31.100 ;
        RECT 78.730 30.650 79.330 31.100 ;
        RECT 70.130 30.450 74.080 30.650 ;
        RECT 75.380 30.450 79.330 30.650 ;
        RECT 79.780 30.450 79.930 38.000 ;
        RECT 80.380 30.450 80.530 38.000 ;
        RECT 80.980 30.450 81.130 38.000 ;
        RECT 81.580 30.450 81.730 38.000 ;
        RECT 82.180 30.450 82.330 38.000 ;
        RECT 82.780 35.150 82.930 38.000 ;
        RECT 83.530 35.600 85.930 38.800 ;
        RECT 89.280 38.650 90.730 38.950 ;
        RECT 86.530 38.450 90.730 38.650 ;
        RECT 98.730 38.950 110.730 39.800 ;
        RECT 98.730 38.900 109.130 38.950 ;
        RECT 98.730 38.650 100.180 38.900 ;
        RECT 100.330 38.800 109.130 38.900 ;
        RECT 98.730 38.450 102.930 38.650 ;
        RECT 86.530 38.300 94.080 38.450 ;
        RECT 95.430 38.300 102.930 38.450 ;
        RECT 86.530 38.000 90.730 38.300 ;
        RECT 86.530 35.150 86.680 38.000 ;
        RECT 87.130 30.450 87.280 38.000 ;
        RECT 87.730 30.450 87.880 38.000 ;
        RECT 88.330 30.450 88.480 38.000 ;
        RECT 88.930 30.450 89.080 38.000 ;
        RECT 89.530 30.450 89.680 38.000 ;
        RECT 90.130 37.850 90.730 38.000 ;
        RECT 98.730 38.000 102.930 38.300 ;
        RECT 98.730 37.850 99.330 38.000 ;
        RECT 90.130 37.700 94.080 37.850 ;
        RECT 95.380 37.700 99.330 37.850 ;
        RECT 90.130 37.250 90.730 37.700 ;
        RECT 98.730 37.250 99.330 37.700 ;
        RECT 90.130 37.100 94.080 37.250 ;
        RECT 95.380 37.100 99.330 37.250 ;
        RECT 90.130 36.650 90.730 37.100 ;
        RECT 98.730 36.650 99.330 37.100 ;
        RECT 90.130 36.500 94.080 36.650 ;
        RECT 95.380 36.500 99.330 36.650 ;
        RECT 90.130 36.050 90.730 36.500 ;
        RECT 98.730 36.050 99.330 36.500 ;
        RECT 90.130 35.900 94.080 36.050 ;
        RECT 95.380 35.900 99.330 36.050 ;
        RECT 90.130 35.450 90.730 35.900 ;
        RECT 98.730 35.450 99.330 35.900 ;
        RECT 90.130 35.300 94.080 35.450 ;
        RECT 95.380 35.300 99.330 35.450 ;
        RECT 90.130 34.850 90.730 35.300 ;
        RECT 98.730 34.850 99.330 35.300 ;
        RECT 90.130 34.700 94.080 34.850 ;
        RECT 95.380 34.700 99.330 34.850 ;
        RECT 90.130 34.250 90.730 34.700 ;
        RECT 98.730 34.250 99.330 34.700 ;
        RECT 90.130 34.100 94.080 34.250 ;
        RECT 95.380 34.100 99.330 34.250 ;
        RECT 90.130 33.650 90.730 34.100 ;
        RECT 98.730 33.650 99.330 34.100 ;
        RECT 90.130 33.500 94.080 33.650 ;
        RECT 95.380 33.500 99.330 33.650 ;
        RECT 90.130 33.050 90.730 33.500 ;
        RECT 98.730 33.050 99.330 33.500 ;
        RECT 90.130 32.900 94.080 33.050 ;
        RECT 95.380 32.900 99.330 33.050 ;
        RECT 90.130 32.450 90.730 32.900 ;
        RECT 98.730 32.450 99.330 32.900 ;
        RECT 90.130 32.300 94.080 32.450 ;
        RECT 95.380 32.300 99.330 32.450 ;
        RECT 90.130 31.850 90.730 32.300 ;
        RECT 98.730 31.850 99.330 32.300 ;
        RECT 90.130 31.700 94.080 31.850 ;
        RECT 95.380 31.700 99.330 31.850 ;
        RECT 90.130 31.250 90.730 31.700 ;
        RECT 98.730 31.250 99.330 31.700 ;
        RECT 90.130 31.100 94.080 31.250 ;
        RECT 95.380 31.100 99.330 31.250 ;
        RECT 90.130 30.650 90.730 31.100 ;
        RECT 98.730 30.650 99.330 31.100 ;
        RECT 90.130 30.450 94.080 30.650 ;
        RECT 95.380 30.450 99.330 30.650 ;
        RECT 99.780 30.450 99.930 38.000 ;
        RECT 100.380 30.450 100.530 38.000 ;
        RECT 100.980 30.450 101.130 38.000 ;
        RECT 101.580 30.450 101.730 38.000 ;
        RECT 102.180 30.450 102.330 38.000 ;
        RECT 102.780 35.150 102.930 38.000 ;
        RECT 103.530 35.600 105.930 38.800 ;
        RECT 109.280 38.650 110.730 38.950 ;
        RECT 106.530 38.450 110.730 38.650 ;
        RECT 118.730 38.900 124.730 39.800 ;
        RECT 118.730 38.650 120.180 38.900 ;
        RECT 120.330 38.800 124.730 38.900 ;
        RECT 118.730 38.450 122.930 38.650 ;
        RECT 106.530 38.300 114.080 38.450 ;
        RECT 115.430 38.300 122.930 38.450 ;
        RECT 106.530 38.000 110.730 38.300 ;
        RECT 106.530 35.150 106.680 38.000 ;
        RECT 107.130 30.450 107.280 38.000 ;
        RECT 107.730 30.450 107.880 38.000 ;
        RECT 108.330 30.450 108.480 38.000 ;
        RECT 108.930 30.450 109.080 38.000 ;
        RECT 109.530 30.450 109.680 38.000 ;
        RECT 110.130 37.850 110.730 38.000 ;
        RECT 118.730 38.000 122.930 38.300 ;
        RECT 118.730 37.850 119.330 38.000 ;
        RECT 110.130 37.700 114.080 37.850 ;
        RECT 115.380 37.700 119.330 37.850 ;
        RECT 110.130 37.250 110.730 37.700 ;
        RECT 118.730 37.250 119.330 37.700 ;
        RECT 110.130 37.100 114.080 37.250 ;
        RECT 115.380 37.100 119.330 37.250 ;
        RECT 110.130 36.650 110.730 37.100 ;
        RECT 118.730 36.650 119.330 37.100 ;
        RECT 110.130 36.500 114.080 36.650 ;
        RECT 115.380 36.500 119.330 36.650 ;
        RECT 110.130 36.050 110.730 36.500 ;
        RECT 118.730 36.050 119.330 36.500 ;
        RECT 110.130 35.900 114.080 36.050 ;
        RECT 115.380 35.900 119.330 36.050 ;
        RECT 110.130 35.450 110.730 35.900 ;
        RECT 118.730 35.450 119.330 35.900 ;
        RECT 110.130 35.300 114.080 35.450 ;
        RECT 115.380 35.300 119.330 35.450 ;
        RECT 110.130 34.850 110.730 35.300 ;
        RECT 118.730 34.850 119.330 35.300 ;
        RECT 110.130 34.700 114.080 34.850 ;
        RECT 115.380 34.700 119.330 34.850 ;
        RECT 110.130 34.250 110.730 34.700 ;
        RECT 118.730 34.250 119.330 34.700 ;
        RECT 110.130 34.100 114.080 34.250 ;
        RECT 115.380 34.100 119.330 34.250 ;
        RECT 110.130 33.650 110.730 34.100 ;
        RECT 118.730 33.650 119.330 34.100 ;
        RECT 110.130 33.500 114.080 33.650 ;
        RECT 115.380 33.500 119.330 33.650 ;
        RECT 110.130 33.050 110.730 33.500 ;
        RECT 118.730 33.050 119.330 33.500 ;
        RECT 110.130 32.900 114.080 33.050 ;
        RECT 115.380 32.900 119.330 33.050 ;
        RECT 110.130 32.450 110.730 32.900 ;
        RECT 118.730 32.450 119.330 32.900 ;
        RECT 110.130 32.300 114.080 32.450 ;
        RECT 115.380 32.300 119.330 32.450 ;
        RECT 110.130 31.850 110.730 32.300 ;
        RECT 118.730 31.850 119.330 32.300 ;
        RECT 110.130 31.700 114.080 31.850 ;
        RECT 115.380 31.700 119.330 31.850 ;
        RECT 110.130 31.250 110.730 31.700 ;
        RECT 118.730 31.250 119.330 31.700 ;
        RECT 110.130 31.100 114.080 31.250 ;
        RECT 115.380 31.100 119.330 31.250 ;
        RECT 110.130 30.650 110.730 31.100 ;
        RECT 118.730 30.650 119.330 31.100 ;
        RECT 110.130 30.450 114.080 30.650 ;
        RECT 115.380 30.450 119.330 30.650 ;
        RECT 119.780 30.450 119.930 38.000 ;
        RECT 120.380 30.450 120.530 38.000 ;
        RECT 120.980 30.450 121.130 38.000 ;
        RECT 121.580 30.450 121.730 38.000 ;
        RECT 122.180 30.450 122.330 38.000 ;
        RECT 122.780 35.150 122.930 38.000 ;
        RECT 123.530 37.310 124.730 38.800 ;
        RECT 123.530 36.035 127.135 37.310 ;
        RECT 123.530 35.600 124.730 36.035 ;
        RECT 2.315 24.445 4.315 26.740 ;
        RECT 4.730 23.320 5.930 24.400 ;
        RECT 2.315 22.045 5.930 23.320 ;
        RECT 4.730 21.200 5.930 22.045 ;
        RECT 6.530 22.000 6.680 24.900 ;
        RECT 7.130 22.000 7.280 29.550 ;
        RECT 7.730 22.000 7.880 29.550 ;
        RECT 8.330 22.000 8.480 29.550 ;
        RECT 8.930 22.000 9.080 29.550 ;
        RECT 9.530 22.000 9.680 29.550 ;
        RECT 10.130 29.350 14.080 29.550 ;
        RECT 15.380 29.350 19.330 29.550 ;
        RECT 10.130 28.900 10.730 29.350 ;
        RECT 18.730 28.900 19.330 29.350 ;
        RECT 10.130 28.750 14.080 28.900 ;
        RECT 15.380 28.750 19.330 28.900 ;
        RECT 10.130 28.300 10.730 28.750 ;
        RECT 18.730 28.300 19.330 28.750 ;
        RECT 10.130 28.150 14.080 28.300 ;
        RECT 15.380 28.150 19.330 28.300 ;
        RECT 10.130 27.700 10.730 28.150 ;
        RECT 18.730 27.700 19.330 28.150 ;
        RECT 10.130 27.550 14.080 27.700 ;
        RECT 15.380 27.550 19.330 27.700 ;
        RECT 10.130 27.100 10.730 27.550 ;
        RECT 18.730 27.100 19.330 27.550 ;
        RECT 10.130 26.950 14.080 27.100 ;
        RECT 15.380 26.950 19.330 27.100 ;
        RECT 10.130 26.500 10.730 26.950 ;
        RECT 18.730 26.500 19.330 26.950 ;
        RECT 10.130 26.350 14.080 26.500 ;
        RECT 15.380 26.350 19.330 26.500 ;
        RECT 10.130 25.900 10.730 26.350 ;
        RECT 18.730 25.900 19.330 26.350 ;
        RECT 10.130 25.750 14.080 25.900 ;
        RECT 15.380 25.750 19.330 25.900 ;
        RECT 10.130 25.300 10.730 25.750 ;
        RECT 18.730 25.300 19.330 25.750 ;
        RECT 10.130 25.150 14.080 25.300 ;
        RECT 15.380 25.150 19.330 25.300 ;
        RECT 10.130 24.700 10.730 25.150 ;
        RECT 18.730 24.700 19.330 25.150 ;
        RECT 10.130 24.550 14.080 24.700 ;
        RECT 15.380 24.550 19.330 24.700 ;
        RECT 10.130 24.100 10.730 24.550 ;
        RECT 18.730 24.100 19.330 24.550 ;
        RECT 10.130 23.950 14.080 24.100 ;
        RECT 15.380 23.950 19.330 24.100 ;
        RECT 10.130 23.500 10.730 23.950 ;
        RECT 18.730 23.500 19.330 23.950 ;
        RECT 10.130 23.350 14.080 23.500 ;
        RECT 15.380 23.350 19.330 23.500 ;
        RECT 10.130 22.900 10.730 23.350 ;
        RECT 18.730 22.900 19.330 23.350 ;
        RECT 10.130 22.750 14.080 22.900 ;
        RECT 15.380 22.750 19.330 22.900 ;
        RECT 10.130 22.300 10.730 22.750 ;
        RECT 18.730 22.300 19.330 22.750 ;
        RECT 10.130 22.150 14.080 22.300 ;
        RECT 15.380 22.150 19.330 22.300 ;
        RECT 10.130 22.000 10.730 22.150 ;
        RECT 6.530 21.700 10.730 22.000 ;
        RECT 18.730 22.000 19.330 22.150 ;
        RECT 19.780 22.000 19.930 29.550 ;
        RECT 20.380 22.000 20.530 29.550 ;
        RECT 20.980 22.000 21.130 29.550 ;
        RECT 21.580 22.000 21.730 29.550 ;
        RECT 22.180 22.000 22.330 29.550 ;
        RECT 22.780 22.000 22.930 24.900 ;
        RECT 18.730 21.700 22.930 22.000 ;
        RECT 6.530 21.550 14.080 21.700 ;
        RECT 15.380 21.550 22.930 21.700 ;
        RECT 6.530 21.350 10.730 21.550 ;
        RECT 4.730 21.050 9.130 21.200 ;
        RECT 9.280 21.050 10.730 21.350 ;
        RECT 4.730 20.150 10.730 21.050 ;
        RECT 18.730 21.350 22.930 21.550 ;
        RECT 18.730 21.050 20.180 21.350 ;
        RECT 23.530 21.200 25.930 24.400 ;
        RECT 26.530 22.000 26.680 24.900 ;
        RECT 27.130 22.000 27.280 29.550 ;
        RECT 27.730 22.000 27.880 29.550 ;
        RECT 28.330 22.000 28.480 29.550 ;
        RECT 28.930 22.000 29.080 29.550 ;
        RECT 29.530 22.000 29.680 29.550 ;
        RECT 30.130 29.350 34.080 29.550 ;
        RECT 35.380 29.350 39.330 29.550 ;
        RECT 30.130 28.900 30.730 29.350 ;
        RECT 38.730 28.900 39.330 29.350 ;
        RECT 30.130 28.750 34.080 28.900 ;
        RECT 35.380 28.750 39.330 28.900 ;
        RECT 30.130 28.300 30.730 28.750 ;
        RECT 38.730 28.300 39.330 28.750 ;
        RECT 30.130 28.150 34.080 28.300 ;
        RECT 35.380 28.150 39.330 28.300 ;
        RECT 30.130 27.700 30.730 28.150 ;
        RECT 38.730 27.700 39.330 28.150 ;
        RECT 30.130 27.550 34.080 27.700 ;
        RECT 35.380 27.550 39.330 27.700 ;
        RECT 30.130 27.100 30.730 27.550 ;
        RECT 38.730 27.100 39.330 27.550 ;
        RECT 30.130 26.950 34.080 27.100 ;
        RECT 35.380 26.950 39.330 27.100 ;
        RECT 30.130 26.500 30.730 26.950 ;
        RECT 38.730 26.500 39.330 26.950 ;
        RECT 30.130 26.350 34.080 26.500 ;
        RECT 35.380 26.350 39.330 26.500 ;
        RECT 30.130 25.900 30.730 26.350 ;
        RECT 38.730 25.900 39.330 26.350 ;
        RECT 30.130 25.750 34.080 25.900 ;
        RECT 35.380 25.750 39.330 25.900 ;
        RECT 30.130 25.300 30.730 25.750 ;
        RECT 38.730 25.300 39.330 25.750 ;
        RECT 30.130 25.150 34.080 25.300 ;
        RECT 35.380 25.150 39.330 25.300 ;
        RECT 30.130 24.700 30.730 25.150 ;
        RECT 38.730 24.700 39.330 25.150 ;
        RECT 30.130 24.550 34.080 24.700 ;
        RECT 35.380 24.550 39.330 24.700 ;
        RECT 30.130 24.100 30.730 24.550 ;
        RECT 38.730 24.100 39.330 24.550 ;
        RECT 30.130 23.950 34.080 24.100 ;
        RECT 35.380 23.950 39.330 24.100 ;
        RECT 30.130 23.500 30.730 23.950 ;
        RECT 38.730 23.500 39.330 23.950 ;
        RECT 30.130 23.350 34.080 23.500 ;
        RECT 35.380 23.350 39.330 23.500 ;
        RECT 30.130 22.900 30.730 23.350 ;
        RECT 38.730 22.900 39.330 23.350 ;
        RECT 30.130 22.750 34.080 22.900 ;
        RECT 35.380 22.750 39.330 22.900 ;
        RECT 30.130 22.300 30.730 22.750 ;
        RECT 38.730 22.300 39.330 22.750 ;
        RECT 30.130 22.150 34.080 22.300 ;
        RECT 35.380 22.150 39.330 22.300 ;
        RECT 30.130 22.000 30.730 22.150 ;
        RECT 26.530 21.700 30.730 22.000 ;
        RECT 38.730 22.000 39.330 22.150 ;
        RECT 39.780 22.000 39.930 29.550 ;
        RECT 40.380 22.000 40.530 29.550 ;
        RECT 40.980 22.000 41.130 29.550 ;
        RECT 41.580 22.000 41.730 29.550 ;
        RECT 42.180 22.000 42.330 29.550 ;
        RECT 42.780 22.000 42.930 24.900 ;
        RECT 38.730 21.700 42.930 22.000 ;
        RECT 26.530 21.550 34.080 21.700 ;
        RECT 35.380 21.550 42.930 21.700 ;
        RECT 26.530 21.350 30.730 21.550 ;
        RECT 20.330 21.050 29.130 21.200 ;
        RECT 29.280 21.050 30.730 21.350 ;
        RECT 18.730 20.150 30.730 21.050 ;
        RECT 38.730 21.350 42.930 21.550 ;
        RECT 38.730 21.050 40.180 21.350 ;
        RECT 43.530 21.200 45.930 24.400 ;
        RECT 46.530 22.000 46.680 24.900 ;
        RECT 47.130 22.000 47.280 29.550 ;
        RECT 47.730 22.000 47.880 29.550 ;
        RECT 48.330 22.000 48.480 29.550 ;
        RECT 48.930 22.000 49.080 29.550 ;
        RECT 49.530 22.000 49.680 29.550 ;
        RECT 50.130 29.350 54.080 29.550 ;
        RECT 55.380 29.350 59.330 29.550 ;
        RECT 50.130 28.900 50.730 29.350 ;
        RECT 58.730 28.900 59.330 29.350 ;
        RECT 50.130 28.750 54.080 28.900 ;
        RECT 55.380 28.750 59.330 28.900 ;
        RECT 50.130 28.300 50.730 28.750 ;
        RECT 58.730 28.300 59.330 28.750 ;
        RECT 50.130 28.150 54.080 28.300 ;
        RECT 55.380 28.150 59.330 28.300 ;
        RECT 50.130 27.700 50.730 28.150 ;
        RECT 58.730 27.700 59.330 28.150 ;
        RECT 50.130 27.550 54.080 27.700 ;
        RECT 55.380 27.550 59.330 27.700 ;
        RECT 50.130 27.100 50.730 27.550 ;
        RECT 58.730 27.100 59.330 27.550 ;
        RECT 50.130 26.950 54.080 27.100 ;
        RECT 55.380 26.950 59.330 27.100 ;
        RECT 50.130 26.500 50.730 26.950 ;
        RECT 58.730 26.500 59.330 26.950 ;
        RECT 50.130 26.350 54.080 26.500 ;
        RECT 55.380 26.350 59.330 26.500 ;
        RECT 50.130 25.900 50.730 26.350 ;
        RECT 58.730 25.900 59.330 26.350 ;
        RECT 50.130 25.750 54.080 25.900 ;
        RECT 55.380 25.750 59.330 25.900 ;
        RECT 50.130 25.300 50.730 25.750 ;
        RECT 58.730 25.300 59.330 25.750 ;
        RECT 50.130 25.150 54.080 25.300 ;
        RECT 55.380 25.150 59.330 25.300 ;
        RECT 50.130 24.700 50.730 25.150 ;
        RECT 58.730 24.700 59.330 25.150 ;
        RECT 50.130 24.550 54.080 24.700 ;
        RECT 55.380 24.550 59.330 24.700 ;
        RECT 50.130 24.100 50.730 24.550 ;
        RECT 58.730 24.100 59.330 24.550 ;
        RECT 50.130 23.950 54.080 24.100 ;
        RECT 55.380 23.950 59.330 24.100 ;
        RECT 50.130 23.500 50.730 23.950 ;
        RECT 58.730 23.500 59.330 23.950 ;
        RECT 50.130 23.350 54.080 23.500 ;
        RECT 55.380 23.350 59.330 23.500 ;
        RECT 50.130 22.900 50.730 23.350 ;
        RECT 58.730 22.900 59.330 23.350 ;
        RECT 50.130 22.750 54.080 22.900 ;
        RECT 55.380 22.750 59.330 22.900 ;
        RECT 50.130 22.300 50.730 22.750 ;
        RECT 58.730 22.300 59.330 22.750 ;
        RECT 50.130 22.150 54.080 22.300 ;
        RECT 55.380 22.150 59.330 22.300 ;
        RECT 50.130 22.000 50.730 22.150 ;
        RECT 46.530 21.700 50.730 22.000 ;
        RECT 58.730 22.000 59.330 22.150 ;
        RECT 59.780 22.000 59.930 29.550 ;
        RECT 60.380 22.000 60.530 29.550 ;
        RECT 60.980 22.000 61.130 29.550 ;
        RECT 61.580 22.000 61.730 29.550 ;
        RECT 62.180 22.000 62.330 29.550 ;
        RECT 62.780 22.000 62.930 24.900 ;
        RECT 58.730 21.700 62.930 22.000 ;
        RECT 46.530 21.550 54.080 21.700 ;
        RECT 55.380 21.550 62.930 21.700 ;
        RECT 46.530 21.350 50.730 21.550 ;
        RECT 40.330 21.050 49.130 21.200 ;
        RECT 49.280 21.050 50.730 21.350 ;
        RECT 38.730 20.150 50.730 21.050 ;
        RECT 58.730 21.350 62.930 21.550 ;
        RECT 58.730 21.050 60.180 21.350 ;
        RECT 63.530 21.200 65.930 24.400 ;
        RECT 66.530 22.000 66.680 24.900 ;
        RECT 67.130 22.000 67.280 29.550 ;
        RECT 67.730 22.000 67.880 29.550 ;
        RECT 68.330 22.000 68.480 29.550 ;
        RECT 68.930 22.000 69.080 29.550 ;
        RECT 69.530 22.000 69.680 29.550 ;
        RECT 70.130 29.350 74.080 29.550 ;
        RECT 75.380 29.350 79.330 29.550 ;
        RECT 70.130 28.900 70.730 29.350 ;
        RECT 78.730 28.900 79.330 29.350 ;
        RECT 70.130 28.750 74.080 28.900 ;
        RECT 75.380 28.750 79.330 28.900 ;
        RECT 70.130 28.300 70.730 28.750 ;
        RECT 78.730 28.300 79.330 28.750 ;
        RECT 70.130 28.150 74.080 28.300 ;
        RECT 75.380 28.150 79.330 28.300 ;
        RECT 70.130 27.700 70.730 28.150 ;
        RECT 78.730 27.700 79.330 28.150 ;
        RECT 70.130 27.550 74.080 27.700 ;
        RECT 75.380 27.550 79.330 27.700 ;
        RECT 70.130 27.100 70.730 27.550 ;
        RECT 78.730 27.100 79.330 27.550 ;
        RECT 70.130 26.950 74.080 27.100 ;
        RECT 75.380 26.950 79.330 27.100 ;
        RECT 70.130 26.500 70.730 26.950 ;
        RECT 78.730 26.500 79.330 26.950 ;
        RECT 70.130 26.350 74.080 26.500 ;
        RECT 75.380 26.350 79.330 26.500 ;
        RECT 70.130 25.900 70.730 26.350 ;
        RECT 78.730 25.900 79.330 26.350 ;
        RECT 70.130 25.750 74.080 25.900 ;
        RECT 75.380 25.750 79.330 25.900 ;
        RECT 70.130 25.300 70.730 25.750 ;
        RECT 78.730 25.300 79.330 25.750 ;
        RECT 70.130 25.150 74.080 25.300 ;
        RECT 75.380 25.150 79.330 25.300 ;
        RECT 70.130 24.700 70.730 25.150 ;
        RECT 78.730 24.700 79.330 25.150 ;
        RECT 70.130 24.550 74.080 24.700 ;
        RECT 75.380 24.550 79.330 24.700 ;
        RECT 70.130 24.100 70.730 24.550 ;
        RECT 78.730 24.100 79.330 24.550 ;
        RECT 70.130 23.950 74.080 24.100 ;
        RECT 75.380 23.950 79.330 24.100 ;
        RECT 70.130 23.500 70.730 23.950 ;
        RECT 78.730 23.500 79.330 23.950 ;
        RECT 70.130 23.350 74.080 23.500 ;
        RECT 75.380 23.350 79.330 23.500 ;
        RECT 70.130 22.900 70.730 23.350 ;
        RECT 78.730 22.900 79.330 23.350 ;
        RECT 70.130 22.750 74.080 22.900 ;
        RECT 75.380 22.750 79.330 22.900 ;
        RECT 70.130 22.300 70.730 22.750 ;
        RECT 78.730 22.300 79.330 22.750 ;
        RECT 70.130 22.150 74.080 22.300 ;
        RECT 75.380 22.150 79.330 22.300 ;
        RECT 70.130 22.000 70.730 22.150 ;
        RECT 66.530 21.700 70.730 22.000 ;
        RECT 78.730 22.000 79.330 22.150 ;
        RECT 79.780 22.000 79.930 29.550 ;
        RECT 80.380 22.000 80.530 29.550 ;
        RECT 80.980 22.000 81.130 29.550 ;
        RECT 81.580 22.000 81.730 29.550 ;
        RECT 82.180 22.000 82.330 29.550 ;
        RECT 82.780 22.000 82.930 24.900 ;
        RECT 78.730 21.700 82.930 22.000 ;
        RECT 66.530 21.550 74.080 21.700 ;
        RECT 75.380 21.550 82.930 21.700 ;
        RECT 66.530 21.350 70.730 21.550 ;
        RECT 60.330 21.050 69.130 21.200 ;
        RECT 69.280 21.050 70.730 21.350 ;
        RECT 58.730 20.150 70.730 21.050 ;
        RECT 78.730 21.350 82.930 21.550 ;
        RECT 78.730 21.050 80.180 21.350 ;
        RECT 83.530 21.200 85.930 24.400 ;
        RECT 86.530 22.000 86.680 24.900 ;
        RECT 87.130 22.000 87.280 29.550 ;
        RECT 87.730 22.000 87.880 29.550 ;
        RECT 88.330 22.000 88.480 29.550 ;
        RECT 88.930 22.000 89.080 29.550 ;
        RECT 89.530 22.000 89.680 29.550 ;
        RECT 90.130 29.350 94.080 29.550 ;
        RECT 95.380 29.350 99.330 29.550 ;
        RECT 90.130 28.900 90.730 29.350 ;
        RECT 98.730 28.900 99.330 29.350 ;
        RECT 90.130 28.750 94.080 28.900 ;
        RECT 95.380 28.750 99.330 28.900 ;
        RECT 90.130 28.300 90.730 28.750 ;
        RECT 98.730 28.300 99.330 28.750 ;
        RECT 90.130 28.150 94.080 28.300 ;
        RECT 95.380 28.150 99.330 28.300 ;
        RECT 90.130 27.700 90.730 28.150 ;
        RECT 98.730 27.700 99.330 28.150 ;
        RECT 90.130 27.550 94.080 27.700 ;
        RECT 95.380 27.550 99.330 27.700 ;
        RECT 90.130 27.100 90.730 27.550 ;
        RECT 98.730 27.100 99.330 27.550 ;
        RECT 90.130 26.950 94.080 27.100 ;
        RECT 95.380 26.950 99.330 27.100 ;
        RECT 90.130 26.500 90.730 26.950 ;
        RECT 98.730 26.500 99.330 26.950 ;
        RECT 90.130 26.350 94.080 26.500 ;
        RECT 95.380 26.350 99.330 26.500 ;
        RECT 90.130 25.900 90.730 26.350 ;
        RECT 98.730 25.900 99.330 26.350 ;
        RECT 90.130 25.750 94.080 25.900 ;
        RECT 95.380 25.750 99.330 25.900 ;
        RECT 90.130 25.300 90.730 25.750 ;
        RECT 98.730 25.300 99.330 25.750 ;
        RECT 90.130 25.150 94.080 25.300 ;
        RECT 95.380 25.150 99.330 25.300 ;
        RECT 90.130 24.700 90.730 25.150 ;
        RECT 98.730 24.700 99.330 25.150 ;
        RECT 90.130 24.550 94.080 24.700 ;
        RECT 95.380 24.550 99.330 24.700 ;
        RECT 90.130 24.100 90.730 24.550 ;
        RECT 98.730 24.100 99.330 24.550 ;
        RECT 90.130 23.950 94.080 24.100 ;
        RECT 95.380 23.950 99.330 24.100 ;
        RECT 90.130 23.500 90.730 23.950 ;
        RECT 98.730 23.500 99.330 23.950 ;
        RECT 90.130 23.350 94.080 23.500 ;
        RECT 95.380 23.350 99.330 23.500 ;
        RECT 90.130 22.900 90.730 23.350 ;
        RECT 98.730 22.900 99.330 23.350 ;
        RECT 90.130 22.750 94.080 22.900 ;
        RECT 95.380 22.750 99.330 22.900 ;
        RECT 90.130 22.300 90.730 22.750 ;
        RECT 98.730 22.300 99.330 22.750 ;
        RECT 90.130 22.150 94.080 22.300 ;
        RECT 95.380 22.150 99.330 22.300 ;
        RECT 90.130 22.000 90.730 22.150 ;
        RECT 86.530 21.700 90.730 22.000 ;
        RECT 98.730 22.000 99.330 22.150 ;
        RECT 99.780 22.000 99.930 29.550 ;
        RECT 100.380 22.000 100.530 29.550 ;
        RECT 100.980 22.000 101.130 29.550 ;
        RECT 101.580 22.000 101.730 29.550 ;
        RECT 102.180 22.000 102.330 29.550 ;
        RECT 102.780 22.000 102.930 24.900 ;
        RECT 98.730 21.700 102.930 22.000 ;
        RECT 86.530 21.550 94.080 21.700 ;
        RECT 95.380 21.550 102.930 21.700 ;
        RECT 86.530 21.350 90.730 21.550 ;
        RECT 80.330 21.050 89.130 21.200 ;
        RECT 89.280 21.050 90.730 21.350 ;
        RECT 78.730 20.150 90.730 21.050 ;
        RECT 98.730 21.350 102.930 21.550 ;
        RECT 98.730 21.050 100.180 21.350 ;
        RECT 103.530 21.200 105.930 24.400 ;
        RECT 106.530 22.000 106.680 24.900 ;
        RECT 107.130 22.000 107.280 29.550 ;
        RECT 107.730 22.000 107.880 29.550 ;
        RECT 108.330 22.000 108.480 29.550 ;
        RECT 108.930 22.000 109.080 29.550 ;
        RECT 109.530 22.000 109.680 29.550 ;
        RECT 110.130 29.350 114.080 29.550 ;
        RECT 115.380 29.350 119.330 29.550 ;
        RECT 110.130 28.900 110.730 29.350 ;
        RECT 118.730 28.900 119.330 29.350 ;
        RECT 110.130 28.750 114.080 28.900 ;
        RECT 115.380 28.750 119.330 28.900 ;
        RECT 110.130 28.300 110.730 28.750 ;
        RECT 118.730 28.300 119.330 28.750 ;
        RECT 110.130 28.150 114.080 28.300 ;
        RECT 115.380 28.150 119.330 28.300 ;
        RECT 110.130 27.700 110.730 28.150 ;
        RECT 118.730 27.700 119.330 28.150 ;
        RECT 110.130 27.550 114.080 27.700 ;
        RECT 115.380 27.550 119.330 27.700 ;
        RECT 110.130 27.100 110.730 27.550 ;
        RECT 118.730 27.100 119.330 27.550 ;
        RECT 110.130 26.950 114.080 27.100 ;
        RECT 115.380 26.950 119.330 27.100 ;
        RECT 110.130 26.500 110.730 26.950 ;
        RECT 118.730 26.500 119.330 26.950 ;
        RECT 110.130 26.350 114.080 26.500 ;
        RECT 115.380 26.350 119.330 26.500 ;
        RECT 110.130 25.900 110.730 26.350 ;
        RECT 118.730 25.900 119.330 26.350 ;
        RECT 110.130 25.750 114.080 25.900 ;
        RECT 115.380 25.750 119.330 25.900 ;
        RECT 110.130 25.300 110.730 25.750 ;
        RECT 118.730 25.300 119.330 25.750 ;
        RECT 110.130 25.150 114.080 25.300 ;
        RECT 115.380 25.150 119.330 25.300 ;
        RECT 110.130 24.700 110.730 25.150 ;
        RECT 118.730 24.700 119.330 25.150 ;
        RECT 110.130 24.550 114.080 24.700 ;
        RECT 115.380 24.550 119.330 24.700 ;
        RECT 110.130 24.100 110.730 24.550 ;
        RECT 118.730 24.100 119.330 24.550 ;
        RECT 110.130 23.950 114.080 24.100 ;
        RECT 115.380 23.950 119.330 24.100 ;
        RECT 110.130 23.500 110.730 23.950 ;
        RECT 118.730 23.500 119.330 23.950 ;
        RECT 110.130 23.350 114.080 23.500 ;
        RECT 115.380 23.350 119.330 23.500 ;
        RECT 110.130 22.900 110.730 23.350 ;
        RECT 118.730 22.900 119.330 23.350 ;
        RECT 110.130 22.750 114.080 22.900 ;
        RECT 115.380 22.750 119.330 22.900 ;
        RECT 110.130 22.300 110.730 22.750 ;
        RECT 118.730 22.300 119.330 22.750 ;
        RECT 110.130 22.150 114.080 22.300 ;
        RECT 115.380 22.150 119.330 22.300 ;
        RECT 110.130 22.000 110.730 22.150 ;
        RECT 106.530 21.700 110.730 22.000 ;
        RECT 118.730 22.000 119.330 22.150 ;
        RECT 119.780 22.000 119.930 29.550 ;
        RECT 120.380 22.000 120.530 29.550 ;
        RECT 120.980 22.000 121.130 29.550 ;
        RECT 121.580 22.000 121.730 29.550 ;
        RECT 122.180 22.000 122.330 29.550 ;
        RECT 122.780 22.000 122.930 24.900 ;
        RECT 118.730 21.700 122.930 22.000 ;
        RECT 106.530 21.550 114.080 21.700 ;
        RECT 115.380 21.550 122.930 21.700 ;
        RECT 106.530 21.350 110.730 21.550 ;
        RECT 100.330 21.050 109.130 21.200 ;
        RECT 109.280 21.050 110.730 21.350 ;
        RECT 98.730 20.150 110.730 21.050 ;
        RECT 118.730 21.350 122.930 21.550 ;
        RECT 123.530 23.095 124.730 24.400 ;
        RECT 123.530 21.820 127.140 23.095 ;
        RECT 118.730 21.050 120.180 21.350 ;
        RECT 123.530 21.200 124.730 21.820 ;
        RECT 120.330 21.050 124.730 21.200 ;
        RECT 118.730 20.150 124.730 21.050 ;
        RECT 4.730 19.850 9.130 20.150 ;
        RECT 20.330 19.850 29.130 20.150 ;
        RECT 40.330 19.850 49.130 20.150 ;
        RECT 60.330 19.850 69.130 20.150 ;
        RECT 80.330 19.850 89.130 20.150 ;
        RECT 100.330 19.850 109.130 20.150 ;
        RECT 4.730 18.950 10.730 19.850 ;
        RECT 20.330 19.800 30.730 19.850 ;
        RECT 40.330 19.800 50.730 19.850 ;
        RECT 60.330 19.800 70.730 19.850 ;
        RECT 80.330 19.800 90.730 19.850 ;
        RECT 100.330 19.800 110.730 19.850 ;
        RECT 120.330 19.800 124.730 20.150 ;
        RECT 4.730 18.800 9.130 18.950 ;
        RECT 4.730 17.765 5.930 18.800 ;
        RECT 9.280 18.650 10.730 18.950 ;
        RECT 2.315 16.490 5.930 17.765 ;
        RECT 4.730 15.600 5.930 16.490 ;
        RECT 6.530 18.450 10.730 18.650 ;
        RECT 18.730 18.950 30.730 19.800 ;
        RECT 18.730 18.900 29.130 18.950 ;
        RECT 18.730 18.650 20.180 18.900 ;
        RECT 20.330 18.800 29.130 18.900 ;
        RECT 18.730 18.450 22.930 18.650 ;
        RECT 6.530 18.300 14.080 18.450 ;
        RECT 15.430 18.300 22.930 18.450 ;
        RECT 6.530 18.000 10.730 18.300 ;
        RECT 2.315 13.255 4.315 15.550 ;
        RECT 6.530 15.150 6.680 18.000 ;
        RECT 7.130 10.450 7.280 18.000 ;
        RECT 7.730 10.450 7.880 18.000 ;
        RECT 8.330 10.450 8.480 18.000 ;
        RECT 8.930 10.450 9.080 18.000 ;
        RECT 9.530 10.450 9.680 18.000 ;
        RECT 10.130 17.850 10.730 18.000 ;
        RECT 18.730 18.000 22.930 18.300 ;
        RECT 18.730 17.850 19.330 18.000 ;
        RECT 10.130 17.700 14.080 17.850 ;
        RECT 15.380 17.700 19.330 17.850 ;
        RECT 10.130 17.250 10.730 17.700 ;
        RECT 18.730 17.250 19.330 17.700 ;
        RECT 10.130 17.100 14.080 17.250 ;
        RECT 15.380 17.100 19.330 17.250 ;
        RECT 10.130 16.650 10.730 17.100 ;
        RECT 18.730 16.650 19.330 17.100 ;
        RECT 10.130 16.500 14.080 16.650 ;
        RECT 15.380 16.500 19.330 16.650 ;
        RECT 10.130 16.050 10.730 16.500 ;
        RECT 18.730 16.050 19.330 16.500 ;
        RECT 10.130 15.900 14.080 16.050 ;
        RECT 15.380 15.900 19.330 16.050 ;
        RECT 10.130 15.450 10.730 15.900 ;
        RECT 18.730 15.450 19.330 15.900 ;
        RECT 10.130 15.300 14.080 15.450 ;
        RECT 15.380 15.300 19.330 15.450 ;
        RECT 10.130 14.850 10.730 15.300 ;
        RECT 18.730 14.850 19.330 15.300 ;
        RECT 10.130 14.700 14.080 14.850 ;
        RECT 15.380 14.700 19.330 14.850 ;
        RECT 10.130 14.250 10.730 14.700 ;
        RECT 18.730 14.250 19.330 14.700 ;
        RECT 10.130 14.100 14.080 14.250 ;
        RECT 15.380 14.100 19.330 14.250 ;
        RECT 10.130 13.650 10.730 14.100 ;
        RECT 18.730 13.650 19.330 14.100 ;
        RECT 10.130 13.500 14.080 13.650 ;
        RECT 15.380 13.500 19.330 13.650 ;
        RECT 10.130 13.050 10.730 13.500 ;
        RECT 18.730 13.050 19.330 13.500 ;
        RECT 10.130 12.900 14.080 13.050 ;
        RECT 15.380 12.900 19.330 13.050 ;
        RECT 10.130 12.450 10.730 12.900 ;
        RECT 18.730 12.450 19.330 12.900 ;
        RECT 10.130 12.300 14.080 12.450 ;
        RECT 15.380 12.300 19.330 12.450 ;
        RECT 10.130 11.850 10.730 12.300 ;
        RECT 18.730 11.850 19.330 12.300 ;
        RECT 10.130 11.700 14.080 11.850 ;
        RECT 15.380 11.700 19.330 11.850 ;
        RECT 10.130 11.250 10.730 11.700 ;
        RECT 18.730 11.250 19.330 11.700 ;
        RECT 10.130 11.100 14.080 11.250 ;
        RECT 15.380 11.100 19.330 11.250 ;
        RECT 10.130 10.650 10.730 11.100 ;
        RECT 18.730 10.650 19.330 11.100 ;
        RECT 10.130 10.450 14.080 10.650 ;
        RECT 15.380 10.450 19.330 10.650 ;
        RECT 19.780 10.450 19.930 18.000 ;
        RECT 20.380 10.450 20.530 18.000 ;
        RECT 20.980 10.450 21.130 18.000 ;
        RECT 21.580 10.450 21.730 18.000 ;
        RECT 22.180 10.450 22.330 18.000 ;
        RECT 22.780 15.150 22.930 18.000 ;
        RECT 23.530 15.600 25.930 18.800 ;
        RECT 29.280 18.650 30.730 18.950 ;
        RECT 26.530 18.450 30.730 18.650 ;
        RECT 38.730 18.950 50.730 19.800 ;
        RECT 38.730 18.900 49.130 18.950 ;
        RECT 38.730 18.650 40.180 18.900 ;
        RECT 40.330 18.800 49.130 18.900 ;
        RECT 38.730 18.450 42.930 18.650 ;
        RECT 26.530 18.300 34.080 18.450 ;
        RECT 35.430 18.300 42.930 18.450 ;
        RECT 26.530 18.000 30.730 18.300 ;
        RECT 26.530 15.150 26.680 18.000 ;
        RECT 27.130 10.450 27.280 18.000 ;
        RECT 27.730 10.450 27.880 18.000 ;
        RECT 28.330 10.450 28.480 18.000 ;
        RECT 28.930 10.450 29.080 18.000 ;
        RECT 29.530 10.450 29.680 18.000 ;
        RECT 30.130 17.850 30.730 18.000 ;
        RECT 38.730 18.000 42.930 18.300 ;
        RECT 38.730 17.850 39.330 18.000 ;
        RECT 30.130 17.700 34.080 17.850 ;
        RECT 35.380 17.700 39.330 17.850 ;
        RECT 30.130 17.250 30.730 17.700 ;
        RECT 38.730 17.250 39.330 17.700 ;
        RECT 30.130 17.100 34.080 17.250 ;
        RECT 35.380 17.100 39.330 17.250 ;
        RECT 30.130 16.650 30.730 17.100 ;
        RECT 38.730 16.650 39.330 17.100 ;
        RECT 30.130 16.500 34.080 16.650 ;
        RECT 35.380 16.500 39.330 16.650 ;
        RECT 30.130 16.050 30.730 16.500 ;
        RECT 38.730 16.050 39.330 16.500 ;
        RECT 30.130 15.900 34.080 16.050 ;
        RECT 35.380 15.900 39.330 16.050 ;
        RECT 30.130 15.450 30.730 15.900 ;
        RECT 38.730 15.450 39.330 15.900 ;
        RECT 30.130 15.300 34.080 15.450 ;
        RECT 35.380 15.300 39.330 15.450 ;
        RECT 30.130 14.850 30.730 15.300 ;
        RECT 38.730 14.850 39.330 15.300 ;
        RECT 30.130 14.700 34.080 14.850 ;
        RECT 35.380 14.700 39.330 14.850 ;
        RECT 30.130 14.250 30.730 14.700 ;
        RECT 38.730 14.250 39.330 14.700 ;
        RECT 30.130 14.100 34.080 14.250 ;
        RECT 35.380 14.100 39.330 14.250 ;
        RECT 30.130 13.650 30.730 14.100 ;
        RECT 38.730 13.650 39.330 14.100 ;
        RECT 30.130 13.500 34.080 13.650 ;
        RECT 35.380 13.500 39.330 13.650 ;
        RECT 30.130 13.050 30.730 13.500 ;
        RECT 38.730 13.050 39.330 13.500 ;
        RECT 30.130 12.900 34.080 13.050 ;
        RECT 35.380 12.900 39.330 13.050 ;
        RECT 30.130 12.450 30.730 12.900 ;
        RECT 38.730 12.450 39.330 12.900 ;
        RECT 30.130 12.300 34.080 12.450 ;
        RECT 35.380 12.300 39.330 12.450 ;
        RECT 30.130 11.850 30.730 12.300 ;
        RECT 38.730 11.850 39.330 12.300 ;
        RECT 30.130 11.700 34.080 11.850 ;
        RECT 35.380 11.700 39.330 11.850 ;
        RECT 30.130 11.250 30.730 11.700 ;
        RECT 38.730 11.250 39.330 11.700 ;
        RECT 30.130 11.100 34.080 11.250 ;
        RECT 35.380 11.100 39.330 11.250 ;
        RECT 30.130 10.650 30.730 11.100 ;
        RECT 38.730 10.650 39.330 11.100 ;
        RECT 30.130 10.450 34.080 10.650 ;
        RECT 35.380 10.450 39.330 10.650 ;
        RECT 39.780 10.450 39.930 18.000 ;
        RECT 40.380 10.450 40.530 18.000 ;
        RECT 40.980 10.450 41.130 18.000 ;
        RECT 41.580 10.450 41.730 18.000 ;
        RECT 42.180 10.450 42.330 18.000 ;
        RECT 42.780 15.150 42.930 18.000 ;
        RECT 43.530 15.600 45.930 18.800 ;
        RECT 49.280 18.650 50.730 18.950 ;
        RECT 46.530 18.450 50.730 18.650 ;
        RECT 58.730 18.950 70.730 19.800 ;
        RECT 58.730 18.900 69.130 18.950 ;
        RECT 58.730 18.650 60.180 18.900 ;
        RECT 60.330 18.800 69.130 18.900 ;
        RECT 58.730 18.450 62.930 18.650 ;
        RECT 46.530 18.300 54.080 18.450 ;
        RECT 55.430 18.300 62.930 18.450 ;
        RECT 46.530 18.000 50.730 18.300 ;
        RECT 46.530 15.150 46.680 18.000 ;
        RECT 47.130 10.450 47.280 18.000 ;
        RECT 47.730 10.450 47.880 18.000 ;
        RECT 48.330 10.450 48.480 18.000 ;
        RECT 48.930 10.450 49.080 18.000 ;
        RECT 49.530 10.450 49.680 18.000 ;
        RECT 50.130 17.850 50.730 18.000 ;
        RECT 58.730 18.000 62.930 18.300 ;
        RECT 58.730 17.850 59.330 18.000 ;
        RECT 50.130 17.700 54.080 17.850 ;
        RECT 55.380 17.700 59.330 17.850 ;
        RECT 50.130 17.250 50.730 17.700 ;
        RECT 58.730 17.250 59.330 17.700 ;
        RECT 50.130 17.100 54.080 17.250 ;
        RECT 55.380 17.100 59.330 17.250 ;
        RECT 50.130 16.650 50.730 17.100 ;
        RECT 58.730 16.650 59.330 17.100 ;
        RECT 50.130 16.500 54.080 16.650 ;
        RECT 55.380 16.500 59.330 16.650 ;
        RECT 50.130 16.050 50.730 16.500 ;
        RECT 58.730 16.050 59.330 16.500 ;
        RECT 50.130 15.900 54.080 16.050 ;
        RECT 55.380 15.900 59.330 16.050 ;
        RECT 50.130 15.450 50.730 15.900 ;
        RECT 58.730 15.450 59.330 15.900 ;
        RECT 50.130 15.300 54.080 15.450 ;
        RECT 55.380 15.300 59.330 15.450 ;
        RECT 50.130 14.850 50.730 15.300 ;
        RECT 58.730 14.850 59.330 15.300 ;
        RECT 50.130 14.700 54.080 14.850 ;
        RECT 55.380 14.700 59.330 14.850 ;
        RECT 50.130 14.250 50.730 14.700 ;
        RECT 58.730 14.250 59.330 14.700 ;
        RECT 50.130 14.100 54.080 14.250 ;
        RECT 55.380 14.100 59.330 14.250 ;
        RECT 50.130 13.650 50.730 14.100 ;
        RECT 58.730 13.650 59.330 14.100 ;
        RECT 50.130 13.500 54.080 13.650 ;
        RECT 55.380 13.500 59.330 13.650 ;
        RECT 50.130 13.050 50.730 13.500 ;
        RECT 58.730 13.050 59.330 13.500 ;
        RECT 50.130 12.900 54.080 13.050 ;
        RECT 55.380 12.900 59.330 13.050 ;
        RECT 50.130 12.450 50.730 12.900 ;
        RECT 58.730 12.450 59.330 12.900 ;
        RECT 50.130 12.300 54.080 12.450 ;
        RECT 55.380 12.300 59.330 12.450 ;
        RECT 50.130 11.850 50.730 12.300 ;
        RECT 58.730 11.850 59.330 12.300 ;
        RECT 50.130 11.700 54.080 11.850 ;
        RECT 55.380 11.700 59.330 11.850 ;
        RECT 50.130 11.250 50.730 11.700 ;
        RECT 58.730 11.250 59.330 11.700 ;
        RECT 50.130 11.100 54.080 11.250 ;
        RECT 55.380 11.100 59.330 11.250 ;
        RECT 50.130 10.650 50.730 11.100 ;
        RECT 58.730 10.650 59.330 11.100 ;
        RECT 50.130 10.450 54.080 10.650 ;
        RECT 55.380 10.450 59.330 10.650 ;
        RECT 59.780 10.450 59.930 18.000 ;
        RECT 60.380 10.450 60.530 18.000 ;
        RECT 60.980 10.450 61.130 18.000 ;
        RECT 61.580 10.450 61.730 18.000 ;
        RECT 62.180 10.450 62.330 18.000 ;
        RECT 62.780 15.150 62.930 18.000 ;
        RECT 63.530 15.600 65.930 18.800 ;
        RECT 69.280 18.650 70.730 18.950 ;
        RECT 66.530 18.450 70.730 18.650 ;
        RECT 78.730 18.950 90.730 19.800 ;
        RECT 78.730 18.900 89.130 18.950 ;
        RECT 78.730 18.650 80.180 18.900 ;
        RECT 80.330 18.800 89.130 18.900 ;
        RECT 78.730 18.450 82.930 18.650 ;
        RECT 66.530 18.300 74.080 18.450 ;
        RECT 75.430 18.300 82.930 18.450 ;
        RECT 66.530 18.000 70.730 18.300 ;
        RECT 66.530 15.150 66.680 18.000 ;
        RECT 67.130 10.450 67.280 18.000 ;
        RECT 67.730 10.450 67.880 18.000 ;
        RECT 68.330 10.450 68.480 18.000 ;
        RECT 68.930 10.450 69.080 18.000 ;
        RECT 69.530 10.450 69.680 18.000 ;
        RECT 70.130 17.850 70.730 18.000 ;
        RECT 78.730 18.000 82.930 18.300 ;
        RECT 78.730 17.850 79.330 18.000 ;
        RECT 70.130 17.700 74.080 17.850 ;
        RECT 75.380 17.700 79.330 17.850 ;
        RECT 70.130 17.250 70.730 17.700 ;
        RECT 78.730 17.250 79.330 17.700 ;
        RECT 70.130 17.100 74.080 17.250 ;
        RECT 75.380 17.100 79.330 17.250 ;
        RECT 70.130 16.650 70.730 17.100 ;
        RECT 78.730 16.650 79.330 17.100 ;
        RECT 70.130 16.500 74.080 16.650 ;
        RECT 75.380 16.500 79.330 16.650 ;
        RECT 70.130 16.050 70.730 16.500 ;
        RECT 78.730 16.050 79.330 16.500 ;
        RECT 70.130 15.900 74.080 16.050 ;
        RECT 75.380 15.900 79.330 16.050 ;
        RECT 70.130 15.450 70.730 15.900 ;
        RECT 78.730 15.450 79.330 15.900 ;
        RECT 70.130 15.300 74.080 15.450 ;
        RECT 75.380 15.300 79.330 15.450 ;
        RECT 70.130 14.850 70.730 15.300 ;
        RECT 78.730 14.850 79.330 15.300 ;
        RECT 70.130 14.700 74.080 14.850 ;
        RECT 75.380 14.700 79.330 14.850 ;
        RECT 70.130 14.250 70.730 14.700 ;
        RECT 78.730 14.250 79.330 14.700 ;
        RECT 70.130 14.100 74.080 14.250 ;
        RECT 75.380 14.100 79.330 14.250 ;
        RECT 70.130 13.650 70.730 14.100 ;
        RECT 78.730 13.650 79.330 14.100 ;
        RECT 70.130 13.500 74.080 13.650 ;
        RECT 75.380 13.500 79.330 13.650 ;
        RECT 70.130 13.050 70.730 13.500 ;
        RECT 78.730 13.050 79.330 13.500 ;
        RECT 70.130 12.900 74.080 13.050 ;
        RECT 75.380 12.900 79.330 13.050 ;
        RECT 70.130 12.450 70.730 12.900 ;
        RECT 78.730 12.450 79.330 12.900 ;
        RECT 70.130 12.300 74.080 12.450 ;
        RECT 75.380 12.300 79.330 12.450 ;
        RECT 70.130 11.850 70.730 12.300 ;
        RECT 78.730 11.850 79.330 12.300 ;
        RECT 70.130 11.700 74.080 11.850 ;
        RECT 75.380 11.700 79.330 11.850 ;
        RECT 70.130 11.250 70.730 11.700 ;
        RECT 78.730 11.250 79.330 11.700 ;
        RECT 70.130 11.100 74.080 11.250 ;
        RECT 75.380 11.100 79.330 11.250 ;
        RECT 70.130 10.650 70.730 11.100 ;
        RECT 78.730 10.650 79.330 11.100 ;
        RECT 70.130 10.450 74.080 10.650 ;
        RECT 75.380 10.450 79.330 10.650 ;
        RECT 79.780 10.450 79.930 18.000 ;
        RECT 80.380 10.450 80.530 18.000 ;
        RECT 80.980 10.450 81.130 18.000 ;
        RECT 81.580 10.450 81.730 18.000 ;
        RECT 82.180 10.450 82.330 18.000 ;
        RECT 82.780 15.150 82.930 18.000 ;
        RECT 83.530 15.600 85.930 18.800 ;
        RECT 89.280 18.650 90.730 18.950 ;
        RECT 86.530 18.450 90.730 18.650 ;
        RECT 98.730 18.950 110.730 19.800 ;
        RECT 98.730 18.900 109.130 18.950 ;
        RECT 98.730 18.650 100.180 18.900 ;
        RECT 100.330 18.800 109.130 18.900 ;
        RECT 98.730 18.450 102.930 18.650 ;
        RECT 86.530 18.300 94.080 18.450 ;
        RECT 95.430 18.300 102.930 18.450 ;
        RECT 86.530 18.000 90.730 18.300 ;
        RECT 86.530 15.150 86.680 18.000 ;
        RECT 87.130 10.450 87.280 18.000 ;
        RECT 87.730 10.450 87.880 18.000 ;
        RECT 88.330 10.450 88.480 18.000 ;
        RECT 88.930 10.450 89.080 18.000 ;
        RECT 89.530 10.450 89.680 18.000 ;
        RECT 90.130 17.850 90.730 18.000 ;
        RECT 98.730 18.000 102.930 18.300 ;
        RECT 98.730 17.850 99.330 18.000 ;
        RECT 90.130 17.700 94.080 17.850 ;
        RECT 95.380 17.700 99.330 17.850 ;
        RECT 90.130 17.250 90.730 17.700 ;
        RECT 98.730 17.250 99.330 17.700 ;
        RECT 90.130 17.100 94.080 17.250 ;
        RECT 95.380 17.100 99.330 17.250 ;
        RECT 90.130 16.650 90.730 17.100 ;
        RECT 98.730 16.650 99.330 17.100 ;
        RECT 90.130 16.500 94.080 16.650 ;
        RECT 95.380 16.500 99.330 16.650 ;
        RECT 90.130 16.050 90.730 16.500 ;
        RECT 98.730 16.050 99.330 16.500 ;
        RECT 90.130 15.900 94.080 16.050 ;
        RECT 95.380 15.900 99.330 16.050 ;
        RECT 90.130 15.450 90.730 15.900 ;
        RECT 98.730 15.450 99.330 15.900 ;
        RECT 90.130 15.300 94.080 15.450 ;
        RECT 95.380 15.300 99.330 15.450 ;
        RECT 90.130 14.850 90.730 15.300 ;
        RECT 98.730 14.850 99.330 15.300 ;
        RECT 90.130 14.700 94.080 14.850 ;
        RECT 95.380 14.700 99.330 14.850 ;
        RECT 90.130 14.250 90.730 14.700 ;
        RECT 98.730 14.250 99.330 14.700 ;
        RECT 90.130 14.100 94.080 14.250 ;
        RECT 95.380 14.100 99.330 14.250 ;
        RECT 90.130 13.650 90.730 14.100 ;
        RECT 98.730 13.650 99.330 14.100 ;
        RECT 90.130 13.500 94.080 13.650 ;
        RECT 95.380 13.500 99.330 13.650 ;
        RECT 90.130 13.050 90.730 13.500 ;
        RECT 98.730 13.050 99.330 13.500 ;
        RECT 90.130 12.900 94.080 13.050 ;
        RECT 95.380 12.900 99.330 13.050 ;
        RECT 90.130 12.450 90.730 12.900 ;
        RECT 98.730 12.450 99.330 12.900 ;
        RECT 90.130 12.300 94.080 12.450 ;
        RECT 95.380 12.300 99.330 12.450 ;
        RECT 90.130 11.850 90.730 12.300 ;
        RECT 98.730 11.850 99.330 12.300 ;
        RECT 90.130 11.700 94.080 11.850 ;
        RECT 95.380 11.700 99.330 11.850 ;
        RECT 90.130 11.250 90.730 11.700 ;
        RECT 98.730 11.250 99.330 11.700 ;
        RECT 90.130 11.100 94.080 11.250 ;
        RECT 95.380 11.100 99.330 11.250 ;
        RECT 90.130 10.650 90.730 11.100 ;
        RECT 98.730 10.650 99.330 11.100 ;
        RECT 90.130 10.450 94.080 10.650 ;
        RECT 95.380 10.450 99.330 10.650 ;
        RECT 99.780 10.450 99.930 18.000 ;
        RECT 100.380 10.450 100.530 18.000 ;
        RECT 100.980 10.450 101.130 18.000 ;
        RECT 101.580 10.450 101.730 18.000 ;
        RECT 102.180 10.450 102.330 18.000 ;
        RECT 102.780 15.150 102.930 18.000 ;
        RECT 103.530 15.600 105.930 18.800 ;
        RECT 109.280 18.650 110.730 18.950 ;
        RECT 106.530 18.450 110.730 18.650 ;
        RECT 118.730 18.900 124.730 19.800 ;
        RECT 118.730 18.650 120.180 18.900 ;
        RECT 120.330 18.800 124.730 18.900 ;
        RECT 118.730 18.450 122.930 18.650 ;
        RECT 106.530 18.300 114.080 18.450 ;
        RECT 115.430 18.300 122.930 18.450 ;
        RECT 106.530 18.000 110.730 18.300 ;
        RECT 106.530 15.150 106.680 18.000 ;
        RECT 107.130 10.450 107.280 18.000 ;
        RECT 107.730 10.450 107.880 18.000 ;
        RECT 108.330 10.450 108.480 18.000 ;
        RECT 108.930 10.450 109.080 18.000 ;
        RECT 109.530 10.450 109.680 18.000 ;
        RECT 110.130 17.850 110.730 18.000 ;
        RECT 118.730 18.000 122.930 18.300 ;
        RECT 118.730 17.850 119.330 18.000 ;
        RECT 110.130 17.700 114.080 17.850 ;
        RECT 115.380 17.700 119.330 17.850 ;
        RECT 110.130 17.250 110.730 17.700 ;
        RECT 118.730 17.250 119.330 17.700 ;
        RECT 110.130 17.100 114.080 17.250 ;
        RECT 115.380 17.100 119.330 17.250 ;
        RECT 110.130 16.650 110.730 17.100 ;
        RECT 118.730 16.650 119.330 17.100 ;
        RECT 110.130 16.500 114.080 16.650 ;
        RECT 115.380 16.500 119.330 16.650 ;
        RECT 110.130 16.050 110.730 16.500 ;
        RECT 118.730 16.050 119.330 16.500 ;
        RECT 110.130 15.900 114.080 16.050 ;
        RECT 115.380 15.900 119.330 16.050 ;
        RECT 110.130 15.450 110.730 15.900 ;
        RECT 118.730 15.450 119.330 15.900 ;
        RECT 110.130 15.300 114.080 15.450 ;
        RECT 115.380 15.300 119.330 15.450 ;
        RECT 110.130 14.850 110.730 15.300 ;
        RECT 118.730 14.850 119.330 15.300 ;
        RECT 110.130 14.700 114.080 14.850 ;
        RECT 115.380 14.700 119.330 14.850 ;
        RECT 110.130 14.250 110.730 14.700 ;
        RECT 118.730 14.250 119.330 14.700 ;
        RECT 110.130 14.100 114.080 14.250 ;
        RECT 115.380 14.100 119.330 14.250 ;
        RECT 110.130 13.650 110.730 14.100 ;
        RECT 118.730 13.650 119.330 14.100 ;
        RECT 110.130 13.500 114.080 13.650 ;
        RECT 115.380 13.500 119.330 13.650 ;
        RECT 110.130 13.050 110.730 13.500 ;
        RECT 118.730 13.050 119.330 13.500 ;
        RECT 110.130 12.900 114.080 13.050 ;
        RECT 115.380 12.900 119.330 13.050 ;
        RECT 110.130 12.450 110.730 12.900 ;
        RECT 118.730 12.450 119.330 12.900 ;
        RECT 110.130 12.300 114.080 12.450 ;
        RECT 115.380 12.300 119.330 12.450 ;
        RECT 110.130 11.850 110.730 12.300 ;
        RECT 118.730 11.850 119.330 12.300 ;
        RECT 110.130 11.700 114.080 11.850 ;
        RECT 115.380 11.700 119.330 11.850 ;
        RECT 110.130 11.250 110.730 11.700 ;
        RECT 118.730 11.250 119.330 11.700 ;
        RECT 110.130 11.100 114.080 11.250 ;
        RECT 115.380 11.100 119.330 11.250 ;
        RECT 110.130 10.650 110.730 11.100 ;
        RECT 118.730 10.650 119.330 11.100 ;
        RECT 110.130 10.450 114.080 10.650 ;
        RECT 115.380 10.450 119.330 10.650 ;
        RECT 119.780 10.450 119.930 18.000 ;
        RECT 120.380 10.450 120.530 18.000 ;
        RECT 120.980 10.450 121.130 18.000 ;
        RECT 121.580 10.450 121.730 18.000 ;
        RECT 122.180 10.450 122.330 18.000 ;
        RECT 122.780 15.150 122.930 18.000 ;
        RECT 123.530 17.310 124.730 18.800 ;
        RECT 123.530 16.035 127.135 17.310 ;
        RECT 123.530 15.600 124.730 16.035 ;
        RECT 2.315 4.450 4.315 6.745 ;
        RECT 4.730 3.650 5.930 4.400 ;
        RECT 2.315 2.375 5.930 3.650 ;
        RECT 4.730 1.200 5.930 2.375 ;
        RECT 6.530 2.000 6.680 4.900 ;
        RECT 7.130 2.000 7.280 9.550 ;
        RECT 7.730 2.000 7.880 9.550 ;
        RECT 8.330 2.000 8.480 9.550 ;
        RECT 8.930 2.000 9.080 9.550 ;
        RECT 9.530 2.000 9.680 9.550 ;
        RECT 10.130 9.350 14.080 9.550 ;
        RECT 15.380 9.350 19.330 9.550 ;
        RECT 10.130 8.900 10.730 9.350 ;
        RECT 18.730 8.900 19.330 9.350 ;
        RECT 10.130 8.750 14.080 8.900 ;
        RECT 15.380 8.750 19.330 8.900 ;
        RECT 10.130 8.300 10.730 8.750 ;
        RECT 18.730 8.300 19.330 8.750 ;
        RECT 10.130 8.150 14.080 8.300 ;
        RECT 15.380 8.150 19.330 8.300 ;
        RECT 10.130 7.700 10.730 8.150 ;
        RECT 18.730 7.700 19.330 8.150 ;
        RECT 10.130 7.550 14.080 7.700 ;
        RECT 15.380 7.550 19.330 7.700 ;
        RECT 10.130 7.100 10.730 7.550 ;
        RECT 18.730 7.100 19.330 7.550 ;
        RECT 10.130 6.950 14.080 7.100 ;
        RECT 15.380 6.950 19.330 7.100 ;
        RECT 10.130 6.500 10.730 6.950 ;
        RECT 18.730 6.500 19.330 6.950 ;
        RECT 10.130 6.350 14.080 6.500 ;
        RECT 15.380 6.350 19.330 6.500 ;
        RECT 10.130 5.900 10.730 6.350 ;
        RECT 18.730 5.900 19.330 6.350 ;
        RECT 10.130 5.750 14.080 5.900 ;
        RECT 15.380 5.750 19.330 5.900 ;
        RECT 10.130 5.300 10.730 5.750 ;
        RECT 18.730 5.300 19.330 5.750 ;
        RECT 10.130 5.150 14.080 5.300 ;
        RECT 15.380 5.150 19.330 5.300 ;
        RECT 10.130 4.700 10.730 5.150 ;
        RECT 18.730 4.700 19.330 5.150 ;
        RECT 10.130 4.550 14.080 4.700 ;
        RECT 15.380 4.550 19.330 4.700 ;
        RECT 10.130 4.100 10.730 4.550 ;
        RECT 18.730 4.100 19.330 4.550 ;
        RECT 10.130 3.950 14.080 4.100 ;
        RECT 15.380 3.950 19.330 4.100 ;
        RECT 10.130 3.500 10.730 3.950 ;
        RECT 18.730 3.500 19.330 3.950 ;
        RECT 10.130 3.350 14.080 3.500 ;
        RECT 15.380 3.350 19.330 3.500 ;
        RECT 10.130 2.900 10.730 3.350 ;
        RECT 18.730 2.900 19.330 3.350 ;
        RECT 10.130 2.750 14.080 2.900 ;
        RECT 15.380 2.750 19.330 2.900 ;
        RECT 10.130 2.300 10.730 2.750 ;
        RECT 18.730 2.300 19.330 2.750 ;
        RECT 10.130 2.150 14.080 2.300 ;
        RECT 15.380 2.150 19.330 2.300 ;
        RECT 10.130 2.000 10.730 2.150 ;
        RECT 6.530 1.700 10.730 2.000 ;
        RECT 18.730 2.000 19.330 2.150 ;
        RECT 19.780 2.000 19.930 9.550 ;
        RECT 20.380 2.000 20.530 9.550 ;
        RECT 20.980 2.000 21.130 9.550 ;
        RECT 21.580 2.000 21.730 9.550 ;
        RECT 22.180 2.000 22.330 9.550 ;
        RECT 22.780 2.000 22.930 4.900 ;
        RECT 18.730 1.700 22.930 2.000 ;
        RECT 6.530 1.550 14.080 1.700 ;
        RECT 15.380 1.550 22.930 1.700 ;
        RECT 6.530 1.350 10.730 1.550 ;
        RECT 4.730 1.050 9.130 1.200 ;
        RECT 9.280 1.050 10.730 1.350 ;
        RECT 4.730 0.150 10.730 1.050 ;
        RECT 18.730 1.350 22.930 1.550 ;
        RECT 18.730 1.050 20.180 1.350 ;
        RECT 23.530 1.200 25.930 4.400 ;
        RECT 26.530 2.000 26.680 4.900 ;
        RECT 27.130 2.000 27.280 9.550 ;
        RECT 27.730 2.000 27.880 9.550 ;
        RECT 28.330 2.000 28.480 9.550 ;
        RECT 28.930 2.000 29.080 9.550 ;
        RECT 29.530 2.000 29.680 9.550 ;
        RECT 30.130 9.350 34.080 9.550 ;
        RECT 35.380 9.350 39.330 9.550 ;
        RECT 30.130 8.900 30.730 9.350 ;
        RECT 38.730 8.900 39.330 9.350 ;
        RECT 30.130 8.750 34.080 8.900 ;
        RECT 35.380 8.750 39.330 8.900 ;
        RECT 30.130 8.300 30.730 8.750 ;
        RECT 38.730 8.300 39.330 8.750 ;
        RECT 30.130 8.150 34.080 8.300 ;
        RECT 35.380 8.150 39.330 8.300 ;
        RECT 30.130 7.700 30.730 8.150 ;
        RECT 38.730 7.700 39.330 8.150 ;
        RECT 30.130 7.550 34.080 7.700 ;
        RECT 35.380 7.550 39.330 7.700 ;
        RECT 30.130 7.100 30.730 7.550 ;
        RECT 38.730 7.100 39.330 7.550 ;
        RECT 30.130 6.950 34.080 7.100 ;
        RECT 35.380 6.950 39.330 7.100 ;
        RECT 30.130 6.500 30.730 6.950 ;
        RECT 38.730 6.500 39.330 6.950 ;
        RECT 30.130 6.350 34.080 6.500 ;
        RECT 35.380 6.350 39.330 6.500 ;
        RECT 30.130 5.900 30.730 6.350 ;
        RECT 38.730 5.900 39.330 6.350 ;
        RECT 30.130 5.750 34.080 5.900 ;
        RECT 35.380 5.750 39.330 5.900 ;
        RECT 30.130 5.300 30.730 5.750 ;
        RECT 38.730 5.300 39.330 5.750 ;
        RECT 30.130 5.150 34.080 5.300 ;
        RECT 35.380 5.150 39.330 5.300 ;
        RECT 30.130 4.700 30.730 5.150 ;
        RECT 38.730 4.700 39.330 5.150 ;
        RECT 30.130 4.550 34.080 4.700 ;
        RECT 35.380 4.550 39.330 4.700 ;
        RECT 30.130 4.100 30.730 4.550 ;
        RECT 38.730 4.100 39.330 4.550 ;
        RECT 30.130 3.950 34.080 4.100 ;
        RECT 35.380 3.950 39.330 4.100 ;
        RECT 30.130 3.500 30.730 3.950 ;
        RECT 38.730 3.500 39.330 3.950 ;
        RECT 30.130 3.350 34.080 3.500 ;
        RECT 35.380 3.350 39.330 3.500 ;
        RECT 30.130 2.900 30.730 3.350 ;
        RECT 38.730 2.900 39.330 3.350 ;
        RECT 30.130 2.750 34.080 2.900 ;
        RECT 35.380 2.750 39.330 2.900 ;
        RECT 30.130 2.300 30.730 2.750 ;
        RECT 38.730 2.300 39.330 2.750 ;
        RECT 30.130 2.150 34.080 2.300 ;
        RECT 35.380 2.150 39.330 2.300 ;
        RECT 30.130 2.000 30.730 2.150 ;
        RECT 26.530 1.700 30.730 2.000 ;
        RECT 38.730 2.000 39.330 2.150 ;
        RECT 39.780 2.000 39.930 9.550 ;
        RECT 40.380 2.000 40.530 9.550 ;
        RECT 40.980 2.000 41.130 9.550 ;
        RECT 41.580 2.000 41.730 9.550 ;
        RECT 42.180 2.000 42.330 9.550 ;
        RECT 42.780 2.000 42.930 4.900 ;
        RECT 38.730 1.700 42.930 2.000 ;
        RECT 26.530 1.550 34.080 1.700 ;
        RECT 35.380 1.550 42.930 1.700 ;
        RECT 26.530 1.350 30.730 1.550 ;
        RECT 20.330 1.050 29.130 1.200 ;
        RECT 29.280 1.050 30.730 1.350 ;
        RECT 18.730 0.150 30.730 1.050 ;
        RECT 38.730 1.350 42.930 1.550 ;
        RECT 38.730 1.050 40.180 1.350 ;
        RECT 43.530 1.200 45.930 4.400 ;
        RECT 46.530 2.000 46.680 4.900 ;
        RECT 47.130 2.000 47.280 9.550 ;
        RECT 47.730 2.000 47.880 9.550 ;
        RECT 48.330 2.000 48.480 9.550 ;
        RECT 48.930 2.000 49.080 9.550 ;
        RECT 49.530 2.000 49.680 9.550 ;
        RECT 50.130 9.350 54.080 9.550 ;
        RECT 55.380 9.350 59.330 9.550 ;
        RECT 50.130 8.900 50.730 9.350 ;
        RECT 58.730 8.900 59.330 9.350 ;
        RECT 50.130 8.750 54.080 8.900 ;
        RECT 55.380 8.750 59.330 8.900 ;
        RECT 50.130 8.300 50.730 8.750 ;
        RECT 58.730 8.300 59.330 8.750 ;
        RECT 50.130 8.150 54.080 8.300 ;
        RECT 55.380 8.150 59.330 8.300 ;
        RECT 50.130 7.700 50.730 8.150 ;
        RECT 58.730 7.700 59.330 8.150 ;
        RECT 50.130 7.550 54.080 7.700 ;
        RECT 55.380 7.550 59.330 7.700 ;
        RECT 50.130 7.100 50.730 7.550 ;
        RECT 58.730 7.100 59.330 7.550 ;
        RECT 50.130 6.950 54.080 7.100 ;
        RECT 55.380 6.950 59.330 7.100 ;
        RECT 50.130 6.500 50.730 6.950 ;
        RECT 58.730 6.500 59.330 6.950 ;
        RECT 50.130 6.350 54.080 6.500 ;
        RECT 55.380 6.350 59.330 6.500 ;
        RECT 50.130 5.900 50.730 6.350 ;
        RECT 58.730 5.900 59.330 6.350 ;
        RECT 50.130 5.750 54.080 5.900 ;
        RECT 55.380 5.750 59.330 5.900 ;
        RECT 50.130 5.300 50.730 5.750 ;
        RECT 58.730 5.300 59.330 5.750 ;
        RECT 50.130 5.150 54.080 5.300 ;
        RECT 55.380 5.150 59.330 5.300 ;
        RECT 50.130 4.700 50.730 5.150 ;
        RECT 58.730 4.700 59.330 5.150 ;
        RECT 50.130 4.550 54.080 4.700 ;
        RECT 55.380 4.550 59.330 4.700 ;
        RECT 50.130 4.100 50.730 4.550 ;
        RECT 58.730 4.100 59.330 4.550 ;
        RECT 50.130 3.950 54.080 4.100 ;
        RECT 55.380 3.950 59.330 4.100 ;
        RECT 50.130 3.500 50.730 3.950 ;
        RECT 58.730 3.500 59.330 3.950 ;
        RECT 50.130 3.350 54.080 3.500 ;
        RECT 55.380 3.350 59.330 3.500 ;
        RECT 50.130 2.900 50.730 3.350 ;
        RECT 58.730 2.900 59.330 3.350 ;
        RECT 50.130 2.750 54.080 2.900 ;
        RECT 55.380 2.750 59.330 2.900 ;
        RECT 50.130 2.300 50.730 2.750 ;
        RECT 58.730 2.300 59.330 2.750 ;
        RECT 50.130 2.150 54.080 2.300 ;
        RECT 55.380 2.150 59.330 2.300 ;
        RECT 50.130 2.000 50.730 2.150 ;
        RECT 46.530 1.700 50.730 2.000 ;
        RECT 58.730 2.000 59.330 2.150 ;
        RECT 59.780 2.000 59.930 9.550 ;
        RECT 60.380 2.000 60.530 9.550 ;
        RECT 60.980 2.000 61.130 9.550 ;
        RECT 61.580 2.000 61.730 9.550 ;
        RECT 62.180 2.000 62.330 9.550 ;
        RECT 62.780 2.000 62.930 4.900 ;
        RECT 58.730 1.700 62.930 2.000 ;
        RECT 46.530 1.550 54.080 1.700 ;
        RECT 55.380 1.550 62.930 1.700 ;
        RECT 46.530 1.350 50.730 1.550 ;
        RECT 40.330 1.050 49.130 1.200 ;
        RECT 49.280 1.050 50.730 1.350 ;
        RECT 38.730 0.150 50.730 1.050 ;
        RECT 58.730 1.350 62.930 1.550 ;
        RECT 58.730 1.050 60.180 1.350 ;
        RECT 63.530 1.200 65.930 4.400 ;
        RECT 66.530 2.000 66.680 4.900 ;
        RECT 67.130 2.000 67.280 9.550 ;
        RECT 67.730 2.000 67.880 9.550 ;
        RECT 68.330 2.000 68.480 9.550 ;
        RECT 68.930 2.000 69.080 9.550 ;
        RECT 69.530 2.000 69.680 9.550 ;
        RECT 70.130 9.350 74.080 9.550 ;
        RECT 75.380 9.350 79.330 9.550 ;
        RECT 70.130 8.900 70.730 9.350 ;
        RECT 78.730 8.900 79.330 9.350 ;
        RECT 70.130 8.750 74.080 8.900 ;
        RECT 75.380 8.750 79.330 8.900 ;
        RECT 70.130 8.300 70.730 8.750 ;
        RECT 78.730 8.300 79.330 8.750 ;
        RECT 70.130 8.150 74.080 8.300 ;
        RECT 75.380 8.150 79.330 8.300 ;
        RECT 70.130 7.700 70.730 8.150 ;
        RECT 78.730 7.700 79.330 8.150 ;
        RECT 70.130 7.550 74.080 7.700 ;
        RECT 75.380 7.550 79.330 7.700 ;
        RECT 70.130 7.100 70.730 7.550 ;
        RECT 78.730 7.100 79.330 7.550 ;
        RECT 70.130 6.950 74.080 7.100 ;
        RECT 75.380 6.950 79.330 7.100 ;
        RECT 70.130 6.500 70.730 6.950 ;
        RECT 78.730 6.500 79.330 6.950 ;
        RECT 70.130 6.350 74.080 6.500 ;
        RECT 75.380 6.350 79.330 6.500 ;
        RECT 70.130 5.900 70.730 6.350 ;
        RECT 78.730 5.900 79.330 6.350 ;
        RECT 70.130 5.750 74.080 5.900 ;
        RECT 75.380 5.750 79.330 5.900 ;
        RECT 70.130 5.300 70.730 5.750 ;
        RECT 78.730 5.300 79.330 5.750 ;
        RECT 70.130 5.150 74.080 5.300 ;
        RECT 75.380 5.150 79.330 5.300 ;
        RECT 70.130 4.700 70.730 5.150 ;
        RECT 78.730 4.700 79.330 5.150 ;
        RECT 70.130 4.550 74.080 4.700 ;
        RECT 75.380 4.550 79.330 4.700 ;
        RECT 70.130 4.100 70.730 4.550 ;
        RECT 78.730 4.100 79.330 4.550 ;
        RECT 70.130 3.950 74.080 4.100 ;
        RECT 75.380 3.950 79.330 4.100 ;
        RECT 70.130 3.500 70.730 3.950 ;
        RECT 78.730 3.500 79.330 3.950 ;
        RECT 70.130 3.350 74.080 3.500 ;
        RECT 75.380 3.350 79.330 3.500 ;
        RECT 70.130 2.900 70.730 3.350 ;
        RECT 78.730 2.900 79.330 3.350 ;
        RECT 70.130 2.750 74.080 2.900 ;
        RECT 75.380 2.750 79.330 2.900 ;
        RECT 70.130 2.300 70.730 2.750 ;
        RECT 78.730 2.300 79.330 2.750 ;
        RECT 70.130 2.150 74.080 2.300 ;
        RECT 75.380 2.150 79.330 2.300 ;
        RECT 70.130 2.000 70.730 2.150 ;
        RECT 66.530 1.700 70.730 2.000 ;
        RECT 78.730 2.000 79.330 2.150 ;
        RECT 79.780 2.000 79.930 9.550 ;
        RECT 80.380 2.000 80.530 9.550 ;
        RECT 80.980 2.000 81.130 9.550 ;
        RECT 81.580 2.000 81.730 9.550 ;
        RECT 82.180 2.000 82.330 9.550 ;
        RECT 82.780 2.000 82.930 4.900 ;
        RECT 78.730 1.700 82.930 2.000 ;
        RECT 66.530 1.550 74.080 1.700 ;
        RECT 75.380 1.550 82.930 1.700 ;
        RECT 66.530 1.350 70.730 1.550 ;
        RECT 60.330 1.050 69.130 1.200 ;
        RECT 69.280 1.050 70.730 1.350 ;
        RECT 58.730 0.150 70.730 1.050 ;
        RECT 78.730 1.350 82.930 1.550 ;
        RECT 78.730 1.050 80.180 1.350 ;
        RECT 83.530 1.200 85.930 4.400 ;
        RECT 86.530 2.000 86.680 4.900 ;
        RECT 87.130 2.000 87.280 9.550 ;
        RECT 87.730 2.000 87.880 9.550 ;
        RECT 88.330 2.000 88.480 9.550 ;
        RECT 88.930 2.000 89.080 9.550 ;
        RECT 89.530 2.000 89.680 9.550 ;
        RECT 90.130 9.350 94.080 9.550 ;
        RECT 95.380 9.350 99.330 9.550 ;
        RECT 90.130 8.900 90.730 9.350 ;
        RECT 98.730 8.900 99.330 9.350 ;
        RECT 90.130 8.750 94.080 8.900 ;
        RECT 95.380 8.750 99.330 8.900 ;
        RECT 90.130 8.300 90.730 8.750 ;
        RECT 98.730 8.300 99.330 8.750 ;
        RECT 90.130 8.150 94.080 8.300 ;
        RECT 95.380 8.150 99.330 8.300 ;
        RECT 90.130 7.700 90.730 8.150 ;
        RECT 98.730 7.700 99.330 8.150 ;
        RECT 90.130 7.550 94.080 7.700 ;
        RECT 95.380 7.550 99.330 7.700 ;
        RECT 90.130 7.100 90.730 7.550 ;
        RECT 98.730 7.100 99.330 7.550 ;
        RECT 90.130 6.950 94.080 7.100 ;
        RECT 95.380 6.950 99.330 7.100 ;
        RECT 90.130 6.500 90.730 6.950 ;
        RECT 98.730 6.500 99.330 6.950 ;
        RECT 90.130 6.350 94.080 6.500 ;
        RECT 95.380 6.350 99.330 6.500 ;
        RECT 90.130 5.900 90.730 6.350 ;
        RECT 98.730 5.900 99.330 6.350 ;
        RECT 90.130 5.750 94.080 5.900 ;
        RECT 95.380 5.750 99.330 5.900 ;
        RECT 90.130 5.300 90.730 5.750 ;
        RECT 98.730 5.300 99.330 5.750 ;
        RECT 90.130 5.150 94.080 5.300 ;
        RECT 95.380 5.150 99.330 5.300 ;
        RECT 90.130 4.700 90.730 5.150 ;
        RECT 98.730 4.700 99.330 5.150 ;
        RECT 90.130 4.550 94.080 4.700 ;
        RECT 95.380 4.550 99.330 4.700 ;
        RECT 90.130 4.100 90.730 4.550 ;
        RECT 98.730 4.100 99.330 4.550 ;
        RECT 90.130 3.950 94.080 4.100 ;
        RECT 95.380 3.950 99.330 4.100 ;
        RECT 90.130 3.500 90.730 3.950 ;
        RECT 98.730 3.500 99.330 3.950 ;
        RECT 90.130 3.350 94.080 3.500 ;
        RECT 95.380 3.350 99.330 3.500 ;
        RECT 90.130 2.900 90.730 3.350 ;
        RECT 98.730 2.900 99.330 3.350 ;
        RECT 90.130 2.750 94.080 2.900 ;
        RECT 95.380 2.750 99.330 2.900 ;
        RECT 90.130 2.300 90.730 2.750 ;
        RECT 98.730 2.300 99.330 2.750 ;
        RECT 90.130 2.150 94.080 2.300 ;
        RECT 95.380 2.150 99.330 2.300 ;
        RECT 90.130 2.000 90.730 2.150 ;
        RECT 86.530 1.700 90.730 2.000 ;
        RECT 98.730 2.000 99.330 2.150 ;
        RECT 99.780 2.000 99.930 9.550 ;
        RECT 100.380 2.000 100.530 9.550 ;
        RECT 100.980 2.000 101.130 9.550 ;
        RECT 101.580 2.000 101.730 9.550 ;
        RECT 102.180 2.000 102.330 9.550 ;
        RECT 102.780 2.000 102.930 4.900 ;
        RECT 98.730 1.700 102.930 2.000 ;
        RECT 86.530 1.550 94.080 1.700 ;
        RECT 95.380 1.550 102.930 1.700 ;
        RECT 86.530 1.350 90.730 1.550 ;
        RECT 80.330 1.050 89.130 1.200 ;
        RECT 89.280 1.050 90.730 1.350 ;
        RECT 78.730 0.150 90.730 1.050 ;
        RECT 98.730 1.350 102.930 1.550 ;
        RECT 98.730 1.050 100.180 1.350 ;
        RECT 103.530 1.200 105.930 4.400 ;
        RECT 106.530 2.000 106.680 4.900 ;
        RECT 107.130 2.000 107.280 9.550 ;
        RECT 107.730 2.000 107.880 9.550 ;
        RECT 108.330 2.000 108.480 9.550 ;
        RECT 108.930 2.000 109.080 9.550 ;
        RECT 109.530 2.000 109.680 9.550 ;
        RECT 110.130 9.350 114.080 9.550 ;
        RECT 115.380 9.350 119.330 9.550 ;
        RECT 110.130 8.900 110.730 9.350 ;
        RECT 118.730 8.900 119.330 9.350 ;
        RECT 110.130 8.750 114.080 8.900 ;
        RECT 115.380 8.750 119.330 8.900 ;
        RECT 110.130 8.300 110.730 8.750 ;
        RECT 118.730 8.300 119.330 8.750 ;
        RECT 110.130 8.150 114.080 8.300 ;
        RECT 115.380 8.150 119.330 8.300 ;
        RECT 110.130 7.700 110.730 8.150 ;
        RECT 118.730 7.700 119.330 8.150 ;
        RECT 110.130 7.550 114.080 7.700 ;
        RECT 115.380 7.550 119.330 7.700 ;
        RECT 110.130 7.100 110.730 7.550 ;
        RECT 118.730 7.100 119.330 7.550 ;
        RECT 110.130 6.950 114.080 7.100 ;
        RECT 115.380 6.950 119.330 7.100 ;
        RECT 110.130 6.500 110.730 6.950 ;
        RECT 118.730 6.500 119.330 6.950 ;
        RECT 110.130 6.350 114.080 6.500 ;
        RECT 115.380 6.350 119.330 6.500 ;
        RECT 110.130 5.900 110.730 6.350 ;
        RECT 118.730 5.900 119.330 6.350 ;
        RECT 110.130 5.750 114.080 5.900 ;
        RECT 115.380 5.750 119.330 5.900 ;
        RECT 110.130 5.300 110.730 5.750 ;
        RECT 118.730 5.300 119.330 5.750 ;
        RECT 110.130 5.150 114.080 5.300 ;
        RECT 115.380 5.150 119.330 5.300 ;
        RECT 110.130 4.700 110.730 5.150 ;
        RECT 118.730 4.700 119.330 5.150 ;
        RECT 110.130 4.550 114.080 4.700 ;
        RECT 115.380 4.550 119.330 4.700 ;
        RECT 110.130 4.100 110.730 4.550 ;
        RECT 118.730 4.100 119.330 4.550 ;
        RECT 110.130 3.950 114.080 4.100 ;
        RECT 115.380 3.950 119.330 4.100 ;
        RECT 110.130 3.500 110.730 3.950 ;
        RECT 118.730 3.500 119.330 3.950 ;
        RECT 110.130 3.350 114.080 3.500 ;
        RECT 115.380 3.350 119.330 3.500 ;
        RECT 110.130 2.900 110.730 3.350 ;
        RECT 118.730 2.900 119.330 3.350 ;
        RECT 110.130 2.750 114.080 2.900 ;
        RECT 115.380 2.750 119.330 2.900 ;
        RECT 110.130 2.300 110.730 2.750 ;
        RECT 118.730 2.300 119.330 2.750 ;
        RECT 110.130 2.150 114.080 2.300 ;
        RECT 115.380 2.150 119.330 2.300 ;
        RECT 110.130 2.000 110.730 2.150 ;
        RECT 106.530 1.700 110.730 2.000 ;
        RECT 118.730 2.000 119.330 2.150 ;
        RECT 119.780 2.000 119.930 9.550 ;
        RECT 120.380 2.000 120.530 9.550 ;
        RECT 120.980 2.000 121.130 9.550 ;
        RECT 121.580 2.000 121.730 9.550 ;
        RECT 122.180 2.000 122.330 9.550 ;
        RECT 122.780 2.000 122.930 4.900 ;
        RECT 118.730 1.700 122.930 2.000 ;
        RECT 106.530 1.550 114.080 1.700 ;
        RECT 115.380 1.550 122.930 1.700 ;
        RECT 106.530 1.350 110.730 1.550 ;
        RECT 100.330 1.050 109.130 1.200 ;
        RECT 109.280 1.050 110.730 1.350 ;
        RECT 98.730 0.150 110.730 1.050 ;
        RECT 118.730 1.350 122.930 1.550 ;
        RECT 123.530 3.095 124.730 4.400 ;
        RECT 123.530 1.820 127.140 3.095 ;
        RECT 118.730 1.050 120.180 1.350 ;
        RECT 123.530 1.200 124.730 1.820 ;
        RECT 120.330 1.050 124.730 1.200 ;
        RECT 118.730 0.150 124.730 1.050 ;
        RECT 4.730 0.000 9.130 0.150 ;
        RECT 20.330 0.000 29.130 0.150 ;
        RECT 40.330 0.000 49.130 0.150 ;
        RECT 60.330 0.000 69.130 0.150 ;
        RECT 80.330 0.000 89.130 0.150 ;
        RECT 100.330 0.000 109.130 0.150 ;
        RECT 120.330 0.000 124.730 0.150 ;
      LAYER via ;
        RECT 4.830 338.900 5.830 339.900 ;
        RECT 6.430 338.900 7.430 339.900 ;
        RECT 8.030 338.900 9.030 339.900 ;
        RECT 4.830 337.300 5.830 338.300 ;
        RECT 2.515 336.880 2.875 337.260 ;
        RECT 3.145 336.880 3.505 337.260 ;
        RECT 3.745 336.880 4.105 337.260 ;
        RECT 2.515 336.290 2.875 336.670 ;
        RECT 3.145 336.290 3.505 336.670 ;
        RECT 3.745 336.290 4.105 336.670 ;
        RECT 4.830 335.700 5.830 336.700 ;
        RECT 20.430 338.900 21.430 339.900 ;
        RECT 22.030 338.900 23.030 339.900 ;
        RECT 23.630 338.900 24.630 339.900 ;
        RECT 24.830 338.900 25.830 339.900 ;
        RECT 26.430 338.900 27.430 339.900 ;
        RECT 28.030 338.900 29.030 339.900 ;
        RECT 2.520 334.920 2.880 335.300 ;
        RECT 3.130 334.920 3.490 335.300 ;
        RECT 3.760 334.920 4.120 335.300 ;
        RECT 2.520 334.185 2.880 334.565 ;
        RECT 3.130 334.185 3.490 334.565 ;
        RECT 3.760 334.185 4.120 334.565 ;
        RECT 2.520 333.500 2.880 333.880 ;
        RECT 3.130 333.500 3.490 333.880 ;
        RECT 3.760 333.500 4.120 333.880 ;
        RECT 23.630 337.300 24.630 338.300 ;
        RECT 24.830 337.300 25.830 338.300 ;
        RECT 23.630 335.700 24.630 336.700 ;
        RECT 24.830 335.700 25.830 336.700 ;
        RECT 40.430 338.900 41.430 339.900 ;
        RECT 42.030 338.900 43.030 339.900 ;
        RECT 43.630 338.900 44.630 339.900 ;
        RECT 44.830 338.900 45.830 339.900 ;
        RECT 46.430 338.900 47.430 339.900 ;
        RECT 48.030 338.900 49.030 339.900 ;
        RECT 43.630 337.300 44.630 338.300 ;
        RECT 44.830 337.300 45.830 338.300 ;
        RECT 43.630 335.700 44.630 336.700 ;
        RECT 44.830 335.700 45.830 336.700 ;
        RECT 60.430 338.900 61.430 339.900 ;
        RECT 62.030 338.900 63.030 339.900 ;
        RECT 63.630 338.900 64.630 339.900 ;
        RECT 64.830 338.900 65.830 339.900 ;
        RECT 66.430 338.900 67.430 339.900 ;
        RECT 68.030 338.900 69.030 339.900 ;
        RECT 63.630 337.300 64.630 338.300 ;
        RECT 64.830 337.300 65.830 338.300 ;
        RECT 63.630 335.700 64.630 336.700 ;
        RECT 64.830 335.700 65.830 336.700 ;
        RECT 80.430 338.900 81.430 339.900 ;
        RECT 82.030 338.900 83.030 339.900 ;
        RECT 83.630 338.900 84.630 339.900 ;
        RECT 84.830 338.900 85.830 339.900 ;
        RECT 86.430 338.900 87.430 339.900 ;
        RECT 88.030 338.900 89.030 339.900 ;
        RECT 83.630 337.300 84.630 338.300 ;
        RECT 84.830 337.300 85.830 338.300 ;
        RECT 83.630 335.700 84.630 336.700 ;
        RECT 84.830 335.700 85.830 336.700 ;
        RECT 100.430 338.900 101.430 339.900 ;
        RECT 102.030 338.900 103.030 339.900 ;
        RECT 103.630 338.900 104.630 339.900 ;
        RECT 104.830 338.900 105.830 339.900 ;
        RECT 106.430 338.900 107.430 339.900 ;
        RECT 108.030 338.900 109.030 339.900 ;
        RECT 103.630 337.300 104.630 338.300 ;
        RECT 104.830 337.300 105.830 338.300 ;
        RECT 103.630 335.700 104.630 336.700 ;
        RECT 104.830 335.700 105.830 336.700 ;
        RECT 120.430 338.900 121.430 339.900 ;
        RECT 122.030 338.900 123.030 339.900 ;
        RECT 123.630 338.900 124.630 339.900 ;
        RECT 123.630 337.300 124.630 338.300 ;
        RECT 125.340 337.080 125.700 337.460 ;
        RECT 125.970 337.080 126.330 337.460 ;
        RECT 126.570 337.080 126.930 337.460 ;
        RECT 123.630 335.700 124.630 336.700 ;
        RECT 125.340 336.490 125.700 336.870 ;
        RECT 125.970 336.490 126.330 336.870 ;
        RECT 126.570 336.490 126.930 336.870 ;
        RECT 2.520 326.120 2.880 326.500 ;
        RECT 3.130 326.120 3.490 326.500 ;
        RECT 3.760 326.120 4.120 326.500 ;
        RECT 2.520 325.385 2.880 325.765 ;
        RECT 3.130 325.385 3.490 325.765 ;
        RECT 3.760 325.385 4.120 325.765 ;
        RECT 2.520 324.700 2.880 325.080 ;
        RECT 3.130 324.700 3.490 325.080 ;
        RECT 3.760 324.700 4.120 325.080 ;
        RECT 2.515 323.515 2.875 323.895 ;
        RECT 3.145 323.515 3.505 323.895 ;
        RECT 3.745 323.515 4.105 323.895 ;
        RECT 2.515 322.925 2.875 323.305 ;
        RECT 3.145 322.925 3.505 323.305 ;
        RECT 3.745 322.925 4.105 323.305 ;
        RECT 4.830 323.300 5.830 324.300 ;
        RECT 4.830 321.700 5.830 322.700 ;
        RECT 4.830 320.100 5.830 321.100 ;
        RECT 6.430 320.100 7.430 321.100 ;
        RECT 8.030 320.100 9.030 321.100 ;
        RECT 23.630 323.300 24.630 324.300 ;
        RECT 24.830 323.300 25.830 324.300 ;
        RECT 23.630 321.700 24.630 322.700 ;
        RECT 24.830 321.700 25.830 322.700 ;
        RECT 4.830 318.900 5.830 319.900 ;
        RECT 6.430 318.900 7.430 319.900 ;
        RECT 8.030 318.900 9.030 319.900 ;
        RECT 20.430 320.100 21.430 321.100 ;
        RECT 22.030 320.100 23.030 321.100 ;
        RECT 23.630 320.100 24.630 321.100 ;
        RECT 24.830 320.100 25.830 321.100 ;
        RECT 26.430 320.100 27.430 321.100 ;
        RECT 28.030 320.100 29.030 321.100 ;
        RECT 43.630 323.300 44.630 324.300 ;
        RECT 44.830 323.300 45.830 324.300 ;
        RECT 43.630 321.700 44.630 322.700 ;
        RECT 44.830 321.700 45.830 322.700 ;
        RECT 4.830 317.300 5.830 318.300 ;
        RECT 2.515 316.870 2.875 317.250 ;
        RECT 3.145 316.870 3.505 317.250 ;
        RECT 3.745 316.870 4.105 317.250 ;
        RECT 2.515 316.280 2.875 316.660 ;
        RECT 3.145 316.280 3.505 316.660 ;
        RECT 3.745 316.280 4.105 316.660 ;
        RECT 4.830 315.700 5.830 316.700 ;
        RECT 20.430 318.900 21.430 319.900 ;
        RECT 22.030 318.900 23.030 319.900 ;
        RECT 23.630 318.900 24.630 319.900 ;
        RECT 24.830 318.900 25.830 319.900 ;
        RECT 26.430 318.900 27.430 319.900 ;
        RECT 28.030 318.900 29.030 319.900 ;
        RECT 40.430 320.100 41.430 321.100 ;
        RECT 42.030 320.100 43.030 321.100 ;
        RECT 43.630 320.100 44.630 321.100 ;
        RECT 44.830 320.100 45.830 321.100 ;
        RECT 46.430 320.100 47.430 321.100 ;
        RECT 48.030 320.100 49.030 321.100 ;
        RECT 63.630 323.300 64.630 324.300 ;
        RECT 64.830 323.300 65.830 324.300 ;
        RECT 63.630 321.700 64.630 322.700 ;
        RECT 64.830 321.700 65.830 322.700 ;
        RECT 2.520 314.920 2.880 315.300 ;
        RECT 3.130 314.920 3.490 315.300 ;
        RECT 3.760 314.920 4.120 315.300 ;
        RECT 2.520 314.185 2.880 314.565 ;
        RECT 3.130 314.185 3.490 314.565 ;
        RECT 3.760 314.185 4.120 314.565 ;
        RECT 2.520 313.500 2.880 313.880 ;
        RECT 3.130 313.500 3.490 313.880 ;
        RECT 3.760 313.500 4.120 313.880 ;
        RECT 23.630 317.300 24.630 318.300 ;
        RECT 24.830 317.300 25.830 318.300 ;
        RECT 23.630 315.700 24.630 316.700 ;
        RECT 24.830 315.700 25.830 316.700 ;
        RECT 40.430 318.900 41.430 319.900 ;
        RECT 42.030 318.900 43.030 319.900 ;
        RECT 43.630 318.900 44.630 319.900 ;
        RECT 44.830 318.900 45.830 319.900 ;
        RECT 46.430 318.900 47.430 319.900 ;
        RECT 48.030 318.900 49.030 319.900 ;
        RECT 60.430 320.100 61.430 321.100 ;
        RECT 62.030 320.100 63.030 321.100 ;
        RECT 63.630 320.100 64.630 321.100 ;
        RECT 64.830 320.100 65.830 321.100 ;
        RECT 66.430 320.100 67.430 321.100 ;
        RECT 68.030 320.100 69.030 321.100 ;
        RECT 83.630 323.300 84.630 324.300 ;
        RECT 84.830 323.300 85.830 324.300 ;
        RECT 83.630 321.700 84.630 322.700 ;
        RECT 84.830 321.700 85.830 322.700 ;
        RECT 43.630 317.300 44.630 318.300 ;
        RECT 44.830 317.300 45.830 318.300 ;
        RECT 43.630 315.700 44.630 316.700 ;
        RECT 44.830 315.700 45.830 316.700 ;
        RECT 60.430 318.900 61.430 319.900 ;
        RECT 62.030 318.900 63.030 319.900 ;
        RECT 63.630 318.900 64.630 319.900 ;
        RECT 64.830 318.900 65.830 319.900 ;
        RECT 66.430 318.900 67.430 319.900 ;
        RECT 68.030 318.900 69.030 319.900 ;
        RECT 80.430 320.100 81.430 321.100 ;
        RECT 82.030 320.100 83.030 321.100 ;
        RECT 83.630 320.100 84.630 321.100 ;
        RECT 84.830 320.100 85.830 321.100 ;
        RECT 86.430 320.100 87.430 321.100 ;
        RECT 88.030 320.100 89.030 321.100 ;
        RECT 103.630 323.300 104.630 324.300 ;
        RECT 104.830 323.300 105.830 324.300 ;
        RECT 103.630 321.700 104.630 322.700 ;
        RECT 104.830 321.700 105.830 322.700 ;
        RECT 63.630 317.300 64.630 318.300 ;
        RECT 64.830 317.300 65.830 318.300 ;
        RECT 63.630 315.700 64.630 316.700 ;
        RECT 64.830 315.700 65.830 316.700 ;
        RECT 80.430 318.900 81.430 319.900 ;
        RECT 82.030 318.900 83.030 319.900 ;
        RECT 83.630 318.900 84.630 319.900 ;
        RECT 84.830 318.900 85.830 319.900 ;
        RECT 86.430 318.900 87.430 319.900 ;
        RECT 88.030 318.900 89.030 319.900 ;
        RECT 100.430 320.100 101.430 321.100 ;
        RECT 102.030 320.100 103.030 321.100 ;
        RECT 103.630 320.100 104.630 321.100 ;
        RECT 104.830 320.100 105.830 321.100 ;
        RECT 106.430 320.100 107.430 321.100 ;
        RECT 108.030 320.100 109.030 321.100 ;
        RECT 123.630 323.300 124.630 324.300 ;
        RECT 125.340 323.095 125.700 323.475 ;
        RECT 125.970 323.095 126.330 323.475 ;
        RECT 126.570 323.095 126.930 323.475 ;
        RECT 123.630 321.700 124.630 322.700 ;
        RECT 125.340 322.505 125.700 322.885 ;
        RECT 125.970 322.505 126.330 322.885 ;
        RECT 126.570 322.505 126.930 322.885 ;
        RECT 83.630 317.300 84.630 318.300 ;
        RECT 84.830 317.300 85.830 318.300 ;
        RECT 83.630 315.700 84.630 316.700 ;
        RECT 84.830 315.700 85.830 316.700 ;
        RECT 100.430 318.900 101.430 319.900 ;
        RECT 102.030 318.900 103.030 319.900 ;
        RECT 103.630 318.900 104.630 319.900 ;
        RECT 104.830 318.900 105.830 319.900 ;
        RECT 106.430 318.900 107.430 319.900 ;
        RECT 108.030 318.900 109.030 319.900 ;
        RECT 120.430 320.100 121.430 321.100 ;
        RECT 122.030 320.100 123.030 321.100 ;
        RECT 123.630 320.100 124.630 321.100 ;
        RECT 103.630 317.300 104.630 318.300 ;
        RECT 104.830 317.300 105.830 318.300 ;
        RECT 103.630 315.700 104.630 316.700 ;
        RECT 104.830 315.700 105.830 316.700 ;
        RECT 120.430 318.900 121.430 319.900 ;
        RECT 122.030 318.900 123.030 319.900 ;
        RECT 123.630 318.900 124.630 319.900 ;
        RECT 123.630 317.300 124.630 318.300 ;
        RECT 125.340 317.080 125.700 317.460 ;
        RECT 125.970 317.080 126.330 317.460 ;
        RECT 126.570 317.080 126.930 317.460 ;
        RECT 123.630 315.700 124.630 316.700 ;
        RECT 125.340 316.490 125.700 316.870 ;
        RECT 125.970 316.490 126.330 316.870 ;
        RECT 126.570 316.490 126.930 316.870 ;
        RECT 2.520 306.125 2.880 306.505 ;
        RECT 3.130 306.125 3.490 306.505 ;
        RECT 3.760 306.125 4.120 306.505 ;
        RECT 2.520 305.390 2.880 305.770 ;
        RECT 3.130 305.390 3.490 305.770 ;
        RECT 3.760 305.390 4.120 305.770 ;
        RECT 2.520 304.705 2.880 305.085 ;
        RECT 3.130 304.705 3.490 305.085 ;
        RECT 3.760 304.705 4.120 305.085 ;
        RECT 2.515 303.170 2.875 303.550 ;
        RECT 3.145 303.170 3.505 303.550 ;
        RECT 3.745 303.170 4.105 303.550 ;
        RECT 4.830 303.300 5.830 304.300 ;
        RECT 2.515 302.580 2.875 302.960 ;
        RECT 3.145 302.580 3.505 302.960 ;
        RECT 3.745 302.580 4.105 302.960 ;
        RECT 4.830 301.700 5.830 302.700 ;
        RECT 4.830 300.100 5.830 301.100 ;
        RECT 6.430 300.100 7.430 301.100 ;
        RECT 8.030 300.100 9.030 301.100 ;
        RECT 23.630 303.300 24.630 304.300 ;
        RECT 24.830 303.300 25.830 304.300 ;
        RECT 23.630 301.700 24.630 302.700 ;
        RECT 24.830 301.700 25.830 302.700 ;
        RECT 4.830 298.900 5.830 299.900 ;
        RECT 6.430 298.900 7.430 299.900 ;
        RECT 8.030 298.900 9.030 299.900 ;
        RECT 20.430 300.100 21.430 301.100 ;
        RECT 22.030 300.100 23.030 301.100 ;
        RECT 23.630 300.100 24.630 301.100 ;
        RECT 24.830 300.100 25.830 301.100 ;
        RECT 26.430 300.100 27.430 301.100 ;
        RECT 28.030 300.100 29.030 301.100 ;
        RECT 43.630 303.300 44.630 304.300 ;
        RECT 44.830 303.300 45.830 304.300 ;
        RECT 43.630 301.700 44.630 302.700 ;
        RECT 44.830 301.700 45.830 302.700 ;
        RECT 2.515 297.280 2.875 297.660 ;
        RECT 3.145 297.280 3.505 297.660 ;
        RECT 3.745 297.280 4.105 297.660 ;
        RECT 4.830 297.300 5.830 298.300 ;
        RECT 2.515 296.690 2.875 297.070 ;
        RECT 3.145 296.690 3.505 297.070 ;
        RECT 3.745 296.690 4.105 297.070 ;
        RECT 4.830 295.700 5.830 296.700 ;
        RECT 20.430 298.900 21.430 299.900 ;
        RECT 22.030 298.900 23.030 299.900 ;
        RECT 23.630 298.900 24.630 299.900 ;
        RECT 24.830 298.900 25.830 299.900 ;
        RECT 26.430 298.900 27.430 299.900 ;
        RECT 28.030 298.900 29.030 299.900 ;
        RECT 40.430 300.100 41.430 301.100 ;
        RECT 42.030 300.100 43.030 301.100 ;
        RECT 43.630 300.100 44.630 301.100 ;
        RECT 44.830 300.100 45.830 301.100 ;
        RECT 46.430 300.100 47.430 301.100 ;
        RECT 48.030 300.100 49.030 301.100 ;
        RECT 63.630 303.300 64.630 304.300 ;
        RECT 64.830 303.300 65.830 304.300 ;
        RECT 63.630 301.700 64.630 302.700 ;
        RECT 64.830 301.700 65.830 302.700 ;
        RECT 2.520 294.920 2.880 295.300 ;
        RECT 3.130 294.920 3.490 295.300 ;
        RECT 3.760 294.920 4.120 295.300 ;
        RECT 2.520 294.185 2.880 294.565 ;
        RECT 3.130 294.185 3.490 294.565 ;
        RECT 3.760 294.185 4.120 294.565 ;
        RECT 2.520 293.500 2.880 293.880 ;
        RECT 3.130 293.500 3.490 293.880 ;
        RECT 3.760 293.500 4.120 293.880 ;
        RECT 23.630 297.300 24.630 298.300 ;
        RECT 24.830 297.300 25.830 298.300 ;
        RECT 23.630 295.700 24.630 296.700 ;
        RECT 24.830 295.700 25.830 296.700 ;
        RECT 40.430 298.900 41.430 299.900 ;
        RECT 42.030 298.900 43.030 299.900 ;
        RECT 43.630 298.900 44.630 299.900 ;
        RECT 44.830 298.900 45.830 299.900 ;
        RECT 46.430 298.900 47.430 299.900 ;
        RECT 48.030 298.900 49.030 299.900 ;
        RECT 60.430 300.100 61.430 301.100 ;
        RECT 62.030 300.100 63.030 301.100 ;
        RECT 63.630 300.100 64.630 301.100 ;
        RECT 64.830 300.100 65.830 301.100 ;
        RECT 66.430 300.100 67.430 301.100 ;
        RECT 68.030 300.100 69.030 301.100 ;
        RECT 83.630 303.300 84.630 304.300 ;
        RECT 84.830 303.300 85.830 304.300 ;
        RECT 83.630 301.700 84.630 302.700 ;
        RECT 84.830 301.700 85.830 302.700 ;
        RECT 43.630 297.300 44.630 298.300 ;
        RECT 44.830 297.300 45.830 298.300 ;
        RECT 43.630 295.700 44.630 296.700 ;
        RECT 44.830 295.700 45.830 296.700 ;
        RECT 60.430 298.900 61.430 299.900 ;
        RECT 62.030 298.900 63.030 299.900 ;
        RECT 63.630 298.900 64.630 299.900 ;
        RECT 64.830 298.900 65.830 299.900 ;
        RECT 66.430 298.900 67.430 299.900 ;
        RECT 68.030 298.900 69.030 299.900 ;
        RECT 80.430 300.100 81.430 301.100 ;
        RECT 82.030 300.100 83.030 301.100 ;
        RECT 83.630 300.100 84.630 301.100 ;
        RECT 84.830 300.100 85.830 301.100 ;
        RECT 86.430 300.100 87.430 301.100 ;
        RECT 88.030 300.100 89.030 301.100 ;
        RECT 103.630 303.300 104.630 304.300 ;
        RECT 104.830 303.300 105.830 304.300 ;
        RECT 103.630 301.700 104.630 302.700 ;
        RECT 104.830 301.700 105.830 302.700 ;
        RECT 63.630 297.300 64.630 298.300 ;
        RECT 64.830 297.300 65.830 298.300 ;
        RECT 63.630 295.700 64.630 296.700 ;
        RECT 64.830 295.700 65.830 296.700 ;
        RECT 80.430 298.900 81.430 299.900 ;
        RECT 82.030 298.900 83.030 299.900 ;
        RECT 83.630 298.900 84.630 299.900 ;
        RECT 84.830 298.900 85.830 299.900 ;
        RECT 86.430 298.900 87.430 299.900 ;
        RECT 88.030 298.900 89.030 299.900 ;
        RECT 100.430 300.100 101.430 301.100 ;
        RECT 102.030 300.100 103.030 301.100 ;
        RECT 103.630 300.100 104.630 301.100 ;
        RECT 104.830 300.100 105.830 301.100 ;
        RECT 106.430 300.100 107.430 301.100 ;
        RECT 108.030 300.100 109.030 301.100 ;
        RECT 123.630 303.300 124.630 304.300 ;
        RECT 125.340 303.095 125.700 303.475 ;
        RECT 125.970 303.095 126.330 303.475 ;
        RECT 126.570 303.095 126.930 303.475 ;
        RECT 123.630 301.700 124.630 302.700 ;
        RECT 125.340 302.505 125.700 302.885 ;
        RECT 125.970 302.505 126.330 302.885 ;
        RECT 126.570 302.505 126.930 302.885 ;
        RECT 83.630 297.300 84.630 298.300 ;
        RECT 84.830 297.300 85.830 298.300 ;
        RECT 83.630 295.700 84.630 296.700 ;
        RECT 84.830 295.700 85.830 296.700 ;
        RECT 100.430 298.900 101.430 299.900 ;
        RECT 102.030 298.900 103.030 299.900 ;
        RECT 103.630 298.900 104.630 299.900 ;
        RECT 104.830 298.900 105.830 299.900 ;
        RECT 106.430 298.900 107.430 299.900 ;
        RECT 108.030 298.900 109.030 299.900 ;
        RECT 120.430 300.100 121.430 301.100 ;
        RECT 122.030 300.100 123.030 301.100 ;
        RECT 123.630 300.100 124.630 301.100 ;
        RECT 103.630 297.300 104.630 298.300 ;
        RECT 104.830 297.300 105.830 298.300 ;
        RECT 103.630 295.700 104.630 296.700 ;
        RECT 104.830 295.700 105.830 296.700 ;
        RECT 120.430 298.900 121.430 299.900 ;
        RECT 122.030 298.900 123.030 299.900 ;
        RECT 123.630 298.900 124.630 299.900 ;
        RECT 123.630 297.300 124.630 298.300 ;
        RECT 125.340 297.080 125.700 297.460 ;
        RECT 125.970 297.080 126.330 297.460 ;
        RECT 126.570 297.080 126.930 297.460 ;
        RECT 123.630 295.700 124.630 296.700 ;
        RECT 125.340 296.490 125.700 296.870 ;
        RECT 125.970 296.490 126.330 296.870 ;
        RECT 126.570 296.490 126.930 296.870 ;
        RECT 2.520 286.125 2.880 286.505 ;
        RECT 3.130 286.125 3.490 286.505 ;
        RECT 3.760 286.125 4.120 286.505 ;
        RECT 2.520 285.390 2.880 285.770 ;
        RECT 3.130 285.390 3.490 285.770 ;
        RECT 3.760 285.390 4.120 285.770 ;
        RECT 2.520 284.705 2.880 285.085 ;
        RECT 3.130 284.705 3.490 285.085 ;
        RECT 3.760 284.705 4.120 285.085 ;
        RECT 2.515 283.040 2.875 283.420 ;
        RECT 3.145 283.040 3.505 283.420 ;
        RECT 3.745 283.040 4.105 283.420 ;
        RECT 4.830 283.300 5.830 284.300 ;
        RECT 2.515 282.450 2.875 282.830 ;
        RECT 3.145 282.450 3.505 282.830 ;
        RECT 3.745 282.450 4.105 282.830 ;
        RECT 4.830 281.700 5.830 282.700 ;
        RECT 4.830 280.100 5.830 281.100 ;
        RECT 6.430 280.100 7.430 281.100 ;
        RECT 8.030 280.100 9.030 281.100 ;
        RECT 23.630 283.300 24.630 284.300 ;
        RECT 24.830 283.300 25.830 284.300 ;
        RECT 23.630 281.700 24.630 282.700 ;
        RECT 24.830 281.700 25.830 282.700 ;
        RECT 4.830 278.900 5.830 279.900 ;
        RECT 6.430 278.900 7.430 279.900 ;
        RECT 8.030 278.900 9.030 279.900 ;
        RECT 20.430 280.100 21.430 281.100 ;
        RECT 22.030 280.100 23.030 281.100 ;
        RECT 23.630 280.100 24.630 281.100 ;
        RECT 24.830 280.100 25.830 281.100 ;
        RECT 26.430 280.100 27.430 281.100 ;
        RECT 28.030 280.100 29.030 281.100 ;
        RECT 43.630 283.300 44.630 284.300 ;
        RECT 44.830 283.300 45.830 284.300 ;
        RECT 43.630 281.700 44.630 282.700 ;
        RECT 44.830 281.700 45.830 282.700 ;
        RECT 2.515 277.025 2.875 277.405 ;
        RECT 3.145 277.025 3.505 277.405 ;
        RECT 3.745 277.025 4.105 277.405 ;
        RECT 4.830 277.300 5.830 278.300 ;
        RECT 2.515 276.435 2.875 276.815 ;
        RECT 3.145 276.435 3.505 276.815 ;
        RECT 3.745 276.435 4.105 276.815 ;
        RECT 4.830 275.700 5.830 276.700 ;
        RECT 20.430 278.900 21.430 279.900 ;
        RECT 22.030 278.900 23.030 279.900 ;
        RECT 23.630 278.900 24.630 279.900 ;
        RECT 24.830 278.900 25.830 279.900 ;
        RECT 26.430 278.900 27.430 279.900 ;
        RECT 28.030 278.900 29.030 279.900 ;
        RECT 40.430 280.100 41.430 281.100 ;
        RECT 42.030 280.100 43.030 281.100 ;
        RECT 43.630 280.100 44.630 281.100 ;
        RECT 44.830 280.100 45.830 281.100 ;
        RECT 46.430 280.100 47.430 281.100 ;
        RECT 48.030 280.100 49.030 281.100 ;
        RECT 63.630 283.300 64.630 284.300 ;
        RECT 64.830 283.300 65.830 284.300 ;
        RECT 63.630 281.700 64.630 282.700 ;
        RECT 64.830 281.700 65.830 282.700 ;
        RECT 2.520 274.920 2.880 275.300 ;
        RECT 3.130 274.920 3.490 275.300 ;
        RECT 3.760 274.920 4.120 275.300 ;
        RECT 2.520 274.185 2.880 274.565 ;
        RECT 3.130 274.185 3.490 274.565 ;
        RECT 3.760 274.185 4.120 274.565 ;
        RECT 2.520 273.500 2.880 273.880 ;
        RECT 3.130 273.500 3.490 273.880 ;
        RECT 3.760 273.500 4.120 273.880 ;
        RECT 23.630 277.300 24.630 278.300 ;
        RECT 24.830 277.300 25.830 278.300 ;
        RECT 23.630 275.700 24.630 276.700 ;
        RECT 24.830 275.700 25.830 276.700 ;
        RECT 40.430 278.900 41.430 279.900 ;
        RECT 42.030 278.900 43.030 279.900 ;
        RECT 43.630 278.900 44.630 279.900 ;
        RECT 44.830 278.900 45.830 279.900 ;
        RECT 46.430 278.900 47.430 279.900 ;
        RECT 48.030 278.900 49.030 279.900 ;
        RECT 60.430 280.100 61.430 281.100 ;
        RECT 62.030 280.100 63.030 281.100 ;
        RECT 63.630 280.100 64.630 281.100 ;
        RECT 64.830 280.100 65.830 281.100 ;
        RECT 66.430 280.100 67.430 281.100 ;
        RECT 68.030 280.100 69.030 281.100 ;
        RECT 83.630 283.300 84.630 284.300 ;
        RECT 84.830 283.300 85.830 284.300 ;
        RECT 83.630 281.700 84.630 282.700 ;
        RECT 84.830 281.700 85.830 282.700 ;
        RECT 43.630 277.300 44.630 278.300 ;
        RECT 44.830 277.300 45.830 278.300 ;
        RECT 43.630 275.700 44.630 276.700 ;
        RECT 44.830 275.700 45.830 276.700 ;
        RECT 60.430 278.900 61.430 279.900 ;
        RECT 62.030 278.900 63.030 279.900 ;
        RECT 63.630 278.900 64.630 279.900 ;
        RECT 64.830 278.900 65.830 279.900 ;
        RECT 66.430 278.900 67.430 279.900 ;
        RECT 68.030 278.900 69.030 279.900 ;
        RECT 80.430 280.100 81.430 281.100 ;
        RECT 82.030 280.100 83.030 281.100 ;
        RECT 83.630 280.100 84.630 281.100 ;
        RECT 84.830 280.100 85.830 281.100 ;
        RECT 86.430 280.100 87.430 281.100 ;
        RECT 88.030 280.100 89.030 281.100 ;
        RECT 103.630 283.300 104.630 284.300 ;
        RECT 104.830 283.300 105.830 284.300 ;
        RECT 103.630 281.700 104.630 282.700 ;
        RECT 104.830 281.700 105.830 282.700 ;
        RECT 63.630 277.300 64.630 278.300 ;
        RECT 64.830 277.300 65.830 278.300 ;
        RECT 63.630 275.700 64.630 276.700 ;
        RECT 64.830 275.700 65.830 276.700 ;
        RECT 80.430 278.900 81.430 279.900 ;
        RECT 82.030 278.900 83.030 279.900 ;
        RECT 83.630 278.900 84.630 279.900 ;
        RECT 84.830 278.900 85.830 279.900 ;
        RECT 86.430 278.900 87.430 279.900 ;
        RECT 88.030 278.900 89.030 279.900 ;
        RECT 100.430 280.100 101.430 281.100 ;
        RECT 102.030 280.100 103.030 281.100 ;
        RECT 103.630 280.100 104.630 281.100 ;
        RECT 104.830 280.100 105.830 281.100 ;
        RECT 106.430 280.100 107.430 281.100 ;
        RECT 108.030 280.100 109.030 281.100 ;
        RECT 123.630 283.300 124.630 284.300 ;
        RECT 125.340 283.095 125.700 283.475 ;
        RECT 125.970 283.095 126.330 283.475 ;
        RECT 126.570 283.095 126.930 283.475 ;
        RECT 123.630 281.700 124.630 282.700 ;
        RECT 125.340 282.505 125.700 282.885 ;
        RECT 125.970 282.505 126.330 282.885 ;
        RECT 126.570 282.505 126.930 282.885 ;
        RECT 83.630 277.300 84.630 278.300 ;
        RECT 84.830 277.300 85.830 278.300 ;
        RECT 83.630 275.700 84.630 276.700 ;
        RECT 84.830 275.700 85.830 276.700 ;
        RECT 100.430 278.900 101.430 279.900 ;
        RECT 102.030 278.900 103.030 279.900 ;
        RECT 103.630 278.900 104.630 279.900 ;
        RECT 104.830 278.900 105.830 279.900 ;
        RECT 106.430 278.900 107.430 279.900 ;
        RECT 108.030 278.900 109.030 279.900 ;
        RECT 120.430 280.100 121.430 281.100 ;
        RECT 122.030 280.100 123.030 281.100 ;
        RECT 123.630 280.100 124.630 281.100 ;
        RECT 103.630 277.300 104.630 278.300 ;
        RECT 104.830 277.300 105.830 278.300 ;
        RECT 103.630 275.700 104.630 276.700 ;
        RECT 104.830 275.700 105.830 276.700 ;
        RECT 120.430 278.900 121.430 279.900 ;
        RECT 122.030 278.900 123.030 279.900 ;
        RECT 123.630 278.900 124.630 279.900 ;
        RECT 123.630 277.300 124.630 278.300 ;
        RECT 125.340 277.350 125.700 277.730 ;
        RECT 125.970 277.350 126.330 277.730 ;
        RECT 126.570 277.350 126.930 277.730 ;
        RECT 125.340 276.760 125.700 277.140 ;
        RECT 125.970 276.760 126.330 277.140 ;
        RECT 126.570 276.760 126.930 277.140 ;
        RECT 123.630 275.700 124.630 276.700 ;
        RECT 2.520 266.115 2.880 266.495 ;
        RECT 3.130 266.115 3.490 266.495 ;
        RECT 3.760 266.115 4.120 266.495 ;
        RECT 2.520 265.380 2.880 265.760 ;
        RECT 3.130 265.380 3.490 265.760 ;
        RECT 3.760 265.380 4.120 265.760 ;
        RECT 2.520 264.695 2.880 265.075 ;
        RECT 3.130 264.695 3.490 265.075 ;
        RECT 3.760 264.695 4.120 265.075 ;
        RECT 2.515 263.140 2.875 263.520 ;
        RECT 3.145 263.140 3.505 263.520 ;
        RECT 3.745 263.140 4.105 263.520 ;
        RECT 4.830 263.300 5.830 264.300 ;
        RECT 2.515 262.550 2.875 262.930 ;
        RECT 3.145 262.550 3.505 262.930 ;
        RECT 3.745 262.550 4.105 262.930 ;
        RECT 4.830 261.700 5.830 262.700 ;
        RECT 4.830 260.100 5.830 261.100 ;
        RECT 6.430 260.100 7.430 261.100 ;
        RECT 8.030 260.100 9.030 261.100 ;
        RECT 23.630 263.300 24.630 264.300 ;
        RECT 24.830 263.300 25.830 264.300 ;
        RECT 23.630 261.700 24.630 262.700 ;
        RECT 24.830 261.700 25.830 262.700 ;
        RECT 4.830 258.900 5.830 259.900 ;
        RECT 6.430 258.900 7.430 259.900 ;
        RECT 8.030 258.900 9.030 259.900 ;
        RECT 20.430 260.100 21.430 261.100 ;
        RECT 22.030 260.100 23.030 261.100 ;
        RECT 23.630 260.100 24.630 261.100 ;
        RECT 24.830 260.100 25.830 261.100 ;
        RECT 26.430 260.100 27.430 261.100 ;
        RECT 28.030 260.100 29.030 261.100 ;
        RECT 43.630 263.300 44.630 264.300 ;
        RECT 44.830 263.300 45.830 264.300 ;
        RECT 43.630 261.700 44.630 262.700 ;
        RECT 44.830 261.700 45.830 262.700 ;
        RECT 2.515 257.105 2.875 257.485 ;
        RECT 3.145 257.105 3.505 257.485 ;
        RECT 3.745 257.105 4.105 257.485 ;
        RECT 4.830 257.300 5.830 258.300 ;
        RECT 2.515 256.515 2.875 256.895 ;
        RECT 3.145 256.515 3.505 256.895 ;
        RECT 3.745 256.515 4.105 256.895 ;
        RECT 4.830 255.700 5.830 256.700 ;
        RECT 20.430 258.900 21.430 259.900 ;
        RECT 22.030 258.900 23.030 259.900 ;
        RECT 23.630 258.900 24.630 259.900 ;
        RECT 24.830 258.900 25.830 259.900 ;
        RECT 26.430 258.900 27.430 259.900 ;
        RECT 28.030 258.900 29.030 259.900 ;
        RECT 40.430 260.100 41.430 261.100 ;
        RECT 42.030 260.100 43.030 261.100 ;
        RECT 43.630 260.100 44.630 261.100 ;
        RECT 44.830 260.100 45.830 261.100 ;
        RECT 46.430 260.100 47.430 261.100 ;
        RECT 48.030 260.100 49.030 261.100 ;
        RECT 63.630 263.300 64.630 264.300 ;
        RECT 64.830 263.300 65.830 264.300 ;
        RECT 63.630 261.700 64.630 262.700 ;
        RECT 64.830 261.700 65.830 262.700 ;
        RECT 2.520 254.920 2.880 255.300 ;
        RECT 3.130 254.920 3.490 255.300 ;
        RECT 3.760 254.920 4.120 255.300 ;
        RECT 2.520 254.185 2.880 254.565 ;
        RECT 3.130 254.185 3.490 254.565 ;
        RECT 3.760 254.185 4.120 254.565 ;
        RECT 2.520 253.500 2.880 253.880 ;
        RECT 3.130 253.500 3.490 253.880 ;
        RECT 3.760 253.500 4.120 253.880 ;
        RECT 23.630 257.300 24.630 258.300 ;
        RECT 24.830 257.300 25.830 258.300 ;
        RECT 23.630 255.700 24.630 256.700 ;
        RECT 24.830 255.700 25.830 256.700 ;
        RECT 40.430 258.900 41.430 259.900 ;
        RECT 42.030 258.900 43.030 259.900 ;
        RECT 43.630 258.900 44.630 259.900 ;
        RECT 44.830 258.900 45.830 259.900 ;
        RECT 46.430 258.900 47.430 259.900 ;
        RECT 48.030 258.900 49.030 259.900 ;
        RECT 60.430 260.100 61.430 261.100 ;
        RECT 62.030 260.100 63.030 261.100 ;
        RECT 63.630 260.100 64.630 261.100 ;
        RECT 64.830 260.100 65.830 261.100 ;
        RECT 66.430 260.100 67.430 261.100 ;
        RECT 68.030 260.100 69.030 261.100 ;
        RECT 83.630 263.300 84.630 264.300 ;
        RECT 84.830 263.300 85.830 264.300 ;
        RECT 83.630 261.700 84.630 262.700 ;
        RECT 84.830 261.700 85.830 262.700 ;
        RECT 43.630 257.300 44.630 258.300 ;
        RECT 44.830 257.300 45.830 258.300 ;
        RECT 43.630 255.700 44.630 256.700 ;
        RECT 44.830 255.700 45.830 256.700 ;
        RECT 60.430 258.900 61.430 259.900 ;
        RECT 62.030 258.900 63.030 259.900 ;
        RECT 63.630 258.900 64.630 259.900 ;
        RECT 64.830 258.900 65.830 259.900 ;
        RECT 66.430 258.900 67.430 259.900 ;
        RECT 68.030 258.900 69.030 259.900 ;
        RECT 80.430 260.100 81.430 261.100 ;
        RECT 82.030 260.100 83.030 261.100 ;
        RECT 83.630 260.100 84.630 261.100 ;
        RECT 84.830 260.100 85.830 261.100 ;
        RECT 86.430 260.100 87.430 261.100 ;
        RECT 88.030 260.100 89.030 261.100 ;
        RECT 103.630 263.300 104.630 264.300 ;
        RECT 104.830 263.300 105.830 264.300 ;
        RECT 103.630 261.700 104.630 262.700 ;
        RECT 104.830 261.700 105.830 262.700 ;
        RECT 63.630 257.300 64.630 258.300 ;
        RECT 64.830 257.300 65.830 258.300 ;
        RECT 63.630 255.700 64.630 256.700 ;
        RECT 64.830 255.700 65.830 256.700 ;
        RECT 80.430 258.900 81.430 259.900 ;
        RECT 82.030 258.900 83.030 259.900 ;
        RECT 83.630 258.900 84.630 259.900 ;
        RECT 84.830 258.900 85.830 259.900 ;
        RECT 86.430 258.900 87.430 259.900 ;
        RECT 88.030 258.900 89.030 259.900 ;
        RECT 100.430 260.100 101.430 261.100 ;
        RECT 102.030 260.100 103.030 261.100 ;
        RECT 103.630 260.100 104.630 261.100 ;
        RECT 104.830 260.100 105.830 261.100 ;
        RECT 106.430 260.100 107.430 261.100 ;
        RECT 108.030 260.100 109.030 261.100 ;
        RECT 123.630 263.300 124.630 264.300 ;
        RECT 125.340 262.770 125.700 263.150 ;
        RECT 125.970 262.770 126.330 263.150 ;
        RECT 126.570 262.770 126.930 263.150 ;
        RECT 123.630 261.700 124.630 262.700 ;
        RECT 125.340 262.180 125.700 262.560 ;
        RECT 125.970 262.180 126.330 262.560 ;
        RECT 126.570 262.180 126.930 262.560 ;
        RECT 83.630 257.300 84.630 258.300 ;
        RECT 84.830 257.300 85.830 258.300 ;
        RECT 83.630 255.700 84.630 256.700 ;
        RECT 84.830 255.700 85.830 256.700 ;
        RECT 100.430 258.900 101.430 259.900 ;
        RECT 102.030 258.900 103.030 259.900 ;
        RECT 103.630 258.900 104.630 259.900 ;
        RECT 104.830 258.900 105.830 259.900 ;
        RECT 106.430 258.900 107.430 259.900 ;
        RECT 108.030 258.900 109.030 259.900 ;
        RECT 120.430 260.100 121.430 261.100 ;
        RECT 122.030 260.100 123.030 261.100 ;
        RECT 123.630 260.100 124.630 261.100 ;
        RECT 103.630 257.300 104.630 258.300 ;
        RECT 104.830 257.300 105.830 258.300 ;
        RECT 103.630 255.700 104.630 256.700 ;
        RECT 104.830 255.700 105.830 256.700 ;
        RECT 120.430 258.900 121.430 259.900 ;
        RECT 122.030 258.900 123.030 259.900 ;
        RECT 123.630 258.900 124.630 259.900 ;
        RECT 123.630 257.300 124.630 258.300 ;
        RECT 125.340 256.855 125.700 257.235 ;
        RECT 125.970 256.855 126.330 257.235 ;
        RECT 126.570 256.855 126.930 257.235 ;
        RECT 123.630 255.700 124.630 256.700 ;
        RECT 125.340 256.265 125.700 256.645 ;
        RECT 125.970 256.265 126.330 256.645 ;
        RECT 126.570 256.265 126.930 256.645 ;
        RECT 2.520 246.125 2.880 246.505 ;
        RECT 3.130 246.125 3.490 246.505 ;
        RECT 3.760 246.125 4.120 246.505 ;
        RECT 2.520 245.390 2.880 245.770 ;
        RECT 3.130 245.390 3.490 245.770 ;
        RECT 3.760 245.390 4.120 245.770 ;
        RECT 2.520 244.705 2.880 245.085 ;
        RECT 3.130 244.705 3.490 245.085 ;
        RECT 3.760 244.705 4.120 245.085 ;
        RECT 2.515 243.275 2.875 243.655 ;
        RECT 3.145 243.275 3.505 243.655 ;
        RECT 3.745 243.275 4.105 243.655 ;
        RECT 4.830 243.300 5.830 244.300 ;
        RECT 2.515 242.685 2.875 243.065 ;
        RECT 3.145 242.685 3.505 243.065 ;
        RECT 3.745 242.685 4.105 243.065 ;
        RECT 4.830 241.700 5.830 242.700 ;
        RECT 4.830 240.100 5.830 241.100 ;
        RECT 6.430 240.100 7.430 241.100 ;
        RECT 8.030 240.100 9.030 241.100 ;
        RECT 23.630 243.300 24.630 244.300 ;
        RECT 24.830 243.300 25.830 244.300 ;
        RECT 23.630 241.700 24.630 242.700 ;
        RECT 24.830 241.700 25.830 242.700 ;
        RECT 4.830 238.900 5.830 239.900 ;
        RECT 6.430 238.900 7.430 239.900 ;
        RECT 8.030 238.900 9.030 239.900 ;
        RECT 20.430 240.100 21.430 241.100 ;
        RECT 22.030 240.100 23.030 241.100 ;
        RECT 23.630 240.100 24.630 241.100 ;
        RECT 24.830 240.100 25.830 241.100 ;
        RECT 26.430 240.100 27.430 241.100 ;
        RECT 28.030 240.100 29.030 241.100 ;
        RECT 43.630 243.300 44.630 244.300 ;
        RECT 44.830 243.300 45.830 244.300 ;
        RECT 43.630 241.700 44.630 242.700 ;
        RECT 44.830 241.700 45.830 242.700 ;
        RECT 2.515 237.340 2.875 237.720 ;
        RECT 3.145 237.340 3.505 237.720 ;
        RECT 3.745 237.340 4.105 237.720 ;
        RECT 4.830 237.300 5.830 238.300 ;
        RECT 2.515 236.750 2.875 237.130 ;
        RECT 3.145 236.750 3.505 237.130 ;
        RECT 3.745 236.750 4.105 237.130 ;
        RECT 4.830 235.700 5.830 236.700 ;
        RECT 20.430 238.900 21.430 239.900 ;
        RECT 22.030 238.900 23.030 239.900 ;
        RECT 23.630 238.900 24.630 239.900 ;
        RECT 24.830 238.900 25.830 239.900 ;
        RECT 26.430 238.900 27.430 239.900 ;
        RECT 28.030 238.900 29.030 239.900 ;
        RECT 40.430 240.100 41.430 241.100 ;
        RECT 42.030 240.100 43.030 241.100 ;
        RECT 43.630 240.100 44.630 241.100 ;
        RECT 44.830 240.100 45.830 241.100 ;
        RECT 46.430 240.100 47.430 241.100 ;
        RECT 48.030 240.100 49.030 241.100 ;
        RECT 63.630 243.300 64.630 244.300 ;
        RECT 64.830 243.300 65.830 244.300 ;
        RECT 63.630 241.700 64.630 242.700 ;
        RECT 64.830 241.700 65.830 242.700 ;
        RECT 2.520 234.920 2.880 235.300 ;
        RECT 3.130 234.920 3.490 235.300 ;
        RECT 3.760 234.920 4.120 235.300 ;
        RECT 2.520 234.185 2.880 234.565 ;
        RECT 3.130 234.185 3.490 234.565 ;
        RECT 3.760 234.185 4.120 234.565 ;
        RECT 2.520 233.500 2.880 233.880 ;
        RECT 3.130 233.500 3.490 233.880 ;
        RECT 3.760 233.500 4.120 233.880 ;
        RECT 23.630 237.300 24.630 238.300 ;
        RECT 24.830 237.300 25.830 238.300 ;
        RECT 23.630 235.700 24.630 236.700 ;
        RECT 24.830 235.700 25.830 236.700 ;
        RECT 40.430 238.900 41.430 239.900 ;
        RECT 42.030 238.900 43.030 239.900 ;
        RECT 43.630 238.900 44.630 239.900 ;
        RECT 44.830 238.900 45.830 239.900 ;
        RECT 46.430 238.900 47.430 239.900 ;
        RECT 48.030 238.900 49.030 239.900 ;
        RECT 60.430 240.100 61.430 241.100 ;
        RECT 62.030 240.100 63.030 241.100 ;
        RECT 63.630 240.100 64.630 241.100 ;
        RECT 64.830 240.100 65.830 241.100 ;
        RECT 66.430 240.100 67.430 241.100 ;
        RECT 68.030 240.100 69.030 241.100 ;
        RECT 83.630 243.300 84.630 244.300 ;
        RECT 84.830 243.300 85.830 244.300 ;
        RECT 83.630 241.700 84.630 242.700 ;
        RECT 84.830 241.700 85.830 242.700 ;
        RECT 43.630 237.300 44.630 238.300 ;
        RECT 44.830 237.300 45.830 238.300 ;
        RECT 43.630 235.700 44.630 236.700 ;
        RECT 44.830 235.700 45.830 236.700 ;
        RECT 60.430 238.900 61.430 239.900 ;
        RECT 62.030 238.900 63.030 239.900 ;
        RECT 63.630 238.900 64.630 239.900 ;
        RECT 64.830 238.900 65.830 239.900 ;
        RECT 66.430 238.900 67.430 239.900 ;
        RECT 68.030 238.900 69.030 239.900 ;
        RECT 80.430 240.100 81.430 241.100 ;
        RECT 82.030 240.100 83.030 241.100 ;
        RECT 83.630 240.100 84.630 241.100 ;
        RECT 84.830 240.100 85.830 241.100 ;
        RECT 86.430 240.100 87.430 241.100 ;
        RECT 88.030 240.100 89.030 241.100 ;
        RECT 103.630 243.300 104.630 244.300 ;
        RECT 104.830 243.300 105.830 244.300 ;
        RECT 103.630 241.700 104.630 242.700 ;
        RECT 104.830 241.700 105.830 242.700 ;
        RECT 63.630 237.300 64.630 238.300 ;
        RECT 64.830 237.300 65.830 238.300 ;
        RECT 63.630 235.700 64.630 236.700 ;
        RECT 64.830 235.700 65.830 236.700 ;
        RECT 80.430 238.900 81.430 239.900 ;
        RECT 82.030 238.900 83.030 239.900 ;
        RECT 83.630 238.900 84.630 239.900 ;
        RECT 84.830 238.900 85.830 239.900 ;
        RECT 86.430 238.900 87.430 239.900 ;
        RECT 88.030 238.900 89.030 239.900 ;
        RECT 100.430 240.100 101.430 241.100 ;
        RECT 102.030 240.100 103.030 241.100 ;
        RECT 103.630 240.100 104.630 241.100 ;
        RECT 104.830 240.100 105.830 241.100 ;
        RECT 106.430 240.100 107.430 241.100 ;
        RECT 108.030 240.100 109.030 241.100 ;
        RECT 123.630 243.300 124.630 244.300 ;
        RECT 123.630 241.700 124.630 242.700 ;
        RECT 125.340 242.495 125.700 242.875 ;
        RECT 125.970 242.495 126.330 242.875 ;
        RECT 126.570 242.495 126.930 242.875 ;
        RECT 125.340 241.905 125.700 242.285 ;
        RECT 125.970 241.905 126.330 242.285 ;
        RECT 126.570 241.905 126.930 242.285 ;
        RECT 83.630 237.300 84.630 238.300 ;
        RECT 84.830 237.300 85.830 238.300 ;
        RECT 83.630 235.700 84.630 236.700 ;
        RECT 84.830 235.700 85.830 236.700 ;
        RECT 100.430 238.900 101.430 239.900 ;
        RECT 102.030 238.900 103.030 239.900 ;
        RECT 103.630 238.900 104.630 239.900 ;
        RECT 104.830 238.900 105.830 239.900 ;
        RECT 106.430 238.900 107.430 239.900 ;
        RECT 108.030 238.900 109.030 239.900 ;
        RECT 120.430 240.100 121.430 241.100 ;
        RECT 122.030 240.100 123.030 241.100 ;
        RECT 123.630 240.100 124.630 241.100 ;
        RECT 103.630 237.300 104.630 238.300 ;
        RECT 104.830 237.300 105.830 238.300 ;
        RECT 103.630 235.700 104.630 236.700 ;
        RECT 104.830 235.700 105.830 236.700 ;
        RECT 120.430 238.900 121.430 239.900 ;
        RECT 122.030 238.900 123.030 239.900 ;
        RECT 123.630 238.900 124.630 239.900 ;
        RECT 123.630 237.300 124.630 238.300 ;
        RECT 125.340 236.820 125.700 237.200 ;
        RECT 125.970 236.820 126.330 237.200 ;
        RECT 126.570 236.820 126.930 237.200 ;
        RECT 123.630 235.700 124.630 236.700 ;
        RECT 125.340 236.230 125.700 236.610 ;
        RECT 125.970 236.230 126.330 236.610 ;
        RECT 126.570 236.230 126.930 236.610 ;
        RECT 2.520 226.125 2.880 226.505 ;
        RECT 3.130 226.125 3.490 226.505 ;
        RECT 3.760 226.125 4.120 226.505 ;
        RECT 2.520 225.390 2.880 225.770 ;
        RECT 3.130 225.390 3.490 225.770 ;
        RECT 3.760 225.390 4.120 225.770 ;
        RECT 2.520 224.705 2.880 225.085 ;
        RECT 3.130 224.705 3.490 225.085 ;
        RECT 3.760 224.705 4.120 225.085 ;
        RECT 2.515 223.230 2.875 223.610 ;
        RECT 3.145 223.230 3.505 223.610 ;
        RECT 3.745 223.230 4.105 223.610 ;
        RECT 4.830 223.300 5.830 224.300 ;
        RECT 2.515 222.640 2.875 223.020 ;
        RECT 3.145 222.640 3.505 223.020 ;
        RECT 3.745 222.640 4.105 223.020 ;
        RECT 4.830 221.700 5.830 222.700 ;
        RECT 4.830 220.100 5.830 221.100 ;
        RECT 6.430 220.100 7.430 221.100 ;
        RECT 8.030 220.100 9.030 221.100 ;
        RECT 23.630 223.300 24.630 224.300 ;
        RECT 24.830 223.300 25.830 224.300 ;
        RECT 23.630 221.700 24.630 222.700 ;
        RECT 24.830 221.700 25.830 222.700 ;
        RECT 4.830 218.900 5.830 219.900 ;
        RECT 6.430 218.900 7.430 219.900 ;
        RECT 8.030 218.900 9.030 219.900 ;
        RECT 20.430 220.100 21.430 221.100 ;
        RECT 22.030 220.100 23.030 221.100 ;
        RECT 23.630 220.100 24.630 221.100 ;
        RECT 24.830 220.100 25.830 221.100 ;
        RECT 26.430 220.100 27.430 221.100 ;
        RECT 28.030 220.100 29.030 221.100 ;
        RECT 43.630 223.300 44.630 224.300 ;
        RECT 44.830 223.300 45.830 224.300 ;
        RECT 43.630 221.700 44.630 222.700 ;
        RECT 44.830 221.700 45.830 222.700 ;
        RECT 2.515 217.465 2.875 217.845 ;
        RECT 3.145 217.465 3.505 217.845 ;
        RECT 3.745 217.465 4.105 217.845 ;
        RECT 4.830 217.300 5.830 218.300 ;
        RECT 2.515 216.875 2.875 217.255 ;
        RECT 3.145 216.875 3.505 217.255 ;
        RECT 3.745 216.875 4.105 217.255 ;
        RECT 4.830 215.700 5.830 216.700 ;
        RECT 20.430 218.900 21.430 219.900 ;
        RECT 22.030 218.900 23.030 219.900 ;
        RECT 23.630 218.900 24.630 219.900 ;
        RECT 24.830 218.900 25.830 219.900 ;
        RECT 26.430 218.900 27.430 219.900 ;
        RECT 28.030 218.900 29.030 219.900 ;
        RECT 40.430 220.100 41.430 221.100 ;
        RECT 42.030 220.100 43.030 221.100 ;
        RECT 43.630 220.100 44.630 221.100 ;
        RECT 44.830 220.100 45.830 221.100 ;
        RECT 46.430 220.100 47.430 221.100 ;
        RECT 48.030 220.100 49.030 221.100 ;
        RECT 63.630 223.300 64.630 224.300 ;
        RECT 64.830 223.300 65.830 224.300 ;
        RECT 63.630 221.700 64.630 222.700 ;
        RECT 64.830 221.700 65.830 222.700 ;
        RECT 2.520 214.920 2.880 215.300 ;
        RECT 3.130 214.920 3.490 215.300 ;
        RECT 3.760 214.920 4.120 215.300 ;
        RECT 2.520 214.185 2.880 214.565 ;
        RECT 3.130 214.185 3.490 214.565 ;
        RECT 3.760 214.185 4.120 214.565 ;
        RECT 2.520 213.500 2.880 213.880 ;
        RECT 3.130 213.500 3.490 213.880 ;
        RECT 3.760 213.500 4.120 213.880 ;
        RECT 23.630 217.300 24.630 218.300 ;
        RECT 24.830 217.300 25.830 218.300 ;
        RECT 23.630 215.700 24.630 216.700 ;
        RECT 24.830 215.700 25.830 216.700 ;
        RECT 40.430 218.900 41.430 219.900 ;
        RECT 42.030 218.900 43.030 219.900 ;
        RECT 43.630 218.900 44.630 219.900 ;
        RECT 44.830 218.900 45.830 219.900 ;
        RECT 46.430 218.900 47.430 219.900 ;
        RECT 48.030 218.900 49.030 219.900 ;
        RECT 60.430 220.100 61.430 221.100 ;
        RECT 62.030 220.100 63.030 221.100 ;
        RECT 63.630 220.100 64.630 221.100 ;
        RECT 64.830 220.100 65.830 221.100 ;
        RECT 66.430 220.100 67.430 221.100 ;
        RECT 68.030 220.100 69.030 221.100 ;
        RECT 83.630 223.300 84.630 224.300 ;
        RECT 84.830 223.300 85.830 224.300 ;
        RECT 83.630 221.700 84.630 222.700 ;
        RECT 84.830 221.700 85.830 222.700 ;
        RECT 43.630 217.300 44.630 218.300 ;
        RECT 44.830 217.300 45.830 218.300 ;
        RECT 43.630 215.700 44.630 216.700 ;
        RECT 44.830 215.700 45.830 216.700 ;
        RECT 60.430 218.900 61.430 219.900 ;
        RECT 62.030 218.900 63.030 219.900 ;
        RECT 63.630 218.900 64.630 219.900 ;
        RECT 64.830 218.900 65.830 219.900 ;
        RECT 66.430 218.900 67.430 219.900 ;
        RECT 68.030 218.900 69.030 219.900 ;
        RECT 80.430 220.100 81.430 221.100 ;
        RECT 82.030 220.100 83.030 221.100 ;
        RECT 83.630 220.100 84.630 221.100 ;
        RECT 84.830 220.100 85.830 221.100 ;
        RECT 86.430 220.100 87.430 221.100 ;
        RECT 88.030 220.100 89.030 221.100 ;
        RECT 103.630 223.300 104.630 224.300 ;
        RECT 104.830 223.300 105.830 224.300 ;
        RECT 103.630 221.700 104.630 222.700 ;
        RECT 104.830 221.700 105.830 222.700 ;
        RECT 63.630 217.300 64.630 218.300 ;
        RECT 64.830 217.300 65.830 218.300 ;
        RECT 63.630 215.700 64.630 216.700 ;
        RECT 64.830 215.700 65.830 216.700 ;
        RECT 80.430 218.900 81.430 219.900 ;
        RECT 82.030 218.900 83.030 219.900 ;
        RECT 83.630 218.900 84.630 219.900 ;
        RECT 84.830 218.900 85.830 219.900 ;
        RECT 86.430 218.900 87.430 219.900 ;
        RECT 88.030 218.900 89.030 219.900 ;
        RECT 100.430 220.100 101.430 221.100 ;
        RECT 102.030 220.100 103.030 221.100 ;
        RECT 103.630 220.100 104.630 221.100 ;
        RECT 104.830 220.100 105.830 221.100 ;
        RECT 106.430 220.100 107.430 221.100 ;
        RECT 108.030 220.100 109.030 221.100 ;
        RECT 123.630 223.300 124.630 224.300 ;
        RECT 125.340 223.025 125.700 223.405 ;
        RECT 125.970 223.025 126.330 223.405 ;
        RECT 126.570 223.025 126.930 223.405 ;
        RECT 123.630 221.700 124.630 222.700 ;
        RECT 125.340 222.435 125.700 222.815 ;
        RECT 125.970 222.435 126.330 222.815 ;
        RECT 126.570 222.435 126.930 222.815 ;
        RECT 83.630 217.300 84.630 218.300 ;
        RECT 84.830 217.300 85.830 218.300 ;
        RECT 83.630 215.700 84.630 216.700 ;
        RECT 84.830 215.700 85.830 216.700 ;
        RECT 100.430 218.900 101.430 219.900 ;
        RECT 102.030 218.900 103.030 219.900 ;
        RECT 103.630 218.900 104.630 219.900 ;
        RECT 104.830 218.900 105.830 219.900 ;
        RECT 106.430 218.900 107.430 219.900 ;
        RECT 108.030 218.900 109.030 219.900 ;
        RECT 120.430 220.100 121.430 221.100 ;
        RECT 122.030 220.100 123.030 221.100 ;
        RECT 123.630 220.100 124.630 221.100 ;
        RECT 103.630 217.300 104.630 218.300 ;
        RECT 104.830 217.300 105.830 218.300 ;
        RECT 103.630 215.700 104.630 216.700 ;
        RECT 104.830 215.700 105.830 216.700 ;
        RECT 120.430 218.900 121.430 219.900 ;
        RECT 122.030 218.900 123.030 219.900 ;
        RECT 123.630 218.900 124.630 219.900 ;
        RECT 123.630 217.300 124.630 218.300 ;
        RECT 125.340 217.260 125.700 217.640 ;
        RECT 125.970 217.260 126.330 217.640 ;
        RECT 126.570 217.260 126.930 217.640 ;
        RECT 123.630 215.700 124.630 216.700 ;
        RECT 125.340 216.670 125.700 217.050 ;
        RECT 125.970 216.670 126.330 217.050 ;
        RECT 126.570 216.670 126.930 217.050 ;
        RECT 2.520 206.120 2.880 206.500 ;
        RECT 3.130 206.120 3.490 206.500 ;
        RECT 3.760 206.120 4.120 206.500 ;
        RECT 2.520 205.385 2.880 205.765 ;
        RECT 3.130 205.385 3.490 205.765 ;
        RECT 3.760 205.385 4.120 205.765 ;
        RECT 2.520 204.700 2.880 205.080 ;
        RECT 3.130 204.700 3.490 205.080 ;
        RECT 3.760 204.700 4.120 205.080 ;
        RECT 4.830 203.300 5.830 204.300 ;
        RECT 2.515 202.165 2.875 202.545 ;
        RECT 3.145 202.165 3.505 202.545 ;
        RECT 3.745 202.165 4.105 202.545 ;
        RECT 2.515 201.575 2.875 201.955 ;
        RECT 3.145 201.575 3.505 201.955 ;
        RECT 3.745 201.575 4.105 201.955 ;
        RECT 4.830 201.700 5.830 202.700 ;
        RECT 4.830 200.100 5.830 201.100 ;
        RECT 6.430 200.100 7.430 201.100 ;
        RECT 8.030 200.100 9.030 201.100 ;
        RECT 23.630 203.300 24.630 204.300 ;
        RECT 24.830 203.300 25.830 204.300 ;
        RECT 23.630 201.700 24.630 202.700 ;
        RECT 24.830 201.700 25.830 202.700 ;
        RECT 20.430 200.100 21.430 201.100 ;
        RECT 22.030 200.100 23.030 201.100 ;
        RECT 23.630 200.100 24.630 201.100 ;
        RECT 24.830 200.100 25.830 201.100 ;
        RECT 26.430 200.100 27.430 201.100 ;
        RECT 28.030 200.100 29.030 201.100 ;
        RECT 43.630 203.300 44.630 204.300 ;
        RECT 44.830 203.300 45.830 204.300 ;
        RECT 43.630 201.700 44.630 202.700 ;
        RECT 44.830 201.700 45.830 202.700 ;
        RECT 40.430 200.100 41.430 201.100 ;
        RECT 42.030 200.100 43.030 201.100 ;
        RECT 43.630 200.100 44.630 201.100 ;
        RECT 44.830 200.100 45.830 201.100 ;
        RECT 46.430 200.100 47.430 201.100 ;
        RECT 48.030 200.100 49.030 201.100 ;
        RECT 63.630 203.300 64.630 204.300 ;
        RECT 64.830 203.300 65.830 204.300 ;
        RECT 63.630 201.700 64.630 202.700 ;
        RECT 64.830 201.700 65.830 202.700 ;
        RECT 60.430 200.100 61.430 201.100 ;
        RECT 62.030 200.100 63.030 201.100 ;
        RECT 63.630 200.100 64.630 201.100 ;
        RECT 64.830 200.100 65.830 201.100 ;
        RECT 66.430 200.100 67.430 201.100 ;
        RECT 68.030 200.100 69.030 201.100 ;
        RECT 83.630 203.300 84.630 204.300 ;
        RECT 84.830 203.300 85.830 204.300 ;
        RECT 83.630 201.700 84.630 202.700 ;
        RECT 84.830 201.700 85.830 202.700 ;
        RECT 80.430 200.100 81.430 201.100 ;
        RECT 82.030 200.100 83.030 201.100 ;
        RECT 83.630 200.100 84.630 201.100 ;
        RECT 84.830 200.100 85.830 201.100 ;
        RECT 86.430 200.100 87.430 201.100 ;
        RECT 88.030 200.100 89.030 201.100 ;
        RECT 103.630 203.300 104.630 204.300 ;
        RECT 104.830 203.300 105.830 204.300 ;
        RECT 103.630 201.700 104.630 202.700 ;
        RECT 104.830 201.700 105.830 202.700 ;
        RECT 100.430 200.100 101.430 201.100 ;
        RECT 102.030 200.100 103.030 201.100 ;
        RECT 103.630 200.100 104.630 201.100 ;
        RECT 104.830 200.100 105.830 201.100 ;
        RECT 106.430 200.100 107.430 201.100 ;
        RECT 108.030 200.100 109.030 201.100 ;
        RECT 123.630 203.300 124.630 204.300 ;
        RECT 123.630 201.700 124.630 202.700 ;
        RECT 125.340 201.680 125.700 202.060 ;
        RECT 125.970 201.680 126.330 202.060 ;
        RECT 126.570 201.680 126.930 202.060 ;
        RECT 120.430 200.100 121.430 201.100 ;
        RECT 122.030 200.100 123.030 201.100 ;
        RECT 123.630 200.100 124.630 201.100 ;
        RECT 125.340 201.090 125.700 201.470 ;
        RECT 125.970 201.090 126.330 201.470 ;
        RECT 126.570 201.090 126.930 201.470 ;
        RECT 2.395 175.260 2.805 175.650 ;
        RECT 2.965 175.260 3.375 175.650 ;
        RECT 3.535 175.260 3.945 175.650 ;
        RECT 42.735 175.560 43.735 176.560 ;
        RECT 44.335 175.560 45.335 176.560 ;
        RECT 45.935 175.560 46.935 176.560 ;
        RECT 42.735 173.960 43.735 174.960 ;
        RECT 42.735 172.360 43.735 173.360 ;
        RECT 58.335 175.560 59.335 176.560 ;
        RECT 59.935 175.560 60.935 176.560 ;
        RECT 61.535 175.560 62.535 176.560 ;
        RECT 62.735 175.560 63.735 176.560 ;
        RECT 64.335 175.560 65.335 176.560 ;
        RECT 65.935 175.560 66.935 176.560 ;
        RECT 2.395 169.820 2.805 170.210 ;
        RECT 2.965 169.820 3.375 170.210 ;
        RECT 3.535 169.820 3.945 170.210 ;
        RECT 61.535 173.960 62.535 174.960 ;
        RECT 62.735 173.960 63.735 174.960 ;
        RECT 61.535 172.360 62.535 173.360 ;
        RECT 62.735 172.360 63.735 173.360 ;
        RECT 78.335 175.560 79.335 176.560 ;
        RECT 79.935 175.560 80.935 176.560 ;
        RECT 81.535 175.560 82.535 176.560 ;
        RECT 82.735 175.560 83.735 176.560 ;
        RECT 84.335 175.560 85.335 176.560 ;
        RECT 85.935 175.560 86.935 176.560 ;
        RECT 81.535 173.960 82.535 174.960 ;
        RECT 82.735 173.960 83.735 174.960 ;
        RECT 81.535 172.360 82.535 173.360 ;
        RECT 82.735 172.360 83.735 173.360 ;
        RECT 98.335 175.560 99.335 176.560 ;
        RECT 99.935 175.560 100.935 176.560 ;
        RECT 101.535 175.560 102.535 176.560 ;
        RECT 102.735 175.560 103.735 176.560 ;
        RECT 104.335 175.560 105.335 176.560 ;
        RECT 105.935 175.560 106.935 176.560 ;
        RECT 101.535 173.960 102.535 174.960 ;
        RECT 102.735 173.960 103.735 174.960 ;
        RECT 101.535 172.360 102.535 173.360 ;
        RECT 102.735 172.360 103.735 173.360 ;
        RECT 118.335 175.560 119.335 176.560 ;
        RECT 119.935 175.560 120.935 176.560 ;
        RECT 121.535 175.560 122.535 176.560 ;
        RECT 121.535 173.960 122.535 174.960 ;
        RECT 125.305 174.460 125.705 174.860 ;
        RECT 125.930 174.460 126.330 174.860 ;
        RECT 126.555 174.460 126.955 174.860 ;
        RECT 125.300 173.860 125.700 174.260 ;
        RECT 125.925 173.860 126.325 174.260 ;
        RECT 126.550 173.860 126.950 174.260 ;
        RECT 121.535 172.360 122.535 173.360 ;
        RECT 125.345 171.580 125.705 171.960 ;
        RECT 125.955 171.580 126.315 171.960 ;
        RECT 126.585 171.580 126.945 171.960 ;
        RECT 125.345 170.845 125.705 171.225 ;
        RECT 125.955 170.845 126.315 171.225 ;
        RECT 126.585 170.845 126.945 171.225 ;
        RECT 125.345 170.160 125.705 170.540 ;
        RECT 125.955 170.160 126.315 170.540 ;
        RECT 126.585 170.160 126.945 170.540 ;
        RECT 2.395 164.380 2.805 164.770 ;
        RECT 2.965 164.380 3.375 164.770 ;
        RECT 3.535 164.380 3.945 164.770 ;
        RECT 42.735 159.960 43.735 160.960 ;
        RECT 42.735 158.360 43.735 159.360 ;
        RECT 42.735 156.760 43.735 157.760 ;
        RECT 44.335 156.760 45.335 157.760 ;
        RECT 45.935 156.760 46.935 157.760 ;
        RECT 61.535 159.960 62.535 160.960 ;
        RECT 62.735 159.960 63.735 160.960 ;
        RECT 61.535 158.360 62.535 159.360 ;
        RECT 62.735 158.360 63.735 159.360 ;
        RECT 58.335 156.760 59.335 157.760 ;
        RECT 59.935 156.760 60.935 157.760 ;
        RECT 61.535 156.760 62.535 157.760 ;
        RECT 62.735 156.760 63.735 157.760 ;
        RECT 64.335 156.760 65.335 157.760 ;
        RECT 65.935 156.760 66.935 157.760 ;
        RECT 81.535 159.960 82.535 160.960 ;
        RECT 82.735 159.960 83.735 160.960 ;
        RECT 81.535 158.360 82.535 159.360 ;
        RECT 82.735 158.360 83.735 159.360 ;
        RECT 78.335 156.760 79.335 157.760 ;
        RECT 79.935 156.760 80.935 157.760 ;
        RECT 81.535 156.760 82.535 157.760 ;
        RECT 82.735 156.760 83.735 157.760 ;
        RECT 84.335 156.760 85.335 157.760 ;
        RECT 85.935 156.760 86.935 157.760 ;
        RECT 101.535 159.960 102.535 160.960 ;
        RECT 102.735 159.960 103.735 160.960 ;
        RECT 101.535 158.360 102.535 159.360 ;
        RECT 102.735 158.360 103.735 159.360 ;
        RECT 125.345 162.780 125.705 163.160 ;
        RECT 125.955 162.780 126.315 163.160 ;
        RECT 126.585 162.780 126.945 163.160 ;
        RECT 125.345 162.045 125.705 162.425 ;
        RECT 125.955 162.045 126.315 162.425 ;
        RECT 126.585 162.045 126.945 162.425 ;
        RECT 125.345 161.360 125.705 161.740 ;
        RECT 125.955 161.360 126.315 161.740 ;
        RECT 126.585 161.360 126.945 161.740 ;
        RECT 98.335 156.760 99.335 157.760 ;
        RECT 99.935 156.760 100.935 157.760 ;
        RECT 101.535 156.760 102.535 157.760 ;
        RECT 102.735 156.760 103.735 157.760 ;
        RECT 104.335 156.760 105.335 157.760 ;
        RECT 105.935 156.760 106.935 157.760 ;
        RECT 121.535 159.960 122.535 160.960 ;
        RECT 121.535 158.360 122.535 159.360 ;
        RECT 125.300 159.185 125.700 159.585 ;
        RECT 125.925 159.185 126.325 159.585 ;
        RECT 126.550 159.185 126.950 159.585 ;
        RECT 125.295 158.585 125.695 158.985 ;
        RECT 125.920 158.585 126.320 158.985 ;
        RECT 126.545 158.585 126.945 158.985 ;
        RECT 118.335 156.760 119.335 157.760 ;
        RECT 119.935 156.760 120.935 157.760 ;
        RECT 121.535 156.760 122.535 157.760 ;
        RECT 2.515 141.130 2.875 141.510 ;
        RECT 3.145 141.130 3.505 141.510 ;
        RECT 3.745 141.130 4.105 141.510 ;
        RECT 125.340 141.130 125.700 141.510 ;
        RECT 125.970 141.130 126.330 141.510 ;
        RECT 126.570 141.130 126.930 141.510 ;
        RECT 2.515 140.540 2.875 140.920 ;
        RECT 3.145 140.540 3.505 140.920 ;
        RECT 3.745 140.540 4.105 140.920 ;
        RECT 125.340 140.540 125.700 140.920 ;
        RECT 125.970 140.540 126.330 140.920 ;
        RECT 126.570 140.540 126.930 140.920 ;
        RECT 4.830 138.900 5.830 139.900 ;
        RECT 6.430 138.900 7.430 139.900 ;
        RECT 8.030 138.900 9.030 139.900 ;
        RECT 2.515 137.220 2.875 137.600 ;
        RECT 3.145 137.220 3.505 137.600 ;
        RECT 3.745 137.220 4.105 137.600 ;
        RECT 4.830 137.300 5.830 138.300 ;
        RECT 2.515 136.630 2.875 137.010 ;
        RECT 3.145 136.630 3.505 137.010 ;
        RECT 3.745 136.630 4.105 137.010 ;
        RECT 4.830 135.700 5.830 136.700 ;
        RECT 20.430 138.900 21.430 139.900 ;
        RECT 22.030 138.900 23.030 139.900 ;
        RECT 23.630 138.900 24.630 139.900 ;
        RECT 24.830 138.900 25.830 139.900 ;
        RECT 26.430 138.900 27.430 139.900 ;
        RECT 28.030 138.900 29.030 139.900 ;
        RECT 2.520 134.925 2.880 135.305 ;
        RECT 3.130 134.925 3.490 135.305 ;
        RECT 3.760 134.925 4.120 135.305 ;
        RECT 2.520 134.190 2.880 134.570 ;
        RECT 3.130 134.190 3.490 134.570 ;
        RECT 3.760 134.190 4.120 134.570 ;
        RECT 2.520 133.505 2.880 133.885 ;
        RECT 3.130 133.505 3.490 133.885 ;
        RECT 3.760 133.505 4.120 133.885 ;
        RECT 23.630 137.300 24.630 138.300 ;
        RECT 24.830 137.300 25.830 138.300 ;
        RECT 23.630 135.700 24.630 136.700 ;
        RECT 24.830 135.700 25.830 136.700 ;
        RECT 40.430 138.900 41.430 139.900 ;
        RECT 42.030 138.900 43.030 139.900 ;
        RECT 43.630 138.900 44.630 139.900 ;
        RECT 44.830 138.900 45.830 139.900 ;
        RECT 46.430 138.900 47.430 139.900 ;
        RECT 48.030 138.900 49.030 139.900 ;
        RECT 43.630 137.300 44.630 138.300 ;
        RECT 44.830 137.300 45.830 138.300 ;
        RECT 43.630 135.700 44.630 136.700 ;
        RECT 44.830 135.700 45.830 136.700 ;
        RECT 60.430 138.900 61.430 139.900 ;
        RECT 62.030 138.900 63.030 139.900 ;
        RECT 63.630 138.900 64.630 139.900 ;
        RECT 64.830 138.900 65.830 139.900 ;
        RECT 66.430 138.900 67.430 139.900 ;
        RECT 68.030 138.900 69.030 139.900 ;
        RECT 63.630 137.300 64.630 138.300 ;
        RECT 64.830 137.300 65.830 138.300 ;
        RECT 63.630 135.700 64.630 136.700 ;
        RECT 64.830 135.700 65.830 136.700 ;
        RECT 80.430 138.900 81.430 139.900 ;
        RECT 82.030 138.900 83.030 139.900 ;
        RECT 83.630 138.900 84.630 139.900 ;
        RECT 84.830 138.900 85.830 139.900 ;
        RECT 86.430 138.900 87.430 139.900 ;
        RECT 88.030 138.900 89.030 139.900 ;
        RECT 83.630 137.300 84.630 138.300 ;
        RECT 84.830 137.300 85.830 138.300 ;
        RECT 83.630 135.700 84.630 136.700 ;
        RECT 84.830 135.700 85.830 136.700 ;
        RECT 100.430 138.900 101.430 139.900 ;
        RECT 102.030 138.900 103.030 139.900 ;
        RECT 103.630 138.900 104.630 139.900 ;
        RECT 104.830 138.900 105.830 139.900 ;
        RECT 106.430 138.900 107.430 139.900 ;
        RECT 108.030 138.900 109.030 139.900 ;
        RECT 103.630 137.300 104.630 138.300 ;
        RECT 104.830 137.300 105.830 138.300 ;
        RECT 103.630 135.700 104.630 136.700 ;
        RECT 104.830 135.700 105.830 136.700 ;
        RECT 120.430 138.900 121.430 139.900 ;
        RECT 122.030 138.900 123.030 139.900 ;
        RECT 123.630 138.900 124.630 139.900 ;
        RECT 123.630 137.300 124.630 138.300 ;
        RECT 125.340 137.220 125.700 137.600 ;
        RECT 125.970 137.220 126.330 137.600 ;
        RECT 126.570 137.220 126.930 137.600 ;
        RECT 123.630 135.700 124.630 136.700 ;
        RECT 125.340 136.630 125.700 137.010 ;
        RECT 125.970 136.630 126.330 137.010 ;
        RECT 126.570 136.630 126.930 137.010 ;
        RECT 2.520 126.090 2.880 126.470 ;
        RECT 3.130 126.090 3.490 126.470 ;
        RECT 3.760 126.090 4.120 126.470 ;
        RECT 2.520 125.355 2.880 125.735 ;
        RECT 3.130 125.355 3.490 125.735 ;
        RECT 3.760 125.355 4.120 125.735 ;
        RECT 2.520 124.670 2.880 125.050 ;
        RECT 3.130 124.670 3.490 125.050 ;
        RECT 3.760 124.670 4.120 125.050 ;
        RECT 4.830 123.300 5.830 124.300 ;
        RECT 2.515 122.660 2.875 123.040 ;
        RECT 3.145 122.660 3.505 123.040 ;
        RECT 3.745 122.660 4.105 123.040 ;
        RECT 2.515 122.070 2.875 122.450 ;
        RECT 3.145 122.070 3.505 122.450 ;
        RECT 3.745 122.070 4.105 122.450 ;
        RECT 4.830 121.700 5.830 122.700 ;
        RECT 4.830 120.100 5.830 121.100 ;
        RECT 6.430 120.100 7.430 121.100 ;
        RECT 8.030 120.100 9.030 121.100 ;
        RECT 23.630 123.300 24.630 124.300 ;
        RECT 24.830 123.300 25.830 124.300 ;
        RECT 23.630 121.700 24.630 122.700 ;
        RECT 24.830 121.700 25.830 122.700 ;
        RECT 4.830 118.900 5.830 119.900 ;
        RECT 6.430 118.900 7.430 119.900 ;
        RECT 8.030 118.900 9.030 119.900 ;
        RECT 20.430 120.100 21.430 121.100 ;
        RECT 22.030 120.100 23.030 121.100 ;
        RECT 23.630 120.100 24.630 121.100 ;
        RECT 24.830 120.100 25.830 121.100 ;
        RECT 26.430 120.100 27.430 121.100 ;
        RECT 28.030 120.100 29.030 121.100 ;
        RECT 43.630 123.300 44.630 124.300 ;
        RECT 44.830 123.300 45.830 124.300 ;
        RECT 43.630 121.700 44.630 122.700 ;
        RECT 44.830 121.700 45.830 122.700 ;
        RECT 2.515 117.640 2.875 118.020 ;
        RECT 3.145 117.640 3.505 118.020 ;
        RECT 3.745 117.640 4.105 118.020 ;
        RECT 2.515 117.050 2.875 117.430 ;
        RECT 3.145 117.050 3.505 117.430 ;
        RECT 3.745 117.050 4.105 117.430 ;
        RECT 4.830 117.300 5.830 118.300 ;
        RECT 4.830 115.700 5.830 116.700 ;
        RECT 20.430 118.900 21.430 119.900 ;
        RECT 22.030 118.900 23.030 119.900 ;
        RECT 23.630 118.900 24.630 119.900 ;
        RECT 24.830 118.900 25.830 119.900 ;
        RECT 26.430 118.900 27.430 119.900 ;
        RECT 28.030 118.900 29.030 119.900 ;
        RECT 40.430 120.100 41.430 121.100 ;
        RECT 42.030 120.100 43.030 121.100 ;
        RECT 43.630 120.100 44.630 121.100 ;
        RECT 44.830 120.100 45.830 121.100 ;
        RECT 46.430 120.100 47.430 121.100 ;
        RECT 48.030 120.100 49.030 121.100 ;
        RECT 63.630 123.300 64.630 124.300 ;
        RECT 64.830 123.300 65.830 124.300 ;
        RECT 63.630 121.700 64.630 122.700 ;
        RECT 64.830 121.700 65.830 122.700 ;
        RECT 2.520 114.920 2.880 115.300 ;
        RECT 3.130 114.920 3.490 115.300 ;
        RECT 3.760 114.920 4.120 115.300 ;
        RECT 2.520 114.185 2.880 114.565 ;
        RECT 3.130 114.185 3.490 114.565 ;
        RECT 3.760 114.185 4.120 114.565 ;
        RECT 2.520 113.500 2.880 113.880 ;
        RECT 3.130 113.500 3.490 113.880 ;
        RECT 3.760 113.500 4.120 113.880 ;
        RECT 23.630 117.300 24.630 118.300 ;
        RECT 24.830 117.300 25.830 118.300 ;
        RECT 23.630 115.700 24.630 116.700 ;
        RECT 24.830 115.700 25.830 116.700 ;
        RECT 40.430 118.900 41.430 119.900 ;
        RECT 42.030 118.900 43.030 119.900 ;
        RECT 43.630 118.900 44.630 119.900 ;
        RECT 44.830 118.900 45.830 119.900 ;
        RECT 46.430 118.900 47.430 119.900 ;
        RECT 48.030 118.900 49.030 119.900 ;
        RECT 60.430 120.100 61.430 121.100 ;
        RECT 62.030 120.100 63.030 121.100 ;
        RECT 63.630 120.100 64.630 121.100 ;
        RECT 64.830 120.100 65.830 121.100 ;
        RECT 66.430 120.100 67.430 121.100 ;
        RECT 68.030 120.100 69.030 121.100 ;
        RECT 83.630 123.300 84.630 124.300 ;
        RECT 84.830 123.300 85.830 124.300 ;
        RECT 83.630 121.700 84.630 122.700 ;
        RECT 84.830 121.700 85.830 122.700 ;
        RECT 43.630 117.300 44.630 118.300 ;
        RECT 44.830 117.300 45.830 118.300 ;
        RECT 43.630 115.700 44.630 116.700 ;
        RECT 44.830 115.700 45.830 116.700 ;
        RECT 60.430 118.900 61.430 119.900 ;
        RECT 62.030 118.900 63.030 119.900 ;
        RECT 63.630 118.900 64.630 119.900 ;
        RECT 64.830 118.900 65.830 119.900 ;
        RECT 66.430 118.900 67.430 119.900 ;
        RECT 68.030 118.900 69.030 119.900 ;
        RECT 80.430 120.100 81.430 121.100 ;
        RECT 82.030 120.100 83.030 121.100 ;
        RECT 83.630 120.100 84.630 121.100 ;
        RECT 84.830 120.100 85.830 121.100 ;
        RECT 86.430 120.100 87.430 121.100 ;
        RECT 88.030 120.100 89.030 121.100 ;
        RECT 103.630 123.300 104.630 124.300 ;
        RECT 104.830 123.300 105.830 124.300 ;
        RECT 103.630 121.700 104.630 122.700 ;
        RECT 104.830 121.700 105.830 122.700 ;
        RECT 63.630 117.300 64.630 118.300 ;
        RECT 64.830 117.300 65.830 118.300 ;
        RECT 63.630 115.700 64.630 116.700 ;
        RECT 64.830 115.700 65.830 116.700 ;
        RECT 80.430 118.900 81.430 119.900 ;
        RECT 82.030 118.900 83.030 119.900 ;
        RECT 83.630 118.900 84.630 119.900 ;
        RECT 84.830 118.900 85.830 119.900 ;
        RECT 86.430 118.900 87.430 119.900 ;
        RECT 88.030 118.900 89.030 119.900 ;
        RECT 100.430 120.100 101.430 121.100 ;
        RECT 102.030 120.100 103.030 121.100 ;
        RECT 103.630 120.100 104.630 121.100 ;
        RECT 104.830 120.100 105.830 121.100 ;
        RECT 106.430 120.100 107.430 121.100 ;
        RECT 108.030 120.100 109.030 121.100 ;
        RECT 123.630 123.300 124.630 124.300 ;
        RECT 123.630 121.700 124.630 122.700 ;
        RECT 125.340 122.415 125.700 122.795 ;
        RECT 125.970 122.415 126.330 122.795 ;
        RECT 126.570 122.415 126.930 122.795 ;
        RECT 125.340 121.825 125.700 122.205 ;
        RECT 125.970 121.825 126.330 122.205 ;
        RECT 126.570 121.825 126.930 122.205 ;
        RECT 83.630 117.300 84.630 118.300 ;
        RECT 84.830 117.300 85.830 118.300 ;
        RECT 83.630 115.700 84.630 116.700 ;
        RECT 84.830 115.700 85.830 116.700 ;
        RECT 100.430 118.900 101.430 119.900 ;
        RECT 102.030 118.900 103.030 119.900 ;
        RECT 103.630 118.900 104.630 119.900 ;
        RECT 104.830 118.900 105.830 119.900 ;
        RECT 106.430 118.900 107.430 119.900 ;
        RECT 108.030 118.900 109.030 119.900 ;
        RECT 120.430 120.100 121.430 121.100 ;
        RECT 122.030 120.100 123.030 121.100 ;
        RECT 123.630 120.100 124.630 121.100 ;
        RECT 103.630 117.300 104.630 118.300 ;
        RECT 104.830 117.300 105.830 118.300 ;
        RECT 103.630 115.700 104.630 116.700 ;
        RECT 104.830 115.700 105.830 116.700 ;
        RECT 120.430 118.900 121.430 119.900 ;
        RECT 122.030 118.900 123.030 119.900 ;
        RECT 123.630 118.900 124.630 119.900 ;
        RECT 123.630 117.300 124.630 118.300 ;
        RECT 125.340 116.830 125.700 117.210 ;
        RECT 125.970 116.830 126.330 117.210 ;
        RECT 126.570 116.830 126.930 117.210 ;
        RECT 123.630 115.700 124.630 116.700 ;
        RECT 125.340 116.240 125.700 116.620 ;
        RECT 125.970 116.240 126.330 116.620 ;
        RECT 126.570 116.240 126.930 116.620 ;
        RECT 2.520 106.120 2.880 106.500 ;
        RECT 3.130 106.120 3.490 106.500 ;
        RECT 3.760 106.120 4.120 106.500 ;
        RECT 2.520 105.385 2.880 105.765 ;
        RECT 3.130 105.385 3.490 105.765 ;
        RECT 3.760 105.385 4.120 105.765 ;
        RECT 2.520 104.700 2.880 105.080 ;
        RECT 3.130 104.700 3.490 105.080 ;
        RECT 3.760 104.700 4.120 105.080 ;
        RECT 4.830 103.300 5.830 104.300 ;
        RECT 2.515 102.750 2.875 103.130 ;
        RECT 3.145 102.750 3.505 103.130 ;
        RECT 3.745 102.750 4.105 103.130 ;
        RECT 2.515 102.160 2.875 102.540 ;
        RECT 3.145 102.160 3.505 102.540 ;
        RECT 3.745 102.160 4.105 102.540 ;
        RECT 4.830 101.700 5.830 102.700 ;
        RECT 4.830 100.100 5.830 101.100 ;
        RECT 6.430 100.100 7.430 101.100 ;
        RECT 8.030 100.100 9.030 101.100 ;
        RECT 23.630 103.300 24.630 104.300 ;
        RECT 24.830 103.300 25.830 104.300 ;
        RECT 23.630 101.700 24.630 102.700 ;
        RECT 24.830 101.700 25.830 102.700 ;
        RECT 4.830 98.900 5.830 99.900 ;
        RECT 6.430 98.900 7.430 99.900 ;
        RECT 8.030 98.900 9.030 99.900 ;
        RECT 20.430 100.100 21.430 101.100 ;
        RECT 22.030 100.100 23.030 101.100 ;
        RECT 23.630 100.100 24.630 101.100 ;
        RECT 24.830 100.100 25.830 101.100 ;
        RECT 26.430 100.100 27.430 101.100 ;
        RECT 28.030 100.100 29.030 101.100 ;
        RECT 43.630 103.300 44.630 104.300 ;
        RECT 44.830 103.300 45.830 104.300 ;
        RECT 43.630 101.700 44.630 102.700 ;
        RECT 44.830 101.700 45.830 102.700 ;
        RECT 2.515 97.340 2.875 97.720 ;
        RECT 3.145 97.340 3.505 97.720 ;
        RECT 3.745 97.340 4.105 97.720 ;
        RECT 4.830 97.300 5.830 98.300 ;
        RECT 2.515 96.750 2.875 97.130 ;
        RECT 3.145 96.750 3.505 97.130 ;
        RECT 3.745 96.750 4.105 97.130 ;
        RECT 4.830 95.700 5.830 96.700 ;
        RECT 20.430 98.900 21.430 99.900 ;
        RECT 22.030 98.900 23.030 99.900 ;
        RECT 23.630 98.900 24.630 99.900 ;
        RECT 24.830 98.900 25.830 99.900 ;
        RECT 26.430 98.900 27.430 99.900 ;
        RECT 28.030 98.900 29.030 99.900 ;
        RECT 40.430 100.100 41.430 101.100 ;
        RECT 42.030 100.100 43.030 101.100 ;
        RECT 43.630 100.100 44.630 101.100 ;
        RECT 44.830 100.100 45.830 101.100 ;
        RECT 46.430 100.100 47.430 101.100 ;
        RECT 48.030 100.100 49.030 101.100 ;
        RECT 63.630 103.300 64.630 104.300 ;
        RECT 64.830 103.300 65.830 104.300 ;
        RECT 63.630 101.700 64.630 102.700 ;
        RECT 64.830 101.700 65.830 102.700 ;
        RECT 2.520 94.920 2.880 95.300 ;
        RECT 3.130 94.920 3.490 95.300 ;
        RECT 3.760 94.920 4.120 95.300 ;
        RECT 2.520 94.185 2.880 94.565 ;
        RECT 3.130 94.185 3.490 94.565 ;
        RECT 3.760 94.185 4.120 94.565 ;
        RECT 2.520 93.500 2.880 93.880 ;
        RECT 3.130 93.500 3.490 93.880 ;
        RECT 3.760 93.500 4.120 93.880 ;
        RECT 23.630 97.300 24.630 98.300 ;
        RECT 24.830 97.300 25.830 98.300 ;
        RECT 23.630 95.700 24.630 96.700 ;
        RECT 24.830 95.700 25.830 96.700 ;
        RECT 40.430 98.900 41.430 99.900 ;
        RECT 42.030 98.900 43.030 99.900 ;
        RECT 43.630 98.900 44.630 99.900 ;
        RECT 44.830 98.900 45.830 99.900 ;
        RECT 46.430 98.900 47.430 99.900 ;
        RECT 48.030 98.900 49.030 99.900 ;
        RECT 60.430 100.100 61.430 101.100 ;
        RECT 62.030 100.100 63.030 101.100 ;
        RECT 63.630 100.100 64.630 101.100 ;
        RECT 64.830 100.100 65.830 101.100 ;
        RECT 66.430 100.100 67.430 101.100 ;
        RECT 68.030 100.100 69.030 101.100 ;
        RECT 83.630 103.300 84.630 104.300 ;
        RECT 84.830 103.300 85.830 104.300 ;
        RECT 83.630 101.700 84.630 102.700 ;
        RECT 84.830 101.700 85.830 102.700 ;
        RECT 43.630 97.300 44.630 98.300 ;
        RECT 44.830 97.300 45.830 98.300 ;
        RECT 43.630 95.700 44.630 96.700 ;
        RECT 44.830 95.700 45.830 96.700 ;
        RECT 60.430 98.900 61.430 99.900 ;
        RECT 62.030 98.900 63.030 99.900 ;
        RECT 63.630 98.900 64.630 99.900 ;
        RECT 64.830 98.900 65.830 99.900 ;
        RECT 66.430 98.900 67.430 99.900 ;
        RECT 68.030 98.900 69.030 99.900 ;
        RECT 80.430 100.100 81.430 101.100 ;
        RECT 82.030 100.100 83.030 101.100 ;
        RECT 83.630 100.100 84.630 101.100 ;
        RECT 84.830 100.100 85.830 101.100 ;
        RECT 86.430 100.100 87.430 101.100 ;
        RECT 88.030 100.100 89.030 101.100 ;
        RECT 103.630 103.300 104.630 104.300 ;
        RECT 104.830 103.300 105.830 104.300 ;
        RECT 103.630 101.700 104.630 102.700 ;
        RECT 104.830 101.700 105.830 102.700 ;
        RECT 63.630 97.300 64.630 98.300 ;
        RECT 64.830 97.300 65.830 98.300 ;
        RECT 63.630 95.700 64.630 96.700 ;
        RECT 64.830 95.700 65.830 96.700 ;
        RECT 80.430 98.900 81.430 99.900 ;
        RECT 82.030 98.900 83.030 99.900 ;
        RECT 83.630 98.900 84.630 99.900 ;
        RECT 84.830 98.900 85.830 99.900 ;
        RECT 86.430 98.900 87.430 99.900 ;
        RECT 88.030 98.900 89.030 99.900 ;
        RECT 100.430 100.100 101.430 101.100 ;
        RECT 102.030 100.100 103.030 101.100 ;
        RECT 103.630 100.100 104.630 101.100 ;
        RECT 104.830 100.100 105.830 101.100 ;
        RECT 106.430 100.100 107.430 101.100 ;
        RECT 108.030 100.100 109.030 101.100 ;
        RECT 123.630 103.300 124.630 104.300 ;
        RECT 123.630 101.700 124.630 102.700 ;
        RECT 125.340 102.615 125.700 102.995 ;
        RECT 125.970 102.615 126.330 102.995 ;
        RECT 126.570 102.615 126.930 102.995 ;
        RECT 125.340 102.025 125.700 102.405 ;
        RECT 125.970 102.025 126.330 102.405 ;
        RECT 126.570 102.025 126.930 102.405 ;
        RECT 83.630 97.300 84.630 98.300 ;
        RECT 84.830 97.300 85.830 98.300 ;
        RECT 83.630 95.700 84.630 96.700 ;
        RECT 84.830 95.700 85.830 96.700 ;
        RECT 100.430 98.900 101.430 99.900 ;
        RECT 102.030 98.900 103.030 99.900 ;
        RECT 103.630 98.900 104.630 99.900 ;
        RECT 104.830 98.900 105.830 99.900 ;
        RECT 106.430 98.900 107.430 99.900 ;
        RECT 108.030 98.900 109.030 99.900 ;
        RECT 120.430 100.100 121.430 101.100 ;
        RECT 122.030 100.100 123.030 101.100 ;
        RECT 123.630 100.100 124.630 101.100 ;
        RECT 103.630 97.300 104.630 98.300 ;
        RECT 104.830 97.300 105.830 98.300 ;
        RECT 103.630 95.700 104.630 96.700 ;
        RECT 104.830 95.700 105.830 96.700 ;
        RECT 120.430 98.900 121.430 99.900 ;
        RECT 122.030 98.900 123.030 99.900 ;
        RECT 123.630 98.900 124.630 99.900 ;
        RECT 123.630 97.300 124.630 98.300 ;
        RECT 125.340 96.740 125.700 97.120 ;
        RECT 125.970 96.740 126.330 97.120 ;
        RECT 126.570 96.740 126.930 97.120 ;
        RECT 123.630 95.700 124.630 96.700 ;
        RECT 125.340 96.150 125.700 96.530 ;
        RECT 125.970 96.150 126.330 96.530 ;
        RECT 126.570 96.150 126.930 96.530 ;
        RECT 2.520 86.125 2.880 86.505 ;
        RECT 3.130 86.125 3.490 86.505 ;
        RECT 3.760 86.125 4.120 86.505 ;
        RECT 2.520 85.390 2.880 85.770 ;
        RECT 3.130 85.390 3.490 85.770 ;
        RECT 3.760 85.390 4.120 85.770 ;
        RECT 2.520 84.705 2.880 85.085 ;
        RECT 3.130 84.705 3.490 85.085 ;
        RECT 3.760 84.705 4.120 85.085 ;
        RECT 2.515 82.965 2.875 83.345 ;
        RECT 3.145 82.965 3.505 83.345 ;
        RECT 3.745 82.965 4.105 83.345 ;
        RECT 4.830 83.300 5.830 84.300 ;
        RECT 2.515 82.375 2.875 82.755 ;
        RECT 3.145 82.375 3.505 82.755 ;
        RECT 3.745 82.375 4.105 82.755 ;
        RECT 4.830 81.700 5.830 82.700 ;
        RECT 4.830 80.100 5.830 81.100 ;
        RECT 6.430 80.100 7.430 81.100 ;
        RECT 8.030 80.100 9.030 81.100 ;
        RECT 23.630 83.300 24.630 84.300 ;
        RECT 24.830 83.300 25.830 84.300 ;
        RECT 23.630 81.700 24.630 82.700 ;
        RECT 24.830 81.700 25.830 82.700 ;
        RECT 4.830 78.900 5.830 79.900 ;
        RECT 6.430 78.900 7.430 79.900 ;
        RECT 8.030 78.900 9.030 79.900 ;
        RECT 20.430 80.100 21.430 81.100 ;
        RECT 22.030 80.100 23.030 81.100 ;
        RECT 23.630 80.100 24.630 81.100 ;
        RECT 24.830 80.100 25.830 81.100 ;
        RECT 26.430 80.100 27.430 81.100 ;
        RECT 28.030 80.100 29.030 81.100 ;
        RECT 43.630 83.300 44.630 84.300 ;
        RECT 44.830 83.300 45.830 84.300 ;
        RECT 43.630 81.700 44.630 82.700 ;
        RECT 44.830 81.700 45.830 82.700 ;
        RECT 2.515 77.460 2.875 77.840 ;
        RECT 3.145 77.460 3.505 77.840 ;
        RECT 3.745 77.460 4.105 77.840 ;
        RECT 4.830 77.300 5.830 78.300 ;
        RECT 2.515 76.870 2.875 77.250 ;
        RECT 3.145 76.870 3.505 77.250 ;
        RECT 3.745 76.870 4.105 77.250 ;
        RECT 4.830 75.700 5.830 76.700 ;
        RECT 20.430 78.900 21.430 79.900 ;
        RECT 22.030 78.900 23.030 79.900 ;
        RECT 23.630 78.900 24.630 79.900 ;
        RECT 24.830 78.900 25.830 79.900 ;
        RECT 26.430 78.900 27.430 79.900 ;
        RECT 28.030 78.900 29.030 79.900 ;
        RECT 40.430 80.100 41.430 81.100 ;
        RECT 42.030 80.100 43.030 81.100 ;
        RECT 43.630 80.100 44.630 81.100 ;
        RECT 44.830 80.100 45.830 81.100 ;
        RECT 46.430 80.100 47.430 81.100 ;
        RECT 48.030 80.100 49.030 81.100 ;
        RECT 63.630 83.300 64.630 84.300 ;
        RECT 64.830 83.300 65.830 84.300 ;
        RECT 63.630 81.700 64.630 82.700 ;
        RECT 64.830 81.700 65.830 82.700 ;
        RECT 2.520 74.920 2.880 75.300 ;
        RECT 3.130 74.920 3.490 75.300 ;
        RECT 3.760 74.920 4.120 75.300 ;
        RECT 2.520 74.185 2.880 74.565 ;
        RECT 3.130 74.185 3.490 74.565 ;
        RECT 3.760 74.185 4.120 74.565 ;
        RECT 2.520 73.500 2.880 73.880 ;
        RECT 3.130 73.500 3.490 73.880 ;
        RECT 3.760 73.500 4.120 73.880 ;
        RECT 23.630 77.300 24.630 78.300 ;
        RECT 24.830 77.300 25.830 78.300 ;
        RECT 23.630 75.700 24.630 76.700 ;
        RECT 24.830 75.700 25.830 76.700 ;
        RECT 40.430 78.900 41.430 79.900 ;
        RECT 42.030 78.900 43.030 79.900 ;
        RECT 43.630 78.900 44.630 79.900 ;
        RECT 44.830 78.900 45.830 79.900 ;
        RECT 46.430 78.900 47.430 79.900 ;
        RECT 48.030 78.900 49.030 79.900 ;
        RECT 60.430 80.100 61.430 81.100 ;
        RECT 62.030 80.100 63.030 81.100 ;
        RECT 63.630 80.100 64.630 81.100 ;
        RECT 64.830 80.100 65.830 81.100 ;
        RECT 66.430 80.100 67.430 81.100 ;
        RECT 68.030 80.100 69.030 81.100 ;
        RECT 83.630 83.300 84.630 84.300 ;
        RECT 84.830 83.300 85.830 84.300 ;
        RECT 83.630 81.700 84.630 82.700 ;
        RECT 84.830 81.700 85.830 82.700 ;
        RECT 43.630 77.300 44.630 78.300 ;
        RECT 44.830 77.300 45.830 78.300 ;
        RECT 43.630 75.700 44.630 76.700 ;
        RECT 44.830 75.700 45.830 76.700 ;
        RECT 60.430 78.900 61.430 79.900 ;
        RECT 62.030 78.900 63.030 79.900 ;
        RECT 63.630 78.900 64.630 79.900 ;
        RECT 64.830 78.900 65.830 79.900 ;
        RECT 66.430 78.900 67.430 79.900 ;
        RECT 68.030 78.900 69.030 79.900 ;
        RECT 80.430 80.100 81.430 81.100 ;
        RECT 82.030 80.100 83.030 81.100 ;
        RECT 83.630 80.100 84.630 81.100 ;
        RECT 84.830 80.100 85.830 81.100 ;
        RECT 86.430 80.100 87.430 81.100 ;
        RECT 88.030 80.100 89.030 81.100 ;
        RECT 103.630 83.300 104.630 84.300 ;
        RECT 104.830 83.300 105.830 84.300 ;
        RECT 103.630 81.700 104.630 82.700 ;
        RECT 104.830 81.700 105.830 82.700 ;
        RECT 63.630 77.300 64.630 78.300 ;
        RECT 64.830 77.300 65.830 78.300 ;
        RECT 63.630 75.700 64.630 76.700 ;
        RECT 64.830 75.700 65.830 76.700 ;
        RECT 80.430 78.900 81.430 79.900 ;
        RECT 82.030 78.900 83.030 79.900 ;
        RECT 83.630 78.900 84.630 79.900 ;
        RECT 84.830 78.900 85.830 79.900 ;
        RECT 86.430 78.900 87.430 79.900 ;
        RECT 88.030 78.900 89.030 79.900 ;
        RECT 100.430 80.100 101.430 81.100 ;
        RECT 102.030 80.100 103.030 81.100 ;
        RECT 103.630 80.100 104.630 81.100 ;
        RECT 104.830 80.100 105.830 81.100 ;
        RECT 106.430 80.100 107.430 81.100 ;
        RECT 108.030 80.100 109.030 81.100 ;
        RECT 123.630 83.300 124.630 84.300 ;
        RECT 123.630 81.700 124.630 82.700 ;
        RECT 125.340 82.535 125.700 82.915 ;
        RECT 125.970 82.535 126.330 82.915 ;
        RECT 126.570 82.535 126.930 82.915 ;
        RECT 125.340 81.945 125.700 82.325 ;
        RECT 125.970 81.945 126.330 82.325 ;
        RECT 126.570 81.945 126.930 82.325 ;
        RECT 83.630 77.300 84.630 78.300 ;
        RECT 84.830 77.300 85.830 78.300 ;
        RECT 83.630 75.700 84.630 76.700 ;
        RECT 84.830 75.700 85.830 76.700 ;
        RECT 100.430 78.900 101.430 79.900 ;
        RECT 102.030 78.900 103.030 79.900 ;
        RECT 103.630 78.900 104.630 79.900 ;
        RECT 104.830 78.900 105.830 79.900 ;
        RECT 106.430 78.900 107.430 79.900 ;
        RECT 108.030 78.900 109.030 79.900 ;
        RECT 120.430 80.100 121.430 81.100 ;
        RECT 122.030 80.100 123.030 81.100 ;
        RECT 123.630 80.100 124.630 81.100 ;
        RECT 103.630 77.300 104.630 78.300 ;
        RECT 104.830 77.300 105.830 78.300 ;
        RECT 103.630 75.700 104.630 76.700 ;
        RECT 104.830 75.700 105.830 76.700 ;
        RECT 120.430 78.900 121.430 79.900 ;
        RECT 122.030 78.900 123.030 79.900 ;
        RECT 123.630 78.900 124.630 79.900 ;
        RECT 123.630 77.300 124.630 78.300 ;
        RECT 123.630 75.700 124.630 76.700 ;
        RECT 125.340 76.680 125.700 77.060 ;
        RECT 125.970 76.680 126.330 77.060 ;
        RECT 126.570 76.680 126.930 77.060 ;
        RECT 125.340 76.090 125.700 76.470 ;
        RECT 125.970 76.090 126.330 76.470 ;
        RECT 126.570 76.090 126.930 76.470 ;
        RECT 2.520 66.120 2.880 66.500 ;
        RECT 3.130 66.120 3.490 66.500 ;
        RECT 3.760 66.120 4.120 66.500 ;
        RECT 2.520 65.385 2.880 65.765 ;
        RECT 3.130 65.385 3.490 65.765 ;
        RECT 3.760 65.385 4.120 65.765 ;
        RECT 2.520 64.700 2.880 65.080 ;
        RECT 3.130 64.700 3.490 65.080 ;
        RECT 3.760 64.700 4.120 65.080 ;
        RECT 2.515 63.130 2.875 63.510 ;
        RECT 3.145 63.130 3.505 63.510 ;
        RECT 3.745 63.130 4.105 63.510 ;
        RECT 4.830 63.300 5.830 64.300 ;
        RECT 2.515 62.540 2.875 62.920 ;
        RECT 3.145 62.540 3.505 62.920 ;
        RECT 3.745 62.540 4.105 62.920 ;
        RECT 4.830 61.700 5.830 62.700 ;
        RECT 4.830 60.100 5.830 61.100 ;
        RECT 6.430 60.100 7.430 61.100 ;
        RECT 8.030 60.100 9.030 61.100 ;
        RECT 23.630 63.300 24.630 64.300 ;
        RECT 24.830 63.300 25.830 64.300 ;
        RECT 23.630 61.700 24.630 62.700 ;
        RECT 24.830 61.700 25.830 62.700 ;
        RECT 4.830 58.900 5.830 59.900 ;
        RECT 6.430 58.900 7.430 59.900 ;
        RECT 8.030 58.900 9.030 59.900 ;
        RECT 20.430 60.100 21.430 61.100 ;
        RECT 22.030 60.100 23.030 61.100 ;
        RECT 23.630 60.100 24.630 61.100 ;
        RECT 24.830 60.100 25.830 61.100 ;
        RECT 26.430 60.100 27.430 61.100 ;
        RECT 28.030 60.100 29.030 61.100 ;
        RECT 43.630 63.300 44.630 64.300 ;
        RECT 44.830 63.300 45.830 64.300 ;
        RECT 43.630 61.700 44.630 62.700 ;
        RECT 44.830 61.700 45.830 62.700 ;
        RECT 2.515 57.050 2.875 57.430 ;
        RECT 3.145 57.050 3.505 57.430 ;
        RECT 3.745 57.050 4.105 57.430 ;
        RECT 4.830 57.300 5.830 58.300 ;
        RECT 2.515 56.460 2.875 56.840 ;
        RECT 3.145 56.460 3.505 56.840 ;
        RECT 3.745 56.460 4.105 56.840 ;
        RECT 4.830 55.700 5.830 56.700 ;
        RECT 20.430 58.900 21.430 59.900 ;
        RECT 22.030 58.900 23.030 59.900 ;
        RECT 23.630 58.900 24.630 59.900 ;
        RECT 24.830 58.900 25.830 59.900 ;
        RECT 26.430 58.900 27.430 59.900 ;
        RECT 28.030 58.900 29.030 59.900 ;
        RECT 40.430 60.100 41.430 61.100 ;
        RECT 42.030 60.100 43.030 61.100 ;
        RECT 43.630 60.100 44.630 61.100 ;
        RECT 44.830 60.100 45.830 61.100 ;
        RECT 46.430 60.100 47.430 61.100 ;
        RECT 48.030 60.100 49.030 61.100 ;
        RECT 63.630 63.300 64.630 64.300 ;
        RECT 64.830 63.300 65.830 64.300 ;
        RECT 63.630 61.700 64.630 62.700 ;
        RECT 64.830 61.700 65.830 62.700 ;
        RECT 2.520 54.920 2.880 55.300 ;
        RECT 3.130 54.920 3.490 55.300 ;
        RECT 3.760 54.920 4.120 55.300 ;
        RECT 2.520 54.185 2.880 54.565 ;
        RECT 3.130 54.185 3.490 54.565 ;
        RECT 3.760 54.185 4.120 54.565 ;
        RECT 2.520 53.500 2.880 53.880 ;
        RECT 3.130 53.500 3.490 53.880 ;
        RECT 3.760 53.500 4.120 53.880 ;
        RECT 23.630 57.300 24.630 58.300 ;
        RECT 24.830 57.300 25.830 58.300 ;
        RECT 23.630 55.700 24.630 56.700 ;
        RECT 24.830 55.700 25.830 56.700 ;
        RECT 40.430 58.900 41.430 59.900 ;
        RECT 42.030 58.900 43.030 59.900 ;
        RECT 43.630 58.900 44.630 59.900 ;
        RECT 44.830 58.900 45.830 59.900 ;
        RECT 46.430 58.900 47.430 59.900 ;
        RECT 48.030 58.900 49.030 59.900 ;
        RECT 60.430 60.100 61.430 61.100 ;
        RECT 62.030 60.100 63.030 61.100 ;
        RECT 63.630 60.100 64.630 61.100 ;
        RECT 64.830 60.100 65.830 61.100 ;
        RECT 66.430 60.100 67.430 61.100 ;
        RECT 68.030 60.100 69.030 61.100 ;
        RECT 83.630 63.300 84.630 64.300 ;
        RECT 84.830 63.300 85.830 64.300 ;
        RECT 83.630 61.700 84.630 62.700 ;
        RECT 84.830 61.700 85.830 62.700 ;
        RECT 43.630 57.300 44.630 58.300 ;
        RECT 44.830 57.300 45.830 58.300 ;
        RECT 43.630 55.700 44.630 56.700 ;
        RECT 44.830 55.700 45.830 56.700 ;
        RECT 60.430 58.900 61.430 59.900 ;
        RECT 62.030 58.900 63.030 59.900 ;
        RECT 63.630 58.900 64.630 59.900 ;
        RECT 64.830 58.900 65.830 59.900 ;
        RECT 66.430 58.900 67.430 59.900 ;
        RECT 68.030 58.900 69.030 59.900 ;
        RECT 80.430 60.100 81.430 61.100 ;
        RECT 82.030 60.100 83.030 61.100 ;
        RECT 83.630 60.100 84.630 61.100 ;
        RECT 84.830 60.100 85.830 61.100 ;
        RECT 86.430 60.100 87.430 61.100 ;
        RECT 88.030 60.100 89.030 61.100 ;
        RECT 103.630 63.300 104.630 64.300 ;
        RECT 104.830 63.300 105.830 64.300 ;
        RECT 103.630 61.700 104.630 62.700 ;
        RECT 104.830 61.700 105.830 62.700 ;
        RECT 63.630 57.300 64.630 58.300 ;
        RECT 64.830 57.300 65.830 58.300 ;
        RECT 63.630 55.700 64.630 56.700 ;
        RECT 64.830 55.700 65.830 56.700 ;
        RECT 80.430 58.900 81.430 59.900 ;
        RECT 82.030 58.900 83.030 59.900 ;
        RECT 83.630 58.900 84.630 59.900 ;
        RECT 84.830 58.900 85.830 59.900 ;
        RECT 86.430 58.900 87.430 59.900 ;
        RECT 88.030 58.900 89.030 59.900 ;
        RECT 100.430 60.100 101.430 61.100 ;
        RECT 102.030 60.100 103.030 61.100 ;
        RECT 103.630 60.100 104.630 61.100 ;
        RECT 104.830 60.100 105.830 61.100 ;
        RECT 106.430 60.100 107.430 61.100 ;
        RECT 108.030 60.100 109.030 61.100 ;
        RECT 123.630 63.300 124.630 64.300 ;
        RECT 125.340 62.875 125.700 63.255 ;
        RECT 125.970 62.875 126.330 63.255 ;
        RECT 126.570 62.875 126.930 63.255 ;
        RECT 123.630 61.700 124.630 62.700 ;
        RECT 125.340 62.285 125.700 62.665 ;
        RECT 125.970 62.285 126.330 62.665 ;
        RECT 126.570 62.285 126.930 62.665 ;
        RECT 83.630 57.300 84.630 58.300 ;
        RECT 84.830 57.300 85.830 58.300 ;
        RECT 83.630 55.700 84.630 56.700 ;
        RECT 84.830 55.700 85.830 56.700 ;
        RECT 100.430 58.900 101.430 59.900 ;
        RECT 102.030 58.900 103.030 59.900 ;
        RECT 103.630 58.900 104.630 59.900 ;
        RECT 104.830 58.900 105.830 59.900 ;
        RECT 106.430 58.900 107.430 59.900 ;
        RECT 108.030 58.900 109.030 59.900 ;
        RECT 120.430 60.100 121.430 61.100 ;
        RECT 122.030 60.100 123.030 61.100 ;
        RECT 123.630 60.100 124.630 61.100 ;
        RECT 103.630 57.300 104.630 58.300 ;
        RECT 104.830 57.300 105.830 58.300 ;
        RECT 103.630 55.700 104.630 56.700 ;
        RECT 104.830 55.700 105.830 56.700 ;
        RECT 120.430 58.900 121.430 59.900 ;
        RECT 122.030 58.900 123.030 59.900 ;
        RECT 123.630 58.900 124.630 59.900 ;
        RECT 123.630 57.300 124.630 58.300 ;
        RECT 125.340 56.805 125.700 57.185 ;
        RECT 125.970 56.805 126.330 57.185 ;
        RECT 126.570 56.805 126.930 57.185 ;
        RECT 123.630 55.700 124.630 56.700 ;
        RECT 125.340 56.215 125.700 56.595 ;
        RECT 125.970 56.215 126.330 56.595 ;
        RECT 126.570 56.215 126.930 56.595 ;
        RECT 2.520 46.120 2.880 46.500 ;
        RECT 3.130 46.120 3.490 46.500 ;
        RECT 3.760 46.120 4.120 46.500 ;
        RECT 2.520 45.385 2.880 45.765 ;
        RECT 3.130 45.385 3.490 45.765 ;
        RECT 3.760 45.385 4.120 45.765 ;
        RECT 2.520 44.700 2.880 45.080 ;
        RECT 3.130 44.700 3.490 45.080 ;
        RECT 3.760 44.700 4.120 45.080 ;
        RECT 4.830 43.300 5.830 44.300 ;
        RECT 2.515 42.725 2.875 43.105 ;
        RECT 3.145 42.725 3.505 43.105 ;
        RECT 3.745 42.725 4.105 43.105 ;
        RECT 2.515 42.135 2.875 42.515 ;
        RECT 3.145 42.135 3.505 42.515 ;
        RECT 3.745 42.135 4.105 42.515 ;
        RECT 4.830 41.700 5.830 42.700 ;
        RECT 4.830 40.100 5.830 41.100 ;
        RECT 6.430 40.100 7.430 41.100 ;
        RECT 8.030 40.100 9.030 41.100 ;
        RECT 23.630 43.300 24.630 44.300 ;
        RECT 24.830 43.300 25.830 44.300 ;
        RECT 23.630 41.700 24.630 42.700 ;
        RECT 24.830 41.700 25.830 42.700 ;
        RECT 4.830 38.900 5.830 39.900 ;
        RECT 6.430 38.900 7.430 39.900 ;
        RECT 8.030 38.900 9.030 39.900 ;
        RECT 20.430 40.100 21.430 41.100 ;
        RECT 22.030 40.100 23.030 41.100 ;
        RECT 23.630 40.100 24.630 41.100 ;
        RECT 24.830 40.100 25.830 41.100 ;
        RECT 26.430 40.100 27.430 41.100 ;
        RECT 28.030 40.100 29.030 41.100 ;
        RECT 43.630 43.300 44.630 44.300 ;
        RECT 44.830 43.300 45.830 44.300 ;
        RECT 43.630 41.700 44.630 42.700 ;
        RECT 44.830 41.700 45.830 42.700 ;
        RECT 2.515 37.115 2.875 37.495 ;
        RECT 3.145 37.115 3.505 37.495 ;
        RECT 3.745 37.115 4.105 37.495 ;
        RECT 4.830 37.300 5.830 38.300 ;
        RECT 2.515 36.525 2.875 36.905 ;
        RECT 3.145 36.525 3.505 36.905 ;
        RECT 3.745 36.525 4.105 36.905 ;
        RECT 4.830 35.700 5.830 36.700 ;
        RECT 20.430 38.900 21.430 39.900 ;
        RECT 22.030 38.900 23.030 39.900 ;
        RECT 23.630 38.900 24.630 39.900 ;
        RECT 24.830 38.900 25.830 39.900 ;
        RECT 26.430 38.900 27.430 39.900 ;
        RECT 28.030 38.900 29.030 39.900 ;
        RECT 40.430 40.100 41.430 41.100 ;
        RECT 42.030 40.100 43.030 41.100 ;
        RECT 43.630 40.100 44.630 41.100 ;
        RECT 44.830 40.100 45.830 41.100 ;
        RECT 46.430 40.100 47.430 41.100 ;
        RECT 48.030 40.100 49.030 41.100 ;
        RECT 63.630 43.300 64.630 44.300 ;
        RECT 64.830 43.300 65.830 44.300 ;
        RECT 63.630 41.700 64.630 42.700 ;
        RECT 64.830 41.700 65.830 42.700 ;
        RECT 2.520 34.925 2.880 35.305 ;
        RECT 3.130 34.925 3.490 35.305 ;
        RECT 3.760 34.925 4.120 35.305 ;
        RECT 2.520 34.190 2.880 34.570 ;
        RECT 3.130 34.190 3.490 34.570 ;
        RECT 3.760 34.190 4.120 34.570 ;
        RECT 2.520 33.505 2.880 33.885 ;
        RECT 3.130 33.505 3.490 33.885 ;
        RECT 3.760 33.505 4.120 33.885 ;
        RECT 23.630 37.300 24.630 38.300 ;
        RECT 24.830 37.300 25.830 38.300 ;
        RECT 23.630 35.700 24.630 36.700 ;
        RECT 24.830 35.700 25.830 36.700 ;
        RECT 40.430 38.900 41.430 39.900 ;
        RECT 42.030 38.900 43.030 39.900 ;
        RECT 43.630 38.900 44.630 39.900 ;
        RECT 44.830 38.900 45.830 39.900 ;
        RECT 46.430 38.900 47.430 39.900 ;
        RECT 48.030 38.900 49.030 39.900 ;
        RECT 60.430 40.100 61.430 41.100 ;
        RECT 62.030 40.100 63.030 41.100 ;
        RECT 63.630 40.100 64.630 41.100 ;
        RECT 64.830 40.100 65.830 41.100 ;
        RECT 66.430 40.100 67.430 41.100 ;
        RECT 68.030 40.100 69.030 41.100 ;
        RECT 83.630 43.300 84.630 44.300 ;
        RECT 84.830 43.300 85.830 44.300 ;
        RECT 83.630 41.700 84.630 42.700 ;
        RECT 84.830 41.700 85.830 42.700 ;
        RECT 43.630 37.300 44.630 38.300 ;
        RECT 44.830 37.300 45.830 38.300 ;
        RECT 43.630 35.700 44.630 36.700 ;
        RECT 44.830 35.700 45.830 36.700 ;
        RECT 60.430 38.900 61.430 39.900 ;
        RECT 62.030 38.900 63.030 39.900 ;
        RECT 63.630 38.900 64.630 39.900 ;
        RECT 64.830 38.900 65.830 39.900 ;
        RECT 66.430 38.900 67.430 39.900 ;
        RECT 68.030 38.900 69.030 39.900 ;
        RECT 80.430 40.100 81.430 41.100 ;
        RECT 82.030 40.100 83.030 41.100 ;
        RECT 83.630 40.100 84.630 41.100 ;
        RECT 84.830 40.100 85.830 41.100 ;
        RECT 86.430 40.100 87.430 41.100 ;
        RECT 88.030 40.100 89.030 41.100 ;
        RECT 103.630 43.300 104.630 44.300 ;
        RECT 104.830 43.300 105.830 44.300 ;
        RECT 103.630 41.700 104.630 42.700 ;
        RECT 104.830 41.700 105.830 42.700 ;
        RECT 63.630 37.300 64.630 38.300 ;
        RECT 64.830 37.300 65.830 38.300 ;
        RECT 63.630 35.700 64.630 36.700 ;
        RECT 64.830 35.700 65.830 36.700 ;
        RECT 80.430 38.900 81.430 39.900 ;
        RECT 82.030 38.900 83.030 39.900 ;
        RECT 83.630 38.900 84.630 39.900 ;
        RECT 84.830 38.900 85.830 39.900 ;
        RECT 86.430 38.900 87.430 39.900 ;
        RECT 88.030 38.900 89.030 39.900 ;
        RECT 100.430 40.100 101.430 41.100 ;
        RECT 102.030 40.100 103.030 41.100 ;
        RECT 103.630 40.100 104.630 41.100 ;
        RECT 104.830 40.100 105.830 41.100 ;
        RECT 106.430 40.100 107.430 41.100 ;
        RECT 108.030 40.100 109.030 41.100 ;
        RECT 123.630 43.300 124.630 44.300 ;
        RECT 123.630 41.700 124.630 42.700 ;
        RECT 125.340 42.590 125.700 42.970 ;
        RECT 125.970 42.590 126.330 42.970 ;
        RECT 126.570 42.590 126.930 42.970 ;
        RECT 125.340 42.000 125.700 42.380 ;
        RECT 125.970 42.000 126.330 42.380 ;
        RECT 126.570 42.000 126.930 42.380 ;
        RECT 83.630 37.300 84.630 38.300 ;
        RECT 84.830 37.300 85.830 38.300 ;
        RECT 83.630 35.700 84.630 36.700 ;
        RECT 84.830 35.700 85.830 36.700 ;
        RECT 100.430 38.900 101.430 39.900 ;
        RECT 102.030 38.900 103.030 39.900 ;
        RECT 103.630 38.900 104.630 39.900 ;
        RECT 104.830 38.900 105.830 39.900 ;
        RECT 106.430 38.900 107.430 39.900 ;
        RECT 108.030 38.900 109.030 39.900 ;
        RECT 120.430 40.100 121.430 41.100 ;
        RECT 122.030 40.100 123.030 41.100 ;
        RECT 123.630 40.100 124.630 41.100 ;
        RECT 103.630 37.300 104.630 38.300 ;
        RECT 104.830 37.300 105.830 38.300 ;
        RECT 103.630 35.700 104.630 36.700 ;
        RECT 104.830 35.700 105.830 36.700 ;
        RECT 120.430 38.900 121.430 39.900 ;
        RECT 122.030 38.900 123.030 39.900 ;
        RECT 123.630 38.900 124.630 39.900 ;
        RECT 123.630 37.300 124.630 38.300 ;
        RECT 125.340 36.805 125.700 37.185 ;
        RECT 125.970 36.805 126.330 37.185 ;
        RECT 126.570 36.805 126.930 37.185 ;
        RECT 123.630 35.700 124.630 36.700 ;
        RECT 125.340 36.215 125.700 36.595 ;
        RECT 125.970 36.215 126.330 36.595 ;
        RECT 126.570 36.215 126.930 36.595 ;
        RECT 2.520 26.115 2.880 26.495 ;
        RECT 3.130 26.115 3.490 26.495 ;
        RECT 3.760 26.115 4.120 26.495 ;
        RECT 2.520 25.380 2.880 25.760 ;
        RECT 3.130 25.380 3.490 25.760 ;
        RECT 3.760 25.380 4.120 25.760 ;
        RECT 2.520 24.695 2.880 25.075 ;
        RECT 3.130 24.695 3.490 25.075 ;
        RECT 3.760 24.695 4.120 25.075 ;
        RECT 4.830 23.300 5.830 24.300 ;
        RECT 2.515 22.815 2.875 23.195 ;
        RECT 3.145 22.815 3.505 23.195 ;
        RECT 3.745 22.815 4.105 23.195 ;
        RECT 2.515 22.225 2.875 22.605 ;
        RECT 3.145 22.225 3.505 22.605 ;
        RECT 3.745 22.225 4.105 22.605 ;
        RECT 4.830 21.700 5.830 22.700 ;
        RECT 4.830 20.100 5.830 21.100 ;
        RECT 6.430 20.100 7.430 21.100 ;
        RECT 8.030 20.100 9.030 21.100 ;
        RECT 23.630 23.300 24.630 24.300 ;
        RECT 24.830 23.300 25.830 24.300 ;
        RECT 23.630 21.700 24.630 22.700 ;
        RECT 24.830 21.700 25.830 22.700 ;
        RECT 4.830 18.900 5.830 19.900 ;
        RECT 6.430 18.900 7.430 19.900 ;
        RECT 8.030 18.900 9.030 19.900 ;
        RECT 20.430 20.100 21.430 21.100 ;
        RECT 22.030 20.100 23.030 21.100 ;
        RECT 23.630 20.100 24.630 21.100 ;
        RECT 24.830 20.100 25.830 21.100 ;
        RECT 26.430 20.100 27.430 21.100 ;
        RECT 28.030 20.100 29.030 21.100 ;
        RECT 43.630 23.300 44.630 24.300 ;
        RECT 44.830 23.300 45.830 24.300 ;
        RECT 43.630 21.700 44.630 22.700 ;
        RECT 44.830 21.700 45.830 22.700 ;
        RECT 2.515 17.260 2.875 17.640 ;
        RECT 3.145 17.260 3.505 17.640 ;
        RECT 3.745 17.260 4.105 17.640 ;
        RECT 4.830 17.300 5.830 18.300 ;
        RECT 2.515 16.670 2.875 17.050 ;
        RECT 3.145 16.670 3.505 17.050 ;
        RECT 3.745 16.670 4.105 17.050 ;
        RECT 4.830 15.700 5.830 16.700 ;
        RECT 20.430 18.900 21.430 19.900 ;
        RECT 22.030 18.900 23.030 19.900 ;
        RECT 23.630 18.900 24.630 19.900 ;
        RECT 24.830 18.900 25.830 19.900 ;
        RECT 26.430 18.900 27.430 19.900 ;
        RECT 28.030 18.900 29.030 19.900 ;
        RECT 40.430 20.100 41.430 21.100 ;
        RECT 42.030 20.100 43.030 21.100 ;
        RECT 43.630 20.100 44.630 21.100 ;
        RECT 44.830 20.100 45.830 21.100 ;
        RECT 46.430 20.100 47.430 21.100 ;
        RECT 48.030 20.100 49.030 21.100 ;
        RECT 63.630 23.300 64.630 24.300 ;
        RECT 64.830 23.300 65.830 24.300 ;
        RECT 63.630 21.700 64.630 22.700 ;
        RECT 64.830 21.700 65.830 22.700 ;
        RECT 2.520 14.925 2.880 15.305 ;
        RECT 3.130 14.925 3.490 15.305 ;
        RECT 3.760 14.925 4.120 15.305 ;
        RECT 2.520 14.190 2.880 14.570 ;
        RECT 3.130 14.190 3.490 14.570 ;
        RECT 3.760 14.190 4.120 14.570 ;
        RECT 2.520 13.505 2.880 13.885 ;
        RECT 3.130 13.505 3.490 13.885 ;
        RECT 3.760 13.505 4.120 13.885 ;
        RECT 23.630 17.300 24.630 18.300 ;
        RECT 24.830 17.300 25.830 18.300 ;
        RECT 23.630 15.700 24.630 16.700 ;
        RECT 24.830 15.700 25.830 16.700 ;
        RECT 40.430 18.900 41.430 19.900 ;
        RECT 42.030 18.900 43.030 19.900 ;
        RECT 43.630 18.900 44.630 19.900 ;
        RECT 44.830 18.900 45.830 19.900 ;
        RECT 46.430 18.900 47.430 19.900 ;
        RECT 48.030 18.900 49.030 19.900 ;
        RECT 60.430 20.100 61.430 21.100 ;
        RECT 62.030 20.100 63.030 21.100 ;
        RECT 63.630 20.100 64.630 21.100 ;
        RECT 64.830 20.100 65.830 21.100 ;
        RECT 66.430 20.100 67.430 21.100 ;
        RECT 68.030 20.100 69.030 21.100 ;
        RECT 83.630 23.300 84.630 24.300 ;
        RECT 84.830 23.300 85.830 24.300 ;
        RECT 83.630 21.700 84.630 22.700 ;
        RECT 84.830 21.700 85.830 22.700 ;
        RECT 43.630 17.300 44.630 18.300 ;
        RECT 44.830 17.300 45.830 18.300 ;
        RECT 43.630 15.700 44.630 16.700 ;
        RECT 44.830 15.700 45.830 16.700 ;
        RECT 60.430 18.900 61.430 19.900 ;
        RECT 62.030 18.900 63.030 19.900 ;
        RECT 63.630 18.900 64.630 19.900 ;
        RECT 64.830 18.900 65.830 19.900 ;
        RECT 66.430 18.900 67.430 19.900 ;
        RECT 68.030 18.900 69.030 19.900 ;
        RECT 80.430 20.100 81.430 21.100 ;
        RECT 82.030 20.100 83.030 21.100 ;
        RECT 83.630 20.100 84.630 21.100 ;
        RECT 84.830 20.100 85.830 21.100 ;
        RECT 86.430 20.100 87.430 21.100 ;
        RECT 88.030 20.100 89.030 21.100 ;
        RECT 103.630 23.300 104.630 24.300 ;
        RECT 104.830 23.300 105.830 24.300 ;
        RECT 103.630 21.700 104.630 22.700 ;
        RECT 104.830 21.700 105.830 22.700 ;
        RECT 63.630 17.300 64.630 18.300 ;
        RECT 64.830 17.300 65.830 18.300 ;
        RECT 63.630 15.700 64.630 16.700 ;
        RECT 64.830 15.700 65.830 16.700 ;
        RECT 80.430 18.900 81.430 19.900 ;
        RECT 82.030 18.900 83.030 19.900 ;
        RECT 83.630 18.900 84.630 19.900 ;
        RECT 84.830 18.900 85.830 19.900 ;
        RECT 86.430 18.900 87.430 19.900 ;
        RECT 88.030 18.900 89.030 19.900 ;
        RECT 100.430 20.100 101.430 21.100 ;
        RECT 102.030 20.100 103.030 21.100 ;
        RECT 103.630 20.100 104.630 21.100 ;
        RECT 104.830 20.100 105.830 21.100 ;
        RECT 106.430 20.100 107.430 21.100 ;
        RECT 108.030 20.100 109.030 21.100 ;
        RECT 123.630 23.300 124.630 24.300 ;
        RECT 123.630 21.700 124.630 22.700 ;
        RECT 125.340 22.590 125.700 22.970 ;
        RECT 125.970 22.590 126.330 22.970 ;
        RECT 126.570 22.590 126.930 22.970 ;
        RECT 125.340 22.000 125.700 22.380 ;
        RECT 125.970 22.000 126.330 22.380 ;
        RECT 126.570 22.000 126.930 22.380 ;
        RECT 83.630 17.300 84.630 18.300 ;
        RECT 84.830 17.300 85.830 18.300 ;
        RECT 83.630 15.700 84.630 16.700 ;
        RECT 84.830 15.700 85.830 16.700 ;
        RECT 100.430 18.900 101.430 19.900 ;
        RECT 102.030 18.900 103.030 19.900 ;
        RECT 103.630 18.900 104.630 19.900 ;
        RECT 104.830 18.900 105.830 19.900 ;
        RECT 106.430 18.900 107.430 19.900 ;
        RECT 108.030 18.900 109.030 19.900 ;
        RECT 120.430 20.100 121.430 21.100 ;
        RECT 122.030 20.100 123.030 21.100 ;
        RECT 123.630 20.100 124.630 21.100 ;
        RECT 103.630 17.300 104.630 18.300 ;
        RECT 104.830 17.300 105.830 18.300 ;
        RECT 103.630 15.700 104.630 16.700 ;
        RECT 104.830 15.700 105.830 16.700 ;
        RECT 120.430 18.900 121.430 19.900 ;
        RECT 122.030 18.900 123.030 19.900 ;
        RECT 123.630 18.900 124.630 19.900 ;
        RECT 123.630 17.300 124.630 18.300 ;
        RECT 125.340 16.805 125.700 17.185 ;
        RECT 125.970 16.805 126.330 17.185 ;
        RECT 126.570 16.805 126.930 17.185 ;
        RECT 123.630 15.700 124.630 16.700 ;
        RECT 125.340 16.215 125.700 16.595 ;
        RECT 125.970 16.215 126.330 16.595 ;
        RECT 126.570 16.215 126.930 16.595 ;
        RECT 2.520 6.120 2.880 6.500 ;
        RECT 3.130 6.120 3.490 6.500 ;
        RECT 3.760 6.120 4.120 6.500 ;
        RECT 2.520 5.385 2.880 5.765 ;
        RECT 3.130 5.385 3.490 5.765 ;
        RECT 3.760 5.385 4.120 5.765 ;
        RECT 2.520 4.700 2.880 5.080 ;
        RECT 3.130 4.700 3.490 5.080 ;
        RECT 3.760 4.700 4.120 5.080 ;
        RECT 2.515 3.145 2.875 3.525 ;
        RECT 3.145 3.145 3.505 3.525 ;
        RECT 3.745 3.145 4.105 3.525 ;
        RECT 4.830 3.300 5.830 4.300 ;
        RECT 2.515 2.555 2.875 2.935 ;
        RECT 3.145 2.555 3.505 2.935 ;
        RECT 3.745 2.555 4.105 2.935 ;
        RECT 4.830 1.700 5.830 2.700 ;
        RECT 4.830 0.100 5.830 1.100 ;
        RECT 6.430 0.100 7.430 1.100 ;
        RECT 8.030 0.100 9.030 1.100 ;
        RECT 23.630 3.300 24.630 4.300 ;
        RECT 24.830 3.300 25.830 4.300 ;
        RECT 23.630 1.700 24.630 2.700 ;
        RECT 24.830 1.700 25.830 2.700 ;
        RECT 20.430 0.100 21.430 1.100 ;
        RECT 22.030 0.100 23.030 1.100 ;
        RECT 23.630 0.100 24.630 1.100 ;
        RECT 24.830 0.100 25.830 1.100 ;
        RECT 26.430 0.100 27.430 1.100 ;
        RECT 28.030 0.100 29.030 1.100 ;
        RECT 43.630 3.300 44.630 4.300 ;
        RECT 44.830 3.300 45.830 4.300 ;
        RECT 43.630 1.700 44.630 2.700 ;
        RECT 44.830 1.700 45.830 2.700 ;
        RECT 40.430 0.100 41.430 1.100 ;
        RECT 42.030 0.100 43.030 1.100 ;
        RECT 43.630 0.100 44.630 1.100 ;
        RECT 44.830 0.100 45.830 1.100 ;
        RECT 46.430 0.100 47.430 1.100 ;
        RECT 48.030 0.100 49.030 1.100 ;
        RECT 63.630 3.300 64.630 4.300 ;
        RECT 64.830 3.300 65.830 4.300 ;
        RECT 63.630 1.700 64.630 2.700 ;
        RECT 64.830 1.700 65.830 2.700 ;
        RECT 60.430 0.100 61.430 1.100 ;
        RECT 62.030 0.100 63.030 1.100 ;
        RECT 63.630 0.100 64.630 1.100 ;
        RECT 64.830 0.100 65.830 1.100 ;
        RECT 66.430 0.100 67.430 1.100 ;
        RECT 68.030 0.100 69.030 1.100 ;
        RECT 83.630 3.300 84.630 4.300 ;
        RECT 84.830 3.300 85.830 4.300 ;
        RECT 83.630 1.700 84.630 2.700 ;
        RECT 84.830 1.700 85.830 2.700 ;
        RECT 80.430 0.100 81.430 1.100 ;
        RECT 82.030 0.100 83.030 1.100 ;
        RECT 83.630 0.100 84.630 1.100 ;
        RECT 84.830 0.100 85.830 1.100 ;
        RECT 86.430 0.100 87.430 1.100 ;
        RECT 88.030 0.100 89.030 1.100 ;
        RECT 103.630 3.300 104.630 4.300 ;
        RECT 104.830 3.300 105.830 4.300 ;
        RECT 103.630 1.700 104.630 2.700 ;
        RECT 104.830 1.700 105.830 2.700 ;
        RECT 100.430 0.100 101.430 1.100 ;
        RECT 102.030 0.100 103.030 1.100 ;
        RECT 103.630 0.100 104.630 1.100 ;
        RECT 104.830 0.100 105.830 1.100 ;
        RECT 106.430 0.100 107.430 1.100 ;
        RECT 108.030 0.100 109.030 1.100 ;
        RECT 123.630 3.300 124.630 4.300 ;
        RECT 123.630 1.700 124.630 2.700 ;
        RECT 125.340 2.590 125.700 2.970 ;
        RECT 125.970 2.590 126.330 2.970 ;
        RECT 126.570 2.590 126.930 2.970 ;
        RECT 125.340 2.000 125.700 2.380 ;
        RECT 125.970 2.000 126.330 2.380 ;
        RECT 126.570 2.000 126.930 2.380 ;
        RECT 120.430 0.100 121.430 1.100 ;
        RECT 122.030 0.100 123.030 1.100 ;
        RECT 123.630 0.100 124.630 1.100 ;
      LAYER met2 ;
        RECT 4.730 338.800 9.130 340.000 ;
        RECT 20.330 338.800 29.130 340.000 ;
        RECT 40.330 338.800 49.130 340.000 ;
        RECT 60.330 338.800 69.130 340.000 ;
        RECT 80.330 338.800 89.130 340.000 ;
        RECT 100.330 338.800 109.130 340.000 ;
        RECT 120.330 338.800 124.730 340.000 ;
        RECT 4.730 337.850 5.940 338.800 ;
        RECT 4.730 337.700 9.880 337.850 ;
        RECT 2.315 336.110 4.320 337.385 ;
        RECT 4.730 337.250 6.330 337.700 ;
        RECT 4.730 337.100 9.880 337.250 ;
        RECT 4.730 336.650 6.330 337.100 ;
        RECT 4.730 336.500 9.880 336.650 ;
        RECT 4.730 336.050 6.330 336.500 ;
        RECT 4.730 335.900 9.880 336.050 ;
        RECT 4.730 335.600 6.330 335.900 ;
        RECT 2.315 333.250 4.315 335.545 ;
        RECT 5.930 335.450 6.330 335.600 ;
        RECT 5.930 335.300 9.880 335.450 ;
        RECT 5.930 334.850 6.330 335.300 ;
        RECT 5.930 334.700 9.880 334.850 ;
        RECT 5.930 334.250 6.330 334.700 ;
        RECT 5.930 334.100 9.880 334.250 ;
        RECT 5.930 333.650 6.330 334.100 ;
        RECT 5.930 333.500 9.880 333.650 ;
        RECT 5.930 333.050 6.330 333.500 ;
        RECT 5.930 332.900 9.880 333.050 ;
        RECT 5.930 332.450 6.330 332.900 ;
        RECT 5.930 332.300 9.880 332.450 ;
        RECT 5.930 331.850 6.330 332.300 ;
        RECT 5.930 331.700 9.880 331.850 ;
        RECT 5.930 331.250 6.330 331.700 ;
        RECT 5.930 331.100 9.880 331.250 ;
        RECT 5.930 330.650 6.330 331.100 ;
        RECT 5.930 330.500 9.880 330.650 ;
        RECT 5.930 330.200 6.330 330.500 ;
        RECT 10.480 330.200 10.630 338.400 ;
        RECT 11.080 330.200 11.230 338.400 ;
        RECT 11.680 330.200 11.830 338.400 ;
        RECT 12.280 330.200 12.430 338.400 ;
        RECT 12.880 330.200 13.030 338.400 ;
        RECT 13.480 330.200 13.630 338.400 ;
        RECT 14.080 330.200 14.230 338.400 ;
        RECT 5.930 329.800 14.230 330.200 ;
        RECT 5.930 329.500 6.330 329.800 ;
        RECT 5.930 329.350 9.880 329.500 ;
        RECT 5.930 328.900 6.330 329.350 ;
        RECT 5.930 328.750 9.880 328.900 ;
        RECT 5.930 328.300 6.330 328.750 ;
        RECT 5.930 328.150 9.880 328.300 ;
        RECT 5.930 327.700 6.330 328.150 ;
        RECT 5.930 327.550 9.880 327.700 ;
        RECT 5.930 327.100 6.330 327.550 ;
        RECT 5.930 326.950 9.880 327.100 ;
        RECT 2.315 324.450 4.315 326.745 ;
        RECT 5.930 326.500 6.330 326.950 ;
        RECT 5.930 326.350 9.880 326.500 ;
        RECT 5.930 325.900 6.330 326.350 ;
        RECT 5.930 325.750 9.880 325.900 ;
        RECT 5.930 325.300 6.330 325.750 ;
        RECT 5.930 325.150 9.880 325.300 ;
        RECT 5.930 324.700 6.330 325.150 ;
        RECT 5.930 324.550 9.880 324.700 ;
        RECT 5.930 324.400 6.330 324.550 ;
        RECT 4.730 324.100 6.330 324.400 ;
        RECT 2.315 322.745 4.320 324.020 ;
        RECT 4.730 323.950 9.880 324.100 ;
        RECT 4.730 323.500 6.330 323.950 ;
        RECT 4.730 323.350 9.880 323.500 ;
        RECT 4.730 322.900 6.330 323.350 ;
        RECT 4.730 322.750 9.880 322.900 ;
        RECT 4.730 322.300 6.330 322.750 ;
        RECT 4.730 322.150 9.880 322.300 ;
        RECT 4.730 321.200 5.930 322.150 ;
        RECT 10.480 321.600 10.630 329.800 ;
        RECT 11.080 321.600 11.230 329.800 ;
        RECT 11.680 321.600 11.830 329.800 ;
        RECT 12.280 321.600 12.430 329.800 ;
        RECT 12.880 321.600 13.030 329.800 ;
        RECT 13.480 321.600 13.630 329.800 ;
        RECT 14.080 321.600 14.230 329.800 ;
        RECT 15.230 330.200 15.380 338.400 ;
        RECT 15.830 330.200 15.980 338.400 ;
        RECT 16.430 330.200 16.580 338.400 ;
        RECT 17.030 330.200 17.180 338.400 ;
        RECT 17.630 330.200 17.780 338.400 ;
        RECT 18.230 330.200 18.380 338.400 ;
        RECT 18.830 330.200 18.980 338.400 ;
        RECT 23.530 337.850 25.940 338.800 ;
        RECT 19.580 337.700 29.880 337.850 ;
        RECT 23.130 337.250 26.330 337.700 ;
        RECT 19.580 337.100 29.880 337.250 ;
        RECT 23.130 336.650 26.330 337.100 ;
        RECT 19.580 336.500 29.880 336.650 ;
        RECT 23.130 336.050 26.330 336.500 ;
        RECT 19.580 335.900 29.880 336.050 ;
        RECT 23.130 335.600 26.330 335.900 ;
        RECT 23.130 335.450 23.530 335.600 ;
        RECT 19.580 335.300 23.530 335.450 ;
        RECT 23.130 334.850 23.530 335.300 ;
        RECT 19.580 334.700 23.530 334.850 ;
        RECT 23.130 334.250 23.530 334.700 ;
        RECT 19.580 334.100 23.530 334.250 ;
        RECT 23.130 333.650 23.530 334.100 ;
        RECT 19.580 333.500 23.530 333.650 ;
        RECT 23.130 333.050 23.530 333.500 ;
        RECT 19.580 332.900 23.530 333.050 ;
        RECT 23.130 332.450 23.530 332.900 ;
        RECT 19.580 332.300 23.530 332.450 ;
        RECT 23.130 331.850 23.530 332.300 ;
        RECT 19.580 331.700 23.530 331.850 ;
        RECT 23.130 331.250 23.530 331.700 ;
        RECT 19.580 331.100 23.530 331.250 ;
        RECT 23.130 330.650 23.530 331.100 ;
        RECT 19.580 330.500 23.530 330.650 ;
        RECT 23.130 330.200 23.530 330.500 ;
        RECT 15.230 329.800 23.530 330.200 ;
        RECT 15.230 321.600 15.380 329.800 ;
        RECT 15.830 321.600 15.980 329.800 ;
        RECT 16.430 321.600 16.580 329.800 ;
        RECT 17.030 321.600 17.180 329.800 ;
        RECT 17.630 321.600 17.780 329.800 ;
        RECT 18.230 321.600 18.380 329.800 ;
        RECT 18.830 321.600 18.980 329.800 ;
        RECT 23.130 329.500 23.530 329.800 ;
        RECT 19.580 329.350 23.530 329.500 ;
        RECT 23.130 328.900 23.530 329.350 ;
        RECT 19.580 328.750 23.530 328.900 ;
        RECT 23.130 328.300 23.530 328.750 ;
        RECT 19.580 328.150 23.530 328.300 ;
        RECT 23.130 327.700 23.530 328.150 ;
        RECT 19.580 327.550 23.530 327.700 ;
        RECT 23.130 327.100 23.530 327.550 ;
        RECT 19.580 326.950 23.530 327.100 ;
        RECT 23.130 326.500 23.530 326.950 ;
        RECT 19.580 326.350 23.530 326.500 ;
        RECT 23.130 325.900 23.530 326.350 ;
        RECT 19.580 325.750 23.530 325.900 ;
        RECT 23.130 325.300 23.530 325.750 ;
        RECT 19.580 325.150 23.530 325.300 ;
        RECT 23.130 324.700 23.530 325.150 ;
        RECT 19.580 324.550 23.530 324.700 ;
        RECT 23.130 324.400 23.530 324.550 ;
        RECT 25.930 335.450 26.330 335.600 ;
        RECT 25.930 335.300 29.880 335.450 ;
        RECT 25.930 334.850 26.330 335.300 ;
        RECT 25.930 334.700 29.880 334.850 ;
        RECT 25.930 334.250 26.330 334.700 ;
        RECT 25.930 334.100 29.880 334.250 ;
        RECT 25.930 333.650 26.330 334.100 ;
        RECT 25.930 333.500 29.880 333.650 ;
        RECT 25.930 333.050 26.330 333.500 ;
        RECT 25.930 332.900 29.880 333.050 ;
        RECT 25.930 332.450 26.330 332.900 ;
        RECT 25.930 332.300 29.880 332.450 ;
        RECT 25.930 331.850 26.330 332.300 ;
        RECT 25.930 331.700 29.880 331.850 ;
        RECT 25.930 331.250 26.330 331.700 ;
        RECT 25.930 331.100 29.880 331.250 ;
        RECT 25.930 330.650 26.330 331.100 ;
        RECT 25.930 330.500 29.880 330.650 ;
        RECT 25.930 330.200 26.330 330.500 ;
        RECT 30.480 330.200 30.630 338.400 ;
        RECT 31.080 330.200 31.230 338.400 ;
        RECT 31.680 330.200 31.830 338.400 ;
        RECT 32.280 330.200 32.430 338.400 ;
        RECT 32.880 330.200 33.030 338.400 ;
        RECT 33.480 330.200 33.630 338.400 ;
        RECT 34.080 330.200 34.230 338.400 ;
        RECT 25.930 329.800 34.230 330.200 ;
        RECT 25.930 329.500 26.330 329.800 ;
        RECT 25.930 329.350 29.880 329.500 ;
        RECT 25.930 328.900 26.330 329.350 ;
        RECT 25.930 328.750 29.880 328.900 ;
        RECT 25.930 328.300 26.330 328.750 ;
        RECT 25.930 328.150 29.880 328.300 ;
        RECT 25.930 327.700 26.330 328.150 ;
        RECT 25.930 327.550 29.880 327.700 ;
        RECT 25.930 327.100 26.330 327.550 ;
        RECT 25.930 326.950 29.880 327.100 ;
        RECT 25.930 326.500 26.330 326.950 ;
        RECT 25.930 326.350 29.880 326.500 ;
        RECT 25.930 325.900 26.330 326.350 ;
        RECT 25.930 325.750 29.880 325.900 ;
        RECT 25.930 325.300 26.330 325.750 ;
        RECT 25.930 325.150 29.880 325.300 ;
        RECT 25.930 324.700 26.330 325.150 ;
        RECT 25.930 324.550 29.880 324.700 ;
        RECT 25.930 324.400 26.330 324.550 ;
        RECT 23.130 324.100 26.330 324.400 ;
        RECT 19.580 323.950 29.880 324.100 ;
        RECT 23.130 323.500 26.330 323.950 ;
        RECT 19.580 323.350 29.880 323.500 ;
        RECT 23.130 322.900 26.330 323.350 ;
        RECT 19.580 322.750 29.880 322.900 ;
        RECT 23.130 322.300 26.330 322.750 ;
        RECT 19.580 322.150 29.880 322.300 ;
        RECT 23.530 321.200 25.930 322.150 ;
        RECT 30.480 321.600 30.630 329.800 ;
        RECT 31.080 321.600 31.230 329.800 ;
        RECT 31.680 321.600 31.830 329.800 ;
        RECT 32.280 321.600 32.430 329.800 ;
        RECT 32.880 321.600 33.030 329.800 ;
        RECT 33.480 321.600 33.630 329.800 ;
        RECT 34.080 321.600 34.230 329.800 ;
        RECT 35.230 330.200 35.380 338.400 ;
        RECT 35.830 330.200 35.980 338.400 ;
        RECT 36.430 330.200 36.580 338.400 ;
        RECT 37.030 330.200 37.180 338.400 ;
        RECT 37.630 330.200 37.780 338.400 ;
        RECT 38.230 330.200 38.380 338.400 ;
        RECT 38.830 330.200 38.980 338.400 ;
        RECT 43.530 337.850 45.940 338.800 ;
        RECT 39.580 337.700 49.880 337.850 ;
        RECT 43.130 337.250 46.330 337.700 ;
        RECT 39.580 337.100 49.880 337.250 ;
        RECT 43.130 336.650 46.330 337.100 ;
        RECT 39.580 336.500 49.880 336.650 ;
        RECT 43.130 336.050 46.330 336.500 ;
        RECT 39.580 335.900 49.880 336.050 ;
        RECT 43.130 335.600 46.330 335.900 ;
        RECT 43.130 335.450 43.530 335.600 ;
        RECT 39.580 335.300 43.530 335.450 ;
        RECT 43.130 334.850 43.530 335.300 ;
        RECT 39.580 334.700 43.530 334.850 ;
        RECT 43.130 334.250 43.530 334.700 ;
        RECT 39.580 334.100 43.530 334.250 ;
        RECT 43.130 333.650 43.530 334.100 ;
        RECT 39.580 333.500 43.530 333.650 ;
        RECT 43.130 333.050 43.530 333.500 ;
        RECT 39.580 332.900 43.530 333.050 ;
        RECT 43.130 332.450 43.530 332.900 ;
        RECT 39.580 332.300 43.530 332.450 ;
        RECT 43.130 331.850 43.530 332.300 ;
        RECT 39.580 331.700 43.530 331.850 ;
        RECT 43.130 331.250 43.530 331.700 ;
        RECT 39.580 331.100 43.530 331.250 ;
        RECT 43.130 330.650 43.530 331.100 ;
        RECT 39.580 330.500 43.530 330.650 ;
        RECT 43.130 330.200 43.530 330.500 ;
        RECT 35.230 329.800 43.530 330.200 ;
        RECT 35.230 321.600 35.380 329.800 ;
        RECT 35.830 321.600 35.980 329.800 ;
        RECT 36.430 321.600 36.580 329.800 ;
        RECT 37.030 321.600 37.180 329.800 ;
        RECT 37.630 321.600 37.780 329.800 ;
        RECT 38.230 321.600 38.380 329.800 ;
        RECT 38.830 321.600 38.980 329.800 ;
        RECT 43.130 329.500 43.530 329.800 ;
        RECT 39.580 329.350 43.530 329.500 ;
        RECT 43.130 328.900 43.530 329.350 ;
        RECT 39.580 328.750 43.530 328.900 ;
        RECT 43.130 328.300 43.530 328.750 ;
        RECT 39.580 328.150 43.530 328.300 ;
        RECT 43.130 327.700 43.530 328.150 ;
        RECT 39.580 327.550 43.530 327.700 ;
        RECT 43.130 327.100 43.530 327.550 ;
        RECT 39.580 326.950 43.530 327.100 ;
        RECT 43.130 326.500 43.530 326.950 ;
        RECT 39.580 326.350 43.530 326.500 ;
        RECT 43.130 325.900 43.530 326.350 ;
        RECT 39.580 325.750 43.530 325.900 ;
        RECT 43.130 325.300 43.530 325.750 ;
        RECT 39.580 325.150 43.530 325.300 ;
        RECT 43.130 324.700 43.530 325.150 ;
        RECT 39.580 324.550 43.530 324.700 ;
        RECT 43.130 324.400 43.530 324.550 ;
        RECT 45.930 335.450 46.330 335.600 ;
        RECT 45.930 335.300 49.880 335.450 ;
        RECT 45.930 334.850 46.330 335.300 ;
        RECT 45.930 334.700 49.880 334.850 ;
        RECT 45.930 334.250 46.330 334.700 ;
        RECT 45.930 334.100 49.880 334.250 ;
        RECT 45.930 333.650 46.330 334.100 ;
        RECT 45.930 333.500 49.880 333.650 ;
        RECT 45.930 333.050 46.330 333.500 ;
        RECT 45.930 332.900 49.880 333.050 ;
        RECT 45.930 332.450 46.330 332.900 ;
        RECT 45.930 332.300 49.880 332.450 ;
        RECT 45.930 331.850 46.330 332.300 ;
        RECT 45.930 331.700 49.880 331.850 ;
        RECT 45.930 331.250 46.330 331.700 ;
        RECT 45.930 331.100 49.880 331.250 ;
        RECT 45.930 330.650 46.330 331.100 ;
        RECT 45.930 330.500 49.880 330.650 ;
        RECT 45.930 330.200 46.330 330.500 ;
        RECT 50.480 330.200 50.630 338.400 ;
        RECT 51.080 330.200 51.230 338.400 ;
        RECT 51.680 330.200 51.830 338.400 ;
        RECT 52.280 330.200 52.430 338.400 ;
        RECT 52.880 330.200 53.030 338.400 ;
        RECT 53.480 330.200 53.630 338.400 ;
        RECT 54.080 330.200 54.230 338.400 ;
        RECT 45.930 329.800 54.230 330.200 ;
        RECT 45.930 329.500 46.330 329.800 ;
        RECT 45.930 329.350 49.880 329.500 ;
        RECT 45.930 328.900 46.330 329.350 ;
        RECT 45.930 328.750 49.880 328.900 ;
        RECT 45.930 328.300 46.330 328.750 ;
        RECT 45.930 328.150 49.880 328.300 ;
        RECT 45.930 327.700 46.330 328.150 ;
        RECT 45.930 327.550 49.880 327.700 ;
        RECT 45.930 327.100 46.330 327.550 ;
        RECT 45.930 326.950 49.880 327.100 ;
        RECT 45.930 326.500 46.330 326.950 ;
        RECT 45.930 326.350 49.880 326.500 ;
        RECT 45.930 325.900 46.330 326.350 ;
        RECT 45.930 325.750 49.880 325.900 ;
        RECT 45.930 325.300 46.330 325.750 ;
        RECT 45.930 325.150 49.880 325.300 ;
        RECT 45.930 324.700 46.330 325.150 ;
        RECT 45.930 324.550 49.880 324.700 ;
        RECT 45.930 324.400 46.330 324.550 ;
        RECT 43.130 324.100 46.330 324.400 ;
        RECT 39.580 323.950 49.880 324.100 ;
        RECT 43.130 323.500 46.330 323.950 ;
        RECT 39.580 323.350 49.880 323.500 ;
        RECT 43.130 322.900 46.330 323.350 ;
        RECT 39.580 322.750 49.880 322.900 ;
        RECT 43.130 322.300 46.330 322.750 ;
        RECT 39.580 322.150 49.880 322.300 ;
        RECT 43.530 321.200 45.930 322.150 ;
        RECT 50.480 321.600 50.630 329.800 ;
        RECT 51.080 321.600 51.230 329.800 ;
        RECT 51.680 321.600 51.830 329.800 ;
        RECT 52.280 321.600 52.430 329.800 ;
        RECT 52.880 321.600 53.030 329.800 ;
        RECT 53.480 321.600 53.630 329.800 ;
        RECT 54.080 321.600 54.230 329.800 ;
        RECT 55.230 330.200 55.380 338.400 ;
        RECT 55.830 330.200 55.980 338.400 ;
        RECT 56.430 330.200 56.580 338.400 ;
        RECT 57.030 330.200 57.180 338.400 ;
        RECT 57.630 330.200 57.780 338.400 ;
        RECT 58.230 330.200 58.380 338.400 ;
        RECT 58.830 330.200 58.980 338.400 ;
        RECT 63.530 337.850 65.940 338.800 ;
        RECT 59.580 337.700 69.880 337.850 ;
        RECT 63.130 337.250 66.330 337.700 ;
        RECT 59.580 337.100 69.880 337.250 ;
        RECT 63.130 336.650 66.330 337.100 ;
        RECT 59.580 336.500 69.880 336.650 ;
        RECT 63.130 336.050 66.330 336.500 ;
        RECT 59.580 335.900 69.880 336.050 ;
        RECT 63.130 335.600 66.330 335.900 ;
        RECT 63.130 335.450 63.530 335.600 ;
        RECT 59.580 335.300 63.530 335.450 ;
        RECT 63.130 334.850 63.530 335.300 ;
        RECT 59.580 334.700 63.530 334.850 ;
        RECT 63.130 334.250 63.530 334.700 ;
        RECT 59.580 334.100 63.530 334.250 ;
        RECT 63.130 333.650 63.530 334.100 ;
        RECT 59.580 333.500 63.530 333.650 ;
        RECT 63.130 333.050 63.530 333.500 ;
        RECT 59.580 332.900 63.530 333.050 ;
        RECT 63.130 332.450 63.530 332.900 ;
        RECT 59.580 332.300 63.530 332.450 ;
        RECT 63.130 331.850 63.530 332.300 ;
        RECT 59.580 331.700 63.530 331.850 ;
        RECT 63.130 331.250 63.530 331.700 ;
        RECT 59.580 331.100 63.530 331.250 ;
        RECT 63.130 330.650 63.530 331.100 ;
        RECT 59.580 330.500 63.530 330.650 ;
        RECT 63.130 330.200 63.530 330.500 ;
        RECT 55.230 329.800 63.530 330.200 ;
        RECT 55.230 321.600 55.380 329.800 ;
        RECT 55.830 321.600 55.980 329.800 ;
        RECT 56.430 321.600 56.580 329.800 ;
        RECT 57.030 321.600 57.180 329.800 ;
        RECT 57.630 321.600 57.780 329.800 ;
        RECT 58.230 321.600 58.380 329.800 ;
        RECT 58.830 321.600 58.980 329.800 ;
        RECT 63.130 329.500 63.530 329.800 ;
        RECT 59.580 329.350 63.530 329.500 ;
        RECT 63.130 328.900 63.530 329.350 ;
        RECT 59.580 328.750 63.530 328.900 ;
        RECT 63.130 328.300 63.530 328.750 ;
        RECT 59.580 328.150 63.530 328.300 ;
        RECT 63.130 327.700 63.530 328.150 ;
        RECT 59.580 327.550 63.530 327.700 ;
        RECT 63.130 327.100 63.530 327.550 ;
        RECT 59.580 326.950 63.530 327.100 ;
        RECT 63.130 326.500 63.530 326.950 ;
        RECT 59.580 326.350 63.530 326.500 ;
        RECT 63.130 325.900 63.530 326.350 ;
        RECT 59.580 325.750 63.530 325.900 ;
        RECT 63.130 325.300 63.530 325.750 ;
        RECT 59.580 325.150 63.530 325.300 ;
        RECT 63.130 324.700 63.530 325.150 ;
        RECT 59.580 324.550 63.530 324.700 ;
        RECT 63.130 324.400 63.530 324.550 ;
        RECT 65.930 335.450 66.330 335.600 ;
        RECT 65.930 335.300 69.880 335.450 ;
        RECT 65.930 334.850 66.330 335.300 ;
        RECT 65.930 334.700 69.880 334.850 ;
        RECT 65.930 334.250 66.330 334.700 ;
        RECT 65.930 334.100 69.880 334.250 ;
        RECT 65.930 333.650 66.330 334.100 ;
        RECT 65.930 333.500 69.880 333.650 ;
        RECT 65.930 333.050 66.330 333.500 ;
        RECT 65.930 332.900 69.880 333.050 ;
        RECT 65.930 332.450 66.330 332.900 ;
        RECT 65.930 332.300 69.880 332.450 ;
        RECT 65.930 331.850 66.330 332.300 ;
        RECT 65.930 331.700 69.880 331.850 ;
        RECT 65.930 331.250 66.330 331.700 ;
        RECT 65.930 331.100 69.880 331.250 ;
        RECT 65.930 330.650 66.330 331.100 ;
        RECT 65.930 330.500 69.880 330.650 ;
        RECT 65.930 330.200 66.330 330.500 ;
        RECT 70.480 330.200 70.630 338.400 ;
        RECT 71.080 330.200 71.230 338.400 ;
        RECT 71.680 330.200 71.830 338.400 ;
        RECT 72.280 330.200 72.430 338.400 ;
        RECT 72.880 330.200 73.030 338.400 ;
        RECT 73.480 330.200 73.630 338.400 ;
        RECT 74.080 330.200 74.230 338.400 ;
        RECT 65.930 329.800 74.230 330.200 ;
        RECT 65.930 329.500 66.330 329.800 ;
        RECT 65.930 329.350 69.880 329.500 ;
        RECT 65.930 328.900 66.330 329.350 ;
        RECT 65.930 328.750 69.880 328.900 ;
        RECT 65.930 328.300 66.330 328.750 ;
        RECT 65.930 328.150 69.880 328.300 ;
        RECT 65.930 327.700 66.330 328.150 ;
        RECT 65.930 327.550 69.880 327.700 ;
        RECT 65.930 327.100 66.330 327.550 ;
        RECT 65.930 326.950 69.880 327.100 ;
        RECT 65.930 326.500 66.330 326.950 ;
        RECT 65.930 326.350 69.880 326.500 ;
        RECT 65.930 325.900 66.330 326.350 ;
        RECT 65.930 325.750 69.880 325.900 ;
        RECT 65.930 325.300 66.330 325.750 ;
        RECT 65.930 325.150 69.880 325.300 ;
        RECT 65.930 324.700 66.330 325.150 ;
        RECT 65.930 324.550 69.880 324.700 ;
        RECT 65.930 324.400 66.330 324.550 ;
        RECT 63.130 324.100 66.330 324.400 ;
        RECT 59.580 323.950 69.880 324.100 ;
        RECT 63.130 323.500 66.330 323.950 ;
        RECT 59.580 323.350 69.880 323.500 ;
        RECT 63.130 322.900 66.330 323.350 ;
        RECT 59.580 322.750 69.880 322.900 ;
        RECT 63.130 322.300 66.330 322.750 ;
        RECT 59.580 322.150 69.880 322.300 ;
        RECT 63.530 321.200 65.930 322.150 ;
        RECT 70.480 321.600 70.630 329.800 ;
        RECT 71.080 321.600 71.230 329.800 ;
        RECT 71.680 321.600 71.830 329.800 ;
        RECT 72.280 321.600 72.430 329.800 ;
        RECT 72.880 321.600 73.030 329.800 ;
        RECT 73.480 321.600 73.630 329.800 ;
        RECT 74.080 321.600 74.230 329.800 ;
        RECT 75.230 330.200 75.380 338.400 ;
        RECT 75.830 330.200 75.980 338.400 ;
        RECT 76.430 330.200 76.580 338.400 ;
        RECT 77.030 330.200 77.180 338.400 ;
        RECT 77.630 330.200 77.780 338.400 ;
        RECT 78.230 330.200 78.380 338.400 ;
        RECT 78.830 330.200 78.980 338.400 ;
        RECT 83.530 337.850 85.940 338.800 ;
        RECT 79.580 337.700 89.880 337.850 ;
        RECT 83.130 337.250 86.330 337.700 ;
        RECT 79.580 337.100 89.880 337.250 ;
        RECT 83.130 336.650 86.330 337.100 ;
        RECT 79.580 336.500 89.880 336.650 ;
        RECT 83.130 336.050 86.330 336.500 ;
        RECT 79.580 335.900 89.880 336.050 ;
        RECT 83.130 335.600 86.330 335.900 ;
        RECT 83.130 335.450 83.530 335.600 ;
        RECT 79.580 335.300 83.530 335.450 ;
        RECT 83.130 334.850 83.530 335.300 ;
        RECT 79.580 334.700 83.530 334.850 ;
        RECT 83.130 334.250 83.530 334.700 ;
        RECT 79.580 334.100 83.530 334.250 ;
        RECT 83.130 333.650 83.530 334.100 ;
        RECT 79.580 333.500 83.530 333.650 ;
        RECT 83.130 333.050 83.530 333.500 ;
        RECT 79.580 332.900 83.530 333.050 ;
        RECT 83.130 332.450 83.530 332.900 ;
        RECT 79.580 332.300 83.530 332.450 ;
        RECT 83.130 331.850 83.530 332.300 ;
        RECT 79.580 331.700 83.530 331.850 ;
        RECT 83.130 331.250 83.530 331.700 ;
        RECT 79.580 331.100 83.530 331.250 ;
        RECT 83.130 330.650 83.530 331.100 ;
        RECT 79.580 330.500 83.530 330.650 ;
        RECT 83.130 330.200 83.530 330.500 ;
        RECT 75.230 329.800 83.530 330.200 ;
        RECT 75.230 321.600 75.380 329.800 ;
        RECT 75.830 321.600 75.980 329.800 ;
        RECT 76.430 321.600 76.580 329.800 ;
        RECT 77.030 321.600 77.180 329.800 ;
        RECT 77.630 321.600 77.780 329.800 ;
        RECT 78.230 321.600 78.380 329.800 ;
        RECT 78.830 321.600 78.980 329.800 ;
        RECT 83.130 329.500 83.530 329.800 ;
        RECT 79.580 329.350 83.530 329.500 ;
        RECT 83.130 328.900 83.530 329.350 ;
        RECT 79.580 328.750 83.530 328.900 ;
        RECT 83.130 328.300 83.530 328.750 ;
        RECT 79.580 328.150 83.530 328.300 ;
        RECT 83.130 327.700 83.530 328.150 ;
        RECT 79.580 327.550 83.530 327.700 ;
        RECT 83.130 327.100 83.530 327.550 ;
        RECT 79.580 326.950 83.530 327.100 ;
        RECT 83.130 326.500 83.530 326.950 ;
        RECT 79.580 326.350 83.530 326.500 ;
        RECT 83.130 325.900 83.530 326.350 ;
        RECT 79.580 325.750 83.530 325.900 ;
        RECT 83.130 325.300 83.530 325.750 ;
        RECT 79.580 325.150 83.530 325.300 ;
        RECT 83.130 324.700 83.530 325.150 ;
        RECT 79.580 324.550 83.530 324.700 ;
        RECT 83.130 324.400 83.530 324.550 ;
        RECT 85.930 335.450 86.330 335.600 ;
        RECT 85.930 335.300 89.880 335.450 ;
        RECT 85.930 334.850 86.330 335.300 ;
        RECT 85.930 334.700 89.880 334.850 ;
        RECT 85.930 334.250 86.330 334.700 ;
        RECT 85.930 334.100 89.880 334.250 ;
        RECT 85.930 333.650 86.330 334.100 ;
        RECT 85.930 333.500 89.880 333.650 ;
        RECT 85.930 333.050 86.330 333.500 ;
        RECT 85.930 332.900 89.880 333.050 ;
        RECT 85.930 332.450 86.330 332.900 ;
        RECT 85.930 332.300 89.880 332.450 ;
        RECT 85.930 331.850 86.330 332.300 ;
        RECT 85.930 331.700 89.880 331.850 ;
        RECT 85.930 331.250 86.330 331.700 ;
        RECT 85.930 331.100 89.880 331.250 ;
        RECT 85.930 330.650 86.330 331.100 ;
        RECT 85.930 330.500 89.880 330.650 ;
        RECT 85.930 330.200 86.330 330.500 ;
        RECT 90.480 330.200 90.630 338.400 ;
        RECT 91.080 330.200 91.230 338.400 ;
        RECT 91.680 330.200 91.830 338.400 ;
        RECT 92.280 330.200 92.430 338.400 ;
        RECT 92.880 330.200 93.030 338.400 ;
        RECT 93.480 330.200 93.630 338.400 ;
        RECT 94.080 330.200 94.230 338.400 ;
        RECT 85.930 329.800 94.230 330.200 ;
        RECT 85.930 329.500 86.330 329.800 ;
        RECT 85.930 329.350 89.880 329.500 ;
        RECT 85.930 328.900 86.330 329.350 ;
        RECT 85.930 328.750 89.880 328.900 ;
        RECT 85.930 328.300 86.330 328.750 ;
        RECT 85.930 328.150 89.880 328.300 ;
        RECT 85.930 327.700 86.330 328.150 ;
        RECT 85.930 327.550 89.880 327.700 ;
        RECT 85.930 327.100 86.330 327.550 ;
        RECT 85.930 326.950 89.880 327.100 ;
        RECT 85.930 326.500 86.330 326.950 ;
        RECT 85.930 326.350 89.880 326.500 ;
        RECT 85.930 325.900 86.330 326.350 ;
        RECT 85.930 325.750 89.880 325.900 ;
        RECT 85.930 325.300 86.330 325.750 ;
        RECT 85.930 325.150 89.880 325.300 ;
        RECT 85.930 324.700 86.330 325.150 ;
        RECT 85.930 324.550 89.880 324.700 ;
        RECT 85.930 324.400 86.330 324.550 ;
        RECT 83.130 324.100 86.330 324.400 ;
        RECT 79.580 323.950 89.880 324.100 ;
        RECT 83.130 323.500 86.330 323.950 ;
        RECT 79.580 323.350 89.880 323.500 ;
        RECT 83.130 322.900 86.330 323.350 ;
        RECT 79.580 322.750 89.880 322.900 ;
        RECT 83.130 322.300 86.330 322.750 ;
        RECT 79.580 322.150 89.880 322.300 ;
        RECT 83.530 321.200 85.930 322.150 ;
        RECT 90.480 321.600 90.630 329.800 ;
        RECT 91.080 321.600 91.230 329.800 ;
        RECT 91.680 321.600 91.830 329.800 ;
        RECT 92.280 321.600 92.430 329.800 ;
        RECT 92.880 321.600 93.030 329.800 ;
        RECT 93.480 321.600 93.630 329.800 ;
        RECT 94.080 321.600 94.230 329.800 ;
        RECT 95.230 330.200 95.380 338.400 ;
        RECT 95.830 330.200 95.980 338.400 ;
        RECT 96.430 330.200 96.580 338.400 ;
        RECT 97.030 330.200 97.180 338.400 ;
        RECT 97.630 330.200 97.780 338.400 ;
        RECT 98.230 330.200 98.380 338.400 ;
        RECT 98.830 330.200 98.980 338.400 ;
        RECT 103.530 337.850 105.940 338.800 ;
        RECT 99.580 337.700 109.880 337.850 ;
        RECT 103.130 337.250 106.330 337.700 ;
        RECT 99.580 337.100 109.880 337.250 ;
        RECT 103.130 336.650 106.330 337.100 ;
        RECT 99.580 336.500 109.880 336.650 ;
        RECT 103.130 336.050 106.330 336.500 ;
        RECT 99.580 335.900 109.880 336.050 ;
        RECT 103.130 335.600 106.330 335.900 ;
        RECT 103.130 335.450 103.530 335.600 ;
        RECT 99.580 335.300 103.530 335.450 ;
        RECT 103.130 334.850 103.530 335.300 ;
        RECT 99.580 334.700 103.530 334.850 ;
        RECT 103.130 334.250 103.530 334.700 ;
        RECT 99.580 334.100 103.530 334.250 ;
        RECT 103.130 333.650 103.530 334.100 ;
        RECT 99.580 333.500 103.530 333.650 ;
        RECT 103.130 333.050 103.530 333.500 ;
        RECT 99.580 332.900 103.530 333.050 ;
        RECT 103.130 332.450 103.530 332.900 ;
        RECT 99.580 332.300 103.530 332.450 ;
        RECT 103.130 331.850 103.530 332.300 ;
        RECT 99.580 331.700 103.530 331.850 ;
        RECT 103.130 331.250 103.530 331.700 ;
        RECT 99.580 331.100 103.530 331.250 ;
        RECT 103.130 330.650 103.530 331.100 ;
        RECT 99.580 330.500 103.530 330.650 ;
        RECT 103.130 330.200 103.530 330.500 ;
        RECT 95.230 329.800 103.530 330.200 ;
        RECT 95.230 321.600 95.380 329.800 ;
        RECT 95.830 321.600 95.980 329.800 ;
        RECT 96.430 321.600 96.580 329.800 ;
        RECT 97.030 321.600 97.180 329.800 ;
        RECT 97.630 321.600 97.780 329.800 ;
        RECT 98.230 321.600 98.380 329.800 ;
        RECT 98.830 321.600 98.980 329.800 ;
        RECT 103.130 329.500 103.530 329.800 ;
        RECT 99.580 329.350 103.530 329.500 ;
        RECT 103.130 328.900 103.530 329.350 ;
        RECT 99.580 328.750 103.530 328.900 ;
        RECT 103.130 328.300 103.530 328.750 ;
        RECT 99.580 328.150 103.530 328.300 ;
        RECT 103.130 327.700 103.530 328.150 ;
        RECT 99.580 327.550 103.530 327.700 ;
        RECT 103.130 327.100 103.530 327.550 ;
        RECT 99.580 326.950 103.530 327.100 ;
        RECT 103.130 326.500 103.530 326.950 ;
        RECT 99.580 326.350 103.530 326.500 ;
        RECT 103.130 325.900 103.530 326.350 ;
        RECT 99.580 325.750 103.530 325.900 ;
        RECT 103.130 325.300 103.530 325.750 ;
        RECT 99.580 325.150 103.530 325.300 ;
        RECT 103.130 324.700 103.530 325.150 ;
        RECT 99.580 324.550 103.530 324.700 ;
        RECT 103.130 324.400 103.530 324.550 ;
        RECT 105.930 335.450 106.330 335.600 ;
        RECT 105.930 335.300 109.880 335.450 ;
        RECT 105.930 334.850 106.330 335.300 ;
        RECT 105.930 334.700 109.880 334.850 ;
        RECT 105.930 334.250 106.330 334.700 ;
        RECT 105.930 334.100 109.880 334.250 ;
        RECT 105.930 333.650 106.330 334.100 ;
        RECT 105.930 333.500 109.880 333.650 ;
        RECT 105.930 333.050 106.330 333.500 ;
        RECT 105.930 332.900 109.880 333.050 ;
        RECT 105.930 332.450 106.330 332.900 ;
        RECT 105.930 332.300 109.880 332.450 ;
        RECT 105.930 331.850 106.330 332.300 ;
        RECT 105.930 331.700 109.880 331.850 ;
        RECT 105.930 331.250 106.330 331.700 ;
        RECT 105.930 331.100 109.880 331.250 ;
        RECT 105.930 330.650 106.330 331.100 ;
        RECT 105.930 330.500 109.880 330.650 ;
        RECT 105.930 330.200 106.330 330.500 ;
        RECT 110.480 330.200 110.630 338.400 ;
        RECT 111.080 330.200 111.230 338.400 ;
        RECT 111.680 330.200 111.830 338.400 ;
        RECT 112.280 330.200 112.430 338.400 ;
        RECT 112.880 330.200 113.030 338.400 ;
        RECT 113.480 330.200 113.630 338.400 ;
        RECT 114.080 330.200 114.230 338.400 ;
        RECT 105.930 329.800 114.230 330.200 ;
        RECT 105.930 329.500 106.330 329.800 ;
        RECT 105.930 329.350 109.880 329.500 ;
        RECT 105.930 328.900 106.330 329.350 ;
        RECT 105.930 328.750 109.880 328.900 ;
        RECT 105.930 328.300 106.330 328.750 ;
        RECT 105.930 328.150 109.880 328.300 ;
        RECT 105.930 327.700 106.330 328.150 ;
        RECT 105.930 327.550 109.880 327.700 ;
        RECT 105.930 327.100 106.330 327.550 ;
        RECT 105.930 326.950 109.880 327.100 ;
        RECT 105.930 326.500 106.330 326.950 ;
        RECT 105.930 326.350 109.880 326.500 ;
        RECT 105.930 325.900 106.330 326.350 ;
        RECT 105.930 325.750 109.880 325.900 ;
        RECT 105.930 325.300 106.330 325.750 ;
        RECT 105.930 325.150 109.880 325.300 ;
        RECT 105.930 324.700 106.330 325.150 ;
        RECT 105.930 324.550 109.880 324.700 ;
        RECT 105.930 324.400 106.330 324.550 ;
        RECT 103.130 324.100 106.330 324.400 ;
        RECT 99.580 323.950 109.880 324.100 ;
        RECT 103.130 323.500 106.330 323.950 ;
        RECT 99.580 323.350 109.880 323.500 ;
        RECT 103.130 322.900 106.330 323.350 ;
        RECT 99.580 322.750 109.880 322.900 ;
        RECT 103.130 322.300 106.330 322.750 ;
        RECT 99.580 322.150 109.880 322.300 ;
        RECT 103.530 321.200 105.930 322.150 ;
        RECT 110.480 321.600 110.630 329.800 ;
        RECT 111.080 321.600 111.230 329.800 ;
        RECT 111.680 321.600 111.830 329.800 ;
        RECT 112.280 321.600 112.430 329.800 ;
        RECT 112.880 321.600 113.030 329.800 ;
        RECT 113.480 321.600 113.630 329.800 ;
        RECT 114.080 321.600 114.230 329.800 ;
        RECT 115.230 330.200 115.380 338.400 ;
        RECT 115.830 330.200 115.980 338.400 ;
        RECT 116.430 330.200 116.580 338.400 ;
        RECT 117.030 330.200 117.180 338.400 ;
        RECT 117.630 330.200 117.780 338.400 ;
        RECT 118.230 330.200 118.380 338.400 ;
        RECT 118.830 330.200 118.980 338.400 ;
        RECT 123.530 337.850 124.730 338.800 ;
        RECT 119.580 337.700 124.730 337.850 ;
        RECT 123.130 337.250 124.730 337.700 ;
        RECT 119.580 337.100 124.730 337.250 ;
        RECT 123.130 336.650 124.730 337.100 ;
        RECT 119.580 336.500 124.730 336.650 ;
        RECT 123.130 336.050 124.730 336.500 ;
        RECT 125.130 336.310 127.130 337.585 ;
        RECT 119.580 335.900 124.730 336.050 ;
        RECT 123.130 335.600 124.730 335.900 ;
        RECT 123.130 335.450 123.530 335.600 ;
        RECT 119.580 335.300 123.530 335.450 ;
        RECT 123.130 334.850 123.530 335.300 ;
        RECT 119.580 334.700 123.530 334.850 ;
        RECT 123.130 334.250 123.530 334.700 ;
        RECT 119.580 334.100 123.530 334.250 ;
        RECT 123.130 333.650 123.530 334.100 ;
        RECT 119.580 333.500 123.530 333.650 ;
        RECT 123.130 333.050 123.530 333.500 ;
        RECT 119.580 332.900 123.530 333.050 ;
        RECT 123.130 332.450 123.530 332.900 ;
        RECT 119.580 332.300 123.530 332.450 ;
        RECT 123.130 331.850 123.530 332.300 ;
        RECT 119.580 331.700 123.530 331.850 ;
        RECT 123.130 331.250 123.530 331.700 ;
        RECT 119.580 331.100 123.530 331.250 ;
        RECT 123.130 330.650 123.530 331.100 ;
        RECT 119.580 330.500 123.530 330.650 ;
        RECT 123.130 330.200 123.530 330.500 ;
        RECT 115.230 329.800 123.530 330.200 ;
        RECT 115.230 321.600 115.380 329.800 ;
        RECT 115.830 321.600 115.980 329.800 ;
        RECT 116.430 321.600 116.580 329.800 ;
        RECT 117.030 321.600 117.180 329.800 ;
        RECT 117.630 321.600 117.780 329.800 ;
        RECT 118.230 321.600 118.380 329.800 ;
        RECT 118.830 321.600 118.980 329.800 ;
        RECT 123.130 329.500 123.530 329.800 ;
        RECT 119.580 329.350 123.530 329.500 ;
        RECT 123.130 328.900 123.530 329.350 ;
        RECT 119.580 328.750 123.530 328.900 ;
        RECT 123.130 328.300 123.530 328.750 ;
        RECT 119.580 328.150 123.530 328.300 ;
        RECT 123.130 327.700 123.530 328.150 ;
        RECT 119.580 327.550 123.530 327.700 ;
        RECT 123.130 327.100 123.530 327.550 ;
        RECT 119.580 326.950 123.530 327.100 ;
        RECT 123.130 326.500 123.530 326.950 ;
        RECT 119.580 326.350 123.530 326.500 ;
        RECT 123.130 325.900 123.530 326.350 ;
        RECT 119.580 325.750 123.530 325.900 ;
        RECT 123.130 325.300 123.530 325.750 ;
        RECT 119.580 325.150 123.530 325.300 ;
        RECT 123.130 324.700 123.530 325.150 ;
        RECT 119.580 324.550 123.530 324.700 ;
        RECT 123.130 324.400 123.530 324.550 ;
        RECT 123.130 324.100 124.730 324.400 ;
        RECT 119.580 323.950 124.730 324.100 ;
        RECT 123.130 323.500 124.730 323.950 ;
        RECT 119.580 323.350 124.730 323.500 ;
        RECT 123.130 322.900 124.730 323.350 ;
        RECT 119.580 322.750 124.730 322.900 ;
        RECT 123.130 322.300 124.730 322.750 ;
        RECT 125.140 322.325 127.140 323.600 ;
        RECT 119.580 322.150 124.730 322.300 ;
        RECT 123.530 321.200 124.730 322.150 ;
        RECT 4.730 318.800 9.130 321.200 ;
        RECT 20.330 318.800 29.130 321.200 ;
        RECT 40.330 318.800 49.130 321.200 ;
        RECT 60.330 318.800 69.130 321.200 ;
        RECT 80.330 318.800 89.130 321.200 ;
        RECT 100.330 318.800 109.130 321.200 ;
        RECT 120.330 318.800 124.730 321.200 ;
        RECT 4.730 317.850 5.940 318.800 ;
        RECT 4.730 317.700 9.880 317.850 ;
        RECT 2.315 316.100 4.320 317.375 ;
        RECT 4.730 317.250 6.330 317.700 ;
        RECT 4.730 317.100 9.880 317.250 ;
        RECT 4.730 316.650 6.330 317.100 ;
        RECT 4.730 316.500 9.880 316.650 ;
        RECT 4.730 316.050 6.330 316.500 ;
        RECT 4.730 315.900 9.880 316.050 ;
        RECT 4.730 315.600 6.330 315.900 ;
        RECT 2.315 313.250 4.315 315.545 ;
        RECT 5.930 315.450 6.330 315.600 ;
        RECT 5.930 315.300 9.880 315.450 ;
        RECT 5.930 314.850 6.330 315.300 ;
        RECT 5.930 314.700 9.880 314.850 ;
        RECT 5.930 314.250 6.330 314.700 ;
        RECT 5.930 314.100 9.880 314.250 ;
        RECT 5.930 313.650 6.330 314.100 ;
        RECT 5.930 313.500 9.880 313.650 ;
        RECT 5.930 313.050 6.330 313.500 ;
        RECT 5.930 312.900 9.880 313.050 ;
        RECT 5.930 312.450 6.330 312.900 ;
        RECT 5.930 312.300 9.880 312.450 ;
        RECT 5.930 311.850 6.330 312.300 ;
        RECT 5.930 311.700 9.880 311.850 ;
        RECT 5.930 311.250 6.330 311.700 ;
        RECT 5.930 311.100 9.880 311.250 ;
        RECT 5.930 310.650 6.330 311.100 ;
        RECT 5.930 310.500 9.880 310.650 ;
        RECT 5.930 310.200 6.330 310.500 ;
        RECT 10.480 310.200 10.630 318.400 ;
        RECT 11.080 310.200 11.230 318.400 ;
        RECT 11.680 310.200 11.830 318.400 ;
        RECT 12.280 310.200 12.430 318.400 ;
        RECT 12.880 310.200 13.030 318.400 ;
        RECT 13.480 310.200 13.630 318.400 ;
        RECT 14.080 310.200 14.230 318.400 ;
        RECT 5.930 309.800 14.230 310.200 ;
        RECT 5.930 309.500 6.330 309.800 ;
        RECT 5.930 309.350 9.880 309.500 ;
        RECT 5.930 308.900 6.330 309.350 ;
        RECT 5.930 308.750 9.880 308.900 ;
        RECT 5.930 308.300 6.330 308.750 ;
        RECT 5.930 308.150 9.880 308.300 ;
        RECT 5.930 307.700 6.330 308.150 ;
        RECT 5.930 307.550 9.880 307.700 ;
        RECT 5.930 307.100 6.330 307.550 ;
        RECT 5.930 306.950 9.880 307.100 ;
        RECT 2.315 304.455 4.315 306.750 ;
        RECT 5.930 306.500 6.330 306.950 ;
        RECT 5.930 306.350 9.880 306.500 ;
        RECT 5.930 305.900 6.330 306.350 ;
        RECT 5.930 305.750 9.880 305.900 ;
        RECT 5.930 305.300 6.330 305.750 ;
        RECT 5.930 305.150 9.880 305.300 ;
        RECT 5.930 304.700 6.330 305.150 ;
        RECT 5.930 304.550 9.880 304.700 ;
        RECT 5.930 304.400 6.330 304.550 ;
        RECT 4.730 304.100 6.330 304.400 ;
        RECT 4.730 303.950 9.880 304.100 ;
        RECT 2.315 302.400 4.320 303.675 ;
        RECT 4.730 303.500 6.330 303.950 ;
        RECT 4.730 303.350 9.880 303.500 ;
        RECT 4.730 302.900 6.330 303.350 ;
        RECT 4.730 302.750 9.880 302.900 ;
        RECT 4.730 302.300 6.330 302.750 ;
        RECT 4.730 302.150 9.880 302.300 ;
        RECT 4.730 301.200 5.930 302.150 ;
        RECT 10.480 301.600 10.630 309.800 ;
        RECT 11.080 301.600 11.230 309.800 ;
        RECT 11.680 301.600 11.830 309.800 ;
        RECT 12.280 301.600 12.430 309.800 ;
        RECT 12.880 301.600 13.030 309.800 ;
        RECT 13.480 301.600 13.630 309.800 ;
        RECT 14.080 301.600 14.230 309.800 ;
        RECT 15.230 310.200 15.380 318.400 ;
        RECT 15.830 310.200 15.980 318.400 ;
        RECT 16.430 310.200 16.580 318.400 ;
        RECT 17.030 310.200 17.180 318.400 ;
        RECT 17.630 310.200 17.780 318.400 ;
        RECT 18.230 310.200 18.380 318.400 ;
        RECT 18.830 310.200 18.980 318.400 ;
        RECT 23.530 317.850 25.940 318.800 ;
        RECT 19.580 317.700 29.880 317.850 ;
        RECT 23.130 317.250 26.330 317.700 ;
        RECT 19.580 317.100 29.880 317.250 ;
        RECT 23.130 316.650 26.330 317.100 ;
        RECT 19.580 316.500 29.880 316.650 ;
        RECT 23.130 316.050 26.330 316.500 ;
        RECT 19.580 315.900 29.880 316.050 ;
        RECT 23.130 315.600 26.330 315.900 ;
        RECT 23.130 315.450 23.530 315.600 ;
        RECT 19.580 315.300 23.530 315.450 ;
        RECT 23.130 314.850 23.530 315.300 ;
        RECT 19.580 314.700 23.530 314.850 ;
        RECT 23.130 314.250 23.530 314.700 ;
        RECT 19.580 314.100 23.530 314.250 ;
        RECT 23.130 313.650 23.530 314.100 ;
        RECT 19.580 313.500 23.530 313.650 ;
        RECT 23.130 313.050 23.530 313.500 ;
        RECT 19.580 312.900 23.530 313.050 ;
        RECT 23.130 312.450 23.530 312.900 ;
        RECT 19.580 312.300 23.530 312.450 ;
        RECT 23.130 311.850 23.530 312.300 ;
        RECT 19.580 311.700 23.530 311.850 ;
        RECT 23.130 311.250 23.530 311.700 ;
        RECT 19.580 311.100 23.530 311.250 ;
        RECT 23.130 310.650 23.530 311.100 ;
        RECT 19.580 310.500 23.530 310.650 ;
        RECT 23.130 310.200 23.530 310.500 ;
        RECT 15.230 309.800 23.530 310.200 ;
        RECT 15.230 301.600 15.380 309.800 ;
        RECT 15.830 301.600 15.980 309.800 ;
        RECT 16.430 301.600 16.580 309.800 ;
        RECT 17.030 301.600 17.180 309.800 ;
        RECT 17.630 301.600 17.780 309.800 ;
        RECT 18.230 301.600 18.380 309.800 ;
        RECT 18.830 301.600 18.980 309.800 ;
        RECT 23.130 309.500 23.530 309.800 ;
        RECT 19.580 309.350 23.530 309.500 ;
        RECT 23.130 308.900 23.530 309.350 ;
        RECT 19.580 308.750 23.530 308.900 ;
        RECT 23.130 308.300 23.530 308.750 ;
        RECT 19.580 308.150 23.530 308.300 ;
        RECT 23.130 307.700 23.530 308.150 ;
        RECT 19.580 307.550 23.530 307.700 ;
        RECT 23.130 307.100 23.530 307.550 ;
        RECT 19.580 306.950 23.530 307.100 ;
        RECT 23.130 306.500 23.530 306.950 ;
        RECT 19.580 306.350 23.530 306.500 ;
        RECT 23.130 305.900 23.530 306.350 ;
        RECT 19.580 305.750 23.530 305.900 ;
        RECT 23.130 305.300 23.530 305.750 ;
        RECT 19.580 305.150 23.530 305.300 ;
        RECT 23.130 304.700 23.530 305.150 ;
        RECT 19.580 304.550 23.530 304.700 ;
        RECT 23.130 304.400 23.530 304.550 ;
        RECT 25.930 315.450 26.330 315.600 ;
        RECT 25.930 315.300 29.880 315.450 ;
        RECT 25.930 314.850 26.330 315.300 ;
        RECT 25.930 314.700 29.880 314.850 ;
        RECT 25.930 314.250 26.330 314.700 ;
        RECT 25.930 314.100 29.880 314.250 ;
        RECT 25.930 313.650 26.330 314.100 ;
        RECT 25.930 313.500 29.880 313.650 ;
        RECT 25.930 313.050 26.330 313.500 ;
        RECT 25.930 312.900 29.880 313.050 ;
        RECT 25.930 312.450 26.330 312.900 ;
        RECT 25.930 312.300 29.880 312.450 ;
        RECT 25.930 311.850 26.330 312.300 ;
        RECT 25.930 311.700 29.880 311.850 ;
        RECT 25.930 311.250 26.330 311.700 ;
        RECT 25.930 311.100 29.880 311.250 ;
        RECT 25.930 310.650 26.330 311.100 ;
        RECT 25.930 310.500 29.880 310.650 ;
        RECT 25.930 310.200 26.330 310.500 ;
        RECT 30.480 310.200 30.630 318.400 ;
        RECT 31.080 310.200 31.230 318.400 ;
        RECT 31.680 310.200 31.830 318.400 ;
        RECT 32.280 310.200 32.430 318.400 ;
        RECT 32.880 310.200 33.030 318.400 ;
        RECT 33.480 310.200 33.630 318.400 ;
        RECT 34.080 310.200 34.230 318.400 ;
        RECT 25.930 309.800 34.230 310.200 ;
        RECT 25.930 309.500 26.330 309.800 ;
        RECT 25.930 309.350 29.880 309.500 ;
        RECT 25.930 308.900 26.330 309.350 ;
        RECT 25.930 308.750 29.880 308.900 ;
        RECT 25.930 308.300 26.330 308.750 ;
        RECT 25.930 308.150 29.880 308.300 ;
        RECT 25.930 307.700 26.330 308.150 ;
        RECT 25.930 307.550 29.880 307.700 ;
        RECT 25.930 307.100 26.330 307.550 ;
        RECT 25.930 306.950 29.880 307.100 ;
        RECT 25.930 306.500 26.330 306.950 ;
        RECT 25.930 306.350 29.880 306.500 ;
        RECT 25.930 305.900 26.330 306.350 ;
        RECT 25.930 305.750 29.880 305.900 ;
        RECT 25.930 305.300 26.330 305.750 ;
        RECT 25.930 305.150 29.880 305.300 ;
        RECT 25.930 304.700 26.330 305.150 ;
        RECT 25.930 304.550 29.880 304.700 ;
        RECT 25.930 304.400 26.330 304.550 ;
        RECT 23.130 304.100 26.330 304.400 ;
        RECT 19.580 303.950 29.880 304.100 ;
        RECT 23.130 303.500 26.330 303.950 ;
        RECT 19.580 303.350 29.880 303.500 ;
        RECT 23.130 302.900 26.330 303.350 ;
        RECT 19.580 302.750 29.880 302.900 ;
        RECT 23.130 302.300 26.330 302.750 ;
        RECT 19.580 302.150 29.880 302.300 ;
        RECT 23.530 301.200 25.930 302.150 ;
        RECT 30.480 301.600 30.630 309.800 ;
        RECT 31.080 301.600 31.230 309.800 ;
        RECT 31.680 301.600 31.830 309.800 ;
        RECT 32.280 301.600 32.430 309.800 ;
        RECT 32.880 301.600 33.030 309.800 ;
        RECT 33.480 301.600 33.630 309.800 ;
        RECT 34.080 301.600 34.230 309.800 ;
        RECT 35.230 310.200 35.380 318.400 ;
        RECT 35.830 310.200 35.980 318.400 ;
        RECT 36.430 310.200 36.580 318.400 ;
        RECT 37.030 310.200 37.180 318.400 ;
        RECT 37.630 310.200 37.780 318.400 ;
        RECT 38.230 310.200 38.380 318.400 ;
        RECT 38.830 310.200 38.980 318.400 ;
        RECT 43.530 317.850 45.940 318.800 ;
        RECT 39.580 317.700 49.880 317.850 ;
        RECT 43.130 317.250 46.330 317.700 ;
        RECT 39.580 317.100 49.880 317.250 ;
        RECT 43.130 316.650 46.330 317.100 ;
        RECT 39.580 316.500 49.880 316.650 ;
        RECT 43.130 316.050 46.330 316.500 ;
        RECT 39.580 315.900 49.880 316.050 ;
        RECT 43.130 315.600 46.330 315.900 ;
        RECT 43.130 315.450 43.530 315.600 ;
        RECT 39.580 315.300 43.530 315.450 ;
        RECT 43.130 314.850 43.530 315.300 ;
        RECT 39.580 314.700 43.530 314.850 ;
        RECT 43.130 314.250 43.530 314.700 ;
        RECT 39.580 314.100 43.530 314.250 ;
        RECT 43.130 313.650 43.530 314.100 ;
        RECT 39.580 313.500 43.530 313.650 ;
        RECT 43.130 313.050 43.530 313.500 ;
        RECT 39.580 312.900 43.530 313.050 ;
        RECT 43.130 312.450 43.530 312.900 ;
        RECT 39.580 312.300 43.530 312.450 ;
        RECT 43.130 311.850 43.530 312.300 ;
        RECT 39.580 311.700 43.530 311.850 ;
        RECT 43.130 311.250 43.530 311.700 ;
        RECT 39.580 311.100 43.530 311.250 ;
        RECT 43.130 310.650 43.530 311.100 ;
        RECT 39.580 310.500 43.530 310.650 ;
        RECT 43.130 310.200 43.530 310.500 ;
        RECT 35.230 309.800 43.530 310.200 ;
        RECT 35.230 301.600 35.380 309.800 ;
        RECT 35.830 301.600 35.980 309.800 ;
        RECT 36.430 301.600 36.580 309.800 ;
        RECT 37.030 301.600 37.180 309.800 ;
        RECT 37.630 301.600 37.780 309.800 ;
        RECT 38.230 301.600 38.380 309.800 ;
        RECT 38.830 301.600 38.980 309.800 ;
        RECT 43.130 309.500 43.530 309.800 ;
        RECT 39.580 309.350 43.530 309.500 ;
        RECT 43.130 308.900 43.530 309.350 ;
        RECT 39.580 308.750 43.530 308.900 ;
        RECT 43.130 308.300 43.530 308.750 ;
        RECT 39.580 308.150 43.530 308.300 ;
        RECT 43.130 307.700 43.530 308.150 ;
        RECT 39.580 307.550 43.530 307.700 ;
        RECT 43.130 307.100 43.530 307.550 ;
        RECT 39.580 306.950 43.530 307.100 ;
        RECT 43.130 306.500 43.530 306.950 ;
        RECT 39.580 306.350 43.530 306.500 ;
        RECT 43.130 305.900 43.530 306.350 ;
        RECT 39.580 305.750 43.530 305.900 ;
        RECT 43.130 305.300 43.530 305.750 ;
        RECT 39.580 305.150 43.530 305.300 ;
        RECT 43.130 304.700 43.530 305.150 ;
        RECT 39.580 304.550 43.530 304.700 ;
        RECT 43.130 304.400 43.530 304.550 ;
        RECT 45.930 315.450 46.330 315.600 ;
        RECT 45.930 315.300 49.880 315.450 ;
        RECT 45.930 314.850 46.330 315.300 ;
        RECT 45.930 314.700 49.880 314.850 ;
        RECT 45.930 314.250 46.330 314.700 ;
        RECT 45.930 314.100 49.880 314.250 ;
        RECT 45.930 313.650 46.330 314.100 ;
        RECT 45.930 313.500 49.880 313.650 ;
        RECT 45.930 313.050 46.330 313.500 ;
        RECT 45.930 312.900 49.880 313.050 ;
        RECT 45.930 312.450 46.330 312.900 ;
        RECT 45.930 312.300 49.880 312.450 ;
        RECT 45.930 311.850 46.330 312.300 ;
        RECT 45.930 311.700 49.880 311.850 ;
        RECT 45.930 311.250 46.330 311.700 ;
        RECT 45.930 311.100 49.880 311.250 ;
        RECT 45.930 310.650 46.330 311.100 ;
        RECT 45.930 310.500 49.880 310.650 ;
        RECT 45.930 310.200 46.330 310.500 ;
        RECT 50.480 310.200 50.630 318.400 ;
        RECT 51.080 310.200 51.230 318.400 ;
        RECT 51.680 310.200 51.830 318.400 ;
        RECT 52.280 310.200 52.430 318.400 ;
        RECT 52.880 310.200 53.030 318.400 ;
        RECT 53.480 310.200 53.630 318.400 ;
        RECT 54.080 310.200 54.230 318.400 ;
        RECT 45.930 309.800 54.230 310.200 ;
        RECT 45.930 309.500 46.330 309.800 ;
        RECT 45.930 309.350 49.880 309.500 ;
        RECT 45.930 308.900 46.330 309.350 ;
        RECT 45.930 308.750 49.880 308.900 ;
        RECT 45.930 308.300 46.330 308.750 ;
        RECT 45.930 308.150 49.880 308.300 ;
        RECT 45.930 307.700 46.330 308.150 ;
        RECT 45.930 307.550 49.880 307.700 ;
        RECT 45.930 307.100 46.330 307.550 ;
        RECT 45.930 306.950 49.880 307.100 ;
        RECT 45.930 306.500 46.330 306.950 ;
        RECT 45.930 306.350 49.880 306.500 ;
        RECT 45.930 305.900 46.330 306.350 ;
        RECT 45.930 305.750 49.880 305.900 ;
        RECT 45.930 305.300 46.330 305.750 ;
        RECT 45.930 305.150 49.880 305.300 ;
        RECT 45.930 304.700 46.330 305.150 ;
        RECT 45.930 304.550 49.880 304.700 ;
        RECT 45.930 304.400 46.330 304.550 ;
        RECT 43.130 304.100 46.330 304.400 ;
        RECT 39.580 303.950 49.880 304.100 ;
        RECT 43.130 303.500 46.330 303.950 ;
        RECT 39.580 303.350 49.880 303.500 ;
        RECT 43.130 302.900 46.330 303.350 ;
        RECT 39.580 302.750 49.880 302.900 ;
        RECT 43.130 302.300 46.330 302.750 ;
        RECT 39.580 302.150 49.880 302.300 ;
        RECT 43.530 301.200 45.930 302.150 ;
        RECT 50.480 301.600 50.630 309.800 ;
        RECT 51.080 301.600 51.230 309.800 ;
        RECT 51.680 301.600 51.830 309.800 ;
        RECT 52.280 301.600 52.430 309.800 ;
        RECT 52.880 301.600 53.030 309.800 ;
        RECT 53.480 301.600 53.630 309.800 ;
        RECT 54.080 301.600 54.230 309.800 ;
        RECT 55.230 310.200 55.380 318.400 ;
        RECT 55.830 310.200 55.980 318.400 ;
        RECT 56.430 310.200 56.580 318.400 ;
        RECT 57.030 310.200 57.180 318.400 ;
        RECT 57.630 310.200 57.780 318.400 ;
        RECT 58.230 310.200 58.380 318.400 ;
        RECT 58.830 310.200 58.980 318.400 ;
        RECT 63.530 317.850 65.940 318.800 ;
        RECT 59.580 317.700 69.880 317.850 ;
        RECT 63.130 317.250 66.330 317.700 ;
        RECT 59.580 317.100 69.880 317.250 ;
        RECT 63.130 316.650 66.330 317.100 ;
        RECT 59.580 316.500 69.880 316.650 ;
        RECT 63.130 316.050 66.330 316.500 ;
        RECT 59.580 315.900 69.880 316.050 ;
        RECT 63.130 315.600 66.330 315.900 ;
        RECT 63.130 315.450 63.530 315.600 ;
        RECT 59.580 315.300 63.530 315.450 ;
        RECT 63.130 314.850 63.530 315.300 ;
        RECT 59.580 314.700 63.530 314.850 ;
        RECT 63.130 314.250 63.530 314.700 ;
        RECT 59.580 314.100 63.530 314.250 ;
        RECT 63.130 313.650 63.530 314.100 ;
        RECT 59.580 313.500 63.530 313.650 ;
        RECT 63.130 313.050 63.530 313.500 ;
        RECT 59.580 312.900 63.530 313.050 ;
        RECT 63.130 312.450 63.530 312.900 ;
        RECT 59.580 312.300 63.530 312.450 ;
        RECT 63.130 311.850 63.530 312.300 ;
        RECT 59.580 311.700 63.530 311.850 ;
        RECT 63.130 311.250 63.530 311.700 ;
        RECT 59.580 311.100 63.530 311.250 ;
        RECT 63.130 310.650 63.530 311.100 ;
        RECT 59.580 310.500 63.530 310.650 ;
        RECT 63.130 310.200 63.530 310.500 ;
        RECT 55.230 309.800 63.530 310.200 ;
        RECT 55.230 301.600 55.380 309.800 ;
        RECT 55.830 301.600 55.980 309.800 ;
        RECT 56.430 301.600 56.580 309.800 ;
        RECT 57.030 301.600 57.180 309.800 ;
        RECT 57.630 301.600 57.780 309.800 ;
        RECT 58.230 301.600 58.380 309.800 ;
        RECT 58.830 301.600 58.980 309.800 ;
        RECT 63.130 309.500 63.530 309.800 ;
        RECT 59.580 309.350 63.530 309.500 ;
        RECT 63.130 308.900 63.530 309.350 ;
        RECT 59.580 308.750 63.530 308.900 ;
        RECT 63.130 308.300 63.530 308.750 ;
        RECT 59.580 308.150 63.530 308.300 ;
        RECT 63.130 307.700 63.530 308.150 ;
        RECT 59.580 307.550 63.530 307.700 ;
        RECT 63.130 307.100 63.530 307.550 ;
        RECT 59.580 306.950 63.530 307.100 ;
        RECT 63.130 306.500 63.530 306.950 ;
        RECT 59.580 306.350 63.530 306.500 ;
        RECT 63.130 305.900 63.530 306.350 ;
        RECT 59.580 305.750 63.530 305.900 ;
        RECT 63.130 305.300 63.530 305.750 ;
        RECT 59.580 305.150 63.530 305.300 ;
        RECT 63.130 304.700 63.530 305.150 ;
        RECT 59.580 304.550 63.530 304.700 ;
        RECT 63.130 304.400 63.530 304.550 ;
        RECT 65.930 315.450 66.330 315.600 ;
        RECT 65.930 315.300 69.880 315.450 ;
        RECT 65.930 314.850 66.330 315.300 ;
        RECT 65.930 314.700 69.880 314.850 ;
        RECT 65.930 314.250 66.330 314.700 ;
        RECT 65.930 314.100 69.880 314.250 ;
        RECT 65.930 313.650 66.330 314.100 ;
        RECT 65.930 313.500 69.880 313.650 ;
        RECT 65.930 313.050 66.330 313.500 ;
        RECT 65.930 312.900 69.880 313.050 ;
        RECT 65.930 312.450 66.330 312.900 ;
        RECT 65.930 312.300 69.880 312.450 ;
        RECT 65.930 311.850 66.330 312.300 ;
        RECT 65.930 311.700 69.880 311.850 ;
        RECT 65.930 311.250 66.330 311.700 ;
        RECT 65.930 311.100 69.880 311.250 ;
        RECT 65.930 310.650 66.330 311.100 ;
        RECT 65.930 310.500 69.880 310.650 ;
        RECT 65.930 310.200 66.330 310.500 ;
        RECT 70.480 310.200 70.630 318.400 ;
        RECT 71.080 310.200 71.230 318.400 ;
        RECT 71.680 310.200 71.830 318.400 ;
        RECT 72.280 310.200 72.430 318.400 ;
        RECT 72.880 310.200 73.030 318.400 ;
        RECT 73.480 310.200 73.630 318.400 ;
        RECT 74.080 310.200 74.230 318.400 ;
        RECT 65.930 309.800 74.230 310.200 ;
        RECT 65.930 309.500 66.330 309.800 ;
        RECT 65.930 309.350 69.880 309.500 ;
        RECT 65.930 308.900 66.330 309.350 ;
        RECT 65.930 308.750 69.880 308.900 ;
        RECT 65.930 308.300 66.330 308.750 ;
        RECT 65.930 308.150 69.880 308.300 ;
        RECT 65.930 307.700 66.330 308.150 ;
        RECT 65.930 307.550 69.880 307.700 ;
        RECT 65.930 307.100 66.330 307.550 ;
        RECT 65.930 306.950 69.880 307.100 ;
        RECT 65.930 306.500 66.330 306.950 ;
        RECT 65.930 306.350 69.880 306.500 ;
        RECT 65.930 305.900 66.330 306.350 ;
        RECT 65.930 305.750 69.880 305.900 ;
        RECT 65.930 305.300 66.330 305.750 ;
        RECT 65.930 305.150 69.880 305.300 ;
        RECT 65.930 304.700 66.330 305.150 ;
        RECT 65.930 304.550 69.880 304.700 ;
        RECT 65.930 304.400 66.330 304.550 ;
        RECT 63.130 304.100 66.330 304.400 ;
        RECT 59.580 303.950 69.880 304.100 ;
        RECT 63.130 303.500 66.330 303.950 ;
        RECT 59.580 303.350 69.880 303.500 ;
        RECT 63.130 302.900 66.330 303.350 ;
        RECT 59.580 302.750 69.880 302.900 ;
        RECT 63.130 302.300 66.330 302.750 ;
        RECT 59.580 302.150 69.880 302.300 ;
        RECT 63.530 301.200 65.930 302.150 ;
        RECT 70.480 301.600 70.630 309.800 ;
        RECT 71.080 301.600 71.230 309.800 ;
        RECT 71.680 301.600 71.830 309.800 ;
        RECT 72.280 301.600 72.430 309.800 ;
        RECT 72.880 301.600 73.030 309.800 ;
        RECT 73.480 301.600 73.630 309.800 ;
        RECT 74.080 301.600 74.230 309.800 ;
        RECT 75.230 310.200 75.380 318.400 ;
        RECT 75.830 310.200 75.980 318.400 ;
        RECT 76.430 310.200 76.580 318.400 ;
        RECT 77.030 310.200 77.180 318.400 ;
        RECT 77.630 310.200 77.780 318.400 ;
        RECT 78.230 310.200 78.380 318.400 ;
        RECT 78.830 310.200 78.980 318.400 ;
        RECT 83.530 317.850 85.940 318.800 ;
        RECT 79.580 317.700 89.880 317.850 ;
        RECT 83.130 317.250 86.330 317.700 ;
        RECT 79.580 317.100 89.880 317.250 ;
        RECT 83.130 316.650 86.330 317.100 ;
        RECT 79.580 316.500 89.880 316.650 ;
        RECT 83.130 316.050 86.330 316.500 ;
        RECT 79.580 315.900 89.880 316.050 ;
        RECT 83.130 315.600 86.330 315.900 ;
        RECT 83.130 315.450 83.530 315.600 ;
        RECT 79.580 315.300 83.530 315.450 ;
        RECT 83.130 314.850 83.530 315.300 ;
        RECT 79.580 314.700 83.530 314.850 ;
        RECT 83.130 314.250 83.530 314.700 ;
        RECT 79.580 314.100 83.530 314.250 ;
        RECT 83.130 313.650 83.530 314.100 ;
        RECT 79.580 313.500 83.530 313.650 ;
        RECT 83.130 313.050 83.530 313.500 ;
        RECT 79.580 312.900 83.530 313.050 ;
        RECT 83.130 312.450 83.530 312.900 ;
        RECT 79.580 312.300 83.530 312.450 ;
        RECT 83.130 311.850 83.530 312.300 ;
        RECT 79.580 311.700 83.530 311.850 ;
        RECT 83.130 311.250 83.530 311.700 ;
        RECT 79.580 311.100 83.530 311.250 ;
        RECT 83.130 310.650 83.530 311.100 ;
        RECT 79.580 310.500 83.530 310.650 ;
        RECT 83.130 310.200 83.530 310.500 ;
        RECT 75.230 309.800 83.530 310.200 ;
        RECT 75.230 301.600 75.380 309.800 ;
        RECT 75.830 301.600 75.980 309.800 ;
        RECT 76.430 301.600 76.580 309.800 ;
        RECT 77.030 301.600 77.180 309.800 ;
        RECT 77.630 301.600 77.780 309.800 ;
        RECT 78.230 301.600 78.380 309.800 ;
        RECT 78.830 301.600 78.980 309.800 ;
        RECT 83.130 309.500 83.530 309.800 ;
        RECT 79.580 309.350 83.530 309.500 ;
        RECT 83.130 308.900 83.530 309.350 ;
        RECT 79.580 308.750 83.530 308.900 ;
        RECT 83.130 308.300 83.530 308.750 ;
        RECT 79.580 308.150 83.530 308.300 ;
        RECT 83.130 307.700 83.530 308.150 ;
        RECT 79.580 307.550 83.530 307.700 ;
        RECT 83.130 307.100 83.530 307.550 ;
        RECT 79.580 306.950 83.530 307.100 ;
        RECT 83.130 306.500 83.530 306.950 ;
        RECT 79.580 306.350 83.530 306.500 ;
        RECT 83.130 305.900 83.530 306.350 ;
        RECT 79.580 305.750 83.530 305.900 ;
        RECT 83.130 305.300 83.530 305.750 ;
        RECT 79.580 305.150 83.530 305.300 ;
        RECT 83.130 304.700 83.530 305.150 ;
        RECT 79.580 304.550 83.530 304.700 ;
        RECT 83.130 304.400 83.530 304.550 ;
        RECT 85.930 315.450 86.330 315.600 ;
        RECT 85.930 315.300 89.880 315.450 ;
        RECT 85.930 314.850 86.330 315.300 ;
        RECT 85.930 314.700 89.880 314.850 ;
        RECT 85.930 314.250 86.330 314.700 ;
        RECT 85.930 314.100 89.880 314.250 ;
        RECT 85.930 313.650 86.330 314.100 ;
        RECT 85.930 313.500 89.880 313.650 ;
        RECT 85.930 313.050 86.330 313.500 ;
        RECT 85.930 312.900 89.880 313.050 ;
        RECT 85.930 312.450 86.330 312.900 ;
        RECT 85.930 312.300 89.880 312.450 ;
        RECT 85.930 311.850 86.330 312.300 ;
        RECT 85.930 311.700 89.880 311.850 ;
        RECT 85.930 311.250 86.330 311.700 ;
        RECT 85.930 311.100 89.880 311.250 ;
        RECT 85.930 310.650 86.330 311.100 ;
        RECT 85.930 310.500 89.880 310.650 ;
        RECT 85.930 310.200 86.330 310.500 ;
        RECT 90.480 310.200 90.630 318.400 ;
        RECT 91.080 310.200 91.230 318.400 ;
        RECT 91.680 310.200 91.830 318.400 ;
        RECT 92.280 310.200 92.430 318.400 ;
        RECT 92.880 310.200 93.030 318.400 ;
        RECT 93.480 310.200 93.630 318.400 ;
        RECT 94.080 310.200 94.230 318.400 ;
        RECT 85.930 309.800 94.230 310.200 ;
        RECT 85.930 309.500 86.330 309.800 ;
        RECT 85.930 309.350 89.880 309.500 ;
        RECT 85.930 308.900 86.330 309.350 ;
        RECT 85.930 308.750 89.880 308.900 ;
        RECT 85.930 308.300 86.330 308.750 ;
        RECT 85.930 308.150 89.880 308.300 ;
        RECT 85.930 307.700 86.330 308.150 ;
        RECT 85.930 307.550 89.880 307.700 ;
        RECT 85.930 307.100 86.330 307.550 ;
        RECT 85.930 306.950 89.880 307.100 ;
        RECT 85.930 306.500 86.330 306.950 ;
        RECT 85.930 306.350 89.880 306.500 ;
        RECT 85.930 305.900 86.330 306.350 ;
        RECT 85.930 305.750 89.880 305.900 ;
        RECT 85.930 305.300 86.330 305.750 ;
        RECT 85.930 305.150 89.880 305.300 ;
        RECT 85.930 304.700 86.330 305.150 ;
        RECT 85.930 304.550 89.880 304.700 ;
        RECT 85.930 304.400 86.330 304.550 ;
        RECT 83.130 304.100 86.330 304.400 ;
        RECT 79.580 303.950 89.880 304.100 ;
        RECT 83.130 303.500 86.330 303.950 ;
        RECT 79.580 303.350 89.880 303.500 ;
        RECT 83.130 302.900 86.330 303.350 ;
        RECT 79.580 302.750 89.880 302.900 ;
        RECT 83.130 302.300 86.330 302.750 ;
        RECT 79.580 302.150 89.880 302.300 ;
        RECT 83.530 301.200 85.930 302.150 ;
        RECT 90.480 301.600 90.630 309.800 ;
        RECT 91.080 301.600 91.230 309.800 ;
        RECT 91.680 301.600 91.830 309.800 ;
        RECT 92.280 301.600 92.430 309.800 ;
        RECT 92.880 301.600 93.030 309.800 ;
        RECT 93.480 301.600 93.630 309.800 ;
        RECT 94.080 301.600 94.230 309.800 ;
        RECT 95.230 310.200 95.380 318.400 ;
        RECT 95.830 310.200 95.980 318.400 ;
        RECT 96.430 310.200 96.580 318.400 ;
        RECT 97.030 310.200 97.180 318.400 ;
        RECT 97.630 310.200 97.780 318.400 ;
        RECT 98.230 310.200 98.380 318.400 ;
        RECT 98.830 310.200 98.980 318.400 ;
        RECT 103.530 317.850 105.940 318.800 ;
        RECT 99.580 317.700 109.880 317.850 ;
        RECT 103.130 317.250 106.330 317.700 ;
        RECT 99.580 317.100 109.880 317.250 ;
        RECT 103.130 316.650 106.330 317.100 ;
        RECT 99.580 316.500 109.880 316.650 ;
        RECT 103.130 316.050 106.330 316.500 ;
        RECT 99.580 315.900 109.880 316.050 ;
        RECT 103.130 315.600 106.330 315.900 ;
        RECT 103.130 315.450 103.530 315.600 ;
        RECT 99.580 315.300 103.530 315.450 ;
        RECT 103.130 314.850 103.530 315.300 ;
        RECT 99.580 314.700 103.530 314.850 ;
        RECT 103.130 314.250 103.530 314.700 ;
        RECT 99.580 314.100 103.530 314.250 ;
        RECT 103.130 313.650 103.530 314.100 ;
        RECT 99.580 313.500 103.530 313.650 ;
        RECT 103.130 313.050 103.530 313.500 ;
        RECT 99.580 312.900 103.530 313.050 ;
        RECT 103.130 312.450 103.530 312.900 ;
        RECT 99.580 312.300 103.530 312.450 ;
        RECT 103.130 311.850 103.530 312.300 ;
        RECT 99.580 311.700 103.530 311.850 ;
        RECT 103.130 311.250 103.530 311.700 ;
        RECT 99.580 311.100 103.530 311.250 ;
        RECT 103.130 310.650 103.530 311.100 ;
        RECT 99.580 310.500 103.530 310.650 ;
        RECT 103.130 310.200 103.530 310.500 ;
        RECT 95.230 309.800 103.530 310.200 ;
        RECT 95.230 301.600 95.380 309.800 ;
        RECT 95.830 301.600 95.980 309.800 ;
        RECT 96.430 301.600 96.580 309.800 ;
        RECT 97.030 301.600 97.180 309.800 ;
        RECT 97.630 301.600 97.780 309.800 ;
        RECT 98.230 301.600 98.380 309.800 ;
        RECT 98.830 301.600 98.980 309.800 ;
        RECT 103.130 309.500 103.530 309.800 ;
        RECT 99.580 309.350 103.530 309.500 ;
        RECT 103.130 308.900 103.530 309.350 ;
        RECT 99.580 308.750 103.530 308.900 ;
        RECT 103.130 308.300 103.530 308.750 ;
        RECT 99.580 308.150 103.530 308.300 ;
        RECT 103.130 307.700 103.530 308.150 ;
        RECT 99.580 307.550 103.530 307.700 ;
        RECT 103.130 307.100 103.530 307.550 ;
        RECT 99.580 306.950 103.530 307.100 ;
        RECT 103.130 306.500 103.530 306.950 ;
        RECT 99.580 306.350 103.530 306.500 ;
        RECT 103.130 305.900 103.530 306.350 ;
        RECT 99.580 305.750 103.530 305.900 ;
        RECT 103.130 305.300 103.530 305.750 ;
        RECT 99.580 305.150 103.530 305.300 ;
        RECT 103.130 304.700 103.530 305.150 ;
        RECT 99.580 304.550 103.530 304.700 ;
        RECT 103.130 304.400 103.530 304.550 ;
        RECT 105.930 315.450 106.330 315.600 ;
        RECT 105.930 315.300 109.880 315.450 ;
        RECT 105.930 314.850 106.330 315.300 ;
        RECT 105.930 314.700 109.880 314.850 ;
        RECT 105.930 314.250 106.330 314.700 ;
        RECT 105.930 314.100 109.880 314.250 ;
        RECT 105.930 313.650 106.330 314.100 ;
        RECT 105.930 313.500 109.880 313.650 ;
        RECT 105.930 313.050 106.330 313.500 ;
        RECT 105.930 312.900 109.880 313.050 ;
        RECT 105.930 312.450 106.330 312.900 ;
        RECT 105.930 312.300 109.880 312.450 ;
        RECT 105.930 311.850 106.330 312.300 ;
        RECT 105.930 311.700 109.880 311.850 ;
        RECT 105.930 311.250 106.330 311.700 ;
        RECT 105.930 311.100 109.880 311.250 ;
        RECT 105.930 310.650 106.330 311.100 ;
        RECT 105.930 310.500 109.880 310.650 ;
        RECT 105.930 310.200 106.330 310.500 ;
        RECT 110.480 310.200 110.630 318.400 ;
        RECT 111.080 310.200 111.230 318.400 ;
        RECT 111.680 310.200 111.830 318.400 ;
        RECT 112.280 310.200 112.430 318.400 ;
        RECT 112.880 310.200 113.030 318.400 ;
        RECT 113.480 310.200 113.630 318.400 ;
        RECT 114.080 310.200 114.230 318.400 ;
        RECT 105.930 309.800 114.230 310.200 ;
        RECT 105.930 309.500 106.330 309.800 ;
        RECT 105.930 309.350 109.880 309.500 ;
        RECT 105.930 308.900 106.330 309.350 ;
        RECT 105.930 308.750 109.880 308.900 ;
        RECT 105.930 308.300 106.330 308.750 ;
        RECT 105.930 308.150 109.880 308.300 ;
        RECT 105.930 307.700 106.330 308.150 ;
        RECT 105.930 307.550 109.880 307.700 ;
        RECT 105.930 307.100 106.330 307.550 ;
        RECT 105.930 306.950 109.880 307.100 ;
        RECT 105.930 306.500 106.330 306.950 ;
        RECT 105.930 306.350 109.880 306.500 ;
        RECT 105.930 305.900 106.330 306.350 ;
        RECT 105.930 305.750 109.880 305.900 ;
        RECT 105.930 305.300 106.330 305.750 ;
        RECT 105.930 305.150 109.880 305.300 ;
        RECT 105.930 304.700 106.330 305.150 ;
        RECT 105.930 304.550 109.880 304.700 ;
        RECT 105.930 304.400 106.330 304.550 ;
        RECT 103.130 304.100 106.330 304.400 ;
        RECT 99.580 303.950 109.880 304.100 ;
        RECT 103.130 303.500 106.330 303.950 ;
        RECT 99.580 303.350 109.880 303.500 ;
        RECT 103.130 302.900 106.330 303.350 ;
        RECT 99.580 302.750 109.880 302.900 ;
        RECT 103.130 302.300 106.330 302.750 ;
        RECT 99.580 302.150 109.880 302.300 ;
        RECT 103.530 301.200 105.930 302.150 ;
        RECT 110.480 301.600 110.630 309.800 ;
        RECT 111.080 301.600 111.230 309.800 ;
        RECT 111.680 301.600 111.830 309.800 ;
        RECT 112.280 301.600 112.430 309.800 ;
        RECT 112.880 301.600 113.030 309.800 ;
        RECT 113.480 301.600 113.630 309.800 ;
        RECT 114.080 301.600 114.230 309.800 ;
        RECT 115.230 310.200 115.380 318.400 ;
        RECT 115.830 310.200 115.980 318.400 ;
        RECT 116.430 310.200 116.580 318.400 ;
        RECT 117.030 310.200 117.180 318.400 ;
        RECT 117.630 310.200 117.780 318.400 ;
        RECT 118.230 310.200 118.380 318.400 ;
        RECT 118.830 310.200 118.980 318.400 ;
        RECT 123.530 317.850 124.730 318.800 ;
        RECT 119.580 317.700 124.730 317.850 ;
        RECT 123.130 317.250 124.730 317.700 ;
        RECT 119.580 317.100 124.730 317.250 ;
        RECT 123.130 316.650 124.730 317.100 ;
        RECT 119.580 316.500 124.730 316.650 ;
        RECT 123.130 316.050 124.730 316.500 ;
        RECT 125.130 316.310 127.130 317.585 ;
        RECT 119.580 315.900 124.730 316.050 ;
        RECT 123.130 315.600 124.730 315.900 ;
        RECT 123.130 315.450 123.530 315.600 ;
        RECT 119.580 315.300 123.530 315.450 ;
        RECT 123.130 314.850 123.530 315.300 ;
        RECT 119.580 314.700 123.530 314.850 ;
        RECT 123.130 314.250 123.530 314.700 ;
        RECT 119.580 314.100 123.530 314.250 ;
        RECT 123.130 313.650 123.530 314.100 ;
        RECT 119.580 313.500 123.530 313.650 ;
        RECT 123.130 313.050 123.530 313.500 ;
        RECT 119.580 312.900 123.530 313.050 ;
        RECT 123.130 312.450 123.530 312.900 ;
        RECT 119.580 312.300 123.530 312.450 ;
        RECT 123.130 311.850 123.530 312.300 ;
        RECT 119.580 311.700 123.530 311.850 ;
        RECT 123.130 311.250 123.530 311.700 ;
        RECT 119.580 311.100 123.530 311.250 ;
        RECT 123.130 310.650 123.530 311.100 ;
        RECT 119.580 310.500 123.530 310.650 ;
        RECT 123.130 310.200 123.530 310.500 ;
        RECT 115.230 309.800 123.530 310.200 ;
        RECT 115.230 301.600 115.380 309.800 ;
        RECT 115.830 301.600 115.980 309.800 ;
        RECT 116.430 301.600 116.580 309.800 ;
        RECT 117.030 301.600 117.180 309.800 ;
        RECT 117.630 301.600 117.780 309.800 ;
        RECT 118.230 301.600 118.380 309.800 ;
        RECT 118.830 301.600 118.980 309.800 ;
        RECT 123.130 309.500 123.530 309.800 ;
        RECT 119.580 309.350 123.530 309.500 ;
        RECT 123.130 308.900 123.530 309.350 ;
        RECT 119.580 308.750 123.530 308.900 ;
        RECT 123.130 308.300 123.530 308.750 ;
        RECT 119.580 308.150 123.530 308.300 ;
        RECT 123.130 307.700 123.530 308.150 ;
        RECT 119.580 307.550 123.530 307.700 ;
        RECT 123.130 307.100 123.530 307.550 ;
        RECT 119.580 306.950 123.530 307.100 ;
        RECT 123.130 306.500 123.530 306.950 ;
        RECT 119.580 306.350 123.530 306.500 ;
        RECT 123.130 305.900 123.530 306.350 ;
        RECT 119.580 305.750 123.530 305.900 ;
        RECT 123.130 305.300 123.530 305.750 ;
        RECT 119.580 305.150 123.530 305.300 ;
        RECT 123.130 304.700 123.530 305.150 ;
        RECT 119.580 304.550 123.530 304.700 ;
        RECT 123.130 304.400 123.530 304.550 ;
        RECT 123.130 304.100 124.730 304.400 ;
        RECT 119.580 303.950 124.730 304.100 ;
        RECT 123.130 303.500 124.730 303.950 ;
        RECT 119.580 303.350 124.730 303.500 ;
        RECT 123.130 302.900 124.730 303.350 ;
        RECT 119.580 302.750 124.730 302.900 ;
        RECT 123.130 302.300 124.730 302.750 ;
        RECT 125.140 302.325 127.140 303.600 ;
        RECT 119.580 302.150 124.730 302.300 ;
        RECT 123.530 301.200 124.730 302.150 ;
        RECT 4.730 298.800 9.130 301.200 ;
        RECT 20.330 298.800 29.130 301.200 ;
        RECT 40.330 298.800 49.130 301.200 ;
        RECT 60.330 298.800 69.130 301.200 ;
        RECT 80.330 298.800 89.130 301.200 ;
        RECT 100.330 298.800 109.130 301.200 ;
        RECT 120.330 298.800 124.730 301.200 ;
        RECT 4.730 297.850 5.940 298.800 ;
        RECT 2.315 296.510 4.320 297.785 ;
        RECT 4.730 297.700 9.880 297.850 ;
        RECT 4.730 297.250 6.330 297.700 ;
        RECT 4.730 297.100 9.880 297.250 ;
        RECT 4.730 296.650 6.330 297.100 ;
        RECT 4.730 296.500 9.880 296.650 ;
        RECT 4.730 296.050 6.330 296.500 ;
        RECT 4.730 295.900 9.880 296.050 ;
        RECT 4.730 295.600 6.330 295.900 ;
        RECT 2.320 295.340 4.320 295.545 ;
        RECT 2.315 293.250 4.320 295.340 ;
        RECT 5.930 295.450 6.330 295.600 ;
        RECT 5.930 295.300 9.880 295.450 ;
        RECT 5.930 294.850 6.330 295.300 ;
        RECT 5.930 294.700 9.880 294.850 ;
        RECT 5.930 294.250 6.330 294.700 ;
        RECT 5.930 294.100 9.880 294.250 ;
        RECT 5.930 293.650 6.330 294.100 ;
        RECT 5.930 293.500 9.880 293.650 ;
        RECT 5.930 293.050 6.330 293.500 ;
        RECT 5.930 292.900 9.880 293.050 ;
        RECT 5.930 292.450 6.330 292.900 ;
        RECT 5.930 292.300 9.880 292.450 ;
        RECT 5.930 291.850 6.330 292.300 ;
        RECT 5.930 291.700 9.880 291.850 ;
        RECT 5.930 291.250 6.330 291.700 ;
        RECT 5.930 291.100 9.880 291.250 ;
        RECT 5.930 290.650 6.330 291.100 ;
        RECT 5.930 290.500 9.880 290.650 ;
        RECT 5.930 290.200 6.330 290.500 ;
        RECT 10.480 290.200 10.630 298.400 ;
        RECT 11.080 290.200 11.230 298.400 ;
        RECT 11.680 290.200 11.830 298.400 ;
        RECT 12.280 290.200 12.430 298.400 ;
        RECT 12.880 290.200 13.030 298.400 ;
        RECT 13.480 290.200 13.630 298.400 ;
        RECT 14.080 290.200 14.230 298.400 ;
        RECT 5.930 289.800 14.230 290.200 ;
        RECT 5.930 289.500 6.330 289.800 ;
        RECT 5.930 289.350 9.880 289.500 ;
        RECT 5.930 288.900 6.330 289.350 ;
        RECT 5.930 288.750 9.880 288.900 ;
        RECT 5.930 288.300 6.330 288.750 ;
        RECT 5.930 288.150 9.880 288.300 ;
        RECT 5.930 287.700 6.330 288.150 ;
        RECT 5.930 287.550 9.880 287.700 ;
        RECT 5.930 287.100 6.330 287.550 ;
        RECT 5.930 286.950 9.880 287.100 ;
        RECT 2.315 284.455 4.315 286.750 ;
        RECT 5.930 286.500 6.330 286.950 ;
        RECT 5.930 286.350 9.880 286.500 ;
        RECT 5.930 285.900 6.330 286.350 ;
        RECT 5.930 285.750 9.880 285.900 ;
        RECT 5.930 285.300 6.330 285.750 ;
        RECT 5.930 285.150 9.880 285.300 ;
        RECT 5.930 284.700 6.330 285.150 ;
        RECT 5.930 284.550 9.880 284.700 ;
        RECT 5.930 284.400 6.330 284.550 ;
        RECT 4.730 284.100 6.330 284.400 ;
        RECT 4.730 283.950 9.880 284.100 ;
        RECT 2.315 282.270 4.330 283.545 ;
        RECT 4.730 283.500 6.330 283.950 ;
        RECT 4.730 283.350 9.880 283.500 ;
        RECT 4.730 282.900 6.330 283.350 ;
        RECT 4.730 282.750 9.880 282.900 ;
        RECT 4.730 282.300 6.330 282.750 ;
        RECT 4.730 282.150 9.880 282.300 ;
        RECT 4.730 281.200 5.930 282.150 ;
        RECT 10.480 281.600 10.630 289.800 ;
        RECT 11.080 281.600 11.230 289.800 ;
        RECT 11.680 281.600 11.830 289.800 ;
        RECT 12.280 281.600 12.430 289.800 ;
        RECT 12.880 281.600 13.030 289.800 ;
        RECT 13.480 281.600 13.630 289.800 ;
        RECT 14.080 281.600 14.230 289.800 ;
        RECT 15.230 290.200 15.380 298.400 ;
        RECT 15.830 290.200 15.980 298.400 ;
        RECT 16.430 290.200 16.580 298.400 ;
        RECT 17.030 290.200 17.180 298.400 ;
        RECT 17.630 290.200 17.780 298.400 ;
        RECT 18.230 290.200 18.380 298.400 ;
        RECT 18.830 290.200 18.980 298.400 ;
        RECT 23.530 297.850 25.940 298.800 ;
        RECT 19.580 297.700 29.880 297.850 ;
        RECT 23.130 297.250 26.330 297.700 ;
        RECT 19.580 297.100 29.880 297.250 ;
        RECT 23.130 296.650 26.330 297.100 ;
        RECT 19.580 296.500 29.880 296.650 ;
        RECT 23.130 296.050 26.330 296.500 ;
        RECT 19.580 295.900 29.880 296.050 ;
        RECT 23.130 295.600 26.330 295.900 ;
        RECT 23.130 295.450 23.530 295.600 ;
        RECT 19.580 295.300 23.530 295.450 ;
        RECT 23.130 294.850 23.530 295.300 ;
        RECT 19.580 294.700 23.530 294.850 ;
        RECT 23.130 294.250 23.530 294.700 ;
        RECT 19.580 294.100 23.530 294.250 ;
        RECT 23.130 293.650 23.530 294.100 ;
        RECT 19.580 293.500 23.530 293.650 ;
        RECT 23.130 293.050 23.530 293.500 ;
        RECT 19.580 292.900 23.530 293.050 ;
        RECT 23.130 292.450 23.530 292.900 ;
        RECT 19.580 292.300 23.530 292.450 ;
        RECT 23.130 291.850 23.530 292.300 ;
        RECT 19.580 291.700 23.530 291.850 ;
        RECT 23.130 291.250 23.530 291.700 ;
        RECT 19.580 291.100 23.530 291.250 ;
        RECT 23.130 290.650 23.530 291.100 ;
        RECT 19.580 290.500 23.530 290.650 ;
        RECT 23.130 290.200 23.530 290.500 ;
        RECT 15.230 289.800 23.530 290.200 ;
        RECT 15.230 281.600 15.380 289.800 ;
        RECT 15.830 281.600 15.980 289.800 ;
        RECT 16.430 281.600 16.580 289.800 ;
        RECT 17.030 281.600 17.180 289.800 ;
        RECT 17.630 281.600 17.780 289.800 ;
        RECT 18.230 281.600 18.380 289.800 ;
        RECT 18.830 281.600 18.980 289.800 ;
        RECT 23.130 289.500 23.530 289.800 ;
        RECT 19.580 289.350 23.530 289.500 ;
        RECT 23.130 288.900 23.530 289.350 ;
        RECT 19.580 288.750 23.530 288.900 ;
        RECT 23.130 288.300 23.530 288.750 ;
        RECT 19.580 288.150 23.530 288.300 ;
        RECT 23.130 287.700 23.530 288.150 ;
        RECT 19.580 287.550 23.530 287.700 ;
        RECT 23.130 287.100 23.530 287.550 ;
        RECT 19.580 286.950 23.530 287.100 ;
        RECT 23.130 286.500 23.530 286.950 ;
        RECT 19.580 286.350 23.530 286.500 ;
        RECT 23.130 285.900 23.530 286.350 ;
        RECT 19.580 285.750 23.530 285.900 ;
        RECT 23.130 285.300 23.530 285.750 ;
        RECT 19.580 285.150 23.530 285.300 ;
        RECT 23.130 284.700 23.530 285.150 ;
        RECT 19.580 284.550 23.530 284.700 ;
        RECT 23.130 284.400 23.530 284.550 ;
        RECT 25.930 295.450 26.330 295.600 ;
        RECT 25.930 295.300 29.880 295.450 ;
        RECT 25.930 294.850 26.330 295.300 ;
        RECT 25.930 294.700 29.880 294.850 ;
        RECT 25.930 294.250 26.330 294.700 ;
        RECT 25.930 294.100 29.880 294.250 ;
        RECT 25.930 293.650 26.330 294.100 ;
        RECT 25.930 293.500 29.880 293.650 ;
        RECT 25.930 293.050 26.330 293.500 ;
        RECT 25.930 292.900 29.880 293.050 ;
        RECT 25.930 292.450 26.330 292.900 ;
        RECT 25.930 292.300 29.880 292.450 ;
        RECT 25.930 291.850 26.330 292.300 ;
        RECT 25.930 291.700 29.880 291.850 ;
        RECT 25.930 291.250 26.330 291.700 ;
        RECT 25.930 291.100 29.880 291.250 ;
        RECT 25.930 290.650 26.330 291.100 ;
        RECT 25.930 290.500 29.880 290.650 ;
        RECT 25.930 290.200 26.330 290.500 ;
        RECT 30.480 290.200 30.630 298.400 ;
        RECT 31.080 290.200 31.230 298.400 ;
        RECT 31.680 290.200 31.830 298.400 ;
        RECT 32.280 290.200 32.430 298.400 ;
        RECT 32.880 290.200 33.030 298.400 ;
        RECT 33.480 290.200 33.630 298.400 ;
        RECT 34.080 290.200 34.230 298.400 ;
        RECT 25.930 289.800 34.230 290.200 ;
        RECT 25.930 289.500 26.330 289.800 ;
        RECT 25.930 289.350 29.880 289.500 ;
        RECT 25.930 288.900 26.330 289.350 ;
        RECT 25.930 288.750 29.880 288.900 ;
        RECT 25.930 288.300 26.330 288.750 ;
        RECT 25.930 288.150 29.880 288.300 ;
        RECT 25.930 287.700 26.330 288.150 ;
        RECT 25.930 287.550 29.880 287.700 ;
        RECT 25.930 287.100 26.330 287.550 ;
        RECT 25.930 286.950 29.880 287.100 ;
        RECT 25.930 286.500 26.330 286.950 ;
        RECT 25.930 286.350 29.880 286.500 ;
        RECT 25.930 285.900 26.330 286.350 ;
        RECT 25.930 285.750 29.880 285.900 ;
        RECT 25.930 285.300 26.330 285.750 ;
        RECT 25.930 285.150 29.880 285.300 ;
        RECT 25.930 284.700 26.330 285.150 ;
        RECT 25.930 284.550 29.880 284.700 ;
        RECT 25.930 284.400 26.330 284.550 ;
        RECT 23.130 284.100 26.330 284.400 ;
        RECT 19.580 283.950 29.880 284.100 ;
        RECT 23.130 283.500 26.330 283.950 ;
        RECT 19.580 283.350 29.880 283.500 ;
        RECT 23.130 282.900 26.330 283.350 ;
        RECT 19.580 282.750 29.880 282.900 ;
        RECT 23.130 282.300 26.330 282.750 ;
        RECT 19.580 282.150 29.880 282.300 ;
        RECT 23.530 281.200 25.930 282.150 ;
        RECT 30.480 281.600 30.630 289.800 ;
        RECT 31.080 281.600 31.230 289.800 ;
        RECT 31.680 281.600 31.830 289.800 ;
        RECT 32.280 281.600 32.430 289.800 ;
        RECT 32.880 281.600 33.030 289.800 ;
        RECT 33.480 281.600 33.630 289.800 ;
        RECT 34.080 281.600 34.230 289.800 ;
        RECT 35.230 290.200 35.380 298.400 ;
        RECT 35.830 290.200 35.980 298.400 ;
        RECT 36.430 290.200 36.580 298.400 ;
        RECT 37.030 290.200 37.180 298.400 ;
        RECT 37.630 290.200 37.780 298.400 ;
        RECT 38.230 290.200 38.380 298.400 ;
        RECT 38.830 290.200 38.980 298.400 ;
        RECT 43.530 297.850 45.940 298.800 ;
        RECT 39.580 297.700 49.880 297.850 ;
        RECT 43.130 297.250 46.330 297.700 ;
        RECT 39.580 297.100 49.880 297.250 ;
        RECT 43.130 296.650 46.330 297.100 ;
        RECT 39.580 296.500 49.880 296.650 ;
        RECT 43.130 296.050 46.330 296.500 ;
        RECT 39.580 295.900 49.880 296.050 ;
        RECT 43.130 295.600 46.330 295.900 ;
        RECT 43.130 295.450 43.530 295.600 ;
        RECT 39.580 295.300 43.530 295.450 ;
        RECT 43.130 294.850 43.530 295.300 ;
        RECT 39.580 294.700 43.530 294.850 ;
        RECT 43.130 294.250 43.530 294.700 ;
        RECT 39.580 294.100 43.530 294.250 ;
        RECT 43.130 293.650 43.530 294.100 ;
        RECT 39.580 293.500 43.530 293.650 ;
        RECT 43.130 293.050 43.530 293.500 ;
        RECT 39.580 292.900 43.530 293.050 ;
        RECT 43.130 292.450 43.530 292.900 ;
        RECT 39.580 292.300 43.530 292.450 ;
        RECT 43.130 291.850 43.530 292.300 ;
        RECT 39.580 291.700 43.530 291.850 ;
        RECT 43.130 291.250 43.530 291.700 ;
        RECT 39.580 291.100 43.530 291.250 ;
        RECT 43.130 290.650 43.530 291.100 ;
        RECT 39.580 290.500 43.530 290.650 ;
        RECT 43.130 290.200 43.530 290.500 ;
        RECT 35.230 289.800 43.530 290.200 ;
        RECT 35.230 281.600 35.380 289.800 ;
        RECT 35.830 281.600 35.980 289.800 ;
        RECT 36.430 281.600 36.580 289.800 ;
        RECT 37.030 281.600 37.180 289.800 ;
        RECT 37.630 281.600 37.780 289.800 ;
        RECT 38.230 281.600 38.380 289.800 ;
        RECT 38.830 281.600 38.980 289.800 ;
        RECT 43.130 289.500 43.530 289.800 ;
        RECT 39.580 289.350 43.530 289.500 ;
        RECT 43.130 288.900 43.530 289.350 ;
        RECT 39.580 288.750 43.530 288.900 ;
        RECT 43.130 288.300 43.530 288.750 ;
        RECT 39.580 288.150 43.530 288.300 ;
        RECT 43.130 287.700 43.530 288.150 ;
        RECT 39.580 287.550 43.530 287.700 ;
        RECT 43.130 287.100 43.530 287.550 ;
        RECT 39.580 286.950 43.530 287.100 ;
        RECT 43.130 286.500 43.530 286.950 ;
        RECT 39.580 286.350 43.530 286.500 ;
        RECT 43.130 285.900 43.530 286.350 ;
        RECT 39.580 285.750 43.530 285.900 ;
        RECT 43.130 285.300 43.530 285.750 ;
        RECT 39.580 285.150 43.530 285.300 ;
        RECT 43.130 284.700 43.530 285.150 ;
        RECT 39.580 284.550 43.530 284.700 ;
        RECT 43.130 284.400 43.530 284.550 ;
        RECT 45.930 295.450 46.330 295.600 ;
        RECT 45.930 295.300 49.880 295.450 ;
        RECT 45.930 294.850 46.330 295.300 ;
        RECT 45.930 294.700 49.880 294.850 ;
        RECT 45.930 294.250 46.330 294.700 ;
        RECT 45.930 294.100 49.880 294.250 ;
        RECT 45.930 293.650 46.330 294.100 ;
        RECT 45.930 293.500 49.880 293.650 ;
        RECT 45.930 293.050 46.330 293.500 ;
        RECT 45.930 292.900 49.880 293.050 ;
        RECT 45.930 292.450 46.330 292.900 ;
        RECT 45.930 292.300 49.880 292.450 ;
        RECT 45.930 291.850 46.330 292.300 ;
        RECT 45.930 291.700 49.880 291.850 ;
        RECT 45.930 291.250 46.330 291.700 ;
        RECT 45.930 291.100 49.880 291.250 ;
        RECT 45.930 290.650 46.330 291.100 ;
        RECT 45.930 290.500 49.880 290.650 ;
        RECT 45.930 290.200 46.330 290.500 ;
        RECT 50.480 290.200 50.630 298.400 ;
        RECT 51.080 290.200 51.230 298.400 ;
        RECT 51.680 290.200 51.830 298.400 ;
        RECT 52.280 290.200 52.430 298.400 ;
        RECT 52.880 290.200 53.030 298.400 ;
        RECT 53.480 290.200 53.630 298.400 ;
        RECT 54.080 290.200 54.230 298.400 ;
        RECT 45.930 289.800 54.230 290.200 ;
        RECT 45.930 289.500 46.330 289.800 ;
        RECT 45.930 289.350 49.880 289.500 ;
        RECT 45.930 288.900 46.330 289.350 ;
        RECT 45.930 288.750 49.880 288.900 ;
        RECT 45.930 288.300 46.330 288.750 ;
        RECT 45.930 288.150 49.880 288.300 ;
        RECT 45.930 287.700 46.330 288.150 ;
        RECT 45.930 287.550 49.880 287.700 ;
        RECT 45.930 287.100 46.330 287.550 ;
        RECT 45.930 286.950 49.880 287.100 ;
        RECT 45.930 286.500 46.330 286.950 ;
        RECT 45.930 286.350 49.880 286.500 ;
        RECT 45.930 285.900 46.330 286.350 ;
        RECT 45.930 285.750 49.880 285.900 ;
        RECT 45.930 285.300 46.330 285.750 ;
        RECT 45.930 285.150 49.880 285.300 ;
        RECT 45.930 284.700 46.330 285.150 ;
        RECT 45.930 284.550 49.880 284.700 ;
        RECT 45.930 284.400 46.330 284.550 ;
        RECT 43.130 284.100 46.330 284.400 ;
        RECT 39.580 283.950 49.880 284.100 ;
        RECT 43.130 283.500 46.330 283.950 ;
        RECT 39.580 283.350 49.880 283.500 ;
        RECT 43.130 282.900 46.330 283.350 ;
        RECT 39.580 282.750 49.880 282.900 ;
        RECT 43.130 282.300 46.330 282.750 ;
        RECT 39.580 282.150 49.880 282.300 ;
        RECT 43.530 281.200 45.930 282.150 ;
        RECT 50.480 281.600 50.630 289.800 ;
        RECT 51.080 281.600 51.230 289.800 ;
        RECT 51.680 281.600 51.830 289.800 ;
        RECT 52.280 281.600 52.430 289.800 ;
        RECT 52.880 281.600 53.030 289.800 ;
        RECT 53.480 281.600 53.630 289.800 ;
        RECT 54.080 281.600 54.230 289.800 ;
        RECT 55.230 290.200 55.380 298.400 ;
        RECT 55.830 290.200 55.980 298.400 ;
        RECT 56.430 290.200 56.580 298.400 ;
        RECT 57.030 290.200 57.180 298.400 ;
        RECT 57.630 290.200 57.780 298.400 ;
        RECT 58.230 290.200 58.380 298.400 ;
        RECT 58.830 290.200 58.980 298.400 ;
        RECT 63.530 297.850 65.940 298.800 ;
        RECT 59.580 297.700 69.880 297.850 ;
        RECT 63.130 297.250 66.330 297.700 ;
        RECT 59.580 297.100 69.880 297.250 ;
        RECT 63.130 296.650 66.330 297.100 ;
        RECT 59.580 296.500 69.880 296.650 ;
        RECT 63.130 296.050 66.330 296.500 ;
        RECT 59.580 295.900 69.880 296.050 ;
        RECT 63.130 295.600 66.330 295.900 ;
        RECT 63.130 295.450 63.530 295.600 ;
        RECT 59.580 295.300 63.530 295.450 ;
        RECT 63.130 294.850 63.530 295.300 ;
        RECT 59.580 294.700 63.530 294.850 ;
        RECT 63.130 294.250 63.530 294.700 ;
        RECT 59.580 294.100 63.530 294.250 ;
        RECT 63.130 293.650 63.530 294.100 ;
        RECT 59.580 293.500 63.530 293.650 ;
        RECT 63.130 293.050 63.530 293.500 ;
        RECT 59.580 292.900 63.530 293.050 ;
        RECT 63.130 292.450 63.530 292.900 ;
        RECT 59.580 292.300 63.530 292.450 ;
        RECT 63.130 291.850 63.530 292.300 ;
        RECT 59.580 291.700 63.530 291.850 ;
        RECT 63.130 291.250 63.530 291.700 ;
        RECT 59.580 291.100 63.530 291.250 ;
        RECT 63.130 290.650 63.530 291.100 ;
        RECT 59.580 290.500 63.530 290.650 ;
        RECT 63.130 290.200 63.530 290.500 ;
        RECT 55.230 289.800 63.530 290.200 ;
        RECT 55.230 281.600 55.380 289.800 ;
        RECT 55.830 281.600 55.980 289.800 ;
        RECT 56.430 281.600 56.580 289.800 ;
        RECT 57.030 281.600 57.180 289.800 ;
        RECT 57.630 281.600 57.780 289.800 ;
        RECT 58.230 281.600 58.380 289.800 ;
        RECT 58.830 281.600 58.980 289.800 ;
        RECT 63.130 289.500 63.530 289.800 ;
        RECT 59.580 289.350 63.530 289.500 ;
        RECT 63.130 288.900 63.530 289.350 ;
        RECT 59.580 288.750 63.530 288.900 ;
        RECT 63.130 288.300 63.530 288.750 ;
        RECT 59.580 288.150 63.530 288.300 ;
        RECT 63.130 287.700 63.530 288.150 ;
        RECT 59.580 287.550 63.530 287.700 ;
        RECT 63.130 287.100 63.530 287.550 ;
        RECT 59.580 286.950 63.530 287.100 ;
        RECT 63.130 286.500 63.530 286.950 ;
        RECT 59.580 286.350 63.530 286.500 ;
        RECT 63.130 285.900 63.530 286.350 ;
        RECT 59.580 285.750 63.530 285.900 ;
        RECT 63.130 285.300 63.530 285.750 ;
        RECT 59.580 285.150 63.530 285.300 ;
        RECT 63.130 284.700 63.530 285.150 ;
        RECT 59.580 284.550 63.530 284.700 ;
        RECT 63.130 284.400 63.530 284.550 ;
        RECT 65.930 295.450 66.330 295.600 ;
        RECT 65.930 295.300 69.880 295.450 ;
        RECT 65.930 294.850 66.330 295.300 ;
        RECT 65.930 294.700 69.880 294.850 ;
        RECT 65.930 294.250 66.330 294.700 ;
        RECT 65.930 294.100 69.880 294.250 ;
        RECT 65.930 293.650 66.330 294.100 ;
        RECT 65.930 293.500 69.880 293.650 ;
        RECT 65.930 293.050 66.330 293.500 ;
        RECT 65.930 292.900 69.880 293.050 ;
        RECT 65.930 292.450 66.330 292.900 ;
        RECT 65.930 292.300 69.880 292.450 ;
        RECT 65.930 291.850 66.330 292.300 ;
        RECT 65.930 291.700 69.880 291.850 ;
        RECT 65.930 291.250 66.330 291.700 ;
        RECT 65.930 291.100 69.880 291.250 ;
        RECT 65.930 290.650 66.330 291.100 ;
        RECT 65.930 290.500 69.880 290.650 ;
        RECT 65.930 290.200 66.330 290.500 ;
        RECT 70.480 290.200 70.630 298.400 ;
        RECT 71.080 290.200 71.230 298.400 ;
        RECT 71.680 290.200 71.830 298.400 ;
        RECT 72.280 290.200 72.430 298.400 ;
        RECT 72.880 290.200 73.030 298.400 ;
        RECT 73.480 290.200 73.630 298.400 ;
        RECT 74.080 290.200 74.230 298.400 ;
        RECT 65.930 289.800 74.230 290.200 ;
        RECT 65.930 289.500 66.330 289.800 ;
        RECT 65.930 289.350 69.880 289.500 ;
        RECT 65.930 288.900 66.330 289.350 ;
        RECT 65.930 288.750 69.880 288.900 ;
        RECT 65.930 288.300 66.330 288.750 ;
        RECT 65.930 288.150 69.880 288.300 ;
        RECT 65.930 287.700 66.330 288.150 ;
        RECT 65.930 287.550 69.880 287.700 ;
        RECT 65.930 287.100 66.330 287.550 ;
        RECT 65.930 286.950 69.880 287.100 ;
        RECT 65.930 286.500 66.330 286.950 ;
        RECT 65.930 286.350 69.880 286.500 ;
        RECT 65.930 285.900 66.330 286.350 ;
        RECT 65.930 285.750 69.880 285.900 ;
        RECT 65.930 285.300 66.330 285.750 ;
        RECT 65.930 285.150 69.880 285.300 ;
        RECT 65.930 284.700 66.330 285.150 ;
        RECT 65.930 284.550 69.880 284.700 ;
        RECT 65.930 284.400 66.330 284.550 ;
        RECT 63.130 284.100 66.330 284.400 ;
        RECT 59.580 283.950 69.880 284.100 ;
        RECT 63.130 283.500 66.330 283.950 ;
        RECT 59.580 283.350 69.880 283.500 ;
        RECT 63.130 282.900 66.330 283.350 ;
        RECT 59.580 282.750 69.880 282.900 ;
        RECT 63.130 282.300 66.330 282.750 ;
        RECT 59.580 282.150 69.880 282.300 ;
        RECT 63.530 281.200 65.930 282.150 ;
        RECT 70.480 281.600 70.630 289.800 ;
        RECT 71.080 281.600 71.230 289.800 ;
        RECT 71.680 281.600 71.830 289.800 ;
        RECT 72.280 281.600 72.430 289.800 ;
        RECT 72.880 281.600 73.030 289.800 ;
        RECT 73.480 281.600 73.630 289.800 ;
        RECT 74.080 281.600 74.230 289.800 ;
        RECT 75.230 290.200 75.380 298.400 ;
        RECT 75.830 290.200 75.980 298.400 ;
        RECT 76.430 290.200 76.580 298.400 ;
        RECT 77.030 290.200 77.180 298.400 ;
        RECT 77.630 290.200 77.780 298.400 ;
        RECT 78.230 290.200 78.380 298.400 ;
        RECT 78.830 290.200 78.980 298.400 ;
        RECT 83.530 297.850 85.940 298.800 ;
        RECT 79.580 297.700 89.880 297.850 ;
        RECT 83.130 297.250 86.330 297.700 ;
        RECT 79.580 297.100 89.880 297.250 ;
        RECT 83.130 296.650 86.330 297.100 ;
        RECT 79.580 296.500 89.880 296.650 ;
        RECT 83.130 296.050 86.330 296.500 ;
        RECT 79.580 295.900 89.880 296.050 ;
        RECT 83.130 295.600 86.330 295.900 ;
        RECT 83.130 295.450 83.530 295.600 ;
        RECT 79.580 295.300 83.530 295.450 ;
        RECT 83.130 294.850 83.530 295.300 ;
        RECT 79.580 294.700 83.530 294.850 ;
        RECT 83.130 294.250 83.530 294.700 ;
        RECT 79.580 294.100 83.530 294.250 ;
        RECT 83.130 293.650 83.530 294.100 ;
        RECT 79.580 293.500 83.530 293.650 ;
        RECT 83.130 293.050 83.530 293.500 ;
        RECT 79.580 292.900 83.530 293.050 ;
        RECT 83.130 292.450 83.530 292.900 ;
        RECT 79.580 292.300 83.530 292.450 ;
        RECT 83.130 291.850 83.530 292.300 ;
        RECT 79.580 291.700 83.530 291.850 ;
        RECT 83.130 291.250 83.530 291.700 ;
        RECT 79.580 291.100 83.530 291.250 ;
        RECT 83.130 290.650 83.530 291.100 ;
        RECT 79.580 290.500 83.530 290.650 ;
        RECT 83.130 290.200 83.530 290.500 ;
        RECT 75.230 289.800 83.530 290.200 ;
        RECT 75.230 281.600 75.380 289.800 ;
        RECT 75.830 281.600 75.980 289.800 ;
        RECT 76.430 281.600 76.580 289.800 ;
        RECT 77.030 281.600 77.180 289.800 ;
        RECT 77.630 281.600 77.780 289.800 ;
        RECT 78.230 281.600 78.380 289.800 ;
        RECT 78.830 281.600 78.980 289.800 ;
        RECT 83.130 289.500 83.530 289.800 ;
        RECT 79.580 289.350 83.530 289.500 ;
        RECT 83.130 288.900 83.530 289.350 ;
        RECT 79.580 288.750 83.530 288.900 ;
        RECT 83.130 288.300 83.530 288.750 ;
        RECT 79.580 288.150 83.530 288.300 ;
        RECT 83.130 287.700 83.530 288.150 ;
        RECT 79.580 287.550 83.530 287.700 ;
        RECT 83.130 287.100 83.530 287.550 ;
        RECT 79.580 286.950 83.530 287.100 ;
        RECT 83.130 286.500 83.530 286.950 ;
        RECT 79.580 286.350 83.530 286.500 ;
        RECT 83.130 285.900 83.530 286.350 ;
        RECT 79.580 285.750 83.530 285.900 ;
        RECT 83.130 285.300 83.530 285.750 ;
        RECT 79.580 285.150 83.530 285.300 ;
        RECT 83.130 284.700 83.530 285.150 ;
        RECT 79.580 284.550 83.530 284.700 ;
        RECT 83.130 284.400 83.530 284.550 ;
        RECT 85.930 295.450 86.330 295.600 ;
        RECT 85.930 295.300 89.880 295.450 ;
        RECT 85.930 294.850 86.330 295.300 ;
        RECT 85.930 294.700 89.880 294.850 ;
        RECT 85.930 294.250 86.330 294.700 ;
        RECT 85.930 294.100 89.880 294.250 ;
        RECT 85.930 293.650 86.330 294.100 ;
        RECT 85.930 293.500 89.880 293.650 ;
        RECT 85.930 293.050 86.330 293.500 ;
        RECT 85.930 292.900 89.880 293.050 ;
        RECT 85.930 292.450 86.330 292.900 ;
        RECT 85.930 292.300 89.880 292.450 ;
        RECT 85.930 291.850 86.330 292.300 ;
        RECT 85.930 291.700 89.880 291.850 ;
        RECT 85.930 291.250 86.330 291.700 ;
        RECT 85.930 291.100 89.880 291.250 ;
        RECT 85.930 290.650 86.330 291.100 ;
        RECT 85.930 290.500 89.880 290.650 ;
        RECT 85.930 290.200 86.330 290.500 ;
        RECT 90.480 290.200 90.630 298.400 ;
        RECT 91.080 290.200 91.230 298.400 ;
        RECT 91.680 290.200 91.830 298.400 ;
        RECT 92.280 290.200 92.430 298.400 ;
        RECT 92.880 290.200 93.030 298.400 ;
        RECT 93.480 290.200 93.630 298.400 ;
        RECT 94.080 290.200 94.230 298.400 ;
        RECT 85.930 289.800 94.230 290.200 ;
        RECT 85.930 289.500 86.330 289.800 ;
        RECT 85.930 289.350 89.880 289.500 ;
        RECT 85.930 288.900 86.330 289.350 ;
        RECT 85.930 288.750 89.880 288.900 ;
        RECT 85.930 288.300 86.330 288.750 ;
        RECT 85.930 288.150 89.880 288.300 ;
        RECT 85.930 287.700 86.330 288.150 ;
        RECT 85.930 287.550 89.880 287.700 ;
        RECT 85.930 287.100 86.330 287.550 ;
        RECT 85.930 286.950 89.880 287.100 ;
        RECT 85.930 286.500 86.330 286.950 ;
        RECT 85.930 286.350 89.880 286.500 ;
        RECT 85.930 285.900 86.330 286.350 ;
        RECT 85.930 285.750 89.880 285.900 ;
        RECT 85.930 285.300 86.330 285.750 ;
        RECT 85.930 285.150 89.880 285.300 ;
        RECT 85.930 284.700 86.330 285.150 ;
        RECT 85.930 284.550 89.880 284.700 ;
        RECT 85.930 284.400 86.330 284.550 ;
        RECT 83.130 284.100 86.330 284.400 ;
        RECT 79.580 283.950 89.880 284.100 ;
        RECT 83.130 283.500 86.330 283.950 ;
        RECT 79.580 283.350 89.880 283.500 ;
        RECT 83.130 282.900 86.330 283.350 ;
        RECT 79.580 282.750 89.880 282.900 ;
        RECT 83.130 282.300 86.330 282.750 ;
        RECT 79.580 282.150 89.880 282.300 ;
        RECT 83.530 281.200 85.930 282.150 ;
        RECT 90.480 281.600 90.630 289.800 ;
        RECT 91.080 281.600 91.230 289.800 ;
        RECT 91.680 281.600 91.830 289.800 ;
        RECT 92.280 281.600 92.430 289.800 ;
        RECT 92.880 281.600 93.030 289.800 ;
        RECT 93.480 281.600 93.630 289.800 ;
        RECT 94.080 281.600 94.230 289.800 ;
        RECT 95.230 290.200 95.380 298.400 ;
        RECT 95.830 290.200 95.980 298.400 ;
        RECT 96.430 290.200 96.580 298.400 ;
        RECT 97.030 290.200 97.180 298.400 ;
        RECT 97.630 290.200 97.780 298.400 ;
        RECT 98.230 290.200 98.380 298.400 ;
        RECT 98.830 290.200 98.980 298.400 ;
        RECT 103.530 297.850 105.940 298.800 ;
        RECT 99.580 297.700 109.880 297.850 ;
        RECT 103.130 297.250 106.330 297.700 ;
        RECT 99.580 297.100 109.880 297.250 ;
        RECT 103.130 296.650 106.330 297.100 ;
        RECT 99.580 296.500 109.880 296.650 ;
        RECT 103.130 296.050 106.330 296.500 ;
        RECT 99.580 295.900 109.880 296.050 ;
        RECT 103.130 295.600 106.330 295.900 ;
        RECT 103.130 295.450 103.530 295.600 ;
        RECT 99.580 295.300 103.530 295.450 ;
        RECT 103.130 294.850 103.530 295.300 ;
        RECT 99.580 294.700 103.530 294.850 ;
        RECT 103.130 294.250 103.530 294.700 ;
        RECT 99.580 294.100 103.530 294.250 ;
        RECT 103.130 293.650 103.530 294.100 ;
        RECT 99.580 293.500 103.530 293.650 ;
        RECT 103.130 293.050 103.530 293.500 ;
        RECT 99.580 292.900 103.530 293.050 ;
        RECT 103.130 292.450 103.530 292.900 ;
        RECT 99.580 292.300 103.530 292.450 ;
        RECT 103.130 291.850 103.530 292.300 ;
        RECT 99.580 291.700 103.530 291.850 ;
        RECT 103.130 291.250 103.530 291.700 ;
        RECT 99.580 291.100 103.530 291.250 ;
        RECT 103.130 290.650 103.530 291.100 ;
        RECT 99.580 290.500 103.530 290.650 ;
        RECT 103.130 290.200 103.530 290.500 ;
        RECT 95.230 289.800 103.530 290.200 ;
        RECT 95.230 281.600 95.380 289.800 ;
        RECT 95.830 281.600 95.980 289.800 ;
        RECT 96.430 281.600 96.580 289.800 ;
        RECT 97.030 281.600 97.180 289.800 ;
        RECT 97.630 281.600 97.780 289.800 ;
        RECT 98.230 281.600 98.380 289.800 ;
        RECT 98.830 281.600 98.980 289.800 ;
        RECT 103.130 289.500 103.530 289.800 ;
        RECT 99.580 289.350 103.530 289.500 ;
        RECT 103.130 288.900 103.530 289.350 ;
        RECT 99.580 288.750 103.530 288.900 ;
        RECT 103.130 288.300 103.530 288.750 ;
        RECT 99.580 288.150 103.530 288.300 ;
        RECT 103.130 287.700 103.530 288.150 ;
        RECT 99.580 287.550 103.530 287.700 ;
        RECT 103.130 287.100 103.530 287.550 ;
        RECT 99.580 286.950 103.530 287.100 ;
        RECT 103.130 286.500 103.530 286.950 ;
        RECT 99.580 286.350 103.530 286.500 ;
        RECT 103.130 285.900 103.530 286.350 ;
        RECT 99.580 285.750 103.530 285.900 ;
        RECT 103.130 285.300 103.530 285.750 ;
        RECT 99.580 285.150 103.530 285.300 ;
        RECT 103.130 284.700 103.530 285.150 ;
        RECT 99.580 284.550 103.530 284.700 ;
        RECT 103.130 284.400 103.530 284.550 ;
        RECT 105.930 295.450 106.330 295.600 ;
        RECT 105.930 295.300 109.880 295.450 ;
        RECT 105.930 294.850 106.330 295.300 ;
        RECT 105.930 294.700 109.880 294.850 ;
        RECT 105.930 294.250 106.330 294.700 ;
        RECT 105.930 294.100 109.880 294.250 ;
        RECT 105.930 293.650 106.330 294.100 ;
        RECT 105.930 293.500 109.880 293.650 ;
        RECT 105.930 293.050 106.330 293.500 ;
        RECT 105.930 292.900 109.880 293.050 ;
        RECT 105.930 292.450 106.330 292.900 ;
        RECT 105.930 292.300 109.880 292.450 ;
        RECT 105.930 291.850 106.330 292.300 ;
        RECT 105.930 291.700 109.880 291.850 ;
        RECT 105.930 291.250 106.330 291.700 ;
        RECT 105.930 291.100 109.880 291.250 ;
        RECT 105.930 290.650 106.330 291.100 ;
        RECT 105.930 290.500 109.880 290.650 ;
        RECT 105.930 290.200 106.330 290.500 ;
        RECT 110.480 290.200 110.630 298.400 ;
        RECT 111.080 290.200 111.230 298.400 ;
        RECT 111.680 290.200 111.830 298.400 ;
        RECT 112.280 290.200 112.430 298.400 ;
        RECT 112.880 290.200 113.030 298.400 ;
        RECT 113.480 290.200 113.630 298.400 ;
        RECT 114.080 290.200 114.230 298.400 ;
        RECT 105.930 289.800 114.230 290.200 ;
        RECT 105.930 289.500 106.330 289.800 ;
        RECT 105.930 289.350 109.880 289.500 ;
        RECT 105.930 288.900 106.330 289.350 ;
        RECT 105.930 288.750 109.880 288.900 ;
        RECT 105.930 288.300 106.330 288.750 ;
        RECT 105.930 288.150 109.880 288.300 ;
        RECT 105.930 287.700 106.330 288.150 ;
        RECT 105.930 287.550 109.880 287.700 ;
        RECT 105.930 287.100 106.330 287.550 ;
        RECT 105.930 286.950 109.880 287.100 ;
        RECT 105.930 286.500 106.330 286.950 ;
        RECT 105.930 286.350 109.880 286.500 ;
        RECT 105.930 285.900 106.330 286.350 ;
        RECT 105.930 285.750 109.880 285.900 ;
        RECT 105.930 285.300 106.330 285.750 ;
        RECT 105.930 285.150 109.880 285.300 ;
        RECT 105.930 284.700 106.330 285.150 ;
        RECT 105.930 284.550 109.880 284.700 ;
        RECT 105.930 284.400 106.330 284.550 ;
        RECT 103.130 284.100 106.330 284.400 ;
        RECT 99.580 283.950 109.880 284.100 ;
        RECT 103.130 283.500 106.330 283.950 ;
        RECT 99.580 283.350 109.880 283.500 ;
        RECT 103.130 282.900 106.330 283.350 ;
        RECT 99.580 282.750 109.880 282.900 ;
        RECT 103.130 282.300 106.330 282.750 ;
        RECT 99.580 282.150 109.880 282.300 ;
        RECT 103.530 281.200 105.930 282.150 ;
        RECT 110.480 281.600 110.630 289.800 ;
        RECT 111.080 281.600 111.230 289.800 ;
        RECT 111.680 281.600 111.830 289.800 ;
        RECT 112.280 281.600 112.430 289.800 ;
        RECT 112.880 281.600 113.030 289.800 ;
        RECT 113.480 281.600 113.630 289.800 ;
        RECT 114.080 281.600 114.230 289.800 ;
        RECT 115.230 290.200 115.380 298.400 ;
        RECT 115.830 290.200 115.980 298.400 ;
        RECT 116.430 290.200 116.580 298.400 ;
        RECT 117.030 290.200 117.180 298.400 ;
        RECT 117.630 290.200 117.780 298.400 ;
        RECT 118.230 290.200 118.380 298.400 ;
        RECT 118.830 290.200 118.980 298.400 ;
        RECT 123.530 297.850 124.730 298.800 ;
        RECT 119.580 297.700 124.730 297.850 ;
        RECT 123.130 297.250 124.730 297.700 ;
        RECT 119.580 297.100 124.730 297.250 ;
        RECT 123.130 296.650 124.730 297.100 ;
        RECT 119.580 296.500 124.730 296.650 ;
        RECT 123.130 296.050 124.730 296.500 ;
        RECT 125.130 296.310 127.130 297.585 ;
        RECT 119.580 295.900 124.730 296.050 ;
        RECT 123.130 295.600 124.730 295.900 ;
        RECT 123.130 295.450 123.530 295.600 ;
        RECT 119.580 295.300 123.530 295.450 ;
        RECT 123.130 294.850 123.530 295.300 ;
        RECT 119.580 294.700 123.530 294.850 ;
        RECT 123.130 294.250 123.530 294.700 ;
        RECT 119.580 294.100 123.530 294.250 ;
        RECT 123.130 293.650 123.530 294.100 ;
        RECT 119.580 293.500 123.530 293.650 ;
        RECT 123.130 293.050 123.530 293.500 ;
        RECT 119.580 292.900 123.530 293.050 ;
        RECT 123.130 292.450 123.530 292.900 ;
        RECT 119.580 292.300 123.530 292.450 ;
        RECT 123.130 291.850 123.530 292.300 ;
        RECT 119.580 291.700 123.530 291.850 ;
        RECT 123.130 291.250 123.530 291.700 ;
        RECT 119.580 291.100 123.530 291.250 ;
        RECT 123.130 290.650 123.530 291.100 ;
        RECT 119.580 290.500 123.530 290.650 ;
        RECT 123.130 290.200 123.530 290.500 ;
        RECT 115.230 289.800 123.530 290.200 ;
        RECT 115.230 281.600 115.380 289.800 ;
        RECT 115.830 281.600 115.980 289.800 ;
        RECT 116.430 281.600 116.580 289.800 ;
        RECT 117.030 281.600 117.180 289.800 ;
        RECT 117.630 281.600 117.780 289.800 ;
        RECT 118.230 281.600 118.380 289.800 ;
        RECT 118.830 281.600 118.980 289.800 ;
        RECT 123.130 289.500 123.530 289.800 ;
        RECT 119.580 289.350 123.530 289.500 ;
        RECT 123.130 288.900 123.530 289.350 ;
        RECT 119.580 288.750 123.530 288.900 ;
        RECT 123.130 288.300 123.530 288.750 ;
        RECT 119.580 288.150 123.530 288.300 ;
        RECT 123.130 287.700 123.530 288.150 ;
        RECT 119.580 287.550 123.530 287.700 ;
        RECT 123.130 287.100 123.530 287.550 ;
        RECT 119.580 286.950 123.530 287.100 ;
        RECT 123.130 286.500 123.530 286.950 ;
        RECT 119.580 286.350 123.530 286.500 ;
        RECT 123.130 285.900 123.530 286.350 ;
        RECT 119.580 285.750 123.530 285.900 ;
        RECT 123.130 285.300 123.530 285.750 ;
        RECT 119.580 285.150 123.530 285.300 ;
        RECT 123.130 284.700 123.530 285.150 ;
        RECT 119.580 284.550 123.530 284.700 ;
        RECT 123.130 284.400 123.530 284.550 ;
        RECT 123.130 284.100 124.730 284.400 ;
        RECT 119.580 283.950 124.730 284.100 ;
        RECT 123.130 283.500 124.730 283.950 ;
        RECT 119.580 283.350 124.730 283.500 ;
        RECT 123.130 282.900 124.730 283.350 ;
        RECT 119.580 282.750 124.730 282.900 ;
        RECT 123.130 282.300 124.730 282.750 ;
        RECT 125.140 282.325 127.140 283.600 ;
        RECT 119.580 282.150 124.730 282.300 ;
        RECT 123.530 281.200 124.730 282.150 ;
        RECT 4.730 278.800 9.130 281.200 ;
        RECT 20.330 278.800 29.130 281.200 ;
        RECT 40.330 278.800 49.130 281.200 ;
        RECT 60.330 278.800 69.130 281.200 ;
        RECT 80.330 278.800 89.130 281.200 ;
        RECT 100.330 278.800 109.130 281.200 ;
        RECT 120.330 278.800 124.730 281.200 ;
        RECT 4.730 277.850 5.940 278.800 ;
        RECT 4.730 277.700 9.880 277.850 ;
        RECT 2.315 276.255 4.320 277.530 ;
        RECT 4.730 277.250 6.330 277.700 ;
        RECT 4.730 277.100 9.880 277.250 ;
        RECT 4.730 276.650 6.330 277.100 ;
        RECT 4.730 276.500 9.880 276.650 ;
        RECT 4.730 276.050 6.330 276.500 ;
        RECT 4.730 275.900 9.880 276.050 ;
        RECT 4.730 275.600 6.330 275.900 ;
        RECT 2.320 275.340 4.320 275.545 ;
        RECT 2.315 273.250 4.320 275.340 ;
        RECT 5.930 275.450 6.330 275.600 ;
        RECT 5.930 275.300 9.880 275.450 ;
        RECT 5.930 274.850 6.330 275.300 ;
        RECT 5.930 274.700 9.880 274.850 ;
        RECT 5.930 274.250 6.330 274.700 ;
        RECT 5.930 274.100 9.880 274.250 ;
        RECT 5.930 273.650 6.330 274.100 ;
        RECT 5.930 273.500 9.880 273.650 ;
        RECT 5.930 273.050 6.330 273.500 ;
        RECT 5.930 272.900 9.880 273.050 ;
        RECT 5.930 272.450 6.330 272.900 ;
        RECT 5.930 272.300 9.880 272.450 ;
        RECT 5.930 271.850 6.330 272.300 ;
        RECT 5.930 271.700 9.880 271.850 ;
        RECT 5.930 271.250 6.330 271.700 ;
        RECT 5.930 271.100 9.880 271.250 ;
        RECT 5.930 270.650 6.330 271.100 ;
        RECT 5.930 270.500 9.880 270.650 ;
        RECT 5.930 270.200 6.330 270.500 ;
        RECT 10.480 270.200 10.630 278.400 ;
        RECT 11.080 270.200 11.230 278.400 ;
        RECT 11.680 270.200 11.830 278.400 ;
        RECT 12.280 270.200 12.430 278.400 ;
        RECT 12.880 270.200 13.030 278.400 ;
        RECT 13.480 270.200 13.630 278.400 ;
        RECT 14.080 270.200 14.230 278.400 ;
        RECT 5.930 269.800 14.230 270.200 ;
        RECT 5.930 269.500 6.330 269.800 ;
        RECT 5.930 269.350 9.880 269.500 ;
        RECT 5.930 268.900 6.330 269.350 ;
        RECT 5.930 268.750 9.880 268.900 ;
        RECT 5.930 268.300 6.330 268.750 ;
        RECT 5.930 268.150 9.880 268.300 ;
        RECT 5.930 267.700 6.330 268.150 ;
        RECT 5.930 267.550 9.880 267.700 ;
        RECT 5.930 267.100 6.330 267.550 ;
        RECT 5.930 266.950 9.880 267.100 ;
        RECT 2.315 264.445 4.315 266.740 ;
        RECT 5.930 266.500 6.330 266.950 ;
        RECT 5.930 266.350 9.880 266.500 ;
        RECT 5.930 265.900 6.330 266.350 ;
        RECT 5.930 265.750 9.880 265.900 ;
        RECT 5.930 265.300 6.330 265.750 ;
        RECT 5.930 265.150 9.880 265.300 ;
        RECT 5.930 264.700 6.330 265.150 ;
        RECT 5.930 264.550 9.880 264.700 ;
        RECT 5.930 264.400 6.330 264.550 ;
        RECT 4.730 264.100 6.330 264.400 ;
        RECT 4.730 263.950 9.880 264.100 ;
        RECT 2.315 262.370 4.320 263.645 ;
        RECT 4.730 263.500 6.330 263.950 ;
        RECT 4.730 263.350 9.880 263.500 ;
        RECT 4.730 262.900 6.330 263.350 ;
        RECT 4.730 262.750 9.880 262.900 ;
        RECT 4.730 262.300 6.330 262.750 ;
        RECT 4.730 262.150 9.880 262.300 ;
        RECT 4.730 261.200 5.930 262.150 ;
        RECT 10.480 261.600 10.630 269.800 ;
        RECT 11.080 261.600 11.230 269.800 ;
        RECT 11.680 261.600 11.830 269.800 ;
        RECT 12.280 261.600 12.430 269.800 ;
        RECT 12.880 261.600 13.030 269.800 ;
        RECT 13.480 261.600 13.630 269.800 ;
        RECT 14.080 261.600 14.230 269.800 ;
        RECT 15.230 270.200 15.380 278.400 ;
        RECT 15.830 270.200 15.980 278.400 ;
        RECT 16.430 270.200 16.580 278.400 ;
        RECT 17.030 270.200 17.180 278.400 ;
        RECT 17.630 270.200 17.780 278.400 ;
        RECT 18.230 270.200 18.380 278.400 ;
        RECT 18.830 270.200 18.980 278.400 ;
        RECT 23.530 277.850 25.940 278.800 ;
        RECT 19.580 277.700 29.880 277.850 ;
        RECT 23.130 277.250 26.330 277.700 ;
        RECT 19.580 277.100 29.880 277.250 ;
        RECT 23.130 276.650 26.330 277.100 ;
        RECT 19.580 276.500 29.880 276.650 ;
        RECT 23.130 276.050 26.330 276.500 ;
        RECT 19.580 275.900 29.880 276.050 ;
        RECT 23.130 275.600 26.330 275.900 ;
        RECT 23.130 275.450 23.530 275.600 ;
        RECT 19.580 275.300 23.530 275.450 ;
        RECT 23.130 274.850 23.530 275.300 ;
        RECT 19.580 274.700 23.530 274.850 ;
        RECT 23.130 274.250 23.530 274.700 ;
        RECT 19.580 274.100 23.530 274.250 ;
        RECT 23.130 273.650 23.530 274.100 ;
        RECT 19.580 273.500 23.530 273.650 ;
        RECT 23.130 273.050 23.530 273.500 ;
        RECT 19.580 272.900 23.530 273.050 ;
        RECT 23.130 272.450 23.530 272.900 ;
        RECT 19.580 272.300 23.530 272.450 ;
        RECT 23.130 271.850 23.530 272.300 ;
        RECT 19.580 271.700 23.530 271.850 ;
        RECT 23.130 271.250 23.530 271.700 ;
        RECT 19.580 271.100 23.530 271.250 ;
        RECT 23.130 270.650 23.530 271.100 ;
        RECT 19.580 270.500 23.530 270.650 ;
        RECT 23.130 270.200 23.530 270.500 ;
        RECT 15.230 269.800 23.530 270.200 ;
        RECT 15.230 261.600 15.380 269.800 ;
        RECT 15.830 261.600 15.980 269.800 ;
        RECT 16.430 261.600 16.580 269.800 ;
        RECT 17.030 261.600 17.180 269.800 ;
        RECT 17.630 261.600 17.780 269.800 ;
        RECT 18.230 261.600 18.380 269.800 ;
        RECT 18.830 261.600 18.980 269.800 ;
        RECT 23.130 269.500 23.530 269.800 ;
        RECT 19.580 269.350 23.530 269.500 ;
        RECT 23.130 268.900 23.530 269.350 ;
        RECT 19.580 268.750 23.530 268.900 ;
        RECT 23.130 268.300 23.530 268.750 ;
        RECT 19.580 268.150 23.530 268.300 ;
        RECT 23.130 267.700 23.530 268.150 ;
        RECT 19.580 267.550 23.530 267.700 ;
        RECT 23.130 267.100 23.530 267.550 ;
        RECT 19.580 266.950 23.530 267.100 ;
        RECT 23.130 266.500 23.530 266.950 ;
        RECT 19.580 266.350 23.530 266.500 ;
        RECT 23.130 265.900 23.530 266.350 ;
        RECT 19.580 265.750 23.530 265.900 ;
        RECT 23.130 265.300 23.530 265.750 ;
        RECT 19.580 265.150 23.530 265.300 ;
        RECT 23.130 264.700 23.530 265.150 ;
        RECT 19.580 264.550 23.530 264.700 ;
        RECT 23.130 264.400 23.530 264.550 ;
        RECT 25.930 275.450 26.330 275.600 ;
        RECT 25.930 275.300 29.880 275.450 ;
        RECT 25.930 274.850 26.330 275.300 ;
        RECT 25.930 274.700 29.880 274.850 ;
        RECT 25.930 274.250 26.330 274.700 ;
        RECT 25.930 274.100 29.880 274.250 ;
        RECT 25.930 273.650 26.330 274.100 ;
        RECT 25.930 273.500 29.880 273.650 ;
        RECT 25.930 273.050 26.330 273.500 ;
        RECT 25.930 272.900 29.880 273.050 ;
        RECT 25.930 272.450 26.330 272.900 ;
        RECT 25.930 272.300 29.880 272.450 ;
        RECT 25.930 271.850 26.330 272.300 ;
        RECT 25.930 271.700 29.880 271.850 ;
        RECT 25.930 271.250 26.330 271.700 ;
        RECT 25.930 271.100 29.880 271.250 ;
        RECT 25.930 270.650 26.330 271.100 ;
        RECT 25.930 270.500 29.880 270.650 ;
        RECT 25.930 270.200 26.330 270.500 ;
        RECT 30.480 270.200 30.630 278.400 ;
        RECT 31.080 270.200 31.230 278.400 ;
        RECT 31.680 270.200 31.830 278.400 ;
        RECT 32.280 270.200 32.430 278.400 ;
        RECT 32.880 270.200 33.030 278.400 ;
        RECT 33.480 270.200 33.630 278.400 ;
        RECT 34.080 270.200 34.230 278.400 ;
        RECT 25.930 269.800 34.230 270.200 ;
        RECT 25.930 269.500 26.330 269.800 ;
        RECT 25.930 269.350 29.880 269.500 ;
        RECT 25.930 268.900 26.330 269.350 ;
        RECT 25.930 268.750 29.880 268.900 ;
        RECT 25.930 268.300 26.330 268.750 ;
        RECT 25.930 268.150 29.880 268.300 ;
        RECT 25.930 267.700 26.330 268.150 ;
        RECT 25.930 267.550 29.880 267.700 ;
        RECT 25.930 267.100 26.330 267.550 ;
        RECT 25.930 266.950 29.880 267.100 ;
        RECT 25.930 266.500 26.330 266.950 ;
        RECT 25.930 266.350 29.880 266.500 ;
        RECT 25.930 265.900 26.330 266.350 ;
        RECT 25.930 265.750 29.880 265.900 ;
        RECT 25.930 265.300 26.330 265.750 ;
        RECT 25.930 265.150 29.880 265.300 ;
        RECT 25.930 264.700 26.330 265.150 ;
        RECT 25.930 264.550 29.880 264.700 ;
        RECT 25.930 264.400 26.330 264.550 ;
        RECT 23.130 264.100 26.330 264.400 ;
        RECT 19.580 263.950 29.880 264.100 ;
        RECT 23.130 263.500 26.330 263.950 ;
        RECT 19.580 263.350 29.880 263.500 ;
        RECT 23.130 262.900 26.330 263.350 ;
        RECT 19.580 262.750 29.880 262.900 ;
        RECT 23.130 262.300 26.330 262.750 ;
        RECT 19.580 262.150 29.880 262.300 ;
        RECT 23.530 261.200 25.930 262.150 ;
        RECT 30.480 261.600 30.630 269.800 ;
        RECT 31.080 261.600 31.230 269.800 ;
        RECT 31.680 261.600 31.830 269.800 ;
        RECT 32.280 261.600 32.430 269.800 ;
        RECT 32.880 261.600 33.030 269.800 ;
        RECT 33.480 261.600 33.630 269.800 ;
        RECT 34.080 261.600 34.230 269.800 ;
        RECT 35.230 270.200 35.380 278.400 ;
        RECT 35.830 270.200 35.980 278.400 ;
        RECT 36.430 270.200 36.580 278.400 ;
        RECT 37.030 270.200 37.180 278.400 ;
        RECT 37.630 270.200 37.780 278.400 ;
        RECT 38.230 270.200 38.380 278.400 ;
        RECT 38.830 270.200 38.980 278.400 ;
        RECT 43.530 277.850 45.940 278.800 ;
        RECT 39.580 277.700 49.880 277.850 ;
        RECT 43.130 277.250 46.330 277.700 ;
        RECT 39.580 277.100 49.880 277.250 ;
        RECT 43.130 276.650 46.330 277.100 ;
        RECT 39.580 276.500 49.880 276.650 ;
        RECT 43.130 276.050 46.330 276.500 ;
        RECT 39.580 275.900 49.880 276.050 ;
        RECT 43.130 275.600 46.330 275.900 ;
        RECT 43.130 275.450 43.530 275.600 ;
        RECT 39.580 275.300 43.530 275.450 ;
        RECT 43.130 274.850 43.530 275.300 ;
        RECT 39.580 274.700 43.530 274.850 ;
        RECT 43.130 274.250 43.530 274.700 ;
        RECT 39.580 274.100 43.530 274.250 ;
        RECT 43.130 273.650 43.530 274.100 ;
        RECT 39.580 273.500 43.530 273.650 ;
        RECT 43.130 273.050 43.530 273.500 ;
        RECT 39.580 272.900 43.530 273.050 ;
        RECT 43.130 272.450 43.530 272.900 ;
        RECT 39.580 272.300 43.530 272.450 ;
        RECT 43.130 271.850 43.530 272.300 ;
        RECT 39.580 271.700 43.530 271.850 ;
        RECT 43.130 271.250 43.530 271.700 ;
        RECT 39.580 271.100 43.530 271.250 ;
        RECT 43.130 270.650 43.530 271.100 ;
        RECT 39.580 270.500 43.530 270.650 ;
        RECT 43.130 270.200 43.530 270.500 ;
        RECT 35.230 269.800 43.530 270.200 ;
        RECT 35.230 261.600 35.380 269.800 ;
        RECT 35.830 261.600 35.980 269.800 ;
        RECT 36.430 261.600 36.580 269.800 ;
        RECT 37.030 261.600 37.180 269.800 ;
        RECT 37.630 261.600 37.780 269.800 ;
        RECT 38.230 261.600 38.380 269.800 ;
        RECT 38.830 261.600 38.980 269.800 ;
        RECT 43.130 269.500 43.530 269.800 ;
        RECT 39.580 269.350 43.530 269.500 ;
        RECT 43.130 268.900 43.530 269.350 ;
        RECT 39.580 268.750 43.530 268.900 ;
        RECT 43.130 268.300 43.530 268.750 ;
        RECT 39.580 268.150 43.530 268.300 ;
        RECT 43.130 267.700 43.530 268.150 ;
        RECT 39.580 267.550 43.530 267.700 ;
        RECT 43.130 267.100 43.530 267.550 ;
        RECT 39.580 266.950 43.530 267.100 ;
        RECT 43.130 266.500 43.530 266.950 ;
        RECT 39.580 266.350 43.530 266.500 ;
        RECT 43.130 265.900 43.530 266.350 ;
        RECT 39.580 265.750 43.530 265.900 ;
        RECT 43.130 265.300 43.530 265.750 ;
        RECT 39.580 265.150 43.530 265.300 ;
        RECT 43.130 264.700 43.530 265.150 ;
        RECT 39.580 264.550 43.530 264.700 ;
        RECT 43.130 264.400 43.530 264.550 ;
        RECT 45.930 275.450 46.330 275.600 ;
        RECT 45.930 275.300 49.880 275.450 ;
        RECT 45.930 274.850 46.330 275.300 ;
        RECT 45.930 274.700 49.880 274.850 ;
        RECT 45.930 274.250 46.330 274.700 ;
        RECT 45.930 274.100 49.880 274.250 ;
        RECT 45.930 273.650 46.330 274.100 ;
        RECT 45.930 273.500 49.880 273.650 ;
        RECT 45.930 273.050 46.330 273.500 ;
        RECT 45.930 272.900 49.880 273.050 ;
        RECT 45.930 272.450 46.330 272.900 ;
        RECT 45.930 272.300 49.880 272.450 ;
        RECT 45.930 271.850 46.330 272.300 ;
        RECT 45.930 271.700 49.880 271.850 ;
        RECT 45.930 271.250 46.330 271.700 ;
        RECT 45.930 271.100 49.880 271.250 ;
        RECT 45.930 270.650 46.330 271.100 ;
        RECT 45.930 270.500 49.880 270.650 ;
        RECT 45.930 270.200 46.330 270.500 ;
        RECT 50.480 270.200 50.630 278.400 ;
        RECT 51.080 270.200 51.230 278.400 ;
        RECT 51.680 270.200 51.830 278.400 ;
        RECT 52.280 270.200 52.430 278.400 ;
        RECT 52.880 270.200 53.030 278.400 ;
        RECT 53.480 270.200 53.630 278.400 ;
        RECT 54.080 270.200 54.230 278.400 ;
        RECT 45.930 269.800 54.230 270.200 ;
        RECT 45.930 269.500 46.330 269.800 ;
        RECT 45.930 269.350 49.880 269.500 ;
        RECT 45.930 268.900 46.330 269.350 ;
        RECT 45.930 268.750 49.880 268.900 ;
        RECT 45.930 268.300 46.330 268.750 ;
        RECT 45.930 268.150 49.880 268.300 ;
        RECT 45.930 267.700 46.330 268.150 ;
        RECT 45.930 267.550 49.880 267.700 ;
        RECT 45.930 267.100 46.330 267.550 ;
        RECT 45.930 266.950 49.880 267.100 ;
        RECT 45.930 266.500 46.330 266.950 ;
        RECT 45.930 266.350 49.880 266.500 ;
        RECT 45.930 265.900 46.330 266.350 ;
        RECT 45.930 265.750 49.880 265.900 ;
        RECT 45.930 265.300 46.330 265.750 ;
        RECT 45.930 265.150 49.880 265.300 ;
        RECT 45.930 264.700 46.330 265.150 ;
        RECT 45.930 264.550 49.880 264.700 ;
        RECT 45.930 264.400 46.330 264.550 ;
        RECT 43.130 264.100 46.330 264.400 ;
        RECT 39.580 263.950 49.880 264.100 ;
        RECT 43.130 263.500 46.330 263.950 ;
        RECT 39.580 263.350 49.880 263.500 ;
        RECT 43.130 262.900 46.330 263.350 ;
        RECT 39.580 262.750 49.880 262.900 ;
        RECT 43.130 262.300 46.330 262.750 ;
        RECT 39.580 262.150 49.880 262.300 ;
        RECT 43.530 261.200 45.930 262.150 ;
        RECT 50.480 261.600 50.630 269.800 ;
        RECT 51.080 261.600 51.230 269.800 ;
        RECT 51.680 261.600 51.830 269.800 ;
        RECT 52.280 261.600 52.430 269.800 ;
        RECT 52.880 261.600 53.030 269.800 ;
        RECT 53.480 261.600 53.630 269.800 ;
        RECT 54.080 261.600 54.230 269.800 ;
        RECT 55.230 270.200 55.380 278.400 ;
        RECT 55.830 270.200 55.980 278.400 ;
        RECT 56.430 270.200 56.580 278.400 ;
        RECT 57.030 270.200 57.180 278.400 ;
        RECT 57.630 270.200 57.780 278.400 ;
        RECT 58.230 270.200 58.380 278.400 ;
        RECT 58.830 270.200 58.980 278.400 ;
        RECT 63.530 277.850 65.940 278.800 ;
        RECT 59.580 277.700 69.880 277.850 ;
        RECT 63.130 277.250 66.330 277.700 ;
        RECT 59.580 277.100 69.880 277.250 ;
        RECT 63.130 276.650 66.330 277.100 ;
        RECT 59.580 276.500 69.880 276.650 ;
        RECT 63.130 276.050 66.330 276.500 ;
        RECT 59.580 275.900 69.880 276.050 ;
        RECT 63.130 275.600 66.330 275.900 ;
        RECT 63.130 275.450 63.530 275.600 ;
        RECT 59.580 275.300 63.530 275.450 ;
        RECT 63.130 274.850 63.530 275.300 ;
        RECT 59.580 274.700 63.530 274.850 ;
        RECT 63.130 274.250 63.530 274.700 ;
        RECT 59.580 274.100 63.530 274.250 ;
        RECT 63.130 273.650 63.530 274.100 ;
        RECT 59.580 273.500 63.530 273.650 ;
        RECT 63.130 273.050 63.530 273.500 ;
        RECT 59.580 272.900 63.530 273.050 ;
        RECT 63.130 272.450 63.530 272.900 ;
        RECT 59.580 272.300 63.530 272.450 ;
        RECT 63.130 271.850 63.530 272.300 ;
        RECT 59.580 271.700 63.530 271.850 ;
        RECT 63.130 271.250 63.530 271.700 ;
        RECT 59.580 271.100 63.530 271.250 ;
        RECT 63.130 270.650 63.530 271.100 ;
        RECT 59.580 270.500 63.530 270.650 ;
        RECT 63.130 270.200 63.530 270.500 ;
        RECT 55.230 269.800 63.530 270.200 ;
        RECT 55.230 261.600 55.380 269.800 ;
        RECT 55.830 261.600 55.980 269.800 ;
        RECT 56.430 261.600 56.580 269.800 ;
        RECT 57.030 261.600 57.180 269.800 ;
        RECT 57.630 261.600 57.780 269.800 ;
        RECT 58.230 261.600 58.380 269.800 ;
        RECT 58.830 261.600 58.980 269.800 ;
        RECT 63.130 269.500 63.530 269.800 ;
        RECT 59.580 269.350 63.530 269.500 ;
        RECT 63.130 268.900 63.530 269.350 ;
        RECT 59.580 268.750 63.530 268.900 ;
        RECT 63.130 268.300 63.530 268.750 ;
        RECT 59.580 268.150 63.530 268.300 ;
        RECT 63.130 267.700 63.530 268.150 ;
        RECT 59.580 267.550 63.530 267.700 ;
        RECT 63.130 267.100 63.530 267.550 ;
        RECT 59.580 266.950 63.530 267.100 ;
        RECT 63.130 266.500 63.530 266.950 ;
        RECT 59.580 266.350 63.530 266.500 ;
        RECT 63.130 265.900 63.530 266.350 ;
        RECT 59.580 265.750 63.530 265.900 ;
        RECT 63.130 265.300 63.530 265.750 ;
        RECT 59.580 265.150 63.530 265.300 ;
        RECT 63.130 264.700 63.530 265.150 ;
        RECT 59.580 264.550 63.530 264.700 ;
        RECT 63.130 264.400 63.530 264.550 ;
        RECT 65.930 275.450 66.330 275.600 ;
        RECT 65.930 275.300 69.880 275.450 ;
        RECT 65.930 274.850 66.330 275.300 ;
        RECT 65.930 274.700 69.880 274.850 ;
        RECT 65.930 274.250 66.330 274.700 ;
        RECT 65.930 274.100 69.880 274.250 ;
        RECT 65.930 273.650 66.330 274.100 ;
        RECT 65.930 273.500 69.880 273.650 ;
        RECT 65.930 273.050 66.330 273.500 ;
        RECT 65.930 272.900 69.880 273.050 ;
        RECT 65.930 272.450 66.330 272.900 ;
        RECT 65.930 272.300 69.880 272.450 ;
        RECT 65.930 271.850 66.330 272.300 ;
        RECT 65.930 271.700 69.880 271.850 ;
        RECT 65.930 271.250 66.330 271.700 ;
        RECT 65.930 271.100 69.880 271.250 ;
        RECT 65.930 270.650 66.330 271.100 ;
        RECT 65.930 270.500 69.880 270.650 ;
        RECT 65.930 270.200 66.330 270.500 ;
        RECT 70.480 270.200 70.630 278.400 ;
        RECT 71.080 270.200 71.230 278.400 ;
        RECT 71.680 270.200 71.830 278.400 ;
        RECT 72.280 270.200 72.430 278.400 ;
        RECT 72.880 270.200 73.030 278.400 ;
        RECT 73.480 270.200 73.630 278.400 ;
        RECT 74.080 270.200 74.230 278.400 ;
        RECT 65.930 269.800 74.230 270.200 ;
        RECT 65.930 269.500 66.330 269.800 ;
        RECT 65.930 269.350 69.880 269.500 ;
        RECT 65.930 268.900 66.330 269.350 ;
        RECT 65.930 268.750 69.880 268.900 ;
        RECT 65.930 268.300 66.330 268.750 ;
        RECT 65.930 268.150 69.880 268.300 ;
        RECT 65.930 267.700 66.330 268.150 ;
        RECT 65.930 267.550 69.880 267.700 ;
        RECT 65.930 267.100 66.330 267.550 ;
        RECT 65.930 266.950 69.880 267.100 ;
        RECT 65.930 266.500 66.330 266.950 ;
        RECT 65.930 266.350 69.880 266.500 ;
        RECT 65.930 265.900 66.330 266.350 ;
        RECT 65.930 265.750 69.880 265.900 ;
        RECT 65.930 265.300 66.330 265.750 ;
        RECT 65.930 265.150 69.880 265.300 ;
        RECT 65.930 264.700 66.330 265.150 ;
        RECT 65.930 264.550 69.880 264.700 ;
        RECT 65.930 264.400 66.330 264.550 ;
        RECT 63.130 264.100 66.330 264.400 ;
        RECT 59.580 263.950 69.880 264.100 ;
        RECT 63.130 263.500 66.330 263.950 ;
        RECT 59.580 263.350 69.880 263.500 ;
        RECT 63.130 262.900 66.330 263.350 ;
        RECT 59.580 262.750 69.880 262.900 ;
        RECT 63.130 262.300 66.330 262.750 ;
        RECT 59.580 262.150 69.880 262.300 ;
        RECT 63.530 261.200 65.930 262.150 ;
        RECT 70.480 261.600 70.630 269.800 ;
        RECT 71.080 261.600 71.230 269.800 ;
        RECT 71.680 261.600 71.830 269.800 ;
        RECT 72.280 261.600 72.430 269.800 ;
        RECT 72.880 261.600 73.030 269.800 ;
        RECT 73.480 261.600 73.630 269.800 ;
        RECT 74.080 261.600 74.230 269.800 ;
        RECT 75.230 270.200 75.380 278.400 ;
        RECT 75.830 270.200 75.980 278.400 ;
        RECT 76.430 270.200 76.580 278.400 ;
        RECT 77.030 270.200 77.180 278.400 ;
        RECT 77.630 270.200 77.780 278.400 ;
        RECT 78.230 270.200 78.380 278.400 ;
        RECT 78.830 270.200 78.980 278.400 ;
        RECT 83.530 277.850 85.940 278.800 ;
        RECT 79.580 277.700 89.880 277.850 ;
        RECT 83.130 277.250 86.330 277.700 ;
        RECT 79.580 277.100 89.880 277.250 ;
        RECT 83.130 276.650 86.330 277.100 ;
        RECT 79.580 276.500 89.880 276.650 ;
        RECT 83.130 276.050 86.330 276.500 ;
        RECT 79.580 275.900 89.880 276.050 ;
        RECT 83.130 275.600 86.330 275.900 ;
        RECT 83.130 275.450 83.530 275.600 ;
        RECT 79.580 275.300 83.530 275.450 ;
        RECT 83.130 274.850 83.530 275.300 ;
        RECT 79.580 274.700 83.530 274.850 ;
        RECT 83.130 274.250 83.530 274.700 ;
        RECT 79.580 274.100 83.530 274.250 ;
        RECT 83.130 273.650 83.530 274.100 ;
        RECT 79.580 273.500 83.530 273.650 ;
        RECT 83.130 273.050 83.530 273.500 ;
        RECT 79.580 272.900 83.530 273.050 ;
        RECT 83.130 272.450 83.530 272.900 ;
        RECT 79.580 272.300 83.530 272.450 ;
        RECT 83.130 271.850 83.530 272.300 ;
        RECT 79.580 271.700 83.530 271.850 ;
        RECT 83.130 271.250 83.530 271.700 ;
        RECT 79.580 271.100 83.530 271.250 ;
        RECT 83.130 270.650 83.530 271.100 ;
        RECT 79.580 270.500 83.530 270.650 ;
        RECT 83.130 270.200 83.530 270.500 ;
        RECT 75.230 269.800 83.530 270.200 ;
        RECT 75.230 261.600 75.380 269.800 ;
        RECT 75.830 261.600 75.980 269.800 ;
        RECT 76.430 261.600 76.580 269.800 ;
        RECT 77.030 261.600 77.180 269.800 ;
        RECT 77.630 261.600 77.780 269.800 ;
        RECT 78.230 261.600 78.380 269.800 ;
        RECT 78.830 261.600 78.980 269.800 ;
        RECT 83.130 269.500 83.530 269.800 ;
        RECT 79.580 269.350 83.530 269.500 ;
        RECT 83.130 268.900 83.530 269.350 ;
        RECT 79.580 268.750 83.530 268.900 ;
        RECT 83.130 268.300 83.530 268.750 ;
        RECT 79.580 268.150 83.530 268.300 ;
        RECT 83.130 267.700 83.530 268.150 ;
        RECT 79.580 267.550 83.530 267.700 ;
        RECT 83.130 267.100 83.530 267.550 ;
        RECT 79.580 266.950 83.530 267.100 ;
        RECT 83.130 266.500 83.530 266.950 ;
        RECT 79.580 266.350 83.530 266.500 ;
        RECT 83.130 265.900 83.530 266.350 ;
        RECT 79.580 265.750 83.530 265.900 ;
        RECT 83.130 265.300 83.530 265.750 ;
        RECT 79.580 265.150 83.530 265.300 ;
        RECT 83.130 264.700 83.530 265.150 ;
        RECT 79.580 264.550 83.530 264.700 ;
        RECT 83.130 264.400 83.530 264.550 ;
        RECT 85.930 275.450 86.330 275.600 ;
        RECT 85.930 275.300 89.880 275.450 ;
        RECT 85.930 274.850 86.330 275.300 ;
        RECT 85.930 274.700 89.880 274.850 ;
        RECT 85.930 274.250 86.330 274.700 ;
        RECT 85.930 274.100 89.880 274.250 ;
        RECT 85.930 273.650 86.330 274.100 ;
        RECT 85.930 273.500 89.880 273.650 ;
        RECT 85.930 273.050 86.330 273.500 ;
        RECT 85.930 272.900 89.880 273.050 ;
        RECT 85.930 272.450 86.330 272.900 ;
        RECT 85.930 272.300 89.880 272.450 ;
        RECT 85.930 271.850 86.330 272.300 ;
        RECT 85.930 271.700 89.880 271.850 ;
        RECT 85.930 271.250 86.330 271.700 ;
        RECT 85.930 271.100 89.880 271.250 ;
        RECT 85.930 270.650 86.330 271.100 ;
        RECT 85.930 270.500 89.880 270.650 ;
        RECT 85.930 270.200 86.330 270.500 ;
        RECT 90.480 270.200 90.630 278.400 ;
        RECT 91.080 270.200 91.230 278.400 ;
        RECT 91.680 270.200 91.830 278.400 ;
        RECT 92.280 270.200 92.430 278.400 ;
        RECT 92.880 270.200 93.030 278.400 ;
        RECT 93.480 270.200 93.630 278.400 ;
        RECT 94.080 270.200 94.230 278.400 ;
        RECT 85.930 269.800 94.230 270.200 ;
        RECT 85.930 269.500 86.330 269.800 ;
        RECT 85.930 269.350 89.880 269.500 ;
        RECT 85.930 268.900 86.330 269.350 ;
        RECT 85.930 268.750 89.880 268.900 ;
        RECT 85.930 268.300 86.330 268.750 ;
        RECT 85.930 268.150 89.880 268.300 ;
        RECT 85.930 267.700 86.330 268.150 ;
        RECT 85.930 267.550 89.880 267.700 ;
        RECT 85.930 267.100 86.330 267.550 ;
        RECT 85.930 266.950 89.880 267.100 ;
        RECT 85.930 266.500 86.330 266.950 ;
        RECT 85.930 266.350 89.880 266.500 ;
        RECT 85.930 265.900 86.330 266.350 ;
        RECT 85.930 265.750 89.880 265.900 ;
        RECT 85.930 265.300 86.330 265.750 ;
        RECT 85.930 265.150 89.880 265.300 ;
        RECT 85.930 264.700 86.330 265.150 ;
        RECT 85.930 264.550 89.880 264.700 ;
        RECT 85.930 264.400 86.330 264.550 ;
        RECT 83.130 264.100 86.330 264.400 ;
        RECT 79.580 263.950 89.880 264.100 ;
        RECT 83.130 263.500 86.330 263.950 ;
        RECT 79.580 263.350 89.880 263.500 ;
        RECT 83.130 262.900 86.330 263.350 ;
        RECT 79.580 262.750 89.880 262.900 ;
        RECT 83.130 262.300 86.330 262.750 ;
        RECT 79.580 262.150 89.880 262.300 ;
        RECT 83.530 261.200 85.930 262.150 ;
        RECT 90.480 261.600 90.630 269.800 ;
        RECT 91.080 261.600 91.230 269.800 ;
        RECT 91.680 261.600 91.830 269.800 ;
        RECT 92.280 261.600 92.430 269.800 ;
        RECT 92.880 261.600 93.030 269.800 ;
        RECT 93.480 261.600 93.630 269.800 ;
        RECT 94.080 261.600 94.230 269.800 ;
        RECT 95.230 270.200 95.380 278.400 ;
        RECT 95.830 270.200 95.980 278.400 ;
        RECT 96.430 270.200 96.580 278.400 ;
        RECT 97.030 270.200 97.180 278.400 ;
        RECT 97.630 270.200 97.780 278.400 ;
        RECT 98.230 270.200 98.380 278.400 ;
        RECT 98.830 270.200 98.980 278.400 ;
        RECT 103.530 277.850 105.940 278.800 ;
        RECT 99.580 277.700 109.880 277.850 ;
        RECT 103.130 277.250 106.330 277.700 ;
        RECT 99.580 277.100 109.880 277.250 ;
        RECT 103.130 276.650 106.330 277.100 ;
        RECT 99.580 276.500 109.880 276.650 ;
        RECT 103.130 276.050 106.330 276.500 ;
        RECT 99.580 275.900 109.880 276.050 ;
        RECT 103.130 275.600 106.330 275.900 ;
        RECT 103.130 275.450 103.530 275.600 ;
        RECT 99.580 275.300 103.530 275.450 ;
        RECT 103.130 274.850 103.530 275.300 ;
        RECT 99.580 274.700 103.530 274.850 ;
        RECT 103.130 274.250 103.530 274.700 ;
        RECT 99.580 274.100 103.530 274.250 ;
        RECT 103.130 273.650 103.530 274.100 ;
        RECT 99.580 273.500 103.530 273.650 ;
        RECT 103.130 273.050 103.530 273.500 ;
        RECT 99.580 272.900 103.530 273.050 ;
        RECT 103.130 272.450 103.530 272.900 ;
        RECT 99.580 272.300 103.530 272.450 ;
        RECT 103.130 271.850 103.530 272.300 ;
        RECT 99.580 271.700 103.530 271.850 ;
        RECT 103.130 271.250 103.530 271.700 ;
        RECT 99.580 271.100 103.530 271.250 ;
        RECT 103.130 270.650 103.530 271.100 ;
        RECT 99.580 270.500 103.530 270.650 ;
        RECT 103.130 270.200 103.530 270.500 ;
        RECT 95.230 269.800 103.530 270.200 ;
        RECT 95.230 261.600 95.380 269.800 ;
        RECT 95.830 261.600 95.980 269.800 ;
        RECT 96.430 261.600 96.580 269.800 ;
        RECT 97.030 261.600 97.180 269.800 ;
        RECT 97.630 261.600 97.780 269.800 ;
        RECT 98.230 261.600 98.380 269.800 ;
        RECT 98.830 261.600 98.980 269.800 ;
        RECT 103.130 269.500 103.530 269.800 ;
        RECT 99.580 269.350 103.530 269.500 ;
        RECT 103.130 268.900 103.530 269.350 ;
        RECT 99.580 268.750 103.530 268.900 ;
        RECT 103.130 268.300 103.530 268.750 ;
        RECT 99.580 268.150 103.530 268.300 ;
        RECT 103.130 267.700 103.530 268.150 ;
        RECT 99.580 267.550 103.530 267.700 ;
        RECT 103.130 267.100 103.530 267.550 ;
        RECT 99.580 266.950 103.530 267.100 ;
        RECT 103.130 266.500 103.530 266.950 ;
        RECT 99.580 266.350 103.530 266.500 ;
        RECT 103.130 265.900 103.530 266.350 ;
        RECT 99.580 265.750 103.530 265.900 ;
        RECT 103.130 265.300 103.530 265.750 ;
        RECT 99.580 265.150 103.530 265.300 ;
        RECT 103.130 264.700 103.530 265.150 ;
        RECT 99.580 264.550 103.530 264.700 ;
        RECT 103.130 264.400 103.530 264.550 ;
        RECT 105.930 275.450 106.330 275.600 ;
        RECT 105.930 275.300 109.880 275.450 ;
        RECT 105.930 274.850 106.330 275.300 ;
        RECT 105.930 274.700 109.880 274.850 ;
        RECT 105.930 274.250 106.330 274.700 ;
        RECT 105.930 274.100 109.880 274.250 ;
        RECT 105.930 273.650 106.330 274.100 ;
        RECT 105.930 273.500 109.880 273.650 ;
        RECT 105.930 273.050 106.330 273.500 ;
        RECT 105.930 272.900 109.880 273.050 ;
        RECT 105.930 272.450 106.330 272.900 ;
        RECT 105.930 272.300 109.880 272.450 ;
        RECT 105.930 271.850 106.330 272.300 ;
        RECT 105.930 271.700 109.880 271.850 ;
        RECT 105.930 271.250 106.330 271.700 ;
        RECT 105.930 271.100 109.880 271.250 ;
        RECT 105.930 270.650 106.330 271.100 ;
        RECT 105.930 270.500 109.880 270.650 ;
        RECT 105.930 270.200 106.330 270.500 ;
        RECT 110.480 270.200 110.630 278.400 ;
        RECT 111.080 270.200 111.230 278.400 ;
        RECT 111.680 270.200 111.830 278.400 ;
        RECT 112.280 270.200 112.430 278.400 ;
        RECT 112.880 270.200 113.030 278.400 ;
        RECT 113.480 270.200 113.630 278.400 ;
        RECT 114.080 270.200 114.230 278.400 ;
        RECT 105.930 269.800 114.230 270.200 ;
        RECT 105.930 269.500 106.330 269.800 ;
        RECT 105.930 269.350 109.880 269.500 ;
        RECT 105.930 268.900 106.330 269.350 ;
        RECT 105.930 268.750 109.880 268.900 ;
        RECT 105.930 268.300 106.330 268.750 ;
        RECT 105.930 268.150 109.880 268.300 ;
        RECT 105.930 267.700 106.330 268.150 ;
        RECT 105.930 267.550 109.880 267.700 ;
        RECT 105.930 267.100 106.330 267.550 ;
        RECT 105.930 266.950 109.880 267.100 ;
        RECT 105.930 266.500 106.330 266.950 ;
        RECT 105.930 266.350 109.880 266.500 ;
        RECT 105.930 265.900 106.330 266.350 ;
        RECT 105.930 265.750 109.880 265.900 ;
        RECT 105.930 265.300 106.330 265.750 ;
        RECT 105.930 265.150 109.880 265.300 ;
        RECT 105.930 264.700 106.330 265.150 ;
        RECT 105.930 264.550 109.880 264.700 ;
        RECT 105.930 264.400 106.330 264.550 ;
        RECT 103.130 264.100 106.330 264.400 ;
        RECT 99.580 263.950 109.880 264.100 ;
        RECT 103.130 263.500 106.330 263.950 ;
        RECT 99.580 263.350 109.880 263.500 ;
        RECT 103.130 262.900 106.330 263.350 ;
        RECT 99.580 262.750 109.880 262.900 ;
        RECT 103.130 262.300 106.330 262.750 ;
        RECT 99.580 262.150 109.880 262.300 ;
        RECT 103.530 261.200 105.930 262.150 ;
        RECT 110.480 261.600 110.630 269.800 ;
        RECT 111.080 261.600 111.230 269.800 ;
        RECT 111.680 261.600 111.830 269.800 ;
        RECT 112.280 261.600 112.430 269.800 ;
        RECT 112.880 261.600 113.030 269.800 ;
        RECT 113.480 261.600 113.630 269.800 ;
        RECT 114.080 261.600 114.230 269.800 ;
        RECT 115.230 270.200 115.380 278.400 ;
        RECT 115.830 270.200 115.980 278.400 ;
        RECT 116.430 270.200 116.580 278.400 ;
        RECT 117.030 270.200 117.180 278.400 ;
        RECT 117.630 270.200 117.780 278.400 ;
        RECT 118.230 270.200 118.380 278.400 ;
        RECT 118.830 270.200 118.980 278.400 ;
        RECT 123.530 277.850 124.730 278.800 ;
        RECT 119.580 277.700 124.730 277.850 ;
        RECT 123.130 277.250 124.730 277.700 ;
        RECT 119.580 277.100 124.730 277.250 ;
        RECT 123.130 276.650 124.730 277.100 ;
        RECT 119.580 276.500 124.730 276.650 ;
        RECT 125.135 276.580 127.135 277.855 ;
        RECT 123.130 276.050 124.730 276.500 ;
        RECT 119.580 275.900 124.730 276.050 ;
        RECT 123.130 275.600 124.730 275.900 ;
        RECT 123.130 275.450 123.530 275.600 ;
        RECT 119.580 275.300 123.530 275.450 ;
        RECT 123.130 274.850 123.530 275.300 ;
        RECT 119.580 274.700 123.530 274.850 ;
        RECT 123.130 274.250 123.530 274.700 ;
        RECT 119.580 274.100 123.530 274.250 ;
        RECT 123.130 273.650 123.530 274.100 ;
        RECT 119.580 273.500 123.530 273.650 ;
        RECT 123.130 273.050 123.530 273.500 ;
        RECT 119.580 272.900 123.530 273.050 ;
        RECT 123.130 272.450 123.530 272.900 ;
        RECT 119.580 272.300 123.530 272.450 ;
        RECT 123.130 271.850 123.530 272.300 ;
        RECT 119.580 271.700 123.530 271.850 ;
        RECT 123.130 271.250 123.530 271.700 ;
        RECT 119.580 271.100 123.530 271.250 ;
        RECT 123.130 270.650 123.530 271.100 ;
        RECT 119.580 270.500 123.530 270.650 ;
        RECT 123.130 270.200 123.530 270.500 ;
        RECT 115.230 269.800 123.530 270.200 ;
        RECT 115.230 261.600 115.380 269.800 ;
        RECT 115.830 261.600 115.980 269.800 ;
        RECT 116.430 261.600 116.580 269.800 ;
        RECT 117.030 261.600 117.180 269.800 ;
        RECT 117.630 261.600 117.780 269.800 ;
        RECT 118.230 261.600 118.380 269.800 ;
        RECT 118.830 261.600 118.980 269.800 ;
        RECT 123.130 269.500 123.530 269.800 ;
        RECT 119.580 269.350 123.530 269.500 ;
        RECT 123.130 268.900 123.530 269.350 ;
        RECT 119.580 268.750 123.530 268.900 ;
        RECT 123.130 268.300 123.530 268.750 ;
        RECT 119.580 268.150 123.530 268.300 ;
        RECT 123.130 267.700 123.530 268.150 ;
        RECT 119.580 267.550 123.530 267.700 ;
        RECT 123.130 267.100 123.530 267.550 ;
        RECT 119.580 266.950 123.530 267.100 ;
        RECT 123.130 266.500 123.530 266.950 ;
        RECT 119.580 266.350 123.530 266.500 ;
        RECT 123.130 265.900 123.530 266.350 ;
        RECT 119.580 265.750 123.530 265.900 ;
        RECT 123.130 265.300 123.530 265.750 ;
        RECT 119.580 265.150 123.530 265.300 ;
        RECT 123.130 264.700 123.530 265.150 ;
        RECT 119.580 264.550 123.530 264.700 ;
        RECT 123.130 264.400 123.530 264.550 ;
        RECT 123.130 264.100 124.730 264.400 ;
        RECT 119.580 263.950 124.730 264.100 ;
        RECT 123.130 263.500 124.730 263.950 ;
        RECT 119.580 263.350 124.730 263.500 ;
        RECT 123.130 262.900 124.730 263.350 ;
        RECT 119.580 262.750 124.730 262.900 ;
        RECT 123.130 262.300 124.730 262.750 ;
        RECT 119.580 262.150 124.730 262.300 ;
        RECT 123.530 261.200 124.730 262.150 ;
        RECT 125.140 262.000 127.140 263.275 ;
        RECT 4.730 258.800 9.130 261.200 ;
        RECT 20.330 258.800 29.130 261.200 ;
        RECT 40.330 258.800 49.130 261.200 ;
        RECT 60.330 258.800 69.130 261.200 ;
        RECT 80.330 258.800 89.130 261.200 ;
        RECT 100.330 258.800 109.130 261.200 ;
        RECT 120.330 258.800 124.730 261.200 ;
        RECT 4.730 257.850 5.940 258.800 ;
        RECT 4.730 257.700 9.880 257.850 ;
        RECT 2.315 256.335 4.330 257.610 ;
        RECT 4.730 257.250 6.330 257.700 ;
        RECT 4.730 257.100 9.880 257.250 ;
        RECT 4.730 256.650 6.330 257.100 ;
        RECT 4.730 256.500 9.880 256.650 ;
        RECT 4.730 256.050 6.330 256.500 ;
        RECT 4.730 255.900 9.880 256.050 ;
        RECT 4.730 255.600 6.330 255.900 ;
        RECT 2.315 253.250 4.315 255.545 ;
        RECT 5.930 255.450 6.330 255.600 ;
        RECT 5.930 255.300 9.880 255.450 ;
        RECT 5.930 254.850 6.330 255.300 ;
        RECT 5.930 254.700 9.880 254.850 ;
        RECT 5.930 254.250 6.330 254.700 ;
        RECT 5.930 254.100 9.880 254.250 ;
        RECT 5.930 253.650 6.330 254.100 ;
        RECT 5.930 253.500 9.880 253.650 ;
        RECT 5.930 253.050 6.330 253.500 ;
        RECT 5.930 252.900 9.880 253.050 ;
        RECT 5.930 252.450 6.330 252.900 ;
        RECT 5.930 252.300 9.880 252.450 ;
        RECT 5.930 251.850 6.330 252.300 ;
        RECT 5.930 251.700 9.880 251.850 ;
        RECT 5.930 251.250 6.330 251.700 ;
        RECT 5.930 251.100 9.880 251.250 ;
        RECT 5.930 250.650 6.330 251.100 ;
        RECT 5.930 250.500 9.880 250.650 ;
        RECT 5.930 250.200 6.330 250.500 ;
        RECT 10.480 250.200 10.630 258.400 ;
        RECT 11.080 250.200 11.230 258.400 ;
        RECT 11.680 250.200 11.830 258.400 ;
        RECT 12.280 250.200 12.430 258.400 ;
        RECT 12.880 250.200 13.030 258.400 ;
        RECT 13.480 250.200 13.630 258.400 ;
        RECT 14.080 250.200 14.230 258.400 ;
        RECT 5.930 249.800 14.230 250.200 ;
        RECT 5.930 249.500 6.330 249.800 ;
        RECT 5.930 249.350 9.880 249.500 ;
        RECT 5.930 248.900 6.330 249.350 ;
        RECT 5.930 248.750 9.880 248.900 ;
        RECT 5.930 248.300 6.330 248.750 ;
        RECT 5.930 248.150 9.880 248.300 ;
        RECT 5.930 247.700 6.330 248.150 ;
        RECT 5.930 247.550 9.880 247.700 ;
        RECT 5.930 247.100 6.330 247.550 ;
        RECT 5.930 246.950 9.880 247.100 ;
        RECT 2.315 244.455 4.315 246.750 ;
        RECT 5.930 246.500 6.330 246.950 ;
        RECT 5.930 246.350 9.880 246.500 ;
        RECT 5.930 245.900 6.330 246.350 ;
        RECT 5.930 245.750 9.880 245.900 ;
        RECT 5.930 245.300 6.330 245.750 ;
        RECT 5.930 245.150 9.880 245.300 ;
        RECT 5.930 244.700 6.330 245.150 ;
        RECT 5.930 244.550 9.880 244.700 ;
        RECT 5.930 244.400 6.330 244.550 ;
        RECT 4.730 244.100 6.330 244.400 ;
        RECT 4.730 243.950 9.880 244.100 ;
        RECT 2.315 242.505 4.320 243.780 ;
        RECT 4.730 243.500 6.330 243.950 ;
        RECT 4.730 243.350 9.880 243.500 ;
        RECT 4.730 242.900 6.330 243.350 ;
        RECT 4.730 242.750 9.880 242.900 ;
        RECT 4.730 242.300 6.330 242.750 ;
        RECT 4.730 242.150 9.880 242.300 ;
        RECT 4.730 241.200 5.930 242.150 ;
        RECT 10.480 241.600 10.630 249.800 ;
        RECT 11.080 241.600 11.230 249.800 ;
        RECT 11.680 241.600 11.830 249.800 ;
        RECT 12.280 241.600 12.430 249.800 ;
        RECT 12.880 241.600 13.030 249.800 ;
        RECT 13.480 241.600 13.630 249.800 ;
        RECT 14.080 241.600 14.230 249.800 ;
        RECT 15.230 250.200 15.380 258.400 ;
        RECT 15.830 250.200 15.980 258.400 ;
        RECT 16.430 250.200 16.580 258.400 ;
        RECT 17.030 250.200 17.180 258.400 ;
        RECT 17.630 250.200 17.780 258.400 ;
        RECT 18.230 250.200 18.380 258.400 ;
        RECT 18.830 250.200 18.980 258.400 ;
        RECT 23.530 257.850 25.940 258.800 ;
        RECT 19.580 257.700 29.880 257.850 ;
        RECT 23.130 257.250 26.330 257.700 ;
        RECT 19.580 257.100 29.880 257.250 ;
        RECT 23.130 256.650 26.330 257.100 ;
        RECT 19.580 256.500 29.880 256.650 ;
        RECT 23.130 256.050 26.330 256.500 ;
        RECT 19.580 255.900 29.880 256.050 ;
        RECT 23.130 255.600 26.330 255.900 ;
        RECT 23.130 255.450 23.530 255.600 ;
        RECT 19.580 255.300 23.530 255.450 ;
        RECT 23.130 254.850 23.530 255.300 ;
        RECT 19.580 254.700 23.530 254.850 ;
        RECT 23.130 254.250 23.530 254.700 ;
        RECT 19.580 254.100 23.530 254.250 ;
        RECT 23.130 253.650 23.530 254.100 ;
        RECT 19.580 253.500 23.530 253.650 ;
        RECT 23.130 253.050 23.530 253.500 ;
        RECT 19.580 252.900 23.530 253.050 ;
        RECT 23.130 252.450 23.530 252.900 ;
        RECT 19.580 252.300 23.530 252.450 ;
        RECT 23.130 251.850 23.530 252.300 ;
        RECT 19.580 251.700 23.530 251.850 ;
        RECT 23.130 251.250 23.530 251.700 ;
        RECT 19.580 251.100 23.530 251.250 ;
        RECT 23.130 250.650 23.530 251.100 ;
        RECT 19.580 250.500 23.530 250.650 ;
        RECT 23.130 250.200 23.530 250.500 ;
        RECT 15.230 249.800 23.530 250.200 ;
        RECT 15.230 241.600 15.380 249.800 ;
        RECT 15.830 241.600 15.980 249.800 ;
        RECT 16.430 241.600 16.580 249.800 ;
        RECT 17.030 241.600 17.180 249.800 ;
        RECT 17.630 241.600 17.780 249.800 ;
        RECT 18.230 241.600 18.380 249.800 ;
        RECT 18.830 241.600 18.980 249.800 ;
        RECT 23.130 249.500 23.530 249.800 ;
        RECT 19.580 249.350 23.530 249.500 ;
        RECT 23.130 248.900 23.530 249.350 ;
        RECT 19.580 248.750 23.530 248.900 ;
        RECT 23.130 248.300 23.530 248.750 ;
        RECT 19.580 248.150 23.530 248.300 ;
        RECT 23.130 247.700 23.530 248.150 ;
        RECT 19.580 247.550 23.530 247.700 ;
        RECT 23.130 247.100 23.530 247.550 ;
        RECT 19.580 246.950 23.530 247.100 ;
        RECT 23.130 246.500 23.530 246.950 ;
        RECT 19.580 246.350 23.530 246.500 ;
        RECT 23.130 245.900 23.530 246.350 ;
        RECT 19.580 245.750 23.530 245.900 ;
        RECT 23.130 245.300 23.530 245.750 ;
        RECT 19.580 245.150 23.530 245.300 ;
        RECT 23.130 244.700 23.530 245.150 ;
        RECT 19.580 244.550 23.530 244.700 ;
        RECT 23.130 244.400 23.530 244.550 ;
        RECT 25.930 255.450 26.330 255.600 ;
        RECT 25.930 255.300 29.880 255.450 ;
        RECT 25.930 254.850 26.330 255.300 ;
        RECT 25.930 254.700 29.880 254.850 ;
        RECT 25.930 254.250 26.330 254.700 ;
        RECT 25.930 254.100 29.880 254.250 ;
        RECT 25.930 253.650 26.330 254.100 ;
        RECT 25.930 253.500 29.880 253.650 ;
        RECT 25.930 253.050 26.330 253.500 ;
        RECT 25.930 252.900 29.880 253.050 ;
        RECT 25.930 252.450 26.330 252.900 ;
        RECT 25.930 252.300 29.880 252.450 ;
        RECT 25.930 251.850 26.330 252.300 ;
        RECT 25.930 251.700 29.880 251.850 ;
        RECT 25.930 251.250 26.330 251.700 ;
        RECT 25.930 251.100 29.880 251.250 ;
        RECT 25.930 250.650 26.330 251.100 ;
        RECT 25.930 250.500 29.880 250.650 ;
        RECT 25.930 250.200 26.330 250.500 ;
        RECT 30.480 250.200 30.630 258.400 ;
        RECT 31.080 250.200 31.230 258.400 ;
        RECT 31.680 250.200 31.830 258.400 ;
        RECT 32.280 250.200 32.430 258.400 ;
        RECT 32.880 250.200 33.030 258.400 ;
        RECT 33.480 250.200 33.630 258.400 ;
        RECT 34.080 250.200 34.230 258.400 ;
        RECT 25.930 249.800 34.230 250.200 ;
        RECT 25.930 249.500 26.330 249.800 ;
        RECT 25.930 249.350 29.880 249.500 ;
        RECT 25.930 248.900 26.330 249.350 ;
        RECT 25.930 248.750 29.880 248.900 ;
        RECT 25.930 248.300 26.330 248.750 ;
        RECT 25.930 248.150 29.880 248.300 ;
        RECT 25.930 247.700 26.330 248.150 ;
        RECT 25.930 247.550 29.880 247.700 ;
        RECT 25.930 247.100 26.330 247.550 ;
        RECT 25.930 246.950 29.880 247.100 ;
        RECT 25.930 246.500 26.330 246.950 ;
        RECT 25.930 246.350 29.880 246.500 ;
        RECT 25.930 245.900 26.330 246.350 ;
        RECT 25.930 245.750 29.880 245.900 ;
        RECT 25.930 245.300 26.330 245.750 ;
        RECT 25.930 245.150 29.880 245.300 ;
        RECT 25.930 244.700 26.330 245.150 ;
        RECT 25.930 244.550 29.880 244.700 ;
        RECT 25.930 244.400 26.330 244.550 ;
        RECT 23.130 244.100 26.330 244.400 ;
        RECT 19.580 243.950 29.880 244.100 ;
        RECT 23.130 243.500 26.330 243.950 ;
        RECT 19.580 243.350 29.880 243.500 ;
        RECT 23.130 242.900 26.330 243.350 ;
        RECT 19.580 242.750 29.880 242.900 ;
        RECT 23.130 242.300 26.330 242.750 ;
        RECT 19.580 242.150 29.880 242.300 ;
        RECT 23.530 241.200 25.930 242.150 ;
        RECT 30.480 241.600 30.630 249.800 ;
        RECT 31.080 241.600 31.230 249.800 ;
        RECT 31.680 241.600 31.830 249.800 ;
        RECT 32.280 241.600 32.430 249.800 ;
        RECT 32.880 241.600 33.030 249.800 ;
        RECT 33.480 241.600 33.630 249.800 ;
        RECT 34.080 241.600 34.230 249.800 ;
        RECT 35.230 250.200 35.380 258.400 ;
        RECT 35.830 250.200 35.980 258.400 ;
        RECT 36.430 250.200 36.580 258.400 ;
        RECT 37.030 250.200 37.180 258.400 ;
        RECT 37.630 250.200 37.780 258.400 ;
        RECT 38.230 250.200 38.380 258.400 ;
        RECT 38.830 250.200 38.980 258.400 ;
        RECT 43.530 257.850 45.940 258.800 ;
        RECT 39.580 257.700 49.880 257.850 ;
        RECT 43.130 257.250 46.330 257.700 ;
        RECT 39.580 257.100 49.880 257.250 ;
        RECT 43.130 256.650 46.330 257.100 ;
        RECT 39.580 256.500 49.880 256.650 ;
        RECT 43.130 256.050 46.330 256.500 ;
        RECT 39.580 255.900 49.880 256.050 ;
        RECT 43.130 255.600 46.330 255.900 ;
        RECT 43.130 255.450 43.530 255.600 ;
        RECT 39.580 255.300 43.530 255.450 ;
        RECT 43.130 254.850 43.530 255.300 ;
        RECT 39.580 254.700 43.530 254.850 ;
        RECT 43.130 254.250 43.530 254.700 ;
        RECT 39.580 254.100 43.530 254.250 ;
        RECT 43.130 253.650 43.530 254.100 ;
        RECT 39.580 253.500 43.530 253.650 ;
        RECT 43.130 253.050 43.530 253.500 ;
        RECT 39.580 252.900 43.530 253.050 ;
        RECT 43.130 252.450 43.530 252.900 ;
        RECT 39.580 252.300 43.530 252.450 ;
        RECT 43.130 251.850 43.530 252.300 ;
        RECT 39.580 251.700 43.530 251.850 ;
        RECT 43.130 251.250 43.530 251.700 ;
        RECT 39.580 251.100 43.530 251.250 ;
        RECT 43.130 250.650 43.530 251.100 ;
        RECT 39.580 250.500 43.530 250.650 ;
        RECT 43.130 250.200 43.530 250.500 ;
        RECT 35.230 249.800 43.530 250.200 ;
        RECT 35.230 241.600 35.380 249.800 ;
        RECT 35.830 241.600 35.980 249.800 ;
        RECT 36.430 241.600 36.580 249.800 ;
        RECT 37.030 241.600 37.180 249.800 ;
        RECT 37.630 241.600 37.780 249.800 ;
        RECT 38.230 241.600 38.380 249.800 ;
        RECT 38.830 241.600 38.980 249.800 ;
        RECT 43.130 249.500 43.530 249.800 ;
        RECT 39.580 249.350 43.530 249.500 ;
        RECT 43.130 248.900 43.530 249.350 ;
        RECT 39.580 248.750 43.530 248.900 ;
        RECT 43.130 248.300 43.530 248.750 ;
        RECT 39.580 248.150 43.530 248.300 ;
        RECT 43.130 247.700 43.530 248.150 ;
        RECT 39.580 247.550 43.530 247.700 ;
        RECT 43.130 247.100 43.530 247.550 ;
        RECT 39.580 246.950 43.530 247.100 ;
        RECT 43.130 246.500 43.530 246.950 ;
        RECT 39.580 246.350 43.530 246.500 ;
        RECT 43.130 245.900 43.530 246.350 ;
        RECT 39.580 245.750 43.530 245.900 ;
        RECT 43.130 245.300 43.530 245.750 ;
        RECT 39.580 245.150 43.530 245.300 ;
        RECT 43.130 244.700 43.530 245.150 ;
        RECT 39.580 244.550 43.530 244.700 ;
        RECT 43.130 244.400 43.530 244.550 ;
        RECT 45.930 255.450 46.330 255.600 ;
        RECT 45.930 255.300 49.880 255.450 ;
        RECT 45.930 254.850 46.330 255.300 ;
        RECT 45.930 254.700 49.880 254.850 ;
        RECT 45.930 254.250 46.330 254.700 ;
        RECT 45.930 254.100 49.880 254.250 ;
        RECT 45.930 253.650 46.330 254.100 ;
        RECT 45.930 253.500 49.880 253.650 ;
        RECT 45.930 253.050 46.330 253.500 ;
        RECT 45.930 252.900 49.880 253.050 ;
        RECT 45.930 252.450 46.330 252.900 ;
        RECT 45.930 252.300 49.880 252.450 ;
        RECT 45.930 251.850 46.330 252.300 ;
        RECT 45.930 251.700 49.880 251.850 ;
        RECT 45.930 251.250 46.330 251.700 ;
        RECT 45.930 251.100 49.880 251.250 ;
        RECT 45.930 250.650 46.330 251.100 ;
        RECT 45.930 250.500 49.880 250.650 ;
        RECT 45.930 250.200 46.330 250.500 ;
        RECT 50.480 250.200 50.630 258.400 ;
        RECT 51.080 250.200 51.230 258.400 ;
        RECT 51.680 250.200 51.830 258.400 ;
        RECT 52.280 250.200 52.430 258.400 ;
        RECT 52.880 250.200 53.030 258.400 ;
        RECT 53.480 250.200 53.630 258.400 ;
        RECT 54.080 250.200 54.230 258.400 ;
        RECT 45.930 249.800 54.230 250.200 ;
        RECT 45.930 249.500 46.330 249.800 ;
        RECT 45.930 249.350 49.880 249.500 ;
        RECT 45.930 248.900 46.330 249.350 ;
        RECT 45.930 248.750 49.880 248.900 ;
        RECT 45.930 248.300 46.330 248.750 ;
        RECT 45.930 248.150 49.880 248.300 ;
        RECT 45.930 247.700 46.330 248.150 ;
        RECT 45.930 247.550 49.880 247.700 ;
        RECT 45.930 247.100 46.330 247.550 ;
        RECT 45.930 246.950 49.880 247.100 ;
        RECT 45.930 246.500 46.330 246.950 ;
        RECT 45.930 246.350 49.880 246.500 ;
        RECT 45.930 245.900 46.330 246.350 ;
        RECT 45.930 245.750 49.880 245.900 ;
        RECT 45.930 245.300 46.330 245.750 ;
        RECT 45.930 245.150 49.880 245.300 ;
        RECT 45.930 244.700 46.330 245.150 ;
        RECT 45.930 244.550 49.880 244.700 ;
        RECT 45.930 244.400 46.330 244.550 ;
        RECT 43.130 244.100 46.330 244.400 ;
        RECT 39.580 243.950 49.880 244.100 ;
        RECT 43.130 243.500 46.330 243.950 ;
        RECT 39.580 243.350 49.880 243.500 ;
        RECT 43.130 242.900 46.330 243.350 ;
        RECT 39.580 242.750 49.880 242.900 ;
        RECT 43.130 242.300 46.330 242.750 ;
        RECT 39.580 242.150 49.880 242.300 ;
        RECT 43.530 241.200 45.930 242.150 ;
        RECT 50.480 241.600 50.630 249.800 ;
        RECT 51.080 241.600 51.230 249.800 ;
        RECT 51.680 241.600 51.830 249.800 ;
        RECT 52.280 241.600 52.430 249.800 ;
        RECT 52.880 241.600 53.030 249.800 ;
        RECT 53.480 241.600 53.630 249.800 ;
        RECT 54.080 241.600 54.230 249.800 ;
        RECT 55.230 250.200 55.380 258.400 ;
        RECT 55.830 250.200 55.980 258.400 ;
        RECT 56.430 250.200 56.580 258.400 ;
        RECT 57.030 250.200 57.180 258.400 ;
        RECT 57.630 250.200 57.780 258.400 ;
        RECT 58.230 250.200 58.380 258.400 ;
        RECT 58.830 250.200 58.980 258.400 ;
        RECT 63.530 257.850 65.940 258.800 ;
        RECT 59.580 257.700 69.880 257.850 ;
        RECT 63.130 257.250 66.330 257.700 ;
        RECT 59.580 257.100 69.880 257.250 ;
        RECT 63.130 256.650 66.330 257.100 ;
        RECT 59.580 256.500 69.880 256.650 ;
        RECT 63.130 256.050 66.330 256.500 ;
        RECT 59.580 255.900 69.880 256.050 ;
        RECT 63.130 255.600 66.330 255.900 ;
        RECT 63.130 255.450 63.530 255.600 ;
        RECT 59.580 255.300 63.530 255.450 ;
        RECT 63.130 254.850 63.530 255.300 ;
        RECT 59.580 254.700 63.530 254.850 ;
        RECT 63.130 254.250 63.530 254.700 ;
        RECT 59.580 254.100 63.530 254.250 ;
        RECT 63.130 253.650 63.530 254.100 ;
        RECT 59.580 253.500 63.530 253.650 ;
        RECT 63.130 253.050 63.530 253.500 ;
        RECT 59.580 252.900 63.530 253.050 ;
        RECT 63.130 252.450 63.530 252.900 ;
        RECT 59.580 252.300 63.530 252.450 ;
        RECT 63.130 251.850 63.530 252.300 ;
        RECT 59.580 251.700 63.530 251.850 ;
        RECT 63.130 251.250 63.530 251.700 ;
        RECT 59.580 251.100 63.530 251.250 ;
        RECT 63.130 250.650 63.530 251.100 ;
        RECT 59.580 250.500 63.530 250.650 ;
        RECT 63.130 250.200 63.530 250.500 ;
        RECT 55.230 249.800 63.530 250.200 ;
        RECT 55.230 241.600 55.380 249.800 ;
        RECT 55.830 241.600 55.980 249.800 ;
        RECT 56.430 241.600 56.580 249.800 ;
        RECT 57.030 241.600 57.180 249.800 ;
        RECT 57.630 241.600 57.780 249.800 ;
        RECT 58.230 241.600 58.380 249.800 ;
        RECT 58.830 241.600 58.980 249.800 ;
        RECT 63.130 249.500 63.530 249.800 ;
        RECT 59.580 249.350 63.530 249.500 ;
        RECT 63.130 248.900 63.530 249.350 ;
        RECT 59.580 248.750 63.530 248.900 ;
        RECT 63.130 248.300 63.530 248.750 ;
        RECT 59.580 248.150 63.530 248.300 ;
        RECT 63.130 247.700 63.530 248.150 ;
        RECT 59.580 247.550 63.530 247.700 ;
        RECT 63.130 247.100 63.530 247.550 ;
        RECT 59.580 246.950 63.530 247.100 ;
        RECT 63.130 246.500 63.530 246.950 ;
        RECT 59.580 246.350 63.530 246.500 ;
        RECT 63.130 245.900 63.530 246.350 ;
        RECT 59.580 245.750 63.530 245.900 ;
        RECT 63.130 245.300 63.530 245.750 ;
        RECT 59.580 245.150 63.530 245.300 ;
        RECT 63.130 244.700 63.530 245.150 ;
        RECT 59.580 244.550 63.530 244.700 ;
        RECT 63.130 244.400 63.530 244.550 ;
        RECT 65.930 255.450 66.330 255.600 ;
        RECT 65.930 255.300 69.880 255.450 ;
        RECT 65.930 254.850 66.330 255.300 ;
        RECT 65.930 254.700 69.880 254.850 ;
        RECT 65.930 254.250 66.330 254.700 ;
        RECT 65.930 254.100 69.880 254.250 ;
        RECT 65.930 253.650 66.330 254.100 ;
        RECT 65.930 253.500 69.880 253.650 ;
        RECT 65.930 253.050 66.330 253.500 ;
        RECT 65.930 252.900 69.880 253.050 ;
        RECT 65.930 252.450 66.330 252.900 ;
        RECT 65.930 252.300 69.880 252.450 ;
        RECT 65.930 251.850 66.330 252.300 ;
        RECT 65.930 251.700 69.880 251.850 ;
        RECT 65.930 251.250 66.330 251.700 ;
        RECT 65.930 251.100 69.880 251.250 ;
        RECT 65.930 250.650 66.330 251.100 ;
        RECT 65.930 250.500 69.880 250.650 ;
        RECT 65.930 250.200 66.330 250.500 ;
        RECT 70.480 250.200 70.630 258.400 ;
        RECT 71.080 250.200 71.230 258.400 ;
        RECT 71.680 250.200 71.830 258.400 ;
        RECT 72.280 250.200 72.430 258.400 ;
        RECT 72.880 250.200 73.030 258.400 ;
        RECT 73.480 250.200 73.630 258.400 ;
        RECT 74.080 250.200 74.230 258.400 ;
        RECT 65.930 249.800 74.230 250.200 ;
        RECT 65.930 249.500 66.330 249.800 ;
        RECT 65.930 249.350 69.880 249.500 ;
        RECT 65.930 248.900 66.330 249.350 ;
        RECT 65.930 248.750 69.880 248.900 ;
        RECT 65.930 248.300 66.330 248.750 ;
        RECT 65.930 248.150 69.880 248.300 ;
        RECT 65.930 247.700 66.330 248.150 ;
        RECT 65.930 247.550 69.880 247.700 ;
        RECT 65.930 247.100 66.330 247.550 ;
        RECT 65.930 246.950 69.880 247.100 ;
        RECT 65.930 246.500 66.330 246.950 ;
        RECT 65.930 246.350 69.880 246.500 ;
        RECT 65.930 245.900 66.330 246.350 ;
        RECT 65.930 245.750 69.880 245.900 ;
        RECT 65.930 245.300 66.330 245.750 ;
        RECT 65.930 245.150 69.880 245.300 ;
        RECT 65.930 244.700 66.330 245.150 ;
        RECT 65.930 244.550 69.880 244.700 ;
        RECT 65.930 244.400 66.330 244.550 ;
        RECT 63.130 244.100 66.330 244.400 ;
        RECT 59.580 243.950 69.880 244.100 ;
        RECT 63.130 243.500 66.330 243.950 ;
        RECT 59.580 243.350 69.880 243.500 ;
        RECT 63.130 242.900 66.330 243.350 ;
        RECT 59.580 242.750 69.880 242.900 ;
        RECT 63.130 242.300 66.330 242.750 ;
        RECT 59.580 242.150 69.880 242.300 ;
        RECT 63.530 241.200 65.930 242.150 ;
        RECT 70.480 241.600 70.630 249.800 ;
        RECT 71.080 241.600 71.230 249.800 ;
        RECT 71.680 241.600 71.830 249.800 ;
        RECT 72.280 241.600 72.430 249.800 ;
        RECT 72.880 241.600 73.030 249.800 ;
        RECT 73.480 241.600 73.630 249.800 ;
        RECT 74.080 241.600 74.230 249.800 ;
        RECT 75.230 250.200 75.380 258.400 ;
        RECT 75.830 250.200 75.980 258.400 ;
        RECT 76.430 250.200 76.580 258.400 ;
        RECT 77.030 250.200 77.180 258.400 ;
        RECT 77.630 250.200 77.780 258.400 ;
        RECT 78.230 250.200 78.380 258.400 ;
        RECT 78.830 250.200 78.980 258.400 ;
        RECT 83.530 257.850 85.940 258.800 ;
        RECT 79.580 257.700 89.880 257.850 ;
        RECT 83.130 257.250 86.330 257.700 ;
        RECT 79.580 257.100 89.880 257.250 ;
        RECT 83.130 256.650 86.330 257.100 ;
        RECT 79.580 256.500 89.880 256.650 ;
        RECT 83.130 256.050 86.330 256.500 ;
        RECT 79.580 255.900 89.880 256.050 ;
        RECT 83.130 255.600 86.330 255.900 ;
        RECT 83.130 255.450 83.530 255.600 ;
        RECT 79.580 255.300 83.530 255.450 ;
        RECT 83.130 254.850 83.530 255.300 ;
        RECT 79.580 254.700 83.530 254.850 ;
        RECT 83.130 254.250 83.530 254.700 ;
        RECT 79.580 254.100 83.530 254.250 ;
        RECT 83.130 253.650 83.530 254.100 ;
        RECT 79.580 253.500 83.530 253.650 ;
        RECT 83.130 253.050 83.530 253.500 ;
        RECT 79.580 252.900 83.530 253.050 ;
        RECT 83.130 252.450 83.530 252.900 ;
        RECT 79.580 252.300 83.530 252.450 ;
        RECT 83.130 251.850 83.530 252.300 ;
        RECT 79.580 251.700 83.530 251.850 ;
        RECT 83.130 251.250 83.530 251.700 ;
        RECT 79.580 251.100 83.530 251.250 ;
        RECT 83.130 250.650 83.530 251.100 ;
        RECT 79.580 250.500 83.530 250.650 ;
        RECT 83.130 250.200 83.530 250.500 ;
        RECT 75.230 249.800 83.530 250.200 ;
        RECT 75.230 241.600 75.380 249.800 ;
        RECT 75.830 241.600 75.980 249.800 ;
        RECT 76.430 241.600 76.580 249.800 ;
        RECT 77.030 241.600 77.180 249.800 ;
        RECT 77.630 241.600 77.780 249.800 ;
        RECT 78.230 241.600 78.380 249.800 ;
        RECT 78.830 241.600 78.980 249.800 ;
        RECT 83.130 249.500 83.530 249.800 ;
        RECT 79.580 249.350 83.530 249.500 ;
        RECT 83.130 248.900 83.530 249.350 ;
        RECT 79.580 248.750 83.530 248.900 ;
        RECT 83.130 248.300 83.530 248.750 ;
        RECT 79.580 248.150 83.530 248.300 ;
        RECT 83.130 247.700 83.530 248.150 ;
        RECT 79.580 247.550 83.530 247.700 ;
        RECT 83.130 247.100 83.530 247.550 ;
        RECT 79.580 246.950 83.530 247.100 ;
        RECT 83.130 246.500 83.530 246.950 ;
        RECT 79.580 246.350 83.530 246.500 ;
        RECT 83.130 245.900 83.530 246.350 ;
        RECT 79.580 245.750 83.530 245.900 ;
        RECT 83.130 245.300 83.530 245.750 ;
        RECT 79.580 245.150 83.530 245.300 ;
        RECT 83.130 244.700 83.530 245.150 ;
        RECT 79.580 244.550 83.530 244.700 ;
        RECT 83.130 244.400 83.530 244.550 ;
        RECT 85.930 255.450 86.330 255.600 ;
        RECT 85.930 255.300 89.880 255.450 ;
        RECT 85.930 254.850 86.330 255.300 ;
        RECT 85.930 254.700 89.880 254.850 ;
        RECT 85.930 254.250 86.330 254.700 ;
        RECT 85.930 254.100 89.880 254.250 ;
        RECT 85.930 253.650 86.330 254.100 ;
        RECT 85.930 253.500 89.880 253.650 ;
        RECT 85.930 253.050 86.330 253.500 ;
        RECT 85.930 252.900 89.880 253.050 ;
        RECT 85.930 252.450 86.330 252.900 ;
        RECT 85.930 252.300 89.880 252.450 ;
        RECT 85.930 251.850 86.330 252.300 ;
        RECT 85.930 251.700 89.880 251.850 ;
        RECT 85.930 251.250 86.330 251.700 ;
        RECT 85.930 251.100 89.880 251.250 ;
        RECT 85.930 250.650 86.330 251.100 ;
        RECT 85.930 250.500 89.880 250.650 ;
        RECT 85.930 250.200 86.330 250.500 ;
        RECT 90.480 250.200 90.630 258.400 ;
        RECT 91.080 250.200 91.230 258.400 ;
        RECT 91.680 250.200 91.830 258.400 ;
        RECT 92.280 250.200 92.430 258.400 ;
        RECT 92.880 250.200 93.030 258.400 ;
        RECT 93.480 250.200 93.630 258.400 ;
        RECT 94.080 250.200 94.230 258.400 ;
        RECT 85.930 249.800 94.230 250.200 ;
        RECT 85.930 249.500 86.330 249.800 ;
        RECT 85.930 249.350 89.880 249.500 ;
        RECT 85.930 248.900 86.330 249.350 ;
        RECT 85.930 248.750 89.880 248.900 ;
        RECT 85.930 248.300 86.330 248.750 ;
        RECT 85.930 248.150 89.880 248.300 ;
        RECT 85.930 247.700 86.330 248.150 ;
        RECT 85.930 247.550 89.880 247.700 ;
        RECT 85.930 247.100 86.330 247.550 ;
        RECT 85.930 246.950 89.880 247.100 ;
        RECT 85.930 246.500 86.330 246.950 ;
        RECT 85.930 246.350 89.880 246.500 ;
        RECT 85.930 245.900 86.330 246.350 ;
        RECT 85.930 245.750 89.880 245.900 ;
        RECT 85.930 245.300 86.330 245.750 ;
        RECT 85.930 245.150 89.880 245.300 ;
        RECT 85.930 244.700 86.330 245.150 ;
        RECT 85.930 244.550 89.880 244.700 ;
        RECT 85.930 244.400 86.330 244.550 ;
        RECT 83.130 244.100 86.330 244.400 ;
        RECT 79.580 243.950 89.880 244.100 ;
        RECT 83.130 243.500 86.330 243.950 ;
        RECT 79.580 243.350 89.880 243.500 ;
        RECT 83.130 242.900 86.330 243.350 ;
        RECT 79.580 242.750 89.880 242.900 ;
        RECT 83.130 242.300 86.330 242.750 ;
        RECT 79.580 242.150 89.880 242.300 ;
        RECT 83.530 241.200 85.930 242.150 ;
        RECT 90.480 241.600 90.630 249.800 ;
        RECT 91.080 241.600 91.230 249.800 ;
        RECT 91.680 241.600 91.830 249.800 ;
        RECT 92.280 241.600 92.430 249.800 ;
        RECT 92.880 241.600 93.030 249.800 ;
        RECT 93.480 241.600 93.630 249.800 ;
        RECT 94.080 241.600 94.230 249.800 ;
        RECT 95.230 250.200 95.380 258.400 ;
        RECT 95.830 250.200 95.980 258.400 ;
        RECT 96.430 250.200 96.580 258.400 ;
        RECT 97.030 250.200 97.180 258.400 ;
        RECT 97.630 250.200 97.780 258.400 ;
        RECT 98.230 250.200 98.380 258.400 ;
        RECT 98.830 250.200 98.980 258.400 ;
        RECT 103.530 257.850 105.940 258.800 ;
        RECT 99.580 257.700 109.880 257.850 ;
        RECT 103.130 257.250 106.330 257.700 ;
        RECT 99.580 257.100 109.880 257.250 ;
        RECT 103.130 256.650 106.330 257.100 ;
        RECT 99.580 256.500 109.880 256.650 ;
        RECT 103.130 256.050 106.330 256.500 ;
        RECT 99.580 255.900 109.880 256.050 ;
        RECT 103.130 255.600 106.330 255.900 ;
        RECT 103.130 255.450 103.530 255.600 ;
        RECT 99.580 255.300 103.530 255.450 ;
        RECT 103.130 254.850 103.530 255.300 ;
        RECT 99.580 254.700 103.530 254.850 ;
        RECT 103.130 254.250 103.530 254.700 ;
        RECT 99.580 254.100 103.530 254.250 ;
        RECT 103.130 253.650 103.530 254.100 ;
        RECT 99.580 253.500 103.530 253.650 ;
        RECT 103.130 253.050 103.530 253.500 ;
        RECT 99.580 252.900 103.530 253.050 ;
        RECT 103.130 252.450 103.530 252.900 ;
        RECT 99.580 252.300 103.530 252.450 ;
        RECT 103.130 251.850 103.530 252.300 ;
        RECT 99.580 251.700 103.530 251.850 ;
        RECT 103.130 251.250 103.530 251.700 ;
        RECT 99.580 251.100 103.530 251.250 ;
        RECT 103.130 250.650 103.530 251.100 ;
        RECT 99.580 250.500 103.530 250.650 ;
        RECT 103.130 250.200 103.530 250.500 ;
        RECT 95.230 249.800 103.530 250.200 ;
        RECT 95.230 241.600 95.380 249.800 ;
        RECT 95.830 241.600 95.980 249.800 ;
        RECT 96.430 241.600 96.580 249.800 ;
        RECT 97.030 241.600 97.180 249.800 ;
        RECT 97.630 241.600 97.780 249.800 ;
        RECT 98.230 241.600 98.380 249.800 ;
        RECT 98.830 241.600 98.980 249.800 ;
        RECT 103.130 249.500 103.530 249.800 ;
        RECT 99.580 249.350 103.530 249.500 ;
        RECT 103.130 248.900 103.530 249.350 ;
        RECT 99.580 248.750 103.530 248.900 ;
        RECT 103.130 248.300 103.530 248.750 ;
        RECT 99.580 248.150 103.530 248.300 ;
        RECT 103.130 247.700 103.530 248.150 ;
        RECT 99.580 247.550 103.530 247.700 ;
        RECT 103.130 247.100 103.530 247.550 ;
        RECT 99.580 246.950 103.530 247.100 ;
        RECT 103.130 246.500 103.530 246.950 ;
        RECT 99.580 246.350 103.530 246.500 ;
        RECT 103.130 245.900 103.530 246.350 ;
        RECT 99.580 245.750 103.530 245.900 ;
        RECT 103.130 245.300 103.530 245.750 ;
        RECT 99.580 245.150 103.530 245.300 ;
        RECT 103.130 244.700 103.530 245.150 ;
        RECT 99.580 244.550 103.530 244.700 ;
        RECT 103.130 244.400 103.530 244.550 ;
        RECT 105.930 255.450 106.330 255.600 ;
        RECT 105.930 255.300 109.880 255.450 ;
        RECT 105.930 254.850 106.330 255.300 ;
        RECT 105.930 254.700 109.880 254.850 ;
        RECT 105.930 254.250 106.330 254.700 ;
        RECT 105.930 254.100 109.880 254.250 ;
        RECT 105.930 253.650 106.330 254.100 ;
        RECT 105.930 253.500 109.880 253.650 ;
        RECT 105.930 253.050 106.330 253.500 ;
        RECT 105.930 252.900 109.880 253.050 ;
        RECT 105.930 252.450 106.330 252.900 ;
        RECT 105.930 252.300 109.880 252.450 ;
        RECT 105.930 251.850 106.330 252.300 ;
        RECT 105.930 251.700 109.880 251.850 ;
        RECT 105.930 251.250 106.330 251.700 ;
        RECT 105.930 251.100 109.880 251.250 ;
        RECT 105.930 250.650 106.330 251.100 ;
        RECT 105.930 250.500 109.880 250.650 ;
        RECT 105.930 250.200 106.330 250.500 ;
        RECT 110.480 250.200 110.630 258.400 ;
        RECT 111.080 250.200 111.230 258.400 ;
        RECT 111.680 250.200 111.830 258.400 ;
        RECT 112.280 250.200 112.430 258.400 ;
        RECT 112.880 250.200 113.030 258.400 ;
        RECT 113.480 250.200 113.630 258.400 ;
        RECT 114.080 250.200 114.230 258.400 ;
        RECT 105.930 249.800 114.230 250.200 ;
        RECT 105.930 249.500 106.330 249.800 ;
        RECT 105.930 249.350 109.880 249.500 ;
        RECT 105.930 248.900 106.330 249.350 ;
        RECT 105.930 248.750 109.880 248.900 ;
        RECT 105.930 248.300 106.330 248.750 ;
        RECT 105.930 248.150 109.880 248.300 ;
        RECT 105.930 247.700 106.330 248.150 ;
        RECT 105.930 247.550 109.880 247.700 ;
        RECT 105.930 247.100 106.330 247.550 ;
        RECT 105.930 246.950 109.880 247.100 ;
        RECT 105.930 246.500 106.330 246.950 ;
        RECT 105.930 246.350 109.880 246.500 ;
        RECT 105.930 245.900 106.330 246.350 ;
        RECT 105.930 245.750 109.880 245.900 ;
        RECT 105.930 245.300 106.330 245.750 ;
        RECT 105.930 245.150 109.880 245.300 ;
        RECT 105.930 244.700 106.330 245.150 ;
        RECT 105.930 244.550 109.880 244.700 ;
        RECT 105.930 244.400 106.330 244.550 ;
        RECT 103.130 244.100 106.330 244.400 ;
        RECT 99.580 243.950 109.880 244.100 ;
        RECT 103.130 243.500 106.330 243.950 ;
        RECT 99.580 243.350 109.880 243.500 ;
        RECT 103.130 242.900 106.330 243.350 ;
        RECT 99.580 242.750 109.880 242.900 ;
        RECT 103.130 242.300 106.330 242.750 ;
        RECT 99.580 242.150 109.880 242.300 ;
        RECT 103.530 241.200 105.930 242.150 ;
        RECT 110.480 241.600 110.630 249.800 ;
        RECT 111.080 241.600 111.230 249.800 ;
        RECT 111.680 241.600 111.830 249.800 ;
        RECT 112.280 241.600 112.430 249.800 ;
        RECT 112.880 241.600 113.030 249.800 ;
        RECT 113.480 241.600 113.630 249.800 ;
        RECT 114.080 241.600 114.230 249.800 ;
        RECT 115.230 250.200 115.380 258.400 ;
        RECT 115.830 250.200 115.980 258.400 ;
        RECT 116.430 250.200 116.580 258.400 ;
        RECT 117.030 250.200 117.180 258.400 ;
        RECT 117.630 250.200 117.780 258.400 ;
        RECT 118.230 250.200 118.380 258.400 ;
        RECT 118.830 250.200 118.980 258.400 ;
        RECT 123.530 257.850 124.730 258.800 ;
        RECT 119.580 257.700 124.730 257.850 ;
        RECT 123.130 257.250 124.730 257.700 ;
        RECT 119.580 257.100 124.730 257.250 ;
        RECT 123.130 256.650 124.730 257.100 ;
        RECT 119.580 256.500 124.730 256.650 ;
        RECT 123.130 256.050 124.730 256.500 ;
        RECT 125.135 256.085 127.135 257.360 ;
        RECT 119.580 255.900 124.730 256.050 ;
        RECT 123.130 255.600 124.730 255.900 ;
        RECT 123.130 255.450 123.530 255.600 ;
        RECT 119.580 255.300 123.530 255.450 ;
        RECT 123.130 254.850 123.530 255.300 ;
        RECT 119.580 254.700 123.530 254.850 ;
        RECT 123.130 254.250 123.530 254.700 ;
        RECT 119.580 254.100 123.530 254.250 ;
        RECT 123.130 253.650 123.530 254.100 ;
        RECT 119.580 253.500 123.530 253.650 ;
        RECT 123.130 253.050 123.530 253.500 ;
        RECT 119.580 252.900 123.530 253.050 ;
        RECT 123.130 252.450 123.530 252.900 ;
        RECT 119.580 252.300 123.530 252.450 ;
        RECT 123.130 251.850 123.530 252.300 ;
        RECT 119.580 251.700 123.530 251.850 ;
        RECT 123.130 251.250 123.530 251.700 ;
        RECT 119.580 251.100 123.530 251.250 ;
        RECT 123.130 250.650 123.530 251.100 ;
        RECT 119.580 250.500 123.530 250.650 ;
        RECT 123.130 250.200 123.530 250.500 ;
        RECT 115.230 249.800 123.530 250.200 ;
        RECT 115.230 241.600 115.380 249.800 ;
        RECT 115.830 241.600 115.980 249.800 ;
        RECT 116.430 241.600 116.580 249.800 ;
        RECT 117.030 241.600 117.180 249.800 ;
        RECT 117.630 241.600 117.780 249.800 ;
        RECT 118.230 241.600 118.380 249.800 ;
        RECT 118.830 241.600 118.980 249.800 ;
        RECT 123.130 249.500 123.530 249.800 ;
        RECT 119.580 249.350 123.530 249.500 ;
        RECT 123.130 248.900 123.530 249.350 ;
        RECT 119.580 248.750 123.530 248.900 ;
        RECT 123.130 248.300 123.530 248.750 ;
        RECT 119.580 248.150 123.530 248.300 ;
        RECT 123.130 247.700 123.530 248.150 ;
        RECT 119.580 247.550 123.530 247.700 ;
        RECT 123.130 247.100 123.530 247.550 ;
        RECT 119.580 246.950 123.530 247.100 ;
        RECT 123.130 246.500 123.530 246.950 ;
        RECT 119.580 246.350 123.530 246.500 ;
        RECT 123.130 245.900 123.530 246.350 ;
        RECT 119.580 245.750 123.530 245.900 ;
        RECT 123.130 245.300 123.530 245.750 ;
        RECT 119.580 245.150 123.530 245.300 ;
        RECT 123.130 244.700 123.530 245.150 ;
        RECT 119.580 244.550 123.530 244.700 ;
        RECT 123.130 244.400 123.530 244.550 ;
        RECT 123.130 244.100 124.730 244.400 ;
        RECT 119.580 243.950 124.730 244.100 ;
        RECT 123.130 243.500 124.730 243.950 ;
        RECT 119.580 243.350 124.730 243.500 ;
        RECT 123.130 242.900 124.730 243.350 ;
        RECT 119.580 242.750 124.730 242.900 ;
        RECT 123.130 242.300 124.730 242.750 ;
        RECT 119.580 242.150 124.730 242.300 ;
        RECT 123.530 241.200 124.730 242.150 ;
        RECT 125.140 241.725 127.140 243.000 ;
        RECT 4.730 238.800 9.130 241.200 ;
        RECT 20.330 238.800 29.130 241.200 ;
        RECT 40.330 238.800 49.130 241.200 ;
        RECT 60.330 238.800 69.130 241.200 ;
        RECT 80.330 238.800 89.130 241.200 ;
        RECT 100.330 238.800 109.130 241.200 ;
        RECT 120.330 238.800 124.730 241.200 ;
        RECT 4.730 237.850 5.940 238.800 ;
        RECT 2.315 236.570 4.320 237.845 ;
        RECT 4.730 237.700 9.880 237.850 ;
        RECT 4.730 237.250 6.330 237.700 ;
        RECT 4.730 237.100 9.880 237.250 ;
        RECT 4.730 236.650 6.330 237.100 ;
        RECT 4.730 236.500 9.880 236.650 ;
        RECT 4.730 236.050 6.330 236.500 ;
        RECT 4.730 235.900 9.880 236.050 ;
        RECT 4.730 235.600 6.330 235.900 ;
        RECT 2.315 233.250 4.315 235.545 ;
        RECT 5.930 235.450 6.330 235.600 ;
        RECT 5.930 235.300 9.880 235.450 ;
        RECT 5.930 234.850 6.330 235.300 ;
        RECT 5.930 234.700 9.880 234.850 ;
        RECT 5.930 234.250 6.330 234.700 ;
        RECT 5.930 234.100 9.880 234.250 ;
        RECT 5.930 233.650 6.330 234.100 ;
        RECT 5.930 233.500 9.880 233.650 ;
        RECT 5.930 233.050 6.330 233.500 ;
        RECT 5.930 232.900 9.880 233.050 ;
        RECT 5.930 232.450 6.330 232.900 ;
        RECT 5.930 232.300 9.880 232.450 ;
        RECT 5.930 231.850 6.330 232.300 ;
        RECT 5.930 231.700 9.880 231.850 ;
        RECT 5.930 231.250 6.330 231.700 ;
        RECT 5.930 231.100 9.880 231.250 ;
        RECT 5.930 230.650 6.330 231.100 ;
        RECT 5.930 230.500 9.880 230.650 ;
        RECT 5.930 230.200 6.330 230.500 ;
        RECT 10.480 230.200 10.630 238.400 ;
        RECT 11.080 230.200 11.230 238.400 ;
        RECT 11.680 230.200 11.830 238.400 ;
        RECT 12.280 230.200 12.430 238.400 ;
        RECT 12.880 230.200 13.030 238.400 ;
        RECT 13.480 230.200 13.630 238.400 ;
        RECT 14.080 230.200 14.230 238.400 ;
        RECT 5.930 229.800 14.230 230.200 ;
        RECT 5.930 229.500 6.330 229.800 ;
        RECT 5.930 229.350 9.880 229.500 ;
        RECT 5.930 228.900 6.330 229.350 ;
        RECT 5.930 228.750 9.880 228.900 ;
        RECT 5.930 228.300 6.330 228.750 ;
        RECT 5.930 228.150 9.880 228.300 ;
        RECT 5.930 227.700 6.330 228.150 ;
        RECT 5.930 227.550 9.880 227.700 ;
        RECT 5.930 227.100 6.330 227.550 ;
        RECT 5.930 226.950 9.880 227.100 ;
        RECT 2.315 224.455 4.315 226.750 ;
        RECT 5.930 226.500 6.330 226.950 ;
        RECT 5.930 226.350 9.880 226.500 ;
        RECT 5.930 225.900 6.330 226.350 ;
        RECT 5.930 225.750 9.880 225.900 ;
        RECT 5.930 225.300 6.330 225.750 ;
        RECT 5.930 225.150 9.880 225.300 ;
        RECT 5.930 224.700 6.330 225.150 ;
        RECT 5.930 224.550 9.880 224.700 ;
        RECT 5.930 224.400 6.330 224.550 ;
        RECT 4.730 224.100 6.330 224.400 ;
        RECT 4.730 223.950 9.880 224.100 ;
        RECT 2.315 222.460 4.320 223.735 ;
        RECT 4.730 223.500 6.330 223.950 ;
        RECT 4.730 223.350 9.880 223.500 ;
        RECT 4.730 222.900 6.330 223.350 ;
        RECT 4.730 222.750 9.880 222.900 ;
        RECT 4.730 222.300 6.330 222.750 ;
        RECT 4.730 222.150 9.880 222.300 ;
        RECT 4.730 221.200 5.930 222.150 ;
        RECT 10.480 221.600 10.630 229.800 ;
        RECT 11.080 221.600 11.230 229.800 ;
        RECT 11.680 221.600 11.830 229.800 ;
        RECT 12.280 221.600 12.430 229.800 ;
        RECT 12.880 221.600 13.030 229.800 ;
        RECT 13.480 221.600 13.630 229.800 ;
        RECT 14.080 221.600 14.230 229.800 ;
        RECT 15.230 230.200 15.380 238.400 ;
        RECT 15.830 230.200 15.980 238.400 ;
        RECT 16.430 230.200 16.580 238.400 ;
        RECT 17.030 230.200 17.180 238.400 ;
        RECT 17.630 230.200 17.780 238.400 ;
        RECT 18.230 230.200 18.380 238.400 ;
        RECT 18.830 230.200 18.980 238.400 ;
        RECT 23.530 237.850 25.940 238.800 ;
        RECT 19.580 237.700 29.880 237.850 ;
        RECT 23.130 237.250 26.330 237.700 ;
        RECT 19.580 237.100 29.880 237.250 ;
        RECT 23.130 236.650 26.330 237.100 ;
        RECT 19.580 236.500 29.880 236.650 ;
        RECT 23.130 236.050 26.330 236.500 ;
        RECT 19.580 235.900 29.880 236.050 ;
        RECT 23.130 235.600 26.330 235.900 ;
        RECT 23.130 235.450 23.530 235.600 ;
        RECT 19.580 235.300 23.530 235.450 ;
        RECT 23.130 234.850 23.530 235.300 ;
        RECT 19.580 234.700 23.530 234.850 ;
        RECT 23.130 234.250 23.530 234.700 ;
        RECT 19.580 234.100 23.530 234.250 ;
        RECT 23.130 233.650 23.530 234.100 ;
        RECT 19.580 233.500 23.530 233.650 ;
        RECT 23.130 233.050 23.530 233.500 ;
        RECT 19.580 232.900 23.530 233.050 ;
        RECT 23.130 232.450 23.530 232.900 ;
        RECT 19.580 232.300 23.530 232.450 ;
        RECT 23.130 231.850 23.530 232.300 ;
        RECT 19.580 231.700 23.530 231.850 ;
        RECT 23.130 231.250 23.530 231.700 ;
        RECT 19.580 231.100 23.530 231.250 ;
        RECT 23.130 230.650 23.530 231.100 ;
        RECT 19.580 230.500 23.530 230.650 ;
        RECT 23.130 230.200 23.530 230.500 ;
        RECT 15.230 229.800 23.530 230.200 ;
        RECT 15.230 221.600 15.380 229.800 ;
        RECT 15.830 221.600 15.980 229.800 ;
        RECT 16.430 221.600 16.580 229.800 ;
        RECT 17.030 221.600 17.180 229.800 ;
        RECT 17.630 221.600 17.780 229.800 ;
        RECT 18.230 221.600 18.380 229.800 ;
        RECT 18.830 221.600 18.980 229.800 ;
        RECT 23.130 229.500 23.530 229.800 ;
        RECT 19.580 229.350 23.530 229.500 ;
        RECT 23.130 228.900 23.530 229.350 ;
        RECT 19.580 228.750 23.530 228.900 ;
        RECT 23.130 228.300 23.530 228.750 ;
        RECT 19.580 228.150 23.530 228.300 ;
        RECT 23.130 227.700 23.530 228.150 ;
        RECT 19.580 227.550 23.530 227.700 ;
        RECT 23.130 227.100 23.530 227.550 ;
        RECT 19.580 226.950 23.530 227.100 ;
        RECT 23.130 226.500 23.530 226.950 ;
        RECT 19.580 226.350 23.530 226.500 ;
        RECT 23.130 225.900 23.530 226.350 ;
        RECT 19.580 225.750 23.530 225.900 ;
        RECT 23.130 225.300 23.530 225.750 ;
        RECT 19.580 225.150 23.530 225.300 ;
        RECT 23.130 224.700 23.530 225.150 ;
        RECT 19.580 224.550 23.530 224.700 ;
        RECT 23.130 224.400 23.530 224.550 ;
        RECT 25.930 235.450 26.330 235.600 ;
        RECT 25.930 235.300 29.880 235.450 ;
        RECT 25.930 234.850 26.330 235.300 ;
        RECT 25.930 234.700 29.880 234.850 ;
        RECT 25.930 234.250 26.330 234.700 ;
        RECT 25.930 234.100 29.880 234.250 ;
        RECT 25.930 233.650 26.330 234.100 ;
        RECT 25.930 233.500 29.880 233.650 ;
        RECT 25.930 233.050 26.330 233.500 ;
        RECT 25.930 232.900 29.880 233.050 ;
        RECT 25.930 232.450 26.330 232.900 ;
        RECT 25.930 232.300 29.880 232.450 ;
        RECT 25.930 231.850 26.330 232.300 ;
        RECT 25.930 231.700 29.880 231.850 ;
        RECT 25.930 231.250 26.330 231.700 ;
        RECT 25.930 231.100 29.880 231.250 ;
        RECT 25.930 230.650 26.330 231.100 ;
        RECT 25.930 230.500 29.880 230.650 ;
        RECT 25.930 230.200 26.330 230.500 ;
        RECT 30.480 230.200 30.630 238.400 ;
        RECT 31.080 230.200 31.230 238.400 ;
        RECT 31.680 230.200 31.830 238.400 ;
        RECT 32.280 230.200 32.430 238.400 ;
        RECT 32.880 230.200 33.030 238.400 ;
        RECT 33.480 230.200 33.630 238.400 ;
        RECT 34.080 230.200 34.230 238.400 ;
        RECT 25.930 229.800 34.230 230.200 ;
        RECT 25.930 229.500 26.330 229.800 ;
        RECT 25.930 229.350 29.880 229.500 ;
        RECT 25.930 228.900 26.330 229.350 ;
        RECT 25.930 228.750 29.880 228.900 ;
        RECT 25.930 228.300 26.330 228.750 ;
        RECT 25.930 228.150 29.880 228.300 ;
        RECT 25.930 227.700 26.330 228.150 ;
        RECT 25.930 227.550 29.880 227.700 ;
        RECT 25.930 227.100 26.330 227.550 ;
        RECT 25.930 226.950 29.880 227.100 ;
        RECT 25.930 226.500 26.330 226.950 ;
        RECT 25.930 226.350 29.880 226.500 ;
        RECT 25.930 225.900 26.330 226.350 ;
        RECT 25.930 225.750 29.880 225.900 ;
        RECT 25.930 225.300 26.330 225.750 ;
        RECT 25.930 225.150 29.880 225.300 ;
        RECT 25.930 224.700 26.330 225.150 ;
        RECT 25.930 224.550 29.880 224.700 ;
        RECT 25.930 224.400 26.330 224.550 ;
        RECT 23.130 224.100 26.330 224.400 ;
        RECT 19.580 223.950 29.880 224.100 ;
        RECT 23.130 223.500 26.330 223.950 ;
        RECT 19.580 223.350 29.880 223.500 ;
        RECT 23.130 222.900 26.330 223.350 ;
        RECT 19.580 222.750 29.880 222.900 ;
        RECT 23.130 222.300 26.330 222.750 ;
        RECT 19.580 222.150 29.880 222.300 ;
        RECT 23.530 221.200 25.930 222.150 ;
        RECT 30.480 221.600 30.630 229.800 ;
        RECT 31.080 221.600 31.230 229.800 ;
        RECT 31.680 221.600 31.830 229.800 ;
        RECT 32.280 221.600 32.430 229.800 ;
        RECT 32.880 221.600 33.030 229.800 ;
        RECT 33.480 221.600 33.630 229.800 ;
        RECT 34.080 221.600 34.230 229.800 ;
        RECT 35.230 230.200 35.380 238.400 ;
        RECT 35.830 230.200 35.980 238.400 ;
        RECT 36.430 230.200 36.580 238.400 ;
        RECT 37.030 230.200 37.180 238.400 ;
        RECT 37.630 230.200 37.780 238.400 ;
        RECT 38.230 230.200 38.380 238.400 ;
        RECT 38.830 230.200 38.980 238.400 ;
        RECT 43.530 237.850 45.940 238.800 ;
        RECT 39.580 237.700 49.880 237.850 ;
        RECT 43.130 237.250 46.330 237.700 ;
        RECT 39.580 237.100 49.880 237.250 ;
        RECT 43.130 236.650 46.330 237.100 ;
        RECT 39.580 236.500 49.880 236.650 ;
        RECT 43.130 236.050 46.330 236.500 ;
        RECT 39.580 235.900 49.880 236.050 ;
        RECT 43.130 235.600 46.330 235.900 ;
        RECT 43.130 235.450 43.530 235.600 ;
        RECT 39.580 235.300 43.530 235.450 ;
        RECT 43.130 234.850 43.530 235.300 ;
        RECT 39.580 234.700 43.530 234.850 ;
        RECT 43.130 234.250 43.530 234.700 ;
        RECT 39.580 234.100 43.530 234.250 ;
        RECT 43.130 233.650 43.530 234.100 ;
        RECT 39.580 233.500 43.530 233.650 ;
        RECT 43.130 233.050 43.530 233.500 ;
        RECT 39.580 232.900 43.530 233.050 ;
        RECT 43.130 232.450 43.530 232.900 ;
        RECT 39.580 232.300 43.530 232.450 ;
        RECT 43.130 231.850 43.530 232.300 ;
        RECT 39.580 231.700 43.530 231.850 ;
        RECT 43.130 231.250 43.530 231.700 ;
        RECT 39.580 231.100 43.530 231.250 ;
        RECT 43.130 230.650 43.530 231.100 ;
        RECT 39.580 230.500 43.530 230.650 ;
        RECT 43.130 230.200 43.530 230.500 ;
        RECT 35.230 229.800 43.530 230.200 ;
        RECT 35.230 221.600 35.380 229.800 ;
        RECT 35.830 221.600 35.980 229.800 ;
        RECT 36.430 221.600 36.580 229.800 ;
        RECT 37.030 221.600 37.180 229.800 ;
        RECT 37.630 221.600 37.780 229.800 ;
        RECT 38.230 221.600 38.380 229.800 ;
        RECT 38.830 221.600 38.980 229.800 ;
        RECT 43.130 229.500 43.530 229.800 ;
        RECT 39.580 229.350 43.530 229.500 ;
        RECT 43.130 228.900 43.530 229.350 ;
        RECT 39.580 228.750 43.530 228.900 ;
        RECT 43.130 228.300 43.530 228.750 ;
        RECT 39.580 228.150 43.530 228.300 ;
        RECT 43.130 227.700 43.530 228.150 ;
        RECT 39.580 227.550 43.530 227.700 ;
        RECT 43.130 227.100 43.530 227.550 ;
        RECT 39.580 226.950 43.530 227.100 ;
        RECT 43.130 226.500 43.530 226.950 ;
        RECT 39.580 226.350 43.530 226.500 ;
        RECT 43.130 225.900 43.530 226.350 ;
        RECT 39.580 225.750 43.530 225.900 ;
        RECT 43.130 225.300 43.530 225.750 ;
        RECT 39.580 225.150 43.530 225.300 ;
        RECT 43.130 224.700 43.530 225.150 ;
        RECT 39.580 224.550 43.530 224.700 ;
        RECT 43.130 224.400 43.530 224.550 ;
        RECT 45.930 235.450 46.330 235.600 ;
        RECT 45.930 235.300 49.880 235.450 ;
        RECT 45.930 234.850 46.330 235.300 ;
        RECT 45.930 234.700 49.880 234.850 ;
        RECT 45.930 234.250 46.330 234.700 ;
        RECT 45.930 234.100 49.880 234.250 ;
        RECT 45.930 233.650 46.330 234.100 ;
        RECT 45.930 233.500 49.880 233.650 ;
        RECT 45.930 233.050 46.330 233.500 ;
        RECT 45.930 232.900 49.880 233.050 ;
        RECT 45.930 232.450 46.330 232.900 ;
        RECT 45.930 232.300 49.880 232.450 ;
        RECT 45.930 231.850 46.330 232.300 ;
        RECT 45.930 231.700 49.880 231.850 ;
        RECT 45.930 231.250 46.330 231.700 ;
        RECT 45.930 231.100 49.880 231.250 ;
        RECT 45.930 230.650 46.330 231.100 ;
        RECT 45.930 230.500 49.880 230.650 ;
        RECT 45.930 230.200 46.330 230.500 ;
        RECT 50.480 230.200 50.630 238.400 ;
        RECT 51.080 230.200 51.230 238.400 ;
        RECT 51.680 230.200 51.830 238.400 ;
        RECT 52.280 230.200 52.430 238.400 ;
        RECT 52.880 230.200 53.030 238.400 ;
        RECT 53.480 230.200 53.630 238.400 ;
        RECT 54.080 230.200 54.230 238.400 ;
        RECT 45.930 229.800 54.230 230.200 ;
        RECT 45.930 229.500 46.330 229.800 ;
        RECT 45.930 229.350 49.880 229.500 ;
        RECT 45.930 228.900 46.330 229.350 ;
        RECT 45.930 228.750 49.880 228.900 ;
        RECT 45.930 228.300 46.330 228.750 ;
        RECT 45.930 228.150 49.880 228.300 ;
        RECT 45.930 227.700 46.330 228.150 ;
        RECT 45.930 227.550 49.880 227.700 ;
        RECT 45.930 227.100 46.330 227.550 ;
        RECT 45.930 226.950 49.880 227.100 ;
        RECT 45.930 226.500 46.330 226.950 ;
        RECT 45.930 226.350 49.880 226.500 ;
        RECT 45.930 225.900 46.330 226.350 ;
        RECT 45.930 225.750 49.880 225.900 ;
        RECT 45.930 225.300 46.330 225.750 ;
        RECT 45.930 225.150 49.880 225.300 ;
        RECT 45.930 224.700 46.330 225.150 ;
        RECT 45.930 224.550 49.880 224.700 ;
        RECT 45.930 224.400 46.330 224.550 ;
        RECT 43.130 224.100 46.330 224.400 ;
        RECT 39.580 223.950 49.880 224.100 ;
        RECT 43.130 223.500 46.330 223.950 ;
        RECT 39.580 223.350 49.880 223.500 ;
        RECT 43.130 222.900 46.330 223.350 ;
        RECT 39.580 222.750 49.880 222.900 ;
        RECT 43.130 222.300 46.330 222.750 ;
        RECT 39.580 222.150 49.880 222.300 ;
        RECT 43.530 221.200 45.930 222.150 ;
        RECT 50.480 221.600 50.630 229.800 ;
        RECT 51.080 221.600 51.230 229.800 ;
        RECT 51.680 221.600 51.830 229.800 ;
        RECT 52.280 221.600 52.430 229.800 ;
        RECT 52.880 221.600 53.030 229.800 ;
        RECT 53.480 221.600 53.630 229.800 ;
        RECT 54.080 221.600 54.230 229.800 ;
        RECT 55.230 230.200 55.380 238.400 ;
        RECT 55.830 230.200 55.980 238.400 ;
        RECT 56.430 230.200 56.580 238.400 ;
        RECT 57.030 230.200 57.180 238.400 ;
        RECT 57.630 230.200 57.780 238.400 ;
        RECT 58.230 230.200 58.380 238.400 ;
        RECT 58.830 230.200 58.980 238.400 ;
        RECT 63.530 237.850 65.940 238.800 ;
        RECT 59.580 237.700 69.880 237.850 ;
        RECT 63.130 237.250 66.330 237.700 ;
        RECT 59.580 237.100 69.880 237.250 ;
        RECT 63.130 236.650 66.330 237.100 ;
        RECT 59.580 236.500 69.880 236.650 ;
        RECT 63.130 236.050 66.330 236.500 ;
        RECT 59.580 235.900 69.880 236.050 ;
        RECT 63.130 235.600 66.330 235.900 ;
        RECT 63.130 235.450 63.530 235.600 ;
        RECT 59.580 235.300 63.530 235.450 ;
        RECT 63.130 234.850 63.530 235.300 ;
        RECT 59.580 234.700 63.530 234.850 ;
        RECT 63.130 234.250 63.530 234.700 ;
        RECT 59.580 234.100 63.530 234.250 ;
        RECT 63.130 233.650 63.530 234.100 ;
        RECT 59.580 233.500 63.530 233.650 ;
        RECT 63.130 233.050 63.530 233.500 ;
        RECT 59.580 232.900 63.530 233.050 ;
        RECT 63.130 232.450 63.530 232.900 ;
        RECT 59.580 232.300 63.530 232.450 ;
        RECT 63.130 231.850 63.530 232.300 ;
        RECT 59.580 231.700 63.530 231.850 ;
        RECT 63.130 231.250 63.530 231.700 ;
        RECT 59.580 231.100 63.530 231.250 ;
        RECT 63.130 230.650 63.530 231.100 ;
        RECT 59.580 230.500 63.530 230.650 ;
        RECT 63.130 230.200 63.530 230.500 ;
        RECT 55.230 229.800 63.530 230.200 ;
        RECT 55.230 221.600 55.380 229.800 ;
        RECT 55.830 221.600 55.980 229.800 ;
        RECT 56.430 221.600 56.580 229.800 ;
        RECT 57.030 221.600 57.180 229.800 ;
        RECT 57.630 221.600 57.780 229.800 ;
        RECT 58.230 221.600 58.380 229.800 ;
        RECT 58.830 221.600 58.980 229.800 ;
        RECT 63.130 229.500 63.530 229.800 ;
        RECT 59.580 229.350 63.530 229.500 ;
        RECT 63.130 228.900 63.530 229.350 ;
        RECT 59.580 228.750 63.530 228.900 ;
        RECT 63.130 228.300 63.530 228.750 ;
        RECT 59.580 228.150 63.530 228.300 ;
        RECT 63.130 227.700 63.530 228.150 ;
        RECT 59.580 227.550 63.530 227.700 ;
        RECT 63.130 227.100 63.530 227.550 ;
        RECT 59.580 226.950 63.530 227.100 ;
        RECT 63.130 226.500 63.530 226.950 ;
        RECT 59.580 226.350 63.530 226.500 ;
        RECT 63.130 225.900 63.530 226.350 ;
        RECT 59.580 225.750 63.530 225.900 ;
        RECT 63.130 225.300 63.530 225.750 ;
        RECT 59.580 225.150 63.530 225.300 ;
        RECT 63.130 224.700 63.530 225.150 ;
        RECT 59.580 224.550 63.530 224.700 ;
        RECT 63.130 224.400 63.530 224.550 ;
        RECT 65.930 235.450 66.330 235.600 ;
        RECT 65.930 235.300 69.880 235.450 ;
        RECT 65.930 234.850 66.330 235.300 ;
        RECT 65.930 234.700 69.880 234.850 ;
        RECT 65.930 234.250 66.330 234.700 ;
        RECT 65.930 234.100 69.880 234.250 ;
        RECT 65.930 233.650 66.330 234.100 ;
        RECT 65.930 233.500 69.880 233.650 ;
        RECT 65.930 233.050 66.330 233.500 ;
        RECT 65.930 232.900 69.880 233.050 ;
        RECT 65.930 232.450 66.330 232.900 ;
        RECT 65.930 232.300 69.880 232.450 ;
        RECT 65.930 231.850 66.330 232.300 ;
        RECT 65.930 231.700 69.880 231.850 ;
        RECT 65.930 231.250 66.330 231.700 ;
        RECT 65.930 231.100 69.880 231.250 ;
        RECT 65.930 230.650 66.330 231.100 ;
        RECT 65.930 230.500 69.880 230.650 ;
        RECT 65.930 230.200 66.330 230.500 ;
        RECT 70.480 230.200 70.630 238.400 ;
        RECT 71.080 230.200 71.230 238.400 ;
        RECT 71.680 230.200 71.830 238.400 ;
        RECT 72.280 230.200 72.430 238.400 ;
        RECT 72.880 230.200 73.030 238.400 ;
        RECT 73.480 230.200 73.630 238.400 ;
        RECT 74.080 230.200 74.230 238.400 ;
        RECT 65.930 229.800 74.230 230.200 ;
        RECT 65.930 229.500 66.330 229.800 ;
        RECT 65.930 229.350 69.880 229.500 ;
        RECT 65.930 228.900 66.330 229.350 ;
        RECT 65.930 228.750 69.880 228.900 ;
        RECT 65.930 228.300 66.330 228.750 ;
        RECT 65.930 228.150 69.880 228.300 ;
        RECT 65.930 227.700 66.330 228.150 ;
        RECT 65.930 227.550 69.880 227.700 ;
        RECT 65.930 227.100 66.330 227.550 ;
        RECT 65.930 226.950 69.880 227.100 ;
        RECT 65.930 226.500 66.330 226.950 ;
        RECT 65.930 226.350 69.880 226.500 ;
        RECT 65.930 225.900 66.330 226.350 ;
        RECT 65.930 225.750 69.880 225.900 ;
        RECT 65.930 225.300 66.330 225.750 ;
        RECT 65.930 225.150 69.880 225.300 ;
        RECT 65.930 224.700 66.330 225.150 ;
        RECT 65.930 224.550 69.880 224.700 ;
        RECT 65.930 224.400 66.330 224.550 ;
        RECT 63.130 224.100 66.330 224.400 ;
        RECT 59.580 223.950 69.880 224.100 ;
        RECT 63.130 223.500 66.330 223.950 ;
        RECT 59.580 223.350 69.880 223.500 ;
        RECT 63.130 222.900 66.330 223.350 ;
        RECT 59.580 222.750 69.880 222.900 ;
        RECT 63.130 222.300 66.330 222.750 ;
        RECT 59.580 222.150 69.880 222.300 ;
        RECT 63.530 221.200 65.930 222.150 ;
        RECT 70.480 221.600 70.630 229.800 ;
        RECT 71.080 221.600 71.230 229.800 ;
        RECT 71.680 221.600 71.830 229.800 ;
        RECT 72.280 221.600 72.430 229.800 ;
        RECT 72.880 221.600 73.030 229.800 ;
        RECT 73.480 221.600 73.630 229.800 ;
        RECT 74.080 221.600 74.230 229.800 ;
        RECT 75.230 230.200 75.380 238.400 ;
        RECT 75.830 230.200 75.980 238.400 ;
        RECT 76.430 230.200 76.580 238.400 ;
        RECT 77.030 230.200 77.180 238.400 ;
        RECT 77.630 230.200 77.780 238.400 ;
        RECT 78.230 230.200 78.380 238.400 ;
        RECT 78.830 230.200 78.980 238.400 ;
        RECT 83.530 237.850 85.940 238.800 ;
        RECT 79.580 237.700 89.880 237.850 ;
        RECT 83.130 237.250 86.330 237.700 ;
        RECT 79.580 237.100 89.880 237.250 ;
        RECT 83.130 236.650 86.330 237.100 ;
        RECT 79.580 236.500 89.880 236.650 ;
        RECT 83.130 236.050 86.330 236.500 ;
        RECT 79.580 235.900 89.880 236.050 ;
        RECT 83.130 235.600 86.330 235.900 ;
        RECT 83.130 235.450 83.530 235.600 ;
        RECT 79.580 235.300 83.530 235.450 ;
        RECT 83.130 234.850 83.530 235.300 ;
        RECT 79.580 234.700 83.530 234.850 ;
        RECT 83.130 234.250 83.530 234.700 ;
        RECT 79.580 234.100 83.530 234.250 ;
        RECT 83.130 233.650 83.530 234.100 ;
        RECT 79.580 233.500 83.530 233.650 ;
        RECT 83.130 233.050 83.530 233.500 ;
        RECT 79.580 232.900 83.530 233.050 ;
        RECT 83.130 232.450 83.530 232.900 ;
        RECT 79.580 232.300 83.530 232.450 ;
        RECT 83.130 231.850 83.530 232.300 ;
        RECT 79.580 231.700 83.530 231.850 ;
        RECT 83.130 231.250 83.530 231.700 ;
        RECT 79.580 231.100 83.530 231.250 ;
        RECT 83.130 230.650 83.530 231.100 ;
        RECT 79.580 230.500 83.530 230.650 ;
        RECT 83.130 230.200 83.530 230.500 ;
        RECT 75.230 229.800 83.530 230.200 ;
        RECT 75.230 221.600 75.380 229.800 ;
        RECT 75.830 221.600 75.980 229.800 ;
        RECT 76.430 221.600 76.580 229.800 ;
        RECT 77.030 221.600 77.180 229.800 ;
        RECT 77.630 221.600 77.780 229.800 ;
        RECT 78.230 221.600 78.380 229.800 ;
        RECT 78.830 221.600 78.980 229.800 ;
        RECT 83.130 229.500 83.530 229.800 ;
        RECT 79.580 229.350 83.530 229.500 ;
        RECT 83.130 228.900 83.530 229.350 ;
        RECT 79.580 228.750 83.530 228.900 ;
        RECT 83.130 228.300 83.530 228.750 ;
        RECT 79.580 228.150 83.530 228.300 ;
        RECT 83.130 227.700 83.530 228.150 ;
        RECT 79.580 227.550 83.530 227.700 ;
        RECT 83.130 227.100 83.530 227.550 ;
        RECT 79.580 226.950 83.530 227.100 ;
        RECT 83.130 226.500 83.530 226.950 ;
        RECT 79.580 226.350 83.530 226.500 ;
        RECT 83.130 225.900 83.530 226.350 ;
        RECT 79.580 225.750 83.530 225.900 ;
        RECT 83.130 225.300 83.530 225.750 ;
        RECT 79.580 225.150 83.530 225.300 ;
        RECT 83.130 224.700 83.530 225.150 ;
        RECT 79.580 224.550 83.530 224.700 ;
        RECT 83.130 224.400 83.530 224.550 ;
        RECT 85.930 235.450 86.330 235.600 ;
        RECT 85.930 235.300 89.880 235.450 ;
        RECT 85.930 234.850 86.330 235.300 ;
        RECT 85.930 234.700 89.880 234.850 ;
        RECT 85.930 234.250 86.330 234.700 ;
        RECT 85.930 234.100 89.880 234.250 ;
        RECT 85.930 233.650 86.330 234.100 ;
        RECT 85.930 233.500 89.880 233.650 ;
        RECT 85.930 233.050 86.330 233.500 ;
        RECT 85.930 232.900 89.880 233.050 ;
        RECT 85.930 232.450 86.330 232.900 ;
        RECT 85.930 232.300 89.880 232.450 ;
        RECT 85.930 231.850 86.330 232.300 ;
        RECT 85.930 231.700 89.880 231.850 ;
        RECT 85.930 231.250 86.330 231.700 ;
        RECT 85.930 231.100 89.880 231.250 ;
        RECT 85.930 230.650 86.330 231.100 ;
        RECT 85.930 230.500 89.880 230.650 ;
        RECT 85.930 230.200 86.330 230.500 ;
        RECT 90.480 230.200 90.630 238.400 ;
        RECT 91.080 230.200 91.230 238.400 ;
        RECT 91.680 230.200 91.830 238.400 ;
        RECT 92.280 230.200 92.430 238.400 ;
        RECT 92.880 230.200 93.030 238.400 ;
        RECT 93.480 230.200 93.630 238.400 ;
        RECT 94.080 230.200 94.230 238.400 ;
        RECT 85.930 229.800 94.230 230.200 ;
        RECT 85.930 229.500 86.330 229.800 ;
        RECT 85.930 229.350 89.880 229.500 ;
        RECT 85.930 228.900 86.330 229.350 ;
        RECT 85.930 228.750 89.880 228.900 ;
        RECT 85.930 228.300 86.330 228.750 ;
        RECT 85.930 228.150 89.880 228.300 ;
        RECT 85.930 227.700 86.330 228.150 ;
        RECT 85.930 227.550 89.880 227.700 ;
        RECT 85.930 227.100 86.330 227.550 ;
        RECT 85.930 226.950 89.880 227.100 ;
        RECT 85.930 226.500 86.330 226.950 ;
        RECT 85.930 226.350 89.880 226.500 ;
        RECT 85.930 225.900 86.330 226.350 ;
        RECT 85.930 225.750 89.880 225.900 ;
        RECT 85.930 225.300 86.330 225.750 ;
        RECT 85.930 225.150 89.880 225.300 ;
        RECT 85.930 224.700 86.330 225.150 ;
        RECT 85.930 224.550 89.880 224.700 ;
        RECT 85.930 224.400 86.330 224.550 ;
        RECT 83.130 224.100 86.330 224.400 ;
        RECT 79.580 223.950 89.880 224.100 ;
        RECT 83.130 223.500 86.330 223.950 ;
        RECT 79.580 223.350 89.880 223.500 ;
        RECT 83.130 222.900 86.330 223.350 ;
        RECT 79.580 222.750 89.880 222.900 ;
        RECT 83.130 222.300 86.330 222.750 ;
        RECT 79.580 222.150 89.880 222.300 ;
        RECT 83.530 221.200 85.930 222.150 ;
        RECT 90.480 221.600 90.630 229.800 ;
        RECT 91.080 221.600 91.230 229.800 ;
        RECT 91.680 221.600 91.830 229.800 ;
        RECT 92.280 221.600 92.430 229.800 ;
        RECT 92.880 221.600 93.030 229.800 ;
        RECT 93.480 221.600 93.630 229.800 ;
        RECT 94.080 221.600 94.230 229.800 ;
        RECT 95.230 230.200 95.380 238.400 ;
        RECT 95.830 230.200 95.980 238.400 ;
        RECT 96.430 230.200 96.580 238.400 ;
        RECT 97.030 230.200 97.180 238.400 ;
        RECT 97.630 230.200 97.780 238.400 ;
        RECT 98.230 230.200 98.380 238.400 ;
        RECT 98.830 230.200 98.980 238.400 ;
        RECT 103.530 237.850 105.940 238.800 ;
        RECT 99.580 237.700 109.880 237.850 ;
        RECT 103.130 237.250 106.330 237.700 ;
        RECT 99.580 237.100 109.880 237.250 ;
        RECT 103.130 236.650 106.330 237.100 ;
        RECT 99.580 236.500 109.880 236.650 ;
        RECT 103.130 236.050 106.330 236.500 ;
        RECT 99.580 235.900 109.880 236.050 ;
        RECT 103.130 235.600 106.330 235.900 ;
        RECT 103.130 235.450 103.530 235.600 ;
        RECT 99.580 235.300 103.530 235.450 ;
        RECT 103.130 234.850 103.530 235.300 ;
        RECT 99.580 234.700 103.530 234.850 ;
        RECT 103.130 234.250 103.530 234.700 ;
        RECT 99.580 234.100 103.530 234.250 ;
        RECT 103.130 233.650 103.530 234.100 ;
        RECT 99.580 233.500 103.530 233.650 ;
        RECT 103.130 233.050 103.530 233.500 ;
        RECT 99.580 232.900 103.530 233.050 ;
        RECT 103.130 232.450 103.530 232.900 ;
        RECT 99.580 232.300 103.530 232.450 ;
        RECT 103.130 231.850 103.530 232.300 ;
        RECT 99.580 231.700 103.530 231.850 ;
        RECT 103.130 231.250 103.530 231.700 ;
        RECT 99.580 231.100 103.530 231.250 ;
        RECT 103.130 230.650 103.530 231.100 ;
        RECT 99.580 230.500 103.530 230.650 ;
        RECT 103.130 230.200 103.530 230.500 ;
        RECT 95.230 229.800 103.530 230.200 ;
        RECT 95.230 221.600 95.380 229.800 ;
        RECT 95.830 221.600 95.980 229.800 ;
        RECT 96.430 221.600 96.580 229.800 ;
        RECT 97.030 221.600 97.180 229.800 ;
        RECT 97.630 221.600 97.780 229.800 ;
        RECT 98.230 221.600 98.380 229.800 ;
        RECT 98.830 221.600 98.980 229.800 ;
        RECT 103.130 229.500 103.530 229.800 ;
        RECT 99.580 229.350 103.530 229.500 ;
        RECT 103.130 228.900 103.530 229.350 ;
        RECT 99.580 228.750 103.530 228.900 ;
        RECT 103.130 228.300 103.530 228.750 ;
        RECT 99.580 228.150 103.530 228.300 ;
        RECT 103.130 227.700 103.530 228.150 ;
        RECT 99.580 227.550 103.530 227.700 ;
        RECT 103.130 227.100 103.530 227.550 ;
        RECT 99.580 226.950 103.530 227.100 ;
        RECT 103.130 226.500 103.530 226.950 ;
        RECT 99.580 226.350 103.530 226.500 ;
        RECT 103.130 225.900 103.530 226.350 ;
        RECT 99.580 225.750 103.530 225.900 ;
        RECT 103.130 225.300 103.530 225.750 ;
        RECT 99.580 225.150 103.530 225.300 ;
        RECT 103.130 224.700 103.530 225.150 ;
        RECT 99.580 224.550 103.530 224.700 ;
        RECT 103.130 224.400 103.530 224.550 ;
        RECT 105.930 235.450 106.330 235.600 ;
        RECT 105.930 235.300 109.880 235.450 ;
        RECT 105.930 234.850 106.330 235.300 ;
        RECT 105.930 234.700 109.880 234.850 ;
        RECT 105.930 234.250 106.330 234.700 ;
        RECT 105.930 234.100 109.880 234.250 ;
        RECT 105.930 233.650 106.330 234.100 ;
        RECT 105.930 233.500 109.880 233.650 ;
        RECT 105.930 233.050 106.330 233.500 ;
        RECT 105.930 232.900 109.880 233.050 ;
        RECT 105.930 232.450 106.330 232.900 ;
        RECT 105.930 232.300 109.880 232.450 ;
        RECT 105.930 231.850 106.330 232.300 ;
        RECT 105.930 231.700 109.880 231.850 ;
        RECT 105.930 231.250 106.330 231.700 ;
        RECT 105.930 231.100 109.880 231.250 ;
        RECT 105.930 230.650 106.330 231.100 ;
        RECT 105.930 230.500 109.880 230.650 ;
        RECT 105.930 230.200 106.330 230.500 ;
        RECT 110.480 230.200 110.630 238.400 ;
        RECT 111.080 230.200 111.230 238.400 ;
        RECT 111.680 230.200 111.830 238.400 ;
        RECT 112.280 230.200 112.430 238.400 ;
        RECT 112.880 230.200 113.030 238.400 ;
        RECT 113.480 230.200 113.630 238.400 ;
        RECT 114.080 230.200 114.230 238.400 ;
        RECT 105.930 229.800 114.230 230.200 ;
        RECT 105.930 229.500 106.330 229.800 ;
        RECT 105.930 229.350 109.880 229.500 ;
        RECT 105.930 228.900 106.330 229.350 ;
        RECT 105.930 228.750 109.880 228.900 ;
        RECT 105.930 228.300 106.330 228.750 ;
        RECT 105.930 228.150 109.880 228.300 ;
        RECT 105.930 227.700 106.330 228.150 ;
        RECT 105.930 227.550 109.880 227.700 ;
        RECT 105.930 227.100 106.330 227.550 ;
        RECT 105.930 226.950 109.880 227.100 ;
        RECT 105.930 226.500 106.330 226.950 ;
        RECT 105.930 226.350 109.880 226.500 ;
        RECT 105.930 225.900 106.330 226.350 ;
        RECT 105.930 225.750 109.880 225.900 ;
        RECT 105.930 225.300 106.330 225.750 ;
        RECT 105.930 225.150 109.880 225.300 ;
        RECT 105.930 224.700 106.330 225.150 ;
        RECT 105.930 224.550 109.880 224.700 ;
        RECT 105.930 224.400 106.330 224.550 ;
        RECT 103.130 224.100 106.330 224.400 ;
        RECT 99.580 223.950 109.880 224.100 ;
        RECT 103.130 223.500 106.330 223.950 ;
        RECT 99.580 223.350 109.880 223.500 ;
        RECT 103.130 222.900 106.330 223.350 ;
        RECT 99.580 222.750 109.880 222.900 ;
        RECT 103.130 222.300 106.330 222.750 ;
        RECT 99.580 222.150 109.880 222.300 ;
        RECT 103.530 221.200 105.930 222.150 ;
        RECT 110.480 221.600 110.630 229.800 ;
        RECT 111.080 221.600 111.230 229.800 ;
        RECT 111.680 221.600 111.830 229.800 ;
        RECT 112.280 221.600 112.430 229.800 ;
        RECT 112.880 221.600 113.030 229.800 ;
        RECT 113.480 221.600 113.630 229.800 ;
        RECT 114.080 221.600 114.230 229.800 ;
        RECT 115.230 230.200 115.380 238.400 ;
        RECT 115.830 230.200 115.980 238.400 ;
        RECT 116.430 230.200 116.580 238.400 ;
        RECT 117.030 230.200 117.180 238.400 ;
        RECT 117.630 230.200 117.780 238.400 ;
        RECT 118.230 230.200 118.380 238.400 ;
        RECT 118.830 230.200 118.980 238.400 ;
        RECT 123.530 237.850 124.730 238.800 ;
        RECT 119.580 237.700 124.730 237.850 ;
        RECT 123.130 237.250 124.730 237.700 ;
        RECT 119.580 237.100 124.730 237.250 ;
        RECT 123.130 236.650 124.730 237.100 ;
        RECT 119.580 236.500 124.730 236.650 ;
        RECT 123.130 236.050 124.730 236.500 ;
        RECT 125.140 236.050 127.140 237.325 ;
        RECT 119.580 235.900 124.730 236.050 ;
        RECT 123.130 235.600 124.730 235.900 ;
        RECT 123.130 235.450 123.530 235.600 ;
        RECT 119.580 235.300 123.530 235.450 ;
        RECT 123.130 234.850 123.530 235.300 ;
        RECT 119.580 234.700 123.530 234.850 ;
        RECT 123.130 234.250 123.530 234.700 ;
        RECT 119.580 234.100 123.530 234.250 ;
        RECT 123.130 233.650 123.530 234.100 ;
        RECT 119.580 233.500 123.530 233.650 ;
        RECT 123.130 233.050 123.530 233.500 ;
        RECT 119.580 232.900 123.530 233.050 ;
        RECT 123.130 232.450 123.530 232.900 ;
        RECT 119.580 232.300 123.530 232.450 ;
        RECT 123.130 231.850 123.530 232.300 ;
        RECT 119.580 231.700 123.530 231.850 ;
        RECT 123.130 231.250 123.530 231.700 ;
        RECT 119.580 231.100 123.530 231.250 ;
        RECT 123.130 230.650 123.530 231.100 ;
        RECT 119.580 230.500 123.530 230.650 ;
        RECT 123.130 230.200 123.530 230.500 ;
        RECT 115.230 229.800 123.530 230.200 ;
        RECT 115.230 221.600 115.380 229.800 ;
        RECT 115.830 221.600 115.980 229.800 ;
        RECT 116.430 221.600 116.580 229.800 ;
        RECT 117.030 221.600 117.180 229.800 ;
        RECT 117.630 221.600 117.780 229.800 ;
        RECT 118.230 221.600 118.380 229.800 ;
        RECT 118.830 221.600 118.980 229.800 ;
        RECT 123.130 229.500 123.530 229.800 ;
        RECT 119.580 229.350 123.530 229.500 ;
        RECT 123.130 228.900 123.530 229.350 ;
        RECT 119.580 228.750 123.530 228.900 ;
        RECT 123.130 228.300 123.530 228.750 ;
        RECT 119.580 228.150 123.530 228.300 ;
        RECT 123.130 227.700 123.530 228.150 ;
        RECT 119.580 227.550 123.530 227.700 ;
        RECT 123.130 227.100 123.530 227.550 ;
        RECT 119.580 226.950 123.530 227.100 ;
        RECT 123.130 226.500 123.530 226.950 ;
        RECT 119.580 226.350 123.530 226.500 ;
        RECT 123.130 225.900 123.530 226.350 ;
        RECT 119.580 225.750 123.530 225.900 ;
        RECT 123.130 225.300 123.530 225.750 ;
        RECT 119.580 225.150 123.530 225.300 ;
        RECT 123.130 224.700 123.530 225.150 ;
        RECT 119.580 224.550 123.530 224.700 ;
        RECT 123.130 224.400 123.530 224.550 ;
        RECT 123.130 224.100 124.730 224.400 ;
        RECT 119.580 223.950 124.730 224.100 ;
        RECT 123.130 223.500 124.730 223.950 ;
        RECT 119.580 223.350 124.730 223.500 ;
        RECT 123.130 222.900 124.730 223.350 ;
        RECT 119.580 222.750 124.730 222.900 ;
        RECT 123.130 222.300 124.730 222.750 ;
        RECT 119.580 222.150 124.730 222.300 ;
        RECT 125.140 222.255 127.140 223.530 ;
        RECT 123.530 221.200 124.730 222.150 ;
        RECT 4.730 218.800 9.130 221.200 ;
        RECT 20.330 218.800 29.130 221.200 ;
        RECT 40.330 218.800 49.130 221.200 ;
        RECT 60.330 218.800 69.130 221.200 ;
        RECT 80.330 218.800 89.130 221.200 ;
        RECT 100.330 218.800 109.130 221.200 ;
        RECT 120.330 218.800 124.730 221.200 ;
        RECT 2.315 216.695 4.320 217.970 ;
        RECT 4.730 217.850 5.940 218.800 ;
        RECT 4.730 217.700 9.880 217.850 ;
        RECT 4.730 217.250 6.330 217.700 ;
        RECT 4.730 217.100 9.880 217.250 ;
        RECT 4.730 216.650 6.330 217.100 ;
        RECT 4.730 216.500 9.880 216.650 ;
        RECT 4.730 216.050 6.330 216.500 ;
        RECT 4.730 215.900 9.880 216.050 ;
        RECT 4.730 215.600 6.330 215.900 ;
        RECT 2.315 213.250 4.315 215.545 ;
        RECT 5.930 215.450 6.330 215.600 ;
        RECT 5.930 215.300 9.880 215.450 ;
        RECT 5.930 214.850 6.330 215.300 ;
        RECT 5.930 214.700 9.880 214.850 ;
        RECT 5.930 214.250 6.330 214.700 ;
        RECT 5.930 214.100 9.880 214.250 ;
        RECT 5.930 213.650 6.330 214.100 ;
        RECT 5.930 213.500 9.880 213.650 ;
        RECT 5.930 213.050 6.330 213.500 ;
        RECT 5.930 212.900 9.880 213.050 ;
        RECT 5.930 212.450 6.330 212.900 ;
        RECT 5.930 212.300 9.880 212.450 ;
        RECT 5.930 211.850 6.330 212.300 ;
        RECT 5.930 211.700 9.880 211.850 ;
        RECT 5.930 211.250 6.330 211.700 ;
        RECT 5.930 211.100 9.880 211.250 ;
        RECT 5.930 210.650 6.330 211.100 ;
        RECT 5.930 210.500 9.880 210.650 ;
        RECT 5.930 210.200 6.330 210.500 ;
        RECT 10.480 210.200 10.630 218.400 ;
        RECT 11.080 210.200 11.230 218.400 ;
        RECT 11.680 210.200 11.830 218.400 ;
        RECT 12.280 210.200 12.430 218.400 ;
        RECT 12.880 210.200 13.030 218.400 ;
        RECT 13.480 210.200 13.630 218.400 ;
        RECT 14.080 210.200 14.230 218.400 ;
        RECT 5.930 209.800 14.230 210.200 ;
        RECT 5.930 209.500 6.330 209.800 ;
        RECT 5.930 209.350 9.880 209.500 ;
        RECT 5.930 208.900 6.330 209.350 ;
        RECT 5.930 208.750 9.880 208.900 ;
        RECT 5.930 208.300 6.330 208.750 ;
        RECT 5.930 208.150 9.880 208.300 ;
        RECT 5.930 207.700 6.330 208.150 ;
        RECT 5.930 207.550 9.880 207.700 ;
        RECT 5.930 207.100 6.330 207.550 ;
        RECT 5.930 206.950 9.880 207.100 ;
        RECT 2.315 204.455 4.315 206.750 ;
        RECT 5.930 206.500 6.330 206.950 ;
        RECT 5.930 206.350 9.880 206.500 ;
        RECT 5.930 205.900 6.330 206.350 ;
        RECT 5.930 205.750 9.880 205.900 ;
        RECT 5.930 205.300 6.330 205.750 ;
        RECT 5.930 205.150 9.880 205.300 ;
        RECT 5.930 204.700 6.330 205.150 ;
        RECT 5.930 204.550 9.880 204.700 ;
        RECT 2.315 204.450 4.180 204.455 ;
        RECT 5.930 204.400 6.330 204.550 ;
        RECT 4.730 204.100 6.330 204.400 ;
        RECT 4.730 203.950 9.880 204.100 ;
        RECT 4.730 203.500 6.330 203.950 ;
        RECT 4.730 203.350 9.880 203.500 ;
        RECT 4.730 202.900 6.330 203.350 ;
        RECT 4.730 202.750 9.880 202.900 ;
        RECT 2.315 201.395 4.315 202.670 ;
        RECT 4.730 202.300 6.330 202.750 ;
        RECT 4.730 202.150 9.880 202.300 ;
        RECT 4.730 201.200 5.930 202.150 ;
        RECT 10.480 201.600 10.630 209.800 ;
        RECT 11.080 201.600 11.230 209.800 ;
        RECT 11.680 201.600 11.830 209.800 ;
        RECT 12.280 201.600 12.430 209.800 ;
        RECT 12.880 201.600 13.030 209.800 ;
        RECT 13.480 201.600 13.630 209.800 ;
        RECT 14.080 201.600 14.230 209.800 ;
        RECT 15.230 210.200 15.380 218.400 ;
        RECT 15.830 210.200 15.980 218.400 ;
        RECT 16.430 210.200 16.580 218.400 ;
        RECT 17.030 210.200 17.180 218.400 ;
        RECT 17.630 210.200 17.780 218.400 ;
        RECT 18.230 210.200 18.380 218.400 ;
        RECT 18.830 210.200 18.980 218.400 ;
        RECT 23.530 217.850 25.940 218.800 ;
        RECT 19.580 217.700 29.880 217.850 ;
        RECT 23.130 217.250 26.330 217.700 ;
        RECT 19.580 217.100 29.880 217.250 ;
        RECT 23.130 216.650 26.330 217.100 ;
        RECT 19.580 216.500 29.880 216.650 ;
        RECT 23.130 216.050 26.330 216.500 ;
        RECT 19.580 215.900 29.880 216.050 ;
        RECT 23.130 215.600 26.330 215.900 ;
        RECT 23.130 215.450 23.530 215.600 ;
        RECT 19.580 215.300 23.530 215.450 ;
        RECT 23.130 214.850 23.530 215.300 ;
        RECT 19.580 214.700 23.530 214.850 ;
        RECT 23.130 214.250 23.530 214.700 ;
        RECT 19.580 214.100 23.530 214.250 ;
        RECT 23.130 213.650 23.530 214.100 ;
        RECT 19.580 213.500 23.530 213.650 ;
        RECT 23.130 213.050 23.530 213.500 ;
        RECT 19.580 212.900 23.530 213.050 ;
        RECT 23.130 212.450 23.530 212.900 ;
        RECT 19.580 212.300 23.530 212.450 ;
        RECT 23.130 211.850 23.530 212.300 ;
        RECT 19.580 211.700 23.530 211.850 ;
        RECT 23.130 211.250 23.530 211.700 ;
        RECT 19.580 211.100 23.530 211.250 ;
        RECT 23.130 210.650 23.530 211.100 ;
        RECT 19.580 210.500 23.530 210.650 ;
        RECT 23.130 210.200 23.530 210.500 ;
        RECT 15.230 209.800 23.530 210.200 ;
        RECT 15.230 201.600 15.380 209.800 ;
        RECT 15.830 201.600 15.980 209.800 ;
        RECT 16.430 201.600 16.580 209.800 ;
        RECT 17.030 201.600 17.180 209.800 ;
        RECT 17.630 201.600 17.780 209.800 ;
        RECT 18.230 201.600 18.380 209.800 ;
        RECT 18.830 201.600 18.980 209.800 ;
        RECT 23.130 209.500 23.530 209.800 ;
        RECT 19.580 209.350 23.530 209.500 ;
        RECT 23.130 208.900 23.530 209.350 ;
        RECT 19.580 208.750 23.530 208.900 ;
        RECT 23.130 208.300 23.530 208.750 ;
        RECT 19.580 208.150 23.530 208.300 ;
        RECT 23.130 207.700 23.530 208.150 ;
        RECT 19.580 207.550 23.530 207.700 ;
        RECT 23.130 207.100 23.530 207.550 ;
        RECT 19.580 206.950 23.530 207.100 ;
        RECT 23.130 206.500 23.530 206.950 ;
        RECT 19.580 206.350 23.530 206.500 ;
        RECT 23.130 205.900 23.530 206.350 ;
        RECT 19.580 205.750 23.530 205.900 ;
        RECT 23.130 205.300 23.530 205.750 ;
        RECT 19.580 205.150 23.530 205.300 ;
        RECT 23.130 204.700 23.530 205.150 ;
        RECT 19.580 204.550 23.530 204.700 ;
        RECT 23.130 204.400 23.530 204.550 ;
        RECT 25.930 215.450 26.330 215.600 ;
        RECT 25.930 215.300 29.880 215.450 ;
        RECT 25.930 214.850 26.330 215.300 ;
        RECT 25.930 214.700 29.880 214.850 ;
        RECT 25.930 214.250 26.330 214.700 ;
        RECT 25.930 214.100 29.880 214.250 ;
        RECT 25.930 213.650 26.330 214.100 ;
        RECT 25.930 213.500 29.880 213.650 ;
        RECT 25.930 213.050 26.330 213.500 ;
        RECT 25.930 212.900 29.880 213.050 ;
        RECT 25.930 212.450 26.330 212.900 ;
        RECT 25.930 212.300 29.880 212.450 ;
        RECT 25.930 211.850 26.330 212.300 ;
        RECT 25.930 211.700 29.880 211.850 ;
        RECT 25.930 211.250 26.330 211.700 ;
        RECT 25.930 211.100 29.880 211.250 ;
        RECT 25.930 210.650 26.330 211.100 ;
        RECT 25.930 210.500 29.880 210.650 ;
        RECT 25.930 210.200 26.330 210.500 ;
        RECT 30.480 210.200 30.630 218.400 ;
        RECT 31.080 210.200 31.230 218.400 ;
        RECT 31.680 210.200 31.830 218.400 ;
        RECT 32.280 210.200 32.430 218.400 ;
        RECT 32.880 210.200 33.030 218.400 ;
        RECT 33.480 210.200 33.630 218.400 ;
        RECT 34.080 210.200 34.230 218.400 ;
        RECT 25.930 209.800 34.230 210.200 ;
        RECT 25.930 209.500 26.330 209.800 ;
        RECT 25.930 209.350 29.880 209.500 ;
        RECT 25.930 208.900 26.330 209.350 ;
        RECT 25.930 208.750 29.880 208.900 ;
        RECT 25.930 208.300 26.330 208.750 ;
        RECT 25.930 208.150 29.880 208.300 ;
        RECT 25.930 207.700 26.330 208.150 ;
        RECT 25.930 207.550 29.880 207.700 ;
        RECT 25.930 207.100 26.330 207.550 ;
        RECT 25.930 206.950 29.880 207.100 ;
        RECT 25.930 206.500 26.330 206.950 ;
        RECT 25.930 206.350 29.880 206.500 ;
        RECT 25.930 205.900 26.330 206.350 ;
        RECT 25.930 205.750 29.880 205.900 ;
        RECT 25.930 205.300 26.330 205.750 ;
        RECT 25.930 205.150 29.880 205.300 ;
        RECT 25.930 204.700 26.330 205.150 ;
        RECT 25.930 204.550 29.880 204.700 ;
        RECT 25.930 204.400 26.330 204.550 ;
        RECT 23.130 204.100 26.330 204.400 ;
        RECT 19.580 203.950 29.880 204.100 ;
        RECT 23.130 203.500 26.330 203.950 ;
        RECT 19.580 203.350 29.880 203.500 ;
        RECT 23.130 202.900 26.330 203.350 ;
        RECT 19.580 202.750 29.880 202.900 ;
        RECT 23.130 202.300 26.330 202.750 ;
        RECT 19.580 202.150 29.880 202.300 ;
        RECT 23.530 201.200 25.930 202.150 ;
        RECT 30.480 201.600 30.630 209.800 ;
        RECT 31.080 201.600 31.230 209.800 ;
        RECT 31.680 201.600 31.830 209.800 ;
        RECT 32.280 201.600 32.430 209.800 ;
        RECT 32.880 201.600 33.030 209.800 ;
        RECT 33.480 201.600 33.630 209.800 ;
        RECT 34.080 201.600 34.230 209.800 ;
        RECT 35.230 210.200 35.380 218.400 ;
        RECT 35.830 210.200 35.980 218.400 ;
        RECT 36.430 210.200 36.580 218.400 ;
        RECT 37.030 210.200 37.180 218.400 ;
        RECT 37.630 210.200 37.780 218.400 ;
        RECT 38.230 210.200 38.380 218.400 ;
        RECT 38.830 210.200 38.980 218.400 ;
        RECT 43.530 217.850 45.940 218.800 ;
        RECT 39.580 217.700 49.880 217.850 ;
        RECT 43.130 217.250 46.330 217.700 ;
        RECT 39.580 217.100 49.880 217.250 ;
        RECT 43.130 216.650 46.330 217.100 ;
        RECT 39.580 216.500 49.880 216.650 ;
        RECT 43.130 216.050 46.330 216.500 ;
        RECT 39.580 215.900 49.880 216.050 ;
        RECT 43.130 215.600 46.330 215.900 ;
        RECT 43.130 215.450 43.530 215.600 ;
        RECT 39.580 215.300 43.530 215.450 ;
        RECT 43.130 214.850 43.530 215.300 ;
        RECT 39.580 214.700 43.530 214.850 ;
        RECT 43.130 214.250 43.530 214.700 ;
        RECT 39.580 214.100 43.530 214.250 ;
        RECT 43.130 213.650 43.530 214.100 ;
        RECT 39.580 213.500 43.530 213.650 ;
        RECT 43.130 213.050 43.530 213.500 ;
        RECT 39.580 212.900 43.530 213.050 ;
        RECT 43.130 212.450 43.530 212.900 ;
        RECT 39.580 212.300 43.530 212.450 ;
        RECT 43.130 211.850 43.530 212.300 ;
        RECT 39.580 211.700 43.530 211.850 ;
        RECT 43.130 211.250 43.530 211.700 ;
        RECT 39.580 211.100 43.530 211.250 ;
        RECT 43.130 210.650 43.530 211.100 ;
        RECT 39.580 210.500 43.530 210.650 ;
        RECT 43.130 210.200 43.530 210.500 ;
        RECT 35.230 209.800 43.530 210.200 ;
        RECT 35.230 201.600 35.380 209.800 ;
        RECT 35.830 201.600 35.980 209.800 ;
        RECT 36.430 201.600 36.580 209.800 ;
        RECT 37.030 201.600 37.180 209.800 ;
        RECT 37.630 201.600 37.780 209.800 ;
        RECT 38.230 201.600 38.380 209.800 ;
        RECT 38.830 201.600 38.980 209.800 ;
        RECT 43.130 209.500 43.530 209.800 ;
        RECT 39.580 209.350 43.530 209.500 ;
        RECT 43.130 208.900 43.530 209.350 ;
        RECT 39.580 208.750 43.530 208.900 ;
        RECT 43.130 208.300 43.530 208.750 ;
        RECT 39.580 208.150 43.530 208.300 ;
        RECT 43.130 207.700 43.530 208.150 ;
        RECT 39.580 207.550 43.530 207.700 ;
        RECT 43.130 207.100 43.530 207.550 ;
        RECT 39.580 206.950 43.530 207.100 ;
        RECT 43.130 206.500 43.530 206.950 ;
        RECT 39.580 206.350 43.530 206.500 ;
        RECT 43.130 205.900 43.530 206.350 ;
        RECT 39.580 205.750 43.530 205.900 ;
        RECT 43.130 205.300 43.530 205.750 ;
        RECT 39.580 205.150 43.530 205.300 ;
        RECT 43.130 204.700 43.530 205.150 ;
        RECT 39.580 204.550 43.530 204.700 ;
        RECT 43.130 204.400 43.530 204.550 ;
        RECT 45.930 215.450 46.330 215.600 ;
        RECT 45.930 215.300 49.880 215.450 ;
        RECT 45.930 214.850 46.330 215.300 ;
        RECT 45.930 214.700 49.880 214.850 ;
        RECT 45.930 214.250 46.330 214.700 ;
        RECT 45.930 214.100 49.880 214.250 ;
        RECT 45.930 213.650 46.330 214.100 ;
        RECT 45.930 213.500 49.880 213.650 ;
        RECT 45.930 213.050 46.330 213.500 ;
        RECT 45.930 212.900 49.880 213.050 ;
        RECT 45.930 212.450 46.330 212.900 ;
        RECT 45.930 212.300 49.880 212.450 ;
        RECT 45.930 211.850 46.330 212.300 ;
        RECT 45.930 211.700 49.880 211.850 ;
        RECT 45.930 211.250 46.330 211.700 ;
        RECT 45.930 211.100 49.880 211.250 ;
        RECT 45.930 210.650 46.330 211.100 ;
        RECT 45.930 210.500 49.880 210.650 ;
        RECT 45.930 210.200 46.330 210.500 ;
        RECT 50.480 210.200 50.630 218.400 ;
        RECT 51.080 210.200 51.230 218.400 ;
        RECT 51.680 210.200 51.830 218.400 ;
        RECT 52.280 210.200 52.430 218.400 ;
        RECT 52.880 210.200 53.030 218.400 ;
        RECT 53.480 210.200 53.630 218.400 ;
        RECT 54.080 210.200 54.230 218.400 ;
        RECT 45.930 209.800 54.230 210.200 ;
        RECT 45.930 209.500 46.330 209.800 ;
        RECT 45.930 209.350 49.880 209.500 ;
        RECT 45.930 208.900 46.330 209.350 ;
        RECT 45.930 208.750 49.880 208.900 ;
        RECT 45.930 208.300 46.330 208.750 ;
        RECT 45.930 208.150 49.880 208.300 ;
        RECT 45.930 207.700 46.330 208.150 ;
        RECT 45.930 207.550 49.880 207.700 ;
        RECT 45.930 207.100 46.330 207.550 ;
        RECT 45.930 206.950 49.880 207.100 ;
        RECT 45.930 206.500 46.330 206.950 ;
        RECT 45.930 206.350 49.880 206.500 ;
        RECT 45.930 205.900 46.330 206.350 ;
        RECT 45.930 205.750 49.880 205.900 ;
        RECT 45.930 205.300 46.330 205.750 ;
        RECT 45.930 205.150 49.880 205.300 ;
        RECT 45.930 204.700 46.330 205.150 ;
        RECT 45.930 204.550 49.880 204.700 ;
        RECT 45.930 204.400 46.330 204.550 ;
        RECT 43.130 204.100 46.330 204.400 ;
        RECT 39.580 203.950 49.880 204.100 ;
        RECT 43.130 203.500 46.330 203.950 ;
        RECT 39.580 203.350 49.880 203.500 ;
        RECT 43.130 202.900 46.330 203.350 ;
        RECT 39.580 202.750 49.880 202.900 ;
        RECT 43.130 202.300 46.330 202.750 ;
        RECT 39.580 202.150 49.880 202.300 ;
        RECT 43.530 201.200 45.930 202.150 ;
        RECT 50.480 201.600 50.630 209.800 ;
        RECT 51.080 201.600 51.230 209.800 ;
        RECT 51.680 201.600 51.830 209.800 ;
        RECT 52.280 201.600 52.430 209.800 ;
        RECT 52.880 201.600 53.030 209.800 ;
        RECT 53.480 201.600 53.630 209.800 ;
        RECT 54.080 201.600 54.230 209.800 ;
        RECT 55.230 210.200 55.380 218.400 ;
        RECT 55.830 210.200 55.980 218.400 ;
        RECT 56.430 210.200 56.580 218.400 ;
        RECT 57.030 210.200 57.180 218.400 ;
        RECT 57.630 210.200 57.780 218.400 ;
        RECT 58.230 210.200 58.380 218.400 ;
        RECT 58.830 210.200 58.980 218.400 ;
        RECT 63.530 217.850 65.940 218.800 ;
        RECT 59.580 217.700 69.880 217.850 ;
        RECT 63.130 217.250 66.330 217.700 ;
        RECT 59.580 217.100 69.880 217.250 ;
        RECT 63.130 216.650 66.330 217.100 ;
        RECT 59.580 216.500 69.880 216.650 ;
        RECT 63.130 216.050 66.330 216.500 ;
        RECT 59.580 215.900 69.880 216.050 ;
        RECT 63.130 215.600 66.330 215.900 ;
        RECT 63.130 215.450 63.530 215.600 ;
        RECT 59.580 215.300 63.530 215.450 ;
        RECT 63.130 214.850 63.530 215.300 ;
        RECT 59.580 214.700 63.530 214.850 ;
        RECT 63.130 214.250 63.530 214.700 ;
        RECT 59.580 214.100 63.530 214.250 ;
        RECT 63.130 213.650 63.530 214.100 ;
        RECT 59.580 213.500 63.530 213.650 ;
        RECT 63.130 213.050 63.530 213.500 ;
        RECT 59.580 212.900 63.530 213.050 ;
        RECT 63.130 212.450 63.530 212.900 ;
        RECT 59.580 212.300 63.530 212.450 ;
        RECT 63.130 211.850 63.530 212.300 ;
        RECT 59.580 211.700 63.530 211.850 ;
        RECT 63.130 211.250 63.530 211.700 ;
        RECT 59.580 211.100 63.530 211.250 ;
        RECT 63.130 210.650 63.530 211.100 ;
        RECT 59.580 210.500 63.530 210.650 ;
        RECT 63.130 210.200 63.530 210.500 ;
        RECT 55.230 209.800 63.530 210.200 ;
        RECT 55.230 201.600 55.380 209.800 ;
        RECT 55.830 201.600 55.980 209.800 ;
        RECT 56.430 201.600 56.580 209.800 ;
        RECT 57.030 201.600 57.180 209.800 ;
        RECT 57.630 201.600 57.780 209.800 ;
        RECT 58.230 201.600 58.380 209.800 ;
        RECT 58.830 201.600 58.980 209.800 ;
        RECT 63.130 209.500 63.530 209.800 ;
        RECT 59.580 209.350 63.530 209.500 ;
        RECT 63.130 208.900 63.530 209.350 ;
        RECT 59.580 208.750 63.530 208.900 ;
        RECT 63.130 208.300 63.530 208.750 ;
        RECT 59.580 208.150 63.530 208.300 ;
        RECT 63.130 207.700 63.530 208.150 ;
        RECT 59.580 207.550 63.530 207.700 ;
        RECT 63.130 207.100 63.530 207.550 ;
        RECT 59.580 206.950 63.530 207.100 ;
        RECT 63.130 206.500 63.530 206.950 ;
        RECT 59.580 206.350 63.530 206.500 ;
        RECT 63.130 205.900 63.530 206.350 ;
        RECT 59.580 205.750 63.530 205.900 ;
        RECT 63.130 205.300 63.530 205.750 ;
        RECT 59.580 205.150 63.530 205.300 ;
        RECT 63.130 204.700 63.530 205.150 ;
        RECT 59.580 204.550 63.530 204.700 ;
        RECT 63.130 204.400 63.530 204.550 ;
        RECT 65.930 215.450 66.330 215.600 ;
        RECT 65.930 215.300 69.880 215.450 ;
        RECT 65.930 214.850 66.330 215.300 ;
        RECT 65.930 214.700 69.880 214.850 ;
        RECT 65.930 214.250 66.330 214.700 ;
        RECT 65.930 214.100 69.880 214.250 ;
        RECT 65.930 213.650 66.330 214.100 ;
        RECT 65.930 213.500 69.880 213.650 ;
        RECT 65.930 213.050 66.330 213.500 ;
        RECT 65.930 212.900 69.880 213.050 ;
        RECT 65.930 212.450 66.330 212.900 ;
        RECT 65.930 212.300 69.880 212.450 ;
        RECT 65.930 211.850 66.330 212.300 ;
        RECT 65.930 211.700 69.880 211.850 ;
        RECT 65.930 211.250 66.330 211.700 ;
        RECT 65.930 211.100 69.880 211.250 ;
        RECT 65.930 210.650 66.330 211.100 ;
        RECT 65.930 210.500 69.880 210.650 ;
        RECT 65.930 210.200 66.330 210.500 ;
        RECT 70.480 210.200 70.630 218.400 ;
        RECT 71.080 210.200 71.230 218.400 ;
        RECT 71.680 210.200 71.830 218.400 ;
        RECT 72.280 210.200 72.430 218.400 ;
        RECT 72.880 210.200 73.030 218.400 ;
        RECT 73.480 210.200 73.630 218.400 ;
        RECT 74.080 210.200 74.230 218.400 ;
        RECT 65.930 209.800 74.230 210.200 ;
        RECT 65.930 209.500 66.330 209.800 ;
        RECT 65.930 209.350 69.880 209.500 ;
        RECT 65.930 208.900 66.330 209.350 ;
        RECT 65.930 208.750 69.880 208.900 ;
        RECT 65.930 208.300 66.330 208.750 ;
        RECT 65.930 208.150 69.880 208.300 ;
        RECT 65.930 207.700 66.330 208.150 ;
        RECT 65.930 207.550 69.880 207.700 ;
        RECT 65.930 207.100 66.330 207.550 ;
        RECT 65.930 206.950 69.880 207.100 ;
        RECT 65.930 206.500 66.330 206.950 ;
        RECT 65.930 206.350 69.880 206.500 ;
        RECT 65.930 205.900 66.330 206.350 ;
        RECT 65.930 205.750 69.880 205.900 ;
        RECT 65.930 205.300 66.330 205.750 ;
        RECT 65.930 205.150 69.880 205.300 ;
        RECT 65.930 204.700 66.330 205.150 ;
        RECT 65.930 204.550 69.880 204.700 ;
        RECT 65.930 204.400 66.330 204.550 ;
        RECT 63.130 204.100 66.330 204.400 ;
        RECT 59.580 203.950 69.880 204.100 ;
        RECT 63.130 203.500 66.330 203.950 ;
        RECT 59.580 203.350 69.880 203.500 ;
        RECT 63.130 202.900 66.330 203.350 ;
        RECT 59.580 202.750 69.880 202.900 ;
        RECT 63.130 202.300 66.330 202.750 ;
        RECT 59.580 202.150 69.880 202.300 ;
        RECT 63.530 201.200 65.930 202.150 ;
        RECT 70.480 201.600 70.630 209.800 ;
        RECT 71.080 201.600 71.230 209.800 ;
        RECT 71.680 201.600 71.830 209.800 ;
        RECT 72.280 201.600 72.430 209.800 ;
        RECT 72.880 201.600 73.030 209.800 ;
        RECT 73.480 201.600 73.630 209.800 ;
        RECT 74.080 201.600 74.230 209.800 ;
        RECT 75.230 210.200 75.380 218.400 ;
        RECT 75.830 210.200 75.980 218.400 ;
        RECT 76.430 210.200 76.580 218.400 ;
        RECT 77.030 210.200 77.180 218.400 ;
        RECT 77.630 210.200 77.780 218.400 ;
        RECT 78.230 210.200 78.380 218.400 ;
        RECT 78.830 210.200 78.980 218.400 ;
        RECT 83.530 217.850 85.940 218.800 ;
        RECT 79.580 217.700 89.880 217.850 ;
        RECT 83.130 217.250 86.330 217.700 ;
        RECT 79.580 217.100 89.880 217.250 ;
        RECT 83.130 216.650 86.330 217.100 ;
        RECT 79.580 216.500 89.880 216.650 ;
        RECT 83.130 216.050 86.330 216.500 ;
        RECT 79.580 215.900 89.880 216.050 ;
        RECT 83.130 215.600 86.330 215.900 ;
        RECT 83.130 215.450 83.530 215.600 ;
        RECT 79.580 215.300 83.530 215.450 ;
        RECT 83.130 214.850 83.530 215.300 ;
        RECT 79.580 214.700 83.530 214.850 ;
        RECT 83.130 214.250 83.530 214.700 ;
        RECT 79.580 214.100 83.530 214.250 ;
        RECT 83.130 213.650 83.530 214.100 ;
        RECT 79.580 213.500 83.530 213.650 ;
        RECT 83.130 213.050 83.530 213.500 ;
        RECT 79.580 212.900 83.530 213.050 ;
        RECT 83.130 212.450 83.530 212.900 ;
        RECT 79.580 212.300 83.530 212.450 ;
        RECT 83.130 211.850 83.530 212.300 ;
        RECT 79.580 211.700 83.530 211.850 ;
        RECT 83.130 211.250 83.530 211.700 ;
        RECT 79.580 211.100 83.530 211.250 ;
        RECT 83.130 210.650 83.530 211.100 ;
        RECT 79.580 210.500 83.530 210.650 ;
        RECT 83.130 210.200 83.530 210.500 ;
        RECT 75.230 209.800 83.530 210.200 ;
        RECT 75.230 201.600 75.380 209.800 ;
        RECT 75.830 201.600 75.980 209.800 ;
        RECT 76.430 201.600 76.580 209.800 ;
        RECT 77.030 201.600 77.180 209.800 ;
        RECT 77.630 201.600 77.780 209.800 ;
        RECT 78.230 201.600 78.380 209.800 ;
        RECT 78.830 201.600 78.980 209.800 ;
        RECT 83.130 209.500 83.530 209.800 ;
        RECT 79.580 209.350 83.530 209.500 ;
        RECT 83.130 208.900 83.530 209.350 ;
        RECT 79.580 208.750 83.530 208.900 ;
        RECT 83.130 208.300 83.530 208.750 ;
        RECT 79.580 208.150 83.530 208.300 ;
        RECT 83.130 207.700 83.530 208.150 ;
        RECT 79.580 207.550 83.530 207.700 ;
        RECT 83.130 207.100 83.530 207.550 ;
        RECT 79.580 206.950 83.530 207.100 ;
        RECT 83.130 206.500 83.530 206.950 ;
        RECT 79.580 206.350 83.530 206.500 ;
        RECT 83.130 205.900 83.530 206.350 ;
        RECT 79.580 205.750 83.530 205.900 ;
        RECT 83.130 205.300 83.530 205.750 ;
        RECT 79.580 205.150 83.530 205.300 ;
        RECT 83.130 204.700 83.530 205.150 ;
        RECT 79.580 204.550 83.530 204.700 ;
        RECT 83.130 204.400 83.530 204.550 ;
        RECT 85.930 215.450 86.330 215.600 ;
        RECT 85.930 215.300 89.880 215.450 ;
        RECT 85.930 214.850 86.330 215.300 ;
        RECT 85.930 214.700 89.880 214.850 ;
        RECT 85.930 214.250 86.330 214.700 ;
        RECT 85.930 214.100 89.880 214.250 ;
        RECT 85.930 213.650 86.330 214.100 ;
        RECT 85.930 213.500 89.880 213.650 ;
        RECT 85.930 213.050 86.330 213.500 ;
        RECT 85.930 212.900 89.880 213.050 ;
        RECT 85.930 212.450 86.330 212.900 ;
        RECT 85.930 212.300 89.880 212.450 ;
        RECT 85.930 211.850 86.330 212.300 ;
        RECT 85.930 211.700 89.880 211.850 ;
        RECT 85.930 211.250 86.330 211.700 ;
        RECT 85.930 211.100 89.880 211.250 ;
        RECT 85.930 210.650 86.330 211.100 ;
        RECT 85.930 210.500 89.880 210.650 ;
        RECT 85.930 210.200 86.330 210.500 ;
        RECT 90.480 210.200 90.630 218.400 ;
        RECT 91.080 210.200 91.230 218.400 ;
        RECT 91.680 210.200 91.830 218.400 ;
        RECT 92.280 210.200 92.430 218.400 ;
        RECT 92.880 210.200 93.030 218.400 ;
        RECT 93.480 210.200 93.630 218.400 ;
        RECT 94.080 210.200 94.230 218.400 ;
        RECT 85.930 209.800 94.230 210.200 ;
        RECT 85.930 209.500 86.330 209.800 ;
        RECT 85.930 209.350 89.880 209.500 ;
        RECT 85.930 208.900 86.330 209.350 ;
        RECT 85.930 208.750 89.880 208.900 ;
        RECT 85.930 208.300 86.330 208.750 ;
        RECT 85.930 208.150 89.880 208.300 ;
        RECT 85.930 207.700 86.330 208.150 ;
        RECT 85.930 207.550 89.880 207.700 ;
        RECT 85.930 207.100 86.330 207.550 ;
        RECT 85.930 206.950 89.880 207.100 ;
        RECT 85.930 206.500 86.330 206.950 ;
        RECT 85.930 206.350 89.880 206.500 ;
        RECT 85.930 205.900 86.330 206.350 ;
        RECT 85.930 205.750 89.880 205.900 ;
        RECT 85.930 205.300 86.330 205.750 ;
        RECT 85.930 205.150 89.880 205.300 ;
        RECT 85.930 204.700 86.330 205.150 ;
        RECT 85.930 204.550 89.880 204.700 ;
        RECT 85.930 204.400 86.330 204.550 ;
        RECT 83.130 204.100 86.330 204.400 ;
        RECT 79.580 203.950 89.880 204.100 ;
        RECT 83.130 203.500 86.330 203.950 ;
        RECT 79.580 203.350 89.880 203.500 ;
        RECT 83.130 202.900 86.330 203.350 ;
        RECT 79.580 202.750 89.880 202.900 ;
        RECT 83.130 202.300 86.330 202.750 ;
        RECT 79.580 202.150 89.880 202.300 ;
        RECT 83.530 201.200 85.930 202.150 ;
        RECT 90.480 201.600 90.630 209.800 ;
        RECT 91.080 201.600 91.230 209.800 ;
        RECT 91.680 201.600 91.830 209.800 ;
        RECT 92.280 201.600 92.430 209.800 ;
        RECT 92.880 201.600 93.030 209.800 ;
        RECT 93.480 201.600 93.630 209.800 ;
        RECT 94.080 201.600 94.230 209.800 ;
        RECT 95.230 210.200 95.380 218.400 ;
        RECT 95.830 210.200 95.980 218.400 ;
        RECT 96.430 210.200 96.580 218.400 ;
        RECT 97.030 210.200 97.180 218.400 ;
        RECT 97.630 210.200 97.780 218.400 ;
        RECT 98.230 210.200 98.380 218.400 ;
        RECT 98.830 210.200 98.980 218.400 ;
        RECT 103.530 217.850 105.940 218.800 ;
        RECT 99.580 217.700 109.880 217.850 ;
        RECT 103.130 217.250 106.330 217.700 ;
        RECT 99.580 217.100 109.880 217.250 ;
        RECT 103.130 216.650 106.330 217.100 ;
        RECT 99.580 216.500 109.880 216.650 ;
        RECT 103.130 216.050 106.330 216.500 ;
        RECT 99.580 215.900 109.880 216.050 ;
        RECT 103.130 215.600 106.330 215.900 ;
        RECT 103.130 215.450 103.530 215.600 ;
        RECT 99.580 215.300 103.530 215.450 ;
        RECT 103.130 214.850 103.530 215.300 ;
        RECT 99.580 214.700 103.530 214.850 ;
        RECT 103.130 214.250 103.530 214.700 ;
        RECT 99.580 214.100 103.530 214.250 ;
        RECT 103.130 213.650 103.530 214.100 ;
        RECT 99.580 213.500 103.530 213.650 ;
        RECT 103.130 213.050 103.530 213.500 ;
        RECT 99.580 212.900 103.530 213.050 ;
        RECT 103.130 212.450 103.530 212.900 ;
        RECT 99.580 212.300 103.530 212.450 ;
        RECT 103.130 211.850 103.530 212.300 ;
        RECT 99.580 211.700 103.530 211.850 ;
        RECT 103.130 211.250 103.530 211.700 ;
        RECT 99.580 211.100 103.530 211.250 ;
        RECT 103.130 210.650 103.530 211.100 ;
        RECT 99.580 210.500 103.530 210.650 ;
        RECT 103.130 210.200 103.530 210.500 ;
        RECT 95.230 209.800 103.530 210.200 ;
        RECT 95.230 201.600 95.380 209.800 ;
        RECT 95.830 201.600 95.980 209.800 ;
        RECT 96.430 201.600 96.580 209.800 ;
        RECT 97.030 201.600 97.180 209.800 ;
        RECT 97.630 201.600 97.780 209.800 ;
        RECT 98.230 201.600 98.380 209.800 ;
        RECT 98.830 201.600 98.980 209.800 ;
        RECT 103.130 209.500 103.530 209.800 ;
        RECT 99.580 209.350 103.530 209.500 ;
        RECT 103.130 208.900 103.530 209.350 ;
        RECT 99.580 208.750 103.530 208.900 ;
        RECT 103.130 208.300 103.530 208.750 ;
        RECT 99.580 208.150 103.530 208.300 ;
        RECT 103.130 207.700 103.530 208.150 ;
        RECT 99.580 207.550 103.530 207.700 ;
        RECT 103.130 207.100 103.530 207.550 ;
        RECT 99.580 206.950 103.530 207.100 ;
        RECT 103.130 206.500 103.530 206.950 ;
        RECT 99.580 206.350 103.530 206.500 ;
        RECT 103.130 205.900 103.530 206.350 ;
        RECT 99.580 205.750 103.530 205.900 ;
        RECT 103.130 205.300 103.530 205.750 ;
        RECT 99.580 205.150 103.530 205.300 ;
        RECT 103.130 204.700 103.530 205.150 ;
        RECT 99.580 204.550 103.530 204.700 ;
        RECT 103.130 204.400 103.530 204.550 ;
        RECT 105.930 215.450 106.330 215.600 ;
        RECT 105.930 215.300 109.880 215.450 ;
        RECT 105.930 214.850 106.330 215.300 ;
        RECT 105.930 214.700 109.880 214.850 ;
        RECT 105.930 214.250 106.330 214.700 ;
        RECT 105.930 214.100 109.880 214.250 ;
        RECT 105.930 213.650 106.330 214.100 ;
        RECT 105.930 213.500 109.880 213.650 ;
        RECT 105.930 213.050 106.330 213.500 ;
        RECT 105.930 212.900 109.880 213.050 ;
        RECT 105.930 212.450 106.330 212.900 ;
        RECT 105.930 212.300 109.880 212.450 ;
        RECT 105.930 211.850 106.330 212.300 ;
        RECT 105.930 211.700 109.880 211.850 ;
        RECT 105.930 211.250 106.330 211.700 ;
        RECT 105.930 211.100 109.880 211.250 ;
        RECT 105.930 210.650 106.330 211.100 ;
        RECT 105.930 210.500 109.880 210.650 ;
        RECT 105.930 210.200 106.330 210.500 ;
        RECT 110.480 210.200 110.630 218.400 ;
        RECT 111.080 210.200 111.230 218.400 ;
        RECT 111.680 210.200 111.830 218.400 ;
        RECT 112.280 210.200 112.430 218.400 ;
        RECT 112.880 210.200 113.030 218.400 ;
        RECT 113.480 210.200 113.630 218.400 ;
        RECT 114.080 210.200 114.230 218.400 ;
        RECT 105.930 209.800 114.230 210.200 ;
        RECT 105.930 209.500 106.330 209.800 ;
        RECT 105.930 209.350 109.880 209.500 ;
        RECT 105.930 208.900 106.330 209.350 ;
        RECT 105.930 208.750 109.880 208.900 ;
        RECT 105.930 208.300 106.330 208.750 ;
        RECT 105.930 208.150 109.880 208.300 ;
        RECT 105.930 207.700 106.330 208.150 ;
        RECT 105.930 207.550 109.880 207.700 ;
        RECT 105.930 207.100 106.330 207.550 ;
        RECT 105.930 206.950 109.880 207.100 ;
        RECT 105.930 206.500 106.330 206.950 ;
        RECT 105.930 206.350 109.880 206.500 ;
        RECT 105.930 205.900 106.330 206.350 ;
        RECT 105.930 205.750 109.880 205.900 ;
        RECT 105.930 205.300 106.330 205.750 ;
        RECT 105.930 205.150 109.880 205.300 ;
        RECT 105.930 204.700 106.330 205.150 ;
        RECT 105.930 204.550 109.880 204.700 ;
        RECT 105.930 204.400 106.330 204.550 ;
        RECT 103.130 204.100 106.330 204.400 ;
        RECT 99.580 203.950 109.880 204.100 ;
        RECT 103.130 203.500 106.330 203.950 ;
        RECT 99.580 203.350 109.880 203.500 ;
        RECT 103.130 202.900 106.330 203.350 ;
        RECT 99.580 202.750 109.880 202.900 ;
        RECT 103.130 202.300 106.330 202.750 ;
        RECT 99.580 202.150 109.880 202.300 ;
        RECT 103.530 201.200 105.930 202.150 ;
        RECT 110.480 201.600 110.630 209.800 ;
        RECT 111.080 201.600 111.230 209.800 ;
        RECT 111.680 201.600 111.830 209.800 ;
        RECT 112.280 201.600 112.430 209.800 ;
        RECT 112.880 201.600 113.030 209.800 ;
        RECT 113.480 201.600 113.630 209.800 ;
        RECT 114.080 201.600 114.230 209.800 ;
        RECT 115.230 210.200 115.380 218.400 ;
        RECT 115.830 210.200 115.980 218.400 ;
        RECT 116.430 210.200 116.580 218.400 ;
        RECT 117.030 210.200 117.180 218.400 ;
        RECT 117.630 210.200 117.780 218.400 ;
        RECT 118.230 210.200 118.380 218.400 ;
        RECT 118.830 210.200 118.980 218.400 ;
        RECT 123.530 217.850 124.730 218.800 ;
        RECT 119.580 217.700 124.730 217.850 ;
        RECT 123.130 217.250 124.730 217.700 ;
        RECT 119.580 217.100 124.730 217.250 ;
        RECT 123.130 216.650 124.730 217.100 ;
        RECT 119.580 216.500 124.730 216.650 ;
        RECT 123.130 216.050 124.730 216.500 ;
        RECT 125.140 216.490 127.140 217.765 ;
        RECT 119.580 215.900 124.730 216.050 ;
        RECT 123.130 215.600 124.730 215.900 ;
        RECT 123.130 215.450 123.530 215.600 ;
        RECT 119.580 215.300 123.530 215.450 ;
        RECT 123.130 214.850 123.530 215.300 ;
        RECT 119.580 214.700 123.530 214.850 ;
        RECT 123.130 214.250 123.530 214.700 ;
        RECT 119.580 214.100 123.530 214.250 ;
        RECT 123.130 213.650 123.530 214.100 ;
        RECT 119.580 213.500 123.530 213.650 ;
        RECT 123.130 213.050 123.530 213.500 ;
        RECT 119.580 212.900 123.530 213.050 ;
        RECT 123.130 212.450 123.530 212.900 ;
        RECT 119.580 212.300 123.530 212.450 ;
        RECT 123.130 211.850 123.530 212.300 ;
        RECT 119.580 211.700 123.530 211.850 ;
        RECT 123.130 211.250 123.530 211.700 ;
        RECT 119.580 211.100 123.530 211.250 ;
        RECT 123.130 210.650 123.530 211.100 ;
        RECT 119.580 210.500 123.530 210.650 ;
        RECT 123.130 210.200 123.530 210.500 ;
        RECT 115.230 209.800 123.530 210.200 ;
        RECT 115.230 201.600 115.380 209.800 ;
        RECT 115.830 201.600 115.980 209.800 ;
        RECT 116.430 201.600 116.580 209.800 ;
        RECT 117.030 201.600 117.180 209.800 ;
        RECT 117.630 201.600 117.780 209.800 ;
        RECT 118.230 201.600 118.380 209.800 ;
        RECT 118.830 201.600 118.980 209.800 ;
        RECT 123.130 209.500 123.530 209.800 ;
        RECT 119.580 209.350 123.530 209.500 ;
        RECT 123.130 208.900 123.530 209.350 ;
        RECT 119.580 208.750 123.530 208.900 ;
        RECT 123.130 208.300 123.530 208.750 ;
        RECT 119.580 208.150 123.530 208.300 ;
        RECT 123.130 207.700 123.530 208.150 ;
        RECT 119.580 207.550 123.530 207.700 ;
        RECT 123.130 207.100 123.530 207.550 ;
        RECT 119.580 206.950 123.530 207.100 ;
        RECT 123.130 206.500 123.530 206.950 ;
        RECT 119.580 206.350 123.530 206.500 ;
        RECT 123.130 205.900 123.530 206.350 ;
        RECT 119.580 205.750 123.530 205.900 ;
        RECT 123.130 205.300 123.530 205.750 ;
        RECT 119.580 205.150 123.530 205.300 ;
        RECT 123.130 204.700 123.530 205.150 ;
        RECT 119.580 204.550 123.530 204.700 ;
        RECT 123.130 204.400 123.530 204.550 ;
        RECT 123.130 204.100 124.730 204.400 ;
        RECT 119.580 203.950 124.730 204.100 ;
        RECT 123.130 203.500 124.730 203.950 ;
        RECT 119.580 203.350 124.730 203.500 ;
        RECT 123.130 202.900 124.730 203.350 ;
        RECT 119.580 202.750 124.730 202.900 ;
        RECT 123.130 202.300 124.730 202.750 ;
        RECT 119.580 202.150 124.730 202.300 ;
        RECT 123.530 201.200 124.730 202.150 ;
        RECT 4.730 200.000 9.130 201.200 ;
        RECT 20.330 200.000 29.130 201.200 ;
        RECT 40.330 200.000 49.130 201.200 ;
        RECT 60.330 200.000 69.130 201.200 ;
        RECT 80.330 200.000 89.130 201.200 ;
        RECT 100.330 200.000 109.130 201.200 ;
        RECT 120.330 200.000 124.730 201.200 ;
        RECT 125.140 200.910 127.140 202.185 ;
        RECT 2.315 175.215 4.025 175.695 ;
        RECT 42.635 175.460 47.035 176.660 ;
        RECT 58.235 175.460 67.035 176.660 ;
        RECT 78.235 175.460 87.035 176.660 ;
        RECT 98.235 175.460 107.035 176.660 ;
        RECT 118.235 175.460 122.635 176.660 ;
        RECT 42.635 174.510 43.845 175.460 ;
        RECT 42.635 174.360 47.785 174.510 ;
        RECT 42.635 173.910 44.235 174.360 ;
        RECT 42.635 173.760 47.785 173.910 ;
        RECT 42.635 173.310 44.235 173.760 ;
        RECT 42.635 173.160 47.785 173.310 ;
        RECT 42.635 172.710 44.235 173.160 ;
        RECT 42.635 172.560 47.785 172.710 ;
        RECT 42.635 172.260 44.235 172.560 ;
        RECT 43.835 172.110 44.235 172.260 ;
        RECT 43.835 171.960 47.785 172.110 ;
        RECT 43.835 171.510 44.235 171.960 ;
        RECT 43.835 171.360 47.785 171.510 ;
        RECT 43.835 170.910 44.235 171.360 ;
        RECT 43.835 170.760 47.785 170.910 ;
        RECT 43.835 170.310 44.235 170.760 ;
        RECT 2.315 169.775 4.025 170.255 ;
        RECT 43.835 170.160 47.785 170.310 ;
        RECT 43.835 169.710 44.235 170.160 ;
        RECT 43.835 169.560 47.785 169.710 ;
        RECT 43.835 169.110 44.235 169.560 ;
        RECT 43.835 168.960 47.785 169.110 ;
        RECT 43.835 168.510 44.235 168.960 ;
        RECT 43.835 168.360 47.785 168.510 ;
        RECT 43.835 167.910 44.235 168.360 ;
        RECT 43.835 167.760 47.785 167.910 ;
        RECT 43.835 167.310 44.235 167.760 ;
        RECT 43.835 167.160 47.785 167.310 ;
        RECT 43.835 166.860 44.235 167.160 ;
        RECT 48.385 166.860 48.535 175.060 ;
        RECT 48.985 166.860 49.135 175.060 ;
        RECT 49.585 166.860 49.735 175.060 ;
        RECT 50.185 166.860 50.335 175.060 ;
        RECT 50.785 166.860 50.935 175.060 ;
        RECT 51.385 166.860 51.535 175.060 ;
        RECT 51.985 166.860 52.135 175.060 ;
        RECT 43.835 166.460 52.135 166.860 ;
        RECT 43.835 166.160 44.235 166.460 ;
        RECT 43.835 166.010 47.785 166.160 ;
        RECT 43.835 165.560 44.235 166.010 ;
        RECT 43.835 165.410 47.785 165.560 ;
        RECT 43.835 164.960 44.235 165.410 ;
        RECT 2.315 164.335 4.025 164.815 ;
        RECT 43.835 164.810 47.785 164.960 ;
        RECT 43.835 164.360 44.235 164.810 ;
        RECT 43.835 164.210 47.785 164.360 ;
        RECT 43.835 163.760 44.235 164.210 ;
        RECT 43.835 163.610 47.785 163.760 ;
        RECT 43.835 163.160 44.235 163.610 ;
        RECT 43.835 163.010 47.785 163.160 ;
        RECT 43.835 162.560 44.235 163.010 ;
        RECT 43.835 162.410 47.785 162.560 ;
        RECT 43.835 161.960 44.235 162.410 ;
        RECT 43.835 161.810 47.785 161.960 ;
        RECT 43.835 161.360 44.235 161.810 ;
        RECT 43.835 161.210 47.785 161.360 ;
        RECT 43.835 161.060 44.235 161.210 ;
        RECT 42.635 160.760 44.235 161.060 ;
        RECT 42.635 160.610 47.785 160.760 ;
        RECT 42.635 160.160 44.235 160.610 ;
        RECT 42.635 160.010 47.785 160.160 ;
        RECT 42.635 159.560 44.235 160.010 ;
        RECT 42.635 159.410 47.785 159.560 ;
        RECT 42.635 158.960 44.235 159.410 ;
        RECT 42.635 158.810 47.785 158.960 ;
        RECT 42.635 157.860 43.835 158.810 ;
        RECT 48.385 158.260 48.535 166.460 ;
        RECT 48.985 158.260 49.135 166.460 ;
        RECT 49.585 158.260 49.735 166.460 ;
        RECT 50.185 158.260 50.335 166.460 ;
        RECT 50.785 158.260 50.935 166.460 ;
        RECT 51.385 158.260 51.535 166.460 ;
        RECT 51.985 158.260 52.135 166.460 ;
        RECT 53.135 166.860 53.285 175.060 ;
        RECT 53.735 166.860 53.885 175.060 ;
        RECT 54.335 166.860 54.485 175.060 ;
        RECT 54.935 166.860 55.085 175.060 ;
        RECT 55.535 166.860 55.685 175.060 ;
        RECT 56.135 166.860 56.285 175.060 ;
        RECT 56.735 166.860 56.885 175.060 ;
        RECT 61.435 174.510 63.845 175.460 ;
        RECT 57.485 174.360 67.785 174.510 ;
        RECT 61.035 173.910 64.235 174.360 ;
        RECT 57.485 173.760 67.785 173.910 ;
        RECT 61.035 173.310 64.235 173.760 ;
        RECT 57.485 173.160 67.785 173.310 ;
        RECT 61.035 172.710 64.235 173.160 ;
        RECT 57.485 172.560 67.785 172.710 ;
        RECT 61.035 172.260 64.235 172.560 ;
        RECT 61.035 172.110 61.435 172.260 ;
        RECT 57.485 171.960 61.435 172.110 ;
        RECT 61.035 171.510 61.435 171.960 ;
        RECT 57.485 171.360 61.435 171.510 ;
        RECT 61.035 170.910 61.435 171.360 ;
        RECT 57.485 170.760 61.435 170.910 ;
        RECT 61.035 170.310 61.435 170.760 ;
        RECT 57.485 170.160 61.435 170.310 ;
        RECT 61.035 169.710 61.435 170.160 ;
        RECT 57.485 169.560 61.435 169.710 ;
        RECT 61.035 169.110 61.435 169.560 ;
        RECT 57.485 168.960 61.435 169.110 ;
        RECT 61.035 168.510 61.435 168.960 ;
        RECT 57.485 168.360 61.435 168.510 ;
        RECT 61.035 167.910 61.435 168.360 ;
        RECT 57.485 167.760 61.435 167.910 ;
        RECT 61.035 167.310 61.435 167.760 ;
        RECT 57.485 167.160 61.435 167.310 ;
        RECT 61.035 166.860 61.435 167.160 ;
        RECT 53.135 166.460 61.435 166.860 ;
        RECT 53.135 158.260 53.285 166.460 ;
        RECT 53.735 158.260 53.885 166.460 ;
        RECT 54.335 158.260 54.485 166.460 ;
        RECT 54.935 158.260 55.085 166.460 ;
        RECT 55.535 158.260 55.685 166.460 ;
        RECT 56.135 158.260 56.285 166.460 ;
        RECT 56.735 158.260 56.885 166.460 ;
        RECT 61.035 166.160 61.435 166.460 ;
        RECT 57.485 166.010 61.435 166.160 ;
        RECT 61.035 165.560 61.435 166.010 ;
        RECT 57.485 165.410 61.435 165.560 ;
        RECT 61.035 164.960 61.435 165.410 ;
        RECT 57.485 164.810 61.435 164.960 ;
        RECT 61.035 164.360 61.435 164.810 ;
        RECT 57.485 164.210 61.435 164.360 ;
        RECT 61.035 163.760 61.435 164.210 ;
        RECT 57.485 163.610 61.435 163.760 ;
        RECT 61.035 163.160 61.435 163.610 ;
        RECT 57.485 163.010 61.435 163.160 ;
        RECT 61.035 162.560 61.435 163.010 ;
        RECT 57.485 162.410 61.435 162.560 ;
        RECT 61.035 161.960 61.435 162.410 ;
        RECT 57.485 161.810 61.435 161.960 ;
        RECT 61.035 161.360 61.435 161.810 ;
        RECT 57.485 161.210 61.435 161.360 ;
        RECT 61.035 161.060 61.435 161.210 ;
        RECT 63.835 172.110 64.235 172.260 ;
        RECT 63.835 171.960 67.785 172.110 ;
        RECT 63.835 171.510 64.235 171.960 ;
        RECT 63.835 171.360 67.785 171.510 ;
        RECT 63.835 170.910 64.235 171.360 ;
        RECT 63.835 170.760 67.785 170.910 ;
        RECT 63.835 170.310 64.235 170.760 ;
        RECT 63.835 170.160 67.785 170.310 ;
        RECT 63.835 169.710 64.235 170.160 ;
        RECT 63.835 169.560 67.785 169.710 ;
        RECT 63.835 169.110 64.235 169.560 ;
        RECT 63.835 168.960 67.785 169.110 ;
        RECT 63.835 168.510 64.235 168.960 ;
        RECT 63.835 168.360 67.785 168.510 ;
        RECT 63.835 167.910 64.235 168.360 ;
        RECT 63.835 167.760 67.785 167.910 ;
        RECT 63.835 167.310 64.235 167.760 ;
        RECT 63.835 167.160 67.785 167.310 ;
        RECT 63.835 166.860 64.235 167.160 ;
        RECT 68.385 166.860 68.535 175.060 ;
        RECT 68.985 166.860 69.135 175.060 ;
        RECT 69.585 166.860 69.735 175.060 ;
        RECT 70.185 166.860 70.335 175.060 ;
        RECT 70.785 166.860 70.935 175.060 ;
        RECT 71.385 166.860 71.535 175.060 ;
        RECT 71.985 166.860 72.135 175.060 ;
        RECT 63.835 166.460 72.135 166.860 ;
        RECT 63.835 166.160 64.235 166.460 ;
        RECT 63.835 166.010 67.785 166.160 ;
        RECT 63.835 165.560 64.235 166.010 ;
        RECT 63.835 165.410 67.785 165.560 ;
        RECT 63.835 164.960 64.235 165.410 ;
        RECT 63.835 164.810 67.785 164.960 ;
        RECT 63.835 164.360 64.235 164.810 ;
        RECT 63.835 164.210 67.785 164.360 ;
        RECT 63.835 163.760 64.235 164.210 ;
        RECT 63.835 163.610 67.785 163.760 ;
        RECT 63.835 163.160 64.235 163.610 ;
        RECT 63.835 163.010 67.785 163.160 ;
        RECT 63.835 162.560 64.235 163.010 ;
        RECT 63.835 162.410 67.785 162.560 ;
        RECT 63.835 161.960 64.235 162.410 ;
        RECT 63.835 161.810 67.785 161.960 ;
        RECT 63.835 161.360 64.235 161.810 ;
        RECT 63.835 161.210 67.785 161.360 ;
        RECT 63.835 161.060 64.235 161.210 ;
        RECT 61.035 160.760 64.235 161.060 ;
        RECT 57.485 160.610 67.785 160.760 ;
        RECT 61.035 160.160 64.235 160.610 ;
        RECT 57.485 160.010 67.785 160.160 ;
        RECT 61.035 159.560 64.235 160.010 ;
        RECT 57.485 159.410 67.785 159.560 ;
        RECT 61.035 158.960 64.235 159.410 ;
        RECT 57.485 158.810 67.785 158.960 ;
        RECT 61.435 157.860 63.835 158.810 ;
        RECT 68.385 158.260 68.535 166.460 ;
        RECT 68.985 158.260 69.135 166.460 ;
        RECT 69.585 158.260 69.735 166.460 ;
        RECT 70.185 158.260 70.335 166.460 ;
        RECT 70.785 158.260 70.935 166.460 ;
        RECT 71.385 158.260 71.535 166.460 ;
        RECT 71.985 158.260 72.135 166.460 ;
        RECT 73.135 166.860 73.285 175.060 ;
        RECT 73.735 166.860 73.885 175.060 ;
        RECT 74.335 166.860 74.485 175.060 ;
        RECT 74.935 166.860 75.085 175.060 ;
        RECT 75.535 166.860 75.685 175.060 ;
        RECT 76.135 166.860 76.285 175.060 ;
        RECT 76.735 166.860 76.885 175.060 ;
        RECT 81.435 174.510 83.845 175.460 ;
        RECT 77.485 174.360 87.785 174.510 ;
        RECT 81.035 173.910 84.235 174.360 ;
        RECT 77.485 173.760 87.785 173.910 ;
        RECT 81.035 173.310 84.235 173.760 ;
        RECT 77.485 173.160 87.785 173.310 ;
        RECT 81.035 172.710 84.235 173.160 ;
        RECT 77.485 172.560 87.785 172.710 ;
        RECT 81.035 172.260 84.235 172.560 ;
        RECT 81.035 172.110 81.435 172.260 ;
        RECT 77.485 171.960 81.435 172.110 ;
        RECT 81.035 171.510 81.435 171.960 ;
        RECT 77.485 171.360 81.435 171.510 ;
        RECT 81.035 170.910 81.435 171.360 ;
        RECT 77.485 170.760 81.435 170.910 ;
        RECT 81.035 170.310 81.435 170.760 ;
        RECT 77.485 170.160 81.435 170.310 ;
        RECT 81.035 169.710 81.435 170.160 ;
        RECT 77.485 169.560 81.435 169.710 ;
        RECT 81.035 169.110 81.435 169.560 ;
        RECT 77.485 168.960 81.435 169.110 ;
        RECT 81.035 168.510 81.435 168.960 ;
        RECT 77.485 168.360 81.435 168.510 ;
        RECT 81.035 167.910 81.435 168.360 ;
        RECT 77.485 167.760 81.435 167.910 ;
        RECT 81.035 167.310 81.435 167.760 ;
        RECT 77.485 167.160 81.435 167.310 ;
        RECT 81.035 166.860 81.435 167.160 ;
        RECT 73.135 166.460 81.435 166.860 ;
        RECT 73.135 158.260 73.285 166.460 ;
        RECT 73.735 158.260 73.885 166.460 ;
        RECT 74.335 158.260 74.485 166.460 ;
        RECT 74.935 158.260 75.085 166.460 ;
        RECT 75.535 158.260 75.685 166.460 ;
        RECT 76.135 158.260 76.285 166.460 ;
        RECT 76.735 158.260 76.885 166.460 ;
        RECT 81.035 166.160 81.435 166.460 ;
        RECT 77.485 166.010 81.435 166.160 ;
        RECT 81.035 165.560 81.435 166.010 ;
        RECT 77.485 165.410 81.435 165.560 ;
        RECT 81.035 164.960 81.435 165.410 ;
        RECT 77.485 164.810 81.435 164.960 ;
        RECT 81.035 164.360 81.435 164.810 ;
        RECT 77.485 164.210 81.435 164.360 ;
        RECT 81.035 163.760 81.435 164.210 ;
        RECT 77.485 163.610 81.435 163.760 ;
        RECT 81.035 163.160 81.435 163.610 ;
        RECT 77.485 163.010 81.435 163.160 ;
        RECT 81.035 162.560 81.435 163.010 ;
        RECT 77.485 162.410 81.435 162.560 ;
        RECT 81.035 161.960 81.435 162.410 ;
        RECT 77.485 161.810 81.435 161.960 ;
        RECT 81.035 161.360 81.435 161.810 ;
        RECT 77.485 161.210 81.435 161.360 ;
        RECT 81.035 161.060 81.435 161.210 ;
        RECT 83.835 172.110 84.235 172.260 ;
        RECT 83.835 171.960 87.785 172.110 ;
        RECT 83.835 171.510 84.235 171.960 ;
        RECT 83.835 171.360 87.785 171.510 ;
        RECT 83.835 170.910 84.235 171.360 ;
        RECT 83.835 170.760 87.785 170.910 ;
        RECT 83.835 170.310 84.235 170.760 ;
        RECT 83.835 170.160 87.785 170.310 ;
        RECT 83.835 169.710 84.235 170.160 ;
        RECT 83.835 169.560 87.785 169.710 ;
        RECT 83.835 169.110 84.235 169.560 ;
        RECT 83.835 168.960 87.785 169.110 ;
        RECT 83.835 168.510 84.235 168.960 ;
        RECT 83.835 168.360 87.785 168.510 ;
        RECT 83.835 167.910 84.235 168.360 ;
        RECT 83.835 167.760 87.785 167.910 ;
        RECT 83.835 167.310 84.235 167.760 ;
        RECT 83.835 167.160 87.785 167.310 ;
        RECT 83.835 166.860 84.235 167.160 ;
        RECT 88.385 166.860 88.535 175.060 ;
        RECT 88.985 166.860 89.135 175.060 ;
        RECT 89.585 166.860 89.735 175.060 ;
        RECT 90.185 166.860 90.335 175.060 ;
        RECT 90.785 166.860 90.935 175.060 ;
        RECT 91.385 166.860 91.535 175.060 ;
        RECT 91.985 166.860 92.135 175.060 ;
        RECT 83.835 166.460 92.135 166.860 ;
        RECT 83.835 166.160 84.235 166.460 ;
        RECT 83.835 166.010 87.785 166.160 ;
        RECT 83.835 165.560 84.235 166.010 ;
        RECT 83.835 165.410 87.785 165.560 ;
        RECT 83.835 164.960 84.235 165.410 ;
        RECT 83.835 164.810 87.785 164.960 ;
        RECT 83.835 164.360 84.235 164.810 ;
        RECT 83.835 164.210 87.785 164.360 ;
        RECT 83.835 163.760 84.235 164.210 ;
        RECT 83.835 163.610 87.785 163.760 ;
        RECT 83.835 163.160 84.235 163.610 ;
        RECT 83.835 163.010 87.785 163.160 ;
        RECT 83.835 162.560 84.235 163.010 ;
        RECT 83.835 162.410 87.785 162.560 ;
        RECT 83.835 161.960 84.235 162.410 ;
        RECT 83.835 161.810 87.785 161.960 ;
        RECT 83.835 161.360 84.235 161.810 ;
        RECT 83.835 161.210 87.785 161.360 ;
        RECT 83.835 161.060 84.235 161.210 ;
        RECT 81.035 160.760 84.235 161.060 ;
        RECT 77.485 160.610 87.785 160.760 ;
        RECT 81.035 160.160 84.235 160.610 ;
        RECT 77.485 160.010 87.785 160.160 ;
        RECT 81.035 159.560 84.235 160.010 ;
        RECT 77.485 159.410 87.785 159.560 ;
        RECT 81.035 158.960 84.235 159.410 ;
        RECT 77.485 158.810 87.785 158.960 ;
        RECT 81.435 157.860 83.835 158.810 ;
        RECT 88.385 158.260 88.535 166.460 ;
        RECT 88.985 158.260 89.135 166.460 ;
        RECT 89.585 158.260 89.735 166.460 ;
        RECT 90.185 158.260 90.335 166.460 ;
        RECT 90.785 158.260 90.935 166.460 ;
        RECT 91.385 158.260 91.535 166.460 ;
        RECT 91.985 158.260 92.135 166.460 ;
        RECT 93.135 166.860 93.285 175.060 ;
        RECT 93.735 166.860 93.885 175.060 ;
        RECT 94.335 166.860 94.485 175.060 ;
        RECT 94.935 166.860 95.085 175.060 ;
        RECT 95.535 166.860 95.685 175.060 ;
        RECT 96.135 166.860 96.285 175.060 ;
        RECT 96.735 166.860 96.885 175.060 ;
        RECT 101.435 174.510 103.845 175.460 ;
        RECT 97.485 174.360 107.785 174.510 ;
        RECT 101.035 173.910 104.235 174.360 ;
        RECT 97.485 173.760 107.785 173.910 ;
        RECT 101.035 173.310 104.235 173.760 ;
        RECT 97.485 173.160 107.785 173.310 ;
        RECT 101.035 172.710 104.235 173.160 ;
        RECT 97.485 172.560 107.785 172.710 ;
        RECT 101.035 172.260 104.235 172.560 ;
        RECT 101.035 172.110 101.435 172.260 ;
        RECT 97.485 171.960 101.435 172.110 ;
        RECT 101.035 171.510 101.435 171.960 ;
        RECT 97.485 171.360 101.435 171.510 ;
        RECT 101.035 170.910 101.435 171.360 ;
        RECT 97.485 170.760 101.435 170.910 ;
        RECT 101.035 170.310 101.435 170.760 ;
        RECT 97.485 170.160 101.435 170.310 ;
        RECT 101.035 169.710 101.435 170.160 ;
        RECT 97.485 169.560 101.435 169.710 ;
        RECT 101.035 169.110 101.435 169.560 ;
        RECT 97.485 168.960 101.435 169.110 ;
        RECT 101.035 168.510 101.435 168.960 ;
        RECT 97.485 168.360 101.435 168.510 ;
        RECT 101.035 167.910 101.435 168.360 ;
        RECT 97.485 167.760 101.435 167.910 ;
        RECT 101.035 167.310 101.435 167.760 ;
        RECT 97.485 167.160 101.435 167.310 ;
        RECT 101.035 166.860 101.435 167.160 ;
        RECT 93.135 166.460 101.435 166.860 ;
        RECT 93.135 158.260 93.285 166.460 ;
        RECT 93.735 158.260 93.885 166.460 ;
        RECT 94.335 158.260 94.485 166.460 ;
        RECT 94.935 158.260 95.085 166.460 ;
        RECT 95.535 158.260 95.685 166.460 ;
        RECT 96.135 158.260 96.285 166.460 ;
        RECT 96.735 158.260 96.885 166.460 ;
        RECT 101.035 166.160 101.435 166.460 ;
        RECT 97.485 166.010 101.435 166.160 ;
        RECT 101.035 165.560 101.435 166.010 ;
        RECT 97.485 165.410 101.435 165.560 ;
        RECT 101.035 164.960 101.435 165.410 ;
        RECT 97.485 164.810 101.435 164.960 ;
        RECT 101.035 164.360 101.435 164.810 ;
        RECT 97.485 164.210 101.435 164.360 ;
        RECT 101.035 163.760 101.435 164.210 ;
        RECT 97.485 163.610 101.435 163.760 ;
        RECT 101.035 163.160 101.435 163.610 ;
        RECT 97.485 163.010 101.435 163.160 ;
        RECT 101.035 162.560 101.435 163.010 ;
        RECT 97.485 162.410 101.435 162.560 ;
        RECT 101.035 161.960 101.435 162.410 ;
        RECT 97.485 161.810 101.435 161.960 ;
        RECT 101.035 161.360 101.435 161.810 ;
        RECT 97.485 161.210 101.435 161.360 ;
        RECT 101.035 161.060 101.435 161.210 ;
        RECT 103.835 172.110 104.235 172.260 ;
        RECT 103.835 171.960 107.785 172.110 ;
        RECT 103.835 171.510 104.235 171.960 ;
        RECT 103.835 171.360 107.785 171.510 ;
        RECT 103.835 170.910 104.235 171.360 ;
        RECT 103.835 170.760 107.785 170.910 ;
        RECT 103.835 170.310 104.235 170.760 ;
        RECT 103.835 170.160 107.785 170.310 ;
        RECT 103.835 169.710 104.235 170.160 ;
        RECT 103.835 169.560 107.785 169.710 ;
        RECT 103.835 169.110 104.235 169.560 ;
        RECT 103.835 168.960 107.785 169.110 ;
        RECT 103.835 168.510 104.235 168.960 ;
        RECT 103.835 168.360 107.785 168.510 ;
        RECT 103.835 167.910 104.235 168.360 ;
        RECT 103.835 167.760 107.785 167.910 ;
        RECT 103.835 167.310 104.235 167.760 ;
        RECT 103.835 167.160 107.785 167.310 ;
        RECT 103.835 166.860 104.235 167.160 ;
        RECT 108.385 166.860 108.535 175.060 ;
        RECT 108.985 166.860 109.135 175.060 ;
        RECT 109.585 166.860 109.735 175.060 ;
        RECT 110.185 166.860 110.335 175.060 ;
        RECT 110.785 166.860 110.935 175.060 ;
        RECT 111.385 166.860 111.535 175.060 ;
        RECT 111.985 166.860 112.135 175.060 ;
        RECT 103.835 166.460 112.135 166.860 ;
        RECT 103.835 166.160 104.235 166.460 ;
        RECT 103.835 166.010 107.785 166.160 ;
        RECT 103.835 165.560 104.235 166.010 ;
        RECT 103.835 165.410 107.785 165.560 ;
        RECT 103.835 164.960 104.235 165.410 ;
        RECT 103.835 164.810 107.785 164.960 ;
        RECT 103.835 164.360 104.235 164.810 ;
        RECT 103.835 164.210 107.785 164.360 ;
        RECT 103.835 163.760 104.235 164.210 ;
        RECT 103.835 163.610 107.785 163.760 ;
        RECT 103.835 163.160 104.235 163.610 ;
        RECT 103.835 163.010 107.785 163.160 ;
        RECT 103.835 162.560 104.235 163.010 ;
        RECT 103.835 162.410 107.785 162.560 ;
        RECT 103.835 161.960 104.235 162.410 ;
        RECT 103.835 161.810 107.785 161.960 ;
        RECT 103.835 161.360 104.235 161.810 ;
        RECT 103.835 161.210 107.785 161.360 ;
        RECT 103.835 161.060 104.235 161.210 ;
        RECT 101.035 160.760 104.235 161.060 ;
        RECT 97.485 160.610 107.785 160.760 ;
        RECT 101.035 160.160 104.235 160.610 ;
        RECT 97.485 160.010 107.785 160.160 ;
        RECT 101.035 159.560 104.235 160.010 ;
        RECT 97.485 159.410 107.785 159.560 ;
        RECT 101.035 158.960 104.235 159.410 ;
        RECT 97.485 158.810 107.785 158.960 ;
        RECT 101.435 157.860 103.835 158.810 ;
        RECT 108.385 158.260 108.535 166.460 ;
        RECT 108.985 158.260 109.135 166.460 ;
        RECT 109.585 158.260 109.735 166.460 ;
        RECT 110.185 158.260 110.335 166.460 ;
        RECT 110.785 158.260 110.935 166.460 ;
        RECT 111.385 158.260 111.535 166.460 ;
        RECT 111.985 158.260 112.135 166.460 ;
        RECT 113.135 166.860 113.285 175.060 ;
        RECT 113.735 166.860 113.885 175.060 ;
        RECT 114.335 166.860 114.485 175.060 ;
        RECT 114.935 166.860 115.085 175.060 ;
        RECT 115.535 166.860 115.685 175.060 ;
        RECT 116.135 166.860 116.285 175.060 ;
        RECT 116.735 166.860 116.885 175.060 ;
        RECT 121.435 174.510 122.635 175.460 ;
        RECT 117.485 174.360 122.635 174.510 ;
        RECT 121.035 173.910 122.635 174.360 ;
        RECT 117.485 173.760 122.635 173.910 ;
        RECT 121.035 173.310 122.635 173.760 ;
        RECT 125.140 173.715 127.140 174.990 ;
        RECT 117.485 173.160 122.635 173.310 ;
        RECT 121.035 172.710 122.635 173.160 ;
        RECT 117.485 172.560 122.635 172.710 ;
        RECT 121.035 172.260 122.635 172.560 ;
        RECT 121.035 172.110 121.435 172.260 ;
        RECT 117.485 171.960 121.435 172.110 ;
        RECT 121.035 171.510 121.435 171.960 ;
        RECT 117.485 171.360 121.435 171.510 ;
        RECT 121.035 170.910 121.435 171.360 ;
        RECT 117.485 170.760 121.435 170.910 ;
        RECT 121.035 170.310 121.435 170.760 ;
        RECT 117.485 170.160 121.435 170.310 ;
        RECT 121.035 169.710 121.435 170.160 ;
        RECT 125.140 169.915 127.140 172.210 ;
        RECT 125.140 169.910 127.005 169.915 ;
        RECT 117.485 169.560 121.435 169.710 ;
        RECT 121.035 169.110 121.435 169.560 ;
        RECT 117.485 168.960 121.435 169.110 ;
        RECT 121.035 168.510 121.435 168.960 ;
        RECT 117.485 168.360 121.435 168.510 ;
        RECT 121.035 167.910 121.435 168.360 ;
        RECT 117.485 167.760 121.435 167.910 ;
        RECT 121.035 167.310 121.435 167.760 ;
        RECT 117.485 167.160 121.435 167.310 ;
        RECT 121.035 166.860 121.435 167.160 ;
        RECT 113.135 166.460 121.435 166.860 ;
        RECT 113.135 158.260 113.285 166.460 ;
        RECT 113.735 158.260 113.885 166.460 ;
        RECT 114.335 158.260 114.485 166.460 ;
        RECT 114.935 158.260 115.085 166.460 ;
        RECT 115.535 158.260 115.685 166.460 ;
        RECT 116.135 158.260 116.285 166.460 ;
        RECT 116.735 158.260 116.885 166.460 ;
        RECT 121.035 166.160 121.435 166.460 ;
        RECT 117.485 166.010 121.435 166.160 ;
        RECT 121.035 165.560 121.435 166.010 ;
        RECT 117.485 165.410 121.435 165.560 ;
        RECT 121.035 164.960 121.435 165.410 ;
        RECT 117.485 164.810 121.435 164.960 ;
        RECT 121.035 164.360 121.435 164.810 ;
        RECT 117.485 164.210 121.435 164.360 ;
        RECT 121.035 163.760 121.435 164.210 ;
        RECT 117.485 163.610 121.435 163.760 ;
        RECT 121.035 163.160 121.435 163.610 ;
        RECT 117.485 163.010 121.435 163.160 ;
        RECT 121.035 162.560 121.435 163.010 ;
        RECT 117.485 162.410 121.435 162.560 ;
        RECT 121.035 161.960 121.435 162.410 ;
        RECT 117.485 161.810 121.435 161.960 ;
        RECT 121.035 161.360 121.435 161.810 ;
        RECT 117.485 161.210 121.435 161.360 ;
        RECT 121.035 161.060 121.435 161.210 ;
        RECT 125.140 161.115 127.140 163.410 ;
        RECT 125.140 161.110 127.005 161.115 ;
        RECT 121.035 160.760 122.635 161.060 ;
        RECT 117.485 160.610 122.635 160.760 ;
        RECT 121.035 160.160 122.635 160.610 ;
        RECT 117.485 160.010 122.635 160.160 ;
        RECT 121.035 159.560 122.635 160.010 ;
        RECT 117.485 159.410 122.635 159.560 ;
        RECT 121.035 158.960 122.635 159.410 ;
        RECT 117.485 158.810 122.635 158.960 ;
        RECT 121.435 157.860 122.635 158.810 ;
        RECT 125.135 158.440 127.135 159.715 ;
        RECT 42.635 156.660 47.035 157.860 ;
        RECT 58.235 156.660 67.035 157.860 ;
        RECT 78.235 156.660 87.035 157.860 ;
        RECT 98.235 156.660 107.035 157.860 ;
        RECT 118.235 156.660 122.635 157.860 ;
        RECT 2.315 140.360 4.330 141.800 ;
        RECT 125.125 140.360 127.140 141.800 ;
        RECT 4.730 138.800 9.130 140.000 ;
        RECT 20.330 138.800 29.130 140.000 ;
        RECT 40.330 138.800 49.130 140.000 ;
        RECT 60.330 138.800 69.130 140.000 ;
        RECT 80.330 138.800 89.130 140.000 ;
        RECT 100.330 138.800 109.130 140.000 ;
        RECT 120.330 138.800 124.730 140.000 ;
        RECT 4.730 137.850 5.940 138.800 ;
        RECT 2.315 136.450 4.315 137.725 ;
        RECT 4.730 137.700 9.880 137.850 ;
        RECT 4.730 137.250 6.330 137.700 ;
        RECT 4.730 137.100 9.880 137.250 ;
        RECT 4.730 136.650 6.330 137.100 ;
        RECT 4.730 136.500 9.880 136.650 ;
        RECT 4.730 136.050 6.330 136.500 ;
        RECT 4.730 135.900 9.880 136.050 ;
        RECT 4.730 135.600 6.330 135.900 ;
        RECT 2.315 133.255 4.315 135.555 ;
        RECT 5.930 135.450 6.330 135.600 ;
        RECT 5.930 135.300 9.880 135.450 ;
        RECT 5.930 134.850 6.330 135.300 ;
        RECT 5.930 134.700 9.880 134.850 ;
        RECT 5.930 134.250 6.330 134.700 ;
        RECT 5.930 134.100 9.880 134.250 ;
        RECT 5.930 133.650 6.330 134.100 ;
        RECT 5.930 133.500 9.880 133.650 ;
        RECT 5.930 133.050 6.330 133.500 ;
        RECT 5.930 132.900 9.880 133.050 ;
        RECT 5.930 132.450 6.330 132.900 ;
        RECT 5.930 132.300 9.880 132.450 ;
        RECT 5.930 131.850 6.330 132.300 ;
        RECT 5.930 131.700 9.880 131.850 ;
        RECT 5.930 131.250 6.330 131.700 ;
        RECT 5.930 131.100 9.880 131.250 ;
        RECT 5.930 130.650 6.330 131.100 ;
        RECT 5.930 130.500 9.880 130.650 ;
        RECT 5.930 130.200 6.330 130.500 ;
        RECT 10.480 130.200 10.630 138.400 ;
        RECT 11.080 130.200 11.230 138.400 ;
        RECT 11.680 130.200 11.830 138.400 ;
        RECT 12.280 130.200 12.430 138.400 ;
        RECT 12.880 130.200 13.030 138.400 ;
        RECT 13.480 130.200 13.630 138.400 ;
        RECT 14.080 130.200 14.230 138.400 ;
        RECT 5.930 129.800 14.230 130.200 ;
        RECT 5.930 129.500 6.330 129.800 ;
        RECT 5.930 129.350 9.880 129.500 ;
        RECT 5.930 128.900 6.330 129.350 ;
        RECT 5.930 128.750 9.880 128.900 ;
        RECT 5.930 128.300 6.330 128.750 ;
        RECT 5.930 128.150 9.880 128.300 ;
        RECT 5.930 127.700 6.330 128.150 ;
        RECT 5.930 127.550 9.880 127.700 ;
        RECT 5.930 127.100 6.330 127.550 ;
        RECT 5.930 126.950 9.880 127.100 ;
        RECT 2.315 124.425 4.315 126.745 ;
        RECT 5.930 126.500 6.330 126.950 ;
        RECT 5.930 126.350 9.880 126.500 ;
        RECT 5.930 125.900 6.330 126.350 ;
        RECT 5.930 125.750 9.880 125.900 ;
        RECT 5.930 125.300 6.330 125.750 ;
        RECT 5.930 125.150 9.880 125.300 ;
        RECT 5.930 124.700 6.330 125.150 ;
        RECT 5.930 124.550 9.880 124.700 ;
        RECT 2.315 124.420 4.310 124.425 ;
        RECT 5.930 124.400 6.330 124.550 ;
        RECT 4.730 124.100 6.330 124.400 ;
        RECT 4.730 123.950 9.880 124.100 ;
        RECT 4.730 123.500 6.330 123.950 ;
        RECT 4.730 123.350 9.880 123.500 ;
        RECT 2.315 121.890 4.315 123.165 ;
        RECT 4.730 122.900 6.330 123.350 ;
        RECT 4.730 122.750 9.880 122.900 ;
        RECT 4.730 122.300 6.330 122.750 ;
        RECT 4.730 122.150 9.880 122.300 ;
        RECT 4.730 121.200 5.930 122.150 ;
        RECT 10.480 121.600 10.630 129.800 ;
        RECT 11.080 121.600 11.230 129.800 ;
        RECT 11.680 121.600 11.830 129.800 ;
        RECT 12.280 121.600 12.430 129.800 ;
        RECT 12.880 121.600 13.030 129.800 ;
        RECT 13.480 121.600 13.630 129.800 ;
        RECT 14.080 121.600 14.230 129.800 ;
        RECT 15.230 130.200 15.380 138.400 ;
        RECT 15.830 130.200 15.980 138.400 ;
        RECT 16.430 130.200 16.580 138.400 ;
        RECT 17.030 130.200 17.180 138.400 ;
        RECT 17.630 130.200 17.780 138.400 ;
        RECT 18.230 130.200 18.380 138.400 ;
        RECT 18.830 130.200 18.980 138.400 ;
        RECT 23.530 137.850 25.940 138.800 ;
        RECT 19.580 137.700 29.880 137.850 ;
        RECT 23.130 137.250 26.330 137.700 ;
        RECT 19.580 137.100 29.880 137.250 ;
        RECT 23.130 136.650 26.330 137.100 ;
        RECT 19.580 136.500 29.880 136.650 ;
        RECT 23.130 136.050 26.330 136.500 ;
        RECT 19.580 135.900 29.880 136.050 ;
        RECT 23.130 135.600 26.330 135.900 ;
        RECT 23.130 135.450 23.530 135.600 ;
        RECT 19.580 135.300 23.530 135.450 ;
        RECT 23.130 134.850 23.530 135.300 ;
        RECT 19.580 134.700 23.530 134.850 ;
        RECT 23.130 134.250 23.530 134.700 ;
        RECT 19.580 134.100 23.530 134.250 ;
        RECT 23.130 133.650 23.530 134.100 ;
        RECT 19.580 133.500 23.530 133.650 ;
        RECT 23.130 133.050 23.530 133.500 ;
        RECT 19.580 132.900 23.530 133.050 ;
        RECT 23.130 132.450 23.530 132.900 ;
        RECT 19.580 132.300 23.530 132.450 ;
        RECT 23.130 131.850 23.530 132.300 ;
        RECT 19.580 131.700 23.530 131.850 ;
        RECT 23.130 131.250 23.530 131.700 ;
        RECT 19.580 131.100 23.530 131.250 ;
        RECT 23.130 130.650 23.530 131.100 ;
        RECT 19.580 130.500 23.530 130.650 ;
        RECT 23.130 130.200 23.530 130.500 ;
        RECT 15.230 129.800 23.530 130.200 ;
        RECT 15.230 121.600 15.380 129.800 ;
        RECT 15.830 121.600 15.980 129.800 ;
        RECT 16.430 121.600 16.580 129.800 ;
        RECT 17.030 121.600 17.180 129.800 ;
        RECT 17.630 121.600 17.780 129.800 ;
        RECT 18.230 121.600 18.380 129.800 ;
        RECT 18.830 121.600 18.980 129.800 ;
        RECT 23.130 129.500 23.530 129.800 ;
        RECT 19.580 129.350 23.530 129.500 ;
        RECT 23.130 128.900 23.530 129.350 ;
        RECT 19.580 128.750 23.530 128.900 ;
        RECT 23.130 128.300 23.530 128.750 ;
        RECT 19.580 128.150 23.530 128.300 ;
        RECT 23.130 127.700 23.530 128.150 ;
        RECT 19.580 127.550 23.530 127.700 ;
        RECT 23.130 127.100 23.530 127.550 ;
        RECT 19.580 126.950 23.530 127.100 ;
        RECT 23.130 126.500 23.530 126.950 ;
        RECT 19.580 126.350 23.530 126.500 ;
        RECT 23.130 125.900 23.530 126.350 ;
        RECT 19.580 125.750 23.530 125.900 ;
        RECT 23.130 125.300 23.530 125.750 ;
        RECT 19.580 125.150 23.530 125.300 ;
        RECT 23.130 124.700 23.530 125.150 ;
        RECT 19.580 124.550 23.530 124.700 ;
        RECT 23.130 124.400 23.530 124.550 ;
        RECT 25.930 135.450 26.330 135.600 ;
        RECT 25.930 135.300 29.880 135.450 ;
        RECT 25.930 134.850 26.330 135.300 ;
        RECT 25.930 134.700 29.880 134.850 ;
        RECT 25.930 134.250 26.330 134.700 ;
        RECT 25.930 134.100 29.880 134.250 ;
        RECT 25.930 133.650 26.330 134.100 ;
        RECT 25.930 133.500 29.880 133.650 ;
        RECT 25.930 133.050 26.330 133.500 ;
        RECT 25.930 132.900 29.880 133.050 ;
        RECT 25.930 132.450 26.330 132.900 ;
        RECT 25.930 132.300 29.880 132.450 ;
        RECT 25.930 131.850 26.330 132.300 ;
        RECT 25.930 131.700 29.880 131.850 ;
        RECT 25.930 131.250 26.330 131.700 ;
        RECT 25.930 131.100 29.880 131.250 ;
        RECT 25.930 130.650 26.330 131.100 ;
        RECT 25.930 130.500 29.880 130.650 ;
        RECT 25.930 130.200 26.330 130.500 ;
        RECT 30.480 130.200 30.630 138.400 ;
        RECT 31.080 130.200 31.230 138.400 ;
        RECT 31.680 130.200 31.830 138.400 ;
        RECT 32.280 130.200 32.430 138.400 ;
        RECT 32.880 130.200 33.030 138.400 ;
        RECT 33.480 130.200 33.630 138.400 ;
        RECT 34.080 130.200 34.230 138.400 ;
        RECT 25.930 129.800 34.230 130.200 ;
        RECT 25.930 129.500 26.330 129.800 ;
        RECT 25.930 129.350 29.880 129.500 ;
        RECT 25.930 128.900 26.330 129.350 ;
        RECT 25.930 128.750 29.880 128.900 ;
        RECT 25.930 128.300 26.330 128.750 ;
        RECT 25.930 128.150 29.880 128.300 ;
        RECT 25.930 127.700 26.330 128.150 ;
        RECT 25.930 127.550 29.880 127.700 ;
        RECT 25.930 127.100 26.330 127.550 ;
        RECT 25.930 126.950 29.880 127.100 ;
        RECT 25.930 126.500 26.330 126.950 ;
        RECT 25.930 126.350 29.880 126.500 ;
        RECT 25.930 125.900 26.330 126.350 ;
        RECT 25.930 125.750 29.880 125.900 ;
        RECT 25.930 125.300 26.330 125.750 ;
        RECT 25.930 125.150 29.880 125.300 ;
        RECT 25.930 124.700 26.330 125.150 ;
        RECT 25.930 124.550 29.880 124.700 ;
        RECT 25.930 124.400 26.330 124.550 ;
        RECT 23.130 124.100 26.330 124.400 ;
        RECT 19.580 123.950 29.880 124.100 ;
        RECT 23.130 123.500 26.330 123.950 ;
        RECT 19.580 123.350 29.880 123.500 ;
        RECT 23.130 122.900 26.330 123.350 ;
        RECT 19.580 122.750 29.880 122.900 ;
        RECT 23.130 122.300 26.330 122.750 ;
        RECT 19.580 122.150 29.880 122.300 ;
        RECT 23.530 121.200 25.930 122.150 ;
        RECT 30.480 121.600 30.630 129.800 ;
        RECT 31.080 121.600 31.230 129.800 ;
        RECT 31.680 121.600 31.830 129.800 ;
        RECT 32.280 121.600 32.430 129.800 ;
        RECT 32.880 121.600 33.030 129.800 ;
        RECT 33.480 121.600 33.630 129.800 ;
        RECT 34.080 121.600 34.230 129.800 ;
        RECT 35.230 130.200 35.380 138.400 ;
        RECT 35.830 130.200 35.980 138.400 ;
        RECT 36.430 130.200 36.580 138.400 ;
        RECT 37.030 130.200 37.180 138.400 ;
        RECT 37.630 130.200 37.780 138.400 ;
        RECT 38.230 130.200 38.380 138.400 ;
        RECT 38.830 130.200 38.980 138.400 ;
        RECT 43.530 137.850 45.940 138.800 ;
        RECT 39.580 137.700 49.880 137.850 ;
        RECT 43.130 137.250 46.330 137.700 ;
        RECT 39.580 137.100 49.880 137.250 ;
        RECT 43.130 136.650 46.330 137.100 ;
        RECT 39.580 136.500 49.880 136.650 ;
        RECT 43.130 136.050 46.330 136.500 ;
        RECT 39.580 135.900 49.880 136.050 ;
        RECT 43.130 135.600 46.330 135.900 ;
        RECT 43.130 135.450 43.530 135.600 ;
        RECT 39.580 135.300 43.530 135.450 ;
        RECT 43.130 134.850 43.530 135.300 ;
        RECT 39.580 134.700 43.530 134.850 ;
        RECT 43.130 134.250 43.530 134.700 ;
        RECT 39.580 134.100 43.530 134.250 ;
        RECT 43.130 133.650 43.530 134.100 ;
        RECT 39.580 133.500 43.530 133.650 ;
        RECT 43.130 133.050 43.530 133.500 ;
        RECT 39.580 132.900 43.530 133.050 ;
        RECT 43.130 132.450 43.530 132.900 ;
        RECT 39.580 132.300 43.530 132.450 ;
        RECT 43.130 131.850 43.530 132.300 ;
        RECT 39.580 131.700 43.530 131.850 ;
        RECT 43.130 131.250 43.530 131.700 ;
        RECT 39.580 131.100 43.530 131.250 ;
        RECT 43.130 130.650 43.530 131.100 ;
        RECT 39.580 130.500 43.530 130.650 ;
        RECT 43.130 130.200 43.530 130.500 ;
        RECT 35.230 129.800 43.530 130.200 ;
        RECT 35.230 121.600 35.380 129.800 ;
        RECT 35.830 121.600 35.980 129.800 ;
        RECT 36.430 121.600 36.580 129.800 ;
        RECT 37.030 121.600 37.180 129.800 ;
        RECT 37.630 121.600 37.780 129.800 ;
        RECT 38.230 121.600 38.380 129.800 ;
        RECT 38.830 121.600 38.980 129.800 ;
        RECT 43.130 129.500 43.530 129.800 ;
        RECT 39.580 129.350 43.530 129.500 ;
        RECT 43.130 128.900 43.530 129.350 ;
        RECT 39.580 128.750 43.530 128.900 ;
        RECT 43.130 128.300 43.530 128.750 ;
        RECT 39.580 128.150 43.530 128.300 ;
        RECT 43.130 127.700 43.530 128.150 ;
        RECT 39.580 127.550 43.530 127.700 ;
        RECT 43.130 127.100 43.530 127.550 ;
        RECT 39.580 126.950 43.530 127.100 ;
        RECT 43.130 126.500 43.530 126.950 ;
        RECT 39.580 126.350 43.530 126.500 ;
        RECT 43.130 125.900 43.530 126.350 ;
        RECT 39.580 125.750 43.530 125.900 ;
        RECT 43.130 125.300 43.530 125.750 ;
        RECT 39.580 125.150 43.530 125.300 ;
        RECT 43.130 124.700 43.530 125.150 ;
        RECT 39.580 124.550 43.530 124.700 ;
        RECT 43.130 124.400 43.530 124.550 ;
        RECT 45.930 135.450 46.330 135.600 ;
        RECT 45.930 135.300 49.880 135.450 ;
        RECT 45.930 134.850 46.330 135.300 ;
        RECT 45.930 134.700 49.880 134.850 ;
        RECT 45.930 134.250 46.330 134.700 ;
        RECT 45.930 134.100 49.880 134.250 ;
        RECT 45.930 133.650 46.330 134.100 ;
        RECT 45.930 133.500 49.880 133.650 ;
        RECT 45.930 133.050 46.330 133.500 ;
        RECT 45.930 132.900 49.880 133.050 ;
        RECT 45.930 132.450 46.330 132.900 ;
        RECT 45.930 132.300 49.880 132.450 ;
        RECT 45.930 131.850 46.330 132.300 ;
        RECT 45.930 131.700 49.880 131.850 ;
        RECT 45.930 131.250 46.330 131.700 ;
        RECT 45.930 131.100 49.880 131.250 ;
        RECT 45.930 130.650 46.330 131.100 ;
        RECT 45.930 130.500 49.880 130.650 ;
        RECT 45.930 130.200 46.330 130.500 ;
        RECT 50.480 130.200 50.630 138.400 ;
        RECT 51.080 130.200 51.230 138.400 ;
        RECT 51.680 130.200 51.830 138.400 ;
        RECT 52.280 130.200 52.430 138.400 ;
        RECT 52.880 130.200 53.030 138.400 ;
        RECT 53.480 130.200 53.630 138.400 ;
        RECT 54.080 130.200 54.230 138.400 ;
        RECT 45.930 129.800 54.230 130.200 ;
        RECT 45.930 129.500 46.330 129.800 ;
        RECT 45.930 129.350 49.880 129.500 ;
        RECT 45.930 128.900 46.330 129.350 ;
        RECT 45.930 128.750 49.880 128.900 ;
        RECT 45.930 128.300 46.330 128.750 ;
        RECT 45.930 128.150 49.880 128.300 ;
        RECT 45.930 127.700 46.330 128.150 ;
        RECT 45.930 127.550 49.880 127.700 ;
        RECT 45.930 127.100 46.330 127.550 ;
        RECT 45.930 126.950 49.880 127.100 ;
        RECT 45.930 126.500 46.330 126.950 ;
        RECT 45.930 126.350 49.880 126.500 ;
        RECT 45.930 125.900 46.330 126.350 ;
        RECT 45.930 125.750 49.880 125.900 ;
        RECT 45.930 125.300 46.330 125.750 ;
        RECT 45.930 125.150 49.880 125.300 ;
        RECT 45.930 124.700 46.330 125.150 ;
        RECT 45.930 124.550 49.880 124.700 ;
        RECT 45.930 124.400 46.330 124.550 ;
        RECT 43.130 124.100 46.330 124.400 ;
        RECT 39.580 123.950 49.880 124.100 ;
        RECT 43.130 123.500 46.330 123.950 ;
        RECT 39.580 123.350 49.880 123.500 ;
        RECT 43.130 122.900 46.330 123.350 ;
        RECT 39.580 122.750 49.880 122.900 ;
        RECT 43.130 122.300 46.330 122.750 ;
        RECT 39.580 122.150 49.880 122.300 ;
        RECT 43.530 121.200 45.930 122.150 ;
        RECT 50.480 121.600 50.630 129.800 ;
        RECT 51.080 121.600 51.230 129.800 ;
        RECT 51.680 121.600 51.830 129.800 ;
        RECT 52.280 121.600 52.430 129.800 ;
        RECT 52.880 121.600 53.030 129.800 ;
        RECT 53.480 121.600 53.630 129.800 ;
        RECT 54.080 121.600 54.230 129.800 ;
        RECT 55.230 130.200 55.380 138.400 ;
        RECT 55.830 130.200 55.980 138.400 ;
        RECT 56.430 130.200 56.580 138.400 ;
        RECT 57.030 130.200 57.180 138.400 ;
        RECT 57.630 130.200 57.780 138.400 ;
        RECT 58.230 130.200 58.380 138.400 ;
        RECT 58.830 130.200 58.980 138.400 ;
        RECT 63.530 137.850 65.940 138.800 ;
        RECT 59.580 137.700 69.880 137.850 ;
        RECT 63.130 137.250 66.330 137.700 ;
        RECT 59.580 137.100 69.880 137.250 ;
        RECT 63.130 136.650 66.330 137.100 ;
        RECT 59.580 136.500 69.880 136.650 ;
        RECT 63.130 136.050 66.330 136.500 ;
        RECT 59.580 135.900 69.880 136.050 ;
        RECT 63.130 135.600 66.330 135.900 ;
        RECT 63.130 135.450 63.530 135.600 ;
        RECT 59.580 135.300 63.530 135.450 ;
        RECT 63.130 134.850 63.530 135.300 ;
        RECT 59.580 134.700 63.530 134.850 ;
        RECT 63.130 134.250 63.530 134.700 ;
        RECT 59.580 134.100 63.530 134.250 ;
        RECT 63.130 133.650 63.530 134.100 ;
        RECT 59.580 133.500 63.530 133.650 ;
        RECT 63.130 133.050 63.530 133.500 ;
        RECT 59.580 132.900 63.530 133.050 ;
        RECT 63.130 132.450 63.530 132.900 ;
        RECT 59.580 132.300 63.530 132.450 ;
        RECT 63.130 131.850 63.530 132.300 ;
        RECT 59.580 131.700 63.530 131.850 ;
        RECT 63.130 131.250 63.530 131.700 ;
        RECT 59.580 131.100 63.530 131.250 ;
        RECT 63.130 130.650 63.530 131.100 ;
        RECT 59.580 130.500 63.530 130.650 ;
        RECT 63.130 130.200 63.530 130.500 ;
        RECT 55.230 129.800 63.530 130.200 ;
        RECT 55.230 121.600 55.380 129.800 ;
        RECT 55.830 121.600 55.980 129.800 ;
        RECT 56.430 121.600 56.580 129.800 ;
        RECT 57.030 121.600 57.180 129.800 ;
        RECT 57.630 121.600 57.780 129.800 ;
        RECT 58.230 121.600 58.380 129.800 ;
        RECT 58.830 121.600 58.980 129.800 ;
        RECT 63.130 129.500 63.530 129.800 ;
        RECT 59.580 129.350 63.530 129.500 ;
        RECT 63.130 128.900 63.530 129.350 ;
        RECT 59.580 128.750 63.530 128.900 ;
        RECT 63.130 128.300 63.530 128.750 ;
        RECT 59.580 128.150 63.530 128.300 ;
        RECT 63.130 127.700 63.530 128.150 ;
        RECT 59.580 127.550 63.530 127.700 ;
        RECT 63.130 127.100 63.530 127.550 ;
        RECT 59.580 126.950 63.530 127.100 ;
        RECT 63.130 126.500 63.530 126.950 ;
        RECT 59.580 126.350 63.530 126.500 ;
        RECT 63.130 125.900 63.530 126.350 ;
        RECT 59.580 125.750 63.530 125.900 ;
        RECT 63.130 125.300 63.530 125.750 ;
        RECT 59.580 125.150 63.530 125.300 ;
        RECT 63.130 124.700 63.530 125.150 ;
        RECT 59.580 124.550 63.530 124.700 ;
        RECT 63.130 124.400 63.530 124.550 ;
        RECT 65.930 135.450 66.330 135.600 ;
        RECT 65.930 135.300 69.880 135.450 ;
        RECT 65.930 134.850 66.330 135.300 ;
        RECT 65.930 134.700 69.880 134.850 ;
        RECT 65.930 134.250 66.330 134.700 ;
        RECT 65.930 134.100 69.880 134.250 ;
        RECT 65.930 133.650 66.330 134.100 ;
        RECT 65.930 133.500 69.880 133.650 ;
        RECT 65.930 133.050 66.330 133.500 ;
        RECT 65.930 132.900 69.880 133.050 ;
        RECT 65.930 132.450 66.330 132.900 ;
        RECT 65.930 132.300 69.880 132.450 ;
        RECT 65.930 131.850 66.330 132.300 ;
        RECT 65.930 131.700 69.880 131.850 ;
        RECT 65.930 131.250 66.330 131.700 ;
        RECT 65.930 131.100 69.880 131.250 ;
        RECT 65.930 130.650 66.330 131.100 ;
        RECT 65.930 130.500 69.880 130.650 ;
        RECT 65.930 130.200 66.330 130.500 ;
        RECT 70.480 130.200 70.630 138.400 ;
        RECT 71.080 130.200 71.230 138.400 ;
        RECT 71.680 130.200 71.830 138.400 ;
        RECT 72.280 130.200 72.430 138.400 ;
        RECT 72.880 130.200 73.030 138.400 ;
        RECT 73.480 130.200 73.630 138.400 ;
        RECT 74.080 130.200 74.230 138.400 ;
        RECT 65.930 129.800 74.230 130.200 ;
        RECT 65.930 129.500 66.330 129.800 ;
        RECT 65.930 129.350 69.880 129.500 ;
        RECT 65.930 128.900 66.330 129.350 ;
        RECT 65.930 128.750 69.880 128.900 ;
        RECT 65.930 128.300 66.330 128.750 ;
        RECT 65.930 128.150 69.880 128.300 ;
        RECT 65.930 127.700 66.330 128.150 ;
        RECT 65.930 127.550 69.880 127.700 ;
        RECT 65.930 127.100 66.330 127.550 ;
        RECT 65.930 126.950 69.880 127.100 ;
        RECT 65.930 126.500 66.330 126.950 ;
        RECT 65.930 126.350 69.880 126.500 ;
        RECT 65.930 125.900 66.330 126.350 ;
        RECT 65.930 125.750 69.880 125.900 ;
        RECT 65.930 125.300 66.330 125.750 ;
        RECT 65.930 125.150 69.880 125.300 ;
        RECT 65.930 124.700 66.330 125.150 ;
        RECT 65.930 124.550 69.880 124.700 ;
        RECT 65.930 124.400 66.330 124.550 ;
        RECT 63.130 124.100 66.330 124.400 ;
        RECT 59.580 123.950 69.880 124.100 ;
        RECT 63.130 123.500 66.330 123.950 ;
        RECT 59.580 123.350 69.880 123.500 ;
        RECT 63.130 122.900 66.330 123.350 ;
        RECT 59.580 122.750 69.880 122.900 ;
        RECT 63.130 122.300 66.330 122.750 ;
        RECT 59.580 122.150 69.880 122.300 ;
        RECT 63.530 121.200 65.930 122.150 ;
        RECT 70.480 121.600 70.630 129.800 ;
        RECT 71.080 121.600 71.230 129.800 ;
        RECT 71.680 121.600 71.830 129.800 ;
        RECT 72.280 121.600 72.430 129.800 ;
        RECT 72.880 121.600 73.030 129.800 ;
        RECT 73.480 121.600 73.630 129.800 ;
        RECT 74.080 121.600 74.230 129.800 ;
        RECT 75.230 130.200 75.380 138.400 ;
        RECT 75.830 130.200 75.980 138.400 ;
        RECT 76.430 130.200 76.580 138.400 ;
        RECT 77.030 130.200 77.180 138.400 ;
        RECT 77.630 130.200 77.780 138.400 ;
        RECT 78.230 130.200 78.380 138.400 ;
        RECT 78.830 130.200 78.980 138.400 ;
        RECT 83.530 137.850 85.940 138.800 ;
        RECT 79.580 137.700 89.880 137.850 ;
        RECT 83.130 137.250 86.330 137.700 ;
        RECT 79.580 137.100 89.880 137.250 ;
        RECT 83.130 136.650 86.330 137.100 ;
        RECT 79.580 136.500 89.880 136.650 ;
        RECT 83.130 136.050 86.330 136.500 ;
        RECT 79.580 135.900 89.880 136.050 ;
        RECT 83.130 135.600 86.330 135.900 ;
        RECT 83.130 135.450 83.530 135.600 ;
        RECT 79.580 135.300 83.530 135.450 ;
        RECT 83.130 134.850 83.530 135.300 ;
        RECT 79.580 134.700 83.530 134.850 ;
        RECT 83.130 134.250 83.530 134.700 ;
        RECT 79.580 134.100 83.530 134.250 ;
        RECT 83.130 133.650 83.530 134.100 ;
        RECT 79.580 133.500 83.530 133.650 ;
        RECT 83.130 133.050 83.530 133.500 ;
        RECT 79.580 132.900 83.530 133.050 ;
        RECT 83.130 132.450 83.530 132.900 ;
        RECT 79.580 132.300 83.530 132.450 ;
        RECT 83.130 131.850 83.530 132.300 ;
        RECT 79.580 131.700 83.530 131.850 ;
        RECT 83.130 131.250 83.530 131.700 ;
        RECT 79.580 131.100 83.530 131.250 ;
        RECT 83.130 130.650 83.530 131.100 ;
        RECT 79.580 130.500 83.530 130.650 ;
        RECT 83.130 130.200 83.530 130.500 ;
        RECT 75.230 129.800 83.530 130.200 ;
        RECT 75.230 121.600 75.380 129.800 ;
        RECT 75.830 121.600 75.980 129.800 ;
        RECT 76.430 121.600 76.580 129.800 ;
        RECT 77.030 121.600 77.180 129.800 ;
        RECT 77.630 121.600 77.780 129.800 ;
        RECT 78.230 121.600 78.380 129.800 ;
        RECT 78.830 121.600 78.980 129.800 ;
        RECT 83.130 129.500 83.530 129.800 ;
        RECT 79.580 129.350 83.530 129.500 ;
        RECT 83.130 128.900 83.530 129.350 ;
        RECT 79.580 128.750 83.530 128.900 ;
        RECT 83.130 128.300 83.530 128.750 ;
        RECT 79.580 128.150 83.530 128.300 ;
        RECT 83.130 127.700 83.530 128.150 ;
        RECT 79.580 127.550 83.530 127.700 ;
        RECT 83.130 127.100 83.530 127.550 ;
        RECT 79.580 126.950 83.530 127.100 ;
        RECT 83.130 126.500 83.530 126.950 ;
        RECT 79.580 126.350 83.530 126.500 ;
        RECT 83.130 125.900 83.530 126.350 ;
        RECT 79.580 125.750 83.530 125.900 ;
        RECT 83.130 125.300 83.530 125.750 ;
        RECT 79.580 125.150 83.530 125.300 ;
        RECT 83.130 124.700 83.530 125.150 ;
        RECT 79.580 124.550 83.530 124.700 ;
        RECT 83.130 124.400 83.530 124.550 ;
        RECT 85.930 135.450 86.330 135.600 ;
        RECT 85.930 135.300 89.880 135.450 ;
        RECT 85.930 134.850 86.330 135.300 ;
        RECT 85.930 134.700 89.880 134.850 ;
        RECT 85.930 134.250 86.330 134.700 ;
        RECT 85.930 134.100 89.880 134.250 ;
        RECT 85.930 133.650 86.330 134.100 ;
        RECT 85.930 133.500 89.880 133.650 ;
        RECT 85.930 133.050 86.330 133.500 ;
        RECT 85.930 132.900 89.880 133.050 ;
        RECT 85.930 132.450 86.330 132.900 ;
        RECT 85.930 132.300 89.880 132.450 ;
        RECT 85.930 131.850 86.330 132.300 ;
        RECT 85.930 131.700 89.880 131.850 ;
        RECT 85.930 131.250 86.330 131.700 ;
        RECT 85.930 131.100 89.880 131.250 ;
        RECT 85.930 130.650 86.330 131.100 ;
        RECT 85.930 130.500 89.880 130.650 ;
        RECT 85.930 130.200 86.330 130.500 ;
        RECT 90.480 130.200 90.630 138.400 ;
        RECT 91.080 130.200 91.230 138.400 ;
        RECT 91.680 130.200 91.830 138.400 ;
        RECT 92.280 130.200 92.430 138.400 ;
        RECT 92.880 130.200 93.030 138.400 ;
        RECT 93.480 130.200 93.630 138.400 ;
        RECT 94.080 130.200 94.230 138.400 ;
        RECT 85.930 129.800 94.230 130.200 ;
        RECT 85.930 129.500 86.330 129.800 ;
        RECT 85.930 129.350 89.880 129.500 ;
        RECT 85.930 128.900 86.330 129.350 ;
        RECT 85.930 128.750 89.880 128.900 ;
        RECT 85.930 128.300 86.330 128.750 ;
        RECT 85.930 128.150 89.880 128.300 ;
        RECT 85.930 127.700 86.330 128.150 ;
        RECT 85.930 127.550 89.880 127.700 ;
        RECT 85.930 127.100 86.330 127.550 ;
        RECT 85.930 126.950 89.880 127.100 ;
        RECT 85.930 126.500 86.330 126.950 ;
        RECT 85.930 126.350 89.880 126.500 ;
        RECT 85.930 125.900 86.330 126.350 ;
        RECT 85.930 125.750 89.880 125.900 ;
        RECT 85.930 125.300 86.330 125.750 ;
        RECT 85.930 125.150 89.880 125.300 ;
        RECT 85.930 124.700 86.330 125.150 ;
        RECT 85.930 124.550 89.880 124.700 ;
        RECT 85.930 124.400 86.330 124.550 ;
        RECT 83.130 124.100 86.330 124.400 ;
        RECT 79.580 123.950 89.880 124.100 ;
        RECT 83.130 123.500 86.330 123.950 ;
        RECT 79.580 123.350 89.880 123.500 ;
        RECT 83.130 122.900 86.330 123.350 ;
        RECT 79.580 122.750 89.880 122.900 ;
        RECT 83.130 122.300 86.330 122.750 ;
        RECT 79.580 122.150 89.880 122.300 ;
        RECT 83.530 121.200 85.930 122.150 ;
        RECT 90.480 121.600 90.630 129.800 ;
        RECT 91.080 121.600 91.230 129.800 ;
        RECT 91.680 121.600 91.830 129.800 ;
        RECT 92.280 121.600 92.430 129.800 ;
        RECT 92.880 121.600 93.030 129.800 ;
        RECT 93.480 121.600 93.630 129.800 ;
        RECT 94.080 121.600 94.230 129.800 ;
        RECT 95.230 130.200 95.380 138.400 ;
        RECT 95.830 130.200 95.980 138.400 ;
        RECT 96.430 130.200 96.580 138.400 ;
        RECT 97.030 130.200 97.180 138.400 ;
        RECT 97.630 130.200 97.780 138.400 ;
        RECT 98.230 130.200 98.380 138.400 ;
        RECT 98.830 130.200 98.980 138.400 ;
        RECT 103.530 137.850 105.940 138.800 ;
        RECT 99.580 137.700 109.880 137.850 ;
        RECT 103.130 137.250 106.330 137.700 ;
        RECT 99.580 137.100 109.880 137.250 ;
        RECT 103.130 136.650 106.330 137.100 ;
        RECT 99.580 136.500 109.880 136.650 ;
        RECT 103.130 136.050 106.330 136.500 ;
        RECT 99.580 135.900 109.880 136.050 ;
        RECT 103.130 135.600 106.330 135.900 ;
        RECT 103.130 135.450 103.530 135.600 ;
        RECT 99.580 135.300 103.530 135.450 ;
        RECT 103.130 134.850 103.530 135.300 ;
        RECT 99.580 134.700 103.530 134.850 ;
        RECT 103.130 134.250 103.530 134.700 ;
        RECT 99.580 134.100 103.530 134.250 ;
        RECT 103.130 133.650 103.530 134.100 ;
        RECT 99.580 133.500 103.530 133.650 ;
        RECT 103.130 133.050 103.530 133.500 ;
        RECT 99.580 132.900 103.530 133.050 ;
        RECT 103.130 132.450 103.530 132.900 ;
        RECT 99.580 132.300 103.530 132.450 ;
        RECT 103.130 131.850 103.530 132.300 ;
        RECT 99.580 131.700 103.530 131.850 ;
        RECT 103.130 131.250 103.530 131.700 ;
        RECT 99.580 131.100 103.530 131.250 ;
        RECT 103.130 130.650 103.530 131.100 ;
        RECT 99.580 130.500 103.530 130.650 ;
        RECT 103.130 130.200 103.530 130.500 ;
        RECT 95.230 129.800 103.530 130.200 ;
        RECT 95.230 121.600 95.380 129.800 ;
        RECT 95.830 121.600 95.980 129.800 ;
        RECT 96.430 121.600 96.580 129.800 ;
        RECT 97.030 121.600 97.180 129.800 ;
        RECT 97.630 121.600 97.780 129.800 ;
        RECT 98.230 121.600 98.380 129.800 ;
        RECT 98.830 121.600 98.980 129.800 ;
        RECT 103.130 129.500 103.530 129.800 ;
        RECT 99.580 129.350 103.530 129.500 ;
        RECT 103.130 128.900 103.530 129.350 ;
        RECT 99.580 128.750 103.530 128.900 ;
        RECT 103.130 128.300 103.530 128.750 ;
        RECT 99.580 128.150 103.530 128.300 ;
        RECT 103.130 127.700 103.530 128.150 ;
        RECT 99.580 127.550 103.530 127.700 ;
        RECT 103.130 127.100 103.530 127.550 ;
        RECT 99.580 126.950 103.530 127.100 ;
        RECT 103.130 126.500 103.530 126.950 ;
        RECT 99.580 126.350 103.530 126.500 ;
        RECT 103.130 125.900 103.530 126.350 ;
        RECT 99.580 125.750 103.530 125.900 ;
        RECT 103.130 125.300 103.530 125.750 ;
        RECT 99.580 125.150 103.530 125.300 ;
        RECT 103.130 124.700 103.530 125.150 ;
        RECT 99.580 124.550 103.530 124.700 ;
        RECT 103.130 124.400 103.530 124.550 ;
        RECT 105.930 135.450 106.330 135.600 ;
        RECT 105.930 135.300 109.880 135.450 ;
        RECT 105.930 134.850 106.330 135.300 ;
        RECT 105.930 134.700 109.880 134.850 ;
        RECT 105.930 134.250 106.330 134.700 ;
        RECT 105.930 134.100 109.880 134.250 ;
        RECT 105.930 133.650 106.330 134.100 ;
        RECT 105.930 133.500 109.880 133.650 ;
        RECT 105.930 133.050 106.330 133.500 ;
        RECT 105.930 132.900 109.880 133.050 ;
        RECT 105.930 132.450 106.330 132.900 ;
        RECT 105.930 132.300 109.880 132.450 ;
        RECT 105.930 131.850 106.330 132.300 ;
        RECT 105.930 131.700 109.880 131.850 ;
        RECT 105.930 131.250 106.330 131.700 ;
        RECT 105.930 131.100 109.880 131.250 ;
        RECT 105.930 130.650 106.330 131.100 ;
        RECT 105.930 130.500 109.880 130.650 ;
        RECT 105.930 130.200 106.330 130.500 ;
        RECT 110.480 130.200 110.630 138.400 ;
        RECT 111.080 130.200 111.230 138.400 ;
        RECT 111.680 130.200 111.830 138.400 ;
        RECT 112.280 130.200 112.430 138.400 ;
        RECT 112.880 130.200 113.030 138.400 ;
        RECT 113.480 130.200 113.630 138.400 ;
        RECT 114.080 130.200 114.230 138.400 ;
        RECT 105.930 129.800 114.230 130.200 ;
        RECT 105.930 129.500 106.330 129.800 ;
        RECT 105.930 129.350 109.880 129.500 ;
        RECT 105.930 128.900 106.330 129.350 ;
        RECT 105.930 128.750 109.880 128.900 ;
        RECT 105.930 128.300 106.330 128.750 ;
        RECT 105.930 128.150 109.880 128.300 ;
        RECT 105.930 127.700 106.330 128.150 ;
        RECT 105.930 127.550 109.880 127.700 ;
        RECT 105.930 127.100 106.330 127.550 ;
        RECT 105.930 126.950 109.880 127.100 ;
        RECT 105.930 126.500 106.330 126.950 ;
        RECT 105.930 126.350 109.880 126.500 ;
        RECT 105.930 125.900 106.330 126.350 ;
        RECT 105.930 125.750 109.880 125.900 ;
        RECT 105.930 125.300 106.330 125.750 ;
        RECT 105.930 125.150 109.880 125.300 ;
        RECT 105.930 124.700 106.330 125.150 ;
        RECT 105.930 124.550 109.880 124.700 ;
        RECT 105.930 124.400 106.330 124.550 ;
        RECT 103.130 124.100 106.330 124.400 ;
        RECT 99.580 123.950 109.880 124.100 ;
        RECT 103.130 123.500 106.330 123.950 ;
        RECT 99.580 123.350 109.880 123.500 ;
        RECT 103.130 122.900 106.330 123.350 ;
        RECT 99.580 122.750 109.880 122.900 ;
        RECT 103.130 122.300 106.330 122.750 ;
        RECT 99.580 122.150 109.880 122.300 ;
        RECT 103.530 121.200 105.930 122.150 ;
        RECT 110.480 121.600 110.630 129.800 ;
        RECT 111.080 121.600 111.230 129.800 ;
        RECT 111.680 121.600 111.830 129.800 ;
        RECT 112.280 121.600 112.430 129.800 ;
        RECT 112.880 121.600 113.030 129.800 ;
        RECT 113.480 121.600 113.630 129.800 ;
        RECT 114.080 121.600 114.230 129.800 ;
        RECT 115.230 130.200 115.380 138.400 ;
        RECT 115.830 130.200 115.980 138.400 ;
        RECT 116.430 130.200 116.580 138.400 ;
        RECT 117.030 130.200 117.180 138.400 ;
        RECT 117.630 130.200 117.780 138.400 ;
        RECT 118.230 130.200 118.380 138.400 ;
        RECT 118.830 130.200 118.980 138.400 ;
        RECT 123.530 137.850 124.730 138.800 ;
        RECT 119.580 137.700 124.730 137.850 ;
        RECT 123.130 137.250 124.730 137.700 ;
        RECT 119.580 137.100 124.730 137.250 ;
        RECT 123.130 136.650 124.730 137.100 ;
        RECT 119.580 136.500 124.730 136.650 ;
        RECT 123.130 136.050 124.730 136.500 ;
        RECT 125.140 136.450 127.140 137.725 ;
        RECT 119.580 135.900 124.730 136.050 ;
        RECT 123.130 135.600 124.730 135.900 ;
        RECT 123.130 135.450 123.530 135.600 ;
        RECT 119.580 135.300 123.530 135.450 ;
        RECT 123.130 134.850 123.530 135.300 ;
        RECT 119.580 134.700 123.530 134.850 ;
        RECT 123.130 134.250 123.530 134.700 ;
        RECT 119.580 134.100 123.530 134.250 ;
        RECT 123.130 133.650 123.530 134.100 ;
        RECT 119.580 133.500 123.530 133.650 ;
        RECT 123.130 133.050 123.530 133.500 ;
        RECT 119.580 132.900 123.530 133.050 ;
        RECT 123.130 132.450 123.530 132.900 ;
        RECT 119.580 132.300 123.530 132.450 ;
        RECT 123.130 131.850 123.530 132.300 ;
        RECT 119.580 131.700 123.530 131.850 ;
        RECT 123.130 131.250 123.530 131.700 ;
        RECT 119.580 131.100 123.530 131.250 ;
        RECT 123.130 130.650 123.530 131.100 ;
        RECT 119.580 130.500 123.530 130.650 ;
        RECT 123.130 130.200 123.530 130.500 ;
        RECT 115.230 129.800 123.530 130.200 ;
        RECT 115.230 121.600 115.380 129.800 ;
        RECT 115.830 121.600 115.980 129.800 ;
        RECT 116.430 121.600 116.580 129.800 ;
        RECT 117.030 121.600 117.180 129.800 ;
        RECT 117.630 121.600 117.780 129.800 ;
        RECT 118.230 121.600 118.380 129.800 ;
        RECT 118.830 121.600 118.980 129.800 ;
        RECT 123.130 129.500 123.530 129.800 ;
        RECT 119.580 129.350 123.530 129.500 ;
        RECT 123.130 128.900 123.530 129.350 ;
        RECT 119.580 128.750 123.530 128.900 ;
        RECT 123.130 128.300 123.530 128.750 ;
        RECT 119.580 128.150 123.530 128.300 ;
        RECT 123.130 127.700 123.530 128.150 ;
        RECT 119.580 127.550 123.530 127.700 ;
        RECT 123.130 127.100 123.530 127.550 ;
        RECT 119.580 126.950 123.530 127.100 ;
        RECT 123.130 126.500 123.530 126.950 ;
        RECT 119.580 126.350 123.530 126.500 ;
        RECT 123.130 125.900 123.530 126.350 ;
        RECT 119.580 125.750 123.530 125.900 ;
        RECT 123.130 125.300 123.530 125.750 ;
        RECT 119.580 125.150 123.530 125.300 ;
        RECT 123.130 124.700 123.530 125.150 ;
        RECT 119.580 124.550 123.530 124.700 ;
        RECT 123.130 124.400 123.530 124.550 ;
        RECT 123.130 124.100 124.730 124.400 ;
        RECT 119.580 123.950 124.730 124.100 ;
        RECT 123.130 123.500 124.730 123.950 ;
        RECT 119.580 123.350 124.730 123.500 ;
        RECT 123.130 122.900 124.730 123.350 ;
        RECT 119.580 122.750 124.730 122.900 ;
        RECT 123.130 122.300 124.730 122.750 ;
        RECT 119.580 122.150 124.730 122.300 ;
        RECT 123.530 121.200 124.730 122.150 ;
        RECT 125.140 121.645 127.140 122.920 ;
        RECT 4.730 118.800 9.130 121.200 ;
        RECT 20.330 118.800 29.130 121.200 ;
        RECT 40.330 118.800 49.130 121.200 ;
        RECT 60.330 118.800 69.130 121.200 ;
        RECT 80.330 118.800 89.130 121.200 ;
        RECT 100.330 118.800 109.130 121.200 ;
        RECT 120.330 118.800 124.730 121.200 ;
        RECT 2.315 116.870 4.315 118.145 ;
        RECT 4.730 117.850 5.940 118.800 ;
        RECT 4.730 117.700 9.880 117.850 ;
        RECT 4.730 117.250 6.330 117.700 ;
        RECT 4.730 117.100 9.880 117.250 ;
        RECT 4.730 116.650 6.330 117.100 ;
        RECT 4.730 116.500 9.880 116.650 ;
        RECT 4.730 116.050 6.330 116.500 ;
        RECT 4.730 115.900 9.880 116.050 ;
        RECT 4.730 115.600 6.330 115.900 ;
        RECT 2.315 113.250 4.315 115.545 ;
        RECT 5.930 115.450 6.330 115.600 ;
        RECT 5.930 115.300 9.880 115.450 ;
        RECT 5.930 114.850 6.330 115.300 ;
        RECT 5.930 114.700 9.880 114.850 ;
        RECT 5.930 114.250 6.330 114.700 ;
        RECT 5.930 114.100 9.880 114.250 ;
        RECT 5.930 113.650 6.330 114.100 ;
        RECT 5.930 113.500 9.880 113.650 ;
        RECT 5.930 113.050 6.330 113.500 ;
        RECT 5.930 112.900 9.880 113.050 ;
        RECT 5.930 112.450 6.330 112.900 ;
        RECT 5.930 112.300 9.880 112.450 ;
        RECT 5.930 111.850 6.330 112.300 ;
        RECT 5.930 111.700 9.880 111.850 ;
        RECT 5.930 111.250 6.330 111.700 ;
        RECT 5.930 111.100 9.880 111.250 ;
        RECT 5.930 110.650 6.330 111.100 ;
        RECT 5.930 110.500 9.880 110.650 ;
        RECT 5.930 110.200 6.330 110.500 ;
        RECT 10.480 110.200 10.630 118.400 ;
        RECT 11.080 110.200 11.230 118.400 ;
        RECT 11.680 110.200 11.830 118.400 ;
        RECT 12.280 110.200 12.430 118.400 ;
        RECT 12.880 110.200 13.030 118.400 ;
        RECT 13.480 110.200 13.630 118.400 ;
        RECT 14.080 110.200 14.230 118.400 ;
        RECT 5.930 109.800 14.230 110.200 ;
        RECT 5.930 109.500 6.330 109.800 ;
        RECT 5.930 109.350 9.880 109.500 ;
        RECT 5.930 108.900 6.330 109.350 ;
        RECT 5.930 108.750 9.880 108.900 ;
        RECT 5.930 108.300 6.330 108.750 ;
        RECT 5.930 108.150 9.880 108.300 ;
        RECT 5.930 107.700 6.330 108.150 ;
        RECT 5.930 107.550 9.880 107.700 ;
        RECT 5.930 107.100 6.330 107.550 ;
        RECT 5.930 106.950 9.880 107.100 ;
        RECT 2.315 104.450 4.315 106.745 ;
        RECT 5.930 106.500 6.330 106.950 ;
        RECT 5.930 106.350 9.880 106.500 ;
        RECT 5.930 105.900 6.330 106.350 ;
        RECT 5.930 105.750 9.880 105.900 ;
        RECT 5.930 105.300 6.330 105.750 ;
        RECT 5.930 105.150 9.880 105.300 ;
        RECT 5.930 104.700 6.330 105.150 ;
        RECT 5.930 104.550 9.880 104.700 ;
        RECT 5.930 104.400 6.330 104.550 ;
        RECT 4.730 104.100 6.330 104.400 ;
        RECT 4.730 103.950 9.880 104.100 ;
        RECT 4.730 103.500 6.330 103.950 ;
        RECT 4.730 103.350 9.880 103.500 ;
        RECT 2.315 101.980 4.320 103.255 ;
        RECT 4.730 102.900 6.330 103.350 ;
        RECT 4.730 102.750 9.880 102.900 ;
        RECT 4.730 102.300 6.330 102.750 ;
        RECT 4.730 102.150 9.880 102.300 ;
        RECT 4.730 101.200 5.930 102.150 ;
        RECT 10.480 101.600 10.630 109.800 ;
        RECT 11.080 101.600 11.230 109.800 ;
        RECT 11.680 101.600 11.830 109.800 ;
        RECT 12.280 101.600 12.430 109.800 ;
        RECT 12.880 101.600 13.030 109.800 ;
        RECT 13.480 101.600 13.630 109.800 ;
        RECT 14.080 101.600 14.230 109.800 ;
        RECT 15.230 110.200 15.380 118.400 ;
        RECT 15.830 110.200 15.980 118.400 ;
        RECT 16.430 110.200 16.580 118.400 ;
        RECT 17.030 110.200 17.180 118.400 ;
        RECT 17.630 110.200 17.780 118.400 ;
        RECT 18.230 110.200 18.380 118.400 ;
        RECT 18.830 110.200 18.980 118.400 ;
        RECT 23.530 117.850 25.940 118.800 ;
        RECT 19.580 117.700 29.880 117.850 ;
        RECT 23.130 117.250 26.330 117.700 ;
        RECT 19.580 117.100 29.880 117.250 ;
        RECT 23.130 116.650 26.330 117.100 ;
        RECT 19.580 116.500 29.880 116.650 ;
        RECT 23.130 116.050 26.330 116.500 ;
        RECT 19.580 115.900 29.880 116.050 ;
        RECT 23.130 115.600 26.330 115.900 ;
        RECT 23.130 115.450 23.530 115.600 ;
        RECT 19.580 115.300 23.530 115.450 ;
        RECT 23.130 114.850 23.530 115.300 ;
        RECT 19.580 114.700 23.530 114.850 ;
        RECT 23.130 114.250 23.530 114.700 ;
        RECT 19.580 114.100 23.530 114.250 ;
        RECT 23.130 113.650 23.530 114.100 ;
        RECT 19.580 113.500 23.530 113.650 ;
        RECT 23.130 113.050 23.530 113.500 ;
        RECT 19.580 112.900 23.530 113.050 ;
        RECT 23.130 112.450 23.530 112.900 ;
        RECT 19.580 112.300 23.530 112.450 ;
        RECT 23.130 111.850 23.530 112.300 ;
        RECT 19.580 111.700 23.530 111.850 ;
        RECT 23.130 111.250 23.530 111.700 ;
        RECT 19.580 111.100 23.530 111.250 ;
        RECT 23.130 110.650 23.530 111.100 ;
        RECT 19.580 110.500 23.530 110.650 ;
        RECT 23.130 110.200 23.530 110.500 ;
        RECT 15.230 109.800 23.530 110.200 ;
        RECT 15.230 101.600 15.380 109.800 ;
        RECT 15.830 101.600 15.980 109.800 ;
        RECT 16.430 101.600 16.580 109.800 ;
        RECT 17.030 101.600 17.180 109.800 ;
        RECT 17.630 101.600 17.780 109.800 ;
        RECT 18.230 101.600 18.380 109.800 ;
        RECT 18.830 101.600 18.980 109.800 ;
        RECT 23.130 109.500 23.530 109.800 ;
        RECT 19.580 109.350 23.530 109.500 ;
        RECT 23.130 108.900 23.530 109.350 ;
        RECT 19.580 108.750 23.530 108.900 ;
        RECT 23.130 108.300 23.530 108.750 ;
        RECT 19.580 108.150 23.530 108.300 ;
        RECT 23.130 107.700 23.530 108.150 ;
        RECT 19.580 107.550 23.530 107.700 ;
        RECT 23.130 107.100 23.530 107.550 ;
        RECT 19.580 106.950 23.530 107.100 ;
        RECT 23.130 106.500 23.530 106.950 ;
        RECT 19.580 106.350 23.530 106.500 ;
        RECT 23.130 105.900 23.530 106.350 ;
        RECT 19.580 105.750 23.530 105.900 ;
        RECT 23.130 105.300 23.530 105.750 ;
        RECT 19.580 105.150 23.530 105.300 ;
        RECT 23.130 104.700 23.530 105.150 ;
        RECT 19.580 104.550 23.530 104.700 ;
        RECT 23.130 104.400 23.530 104.550 ;
        RECT 25.930 115.450 26.330 115.600 ;
        RECT 25.930 115.300 29.880 115.450 ;
        RECT 25.930 114.850 26.330 115.300 ;
        RECT 25.930 114.700 29.880 114.850 ;
        RECT 25.930 114.250 26.330 114.700 ;
        RECT 25.930 114.100 29.880 114.250 ;
        RECT 25.930 113.650 26.330 114.100 ;
        RECT 25.930 113.500 29.880 113.650 ;
        RECT 25.930 113.050 26.330 113.500 ;
        RECT 25.930 112.900 29.880 113.050 ;
        RECT 25.930 112.450 26.330 112.900 ;
        RECT 25.930 112.300 29.880 112.450 ;
        RECT 25.930 111.850 26.330 112.300 ;
        RECT 25.930 111.700 29.880 111.850 ;
        RECT 25.930 111.250 26.330 111.700 ;
        RECT 25.930 111.100 29.880 111.250 ;
        RECT 25.930 110.650 26.330 111.100 ;
        RECT 25.930 110.500 29.880 110.650 ;
        RECT 25.930 110.200 26.330 110.500 ;
        RECT 30.480 110.200 30.630 118.400 ;
        RECT 31.080 110.200 31.230 118.400 ;
        RECT 31.680 110.200 31.830 118.400 ;
        RECT 32.280 110.200 32.430 118.400 ;
        RECT 32.880 110.200 33.030 118.400 ;
        RECT 33.480 110.200 33.630 118.400 ;
        RECT 34.080 110.200 34.230 118.400 ;
        RECT 25.930 109.800 34.230 110.200 ;
        RECT 25.930 109.500 26.330 109.800 ;
        RECT 25.930 109.350 29.880 109.500 ;
        RECT 25.930 108.900 26.330 109.350 ;
        RECT 25.930 108.750 29.880 108.900 ;
        RECT 25.930 108.300 26.330 108.750 ;
        RECT 25.930 108.150 29.880 108.300 ;
        RECT 25.930 107.700 26.330 108.150 ;
        RECT 25.930 107.550 29.880 107.700 ;
        RECT 25.930 107.100 26.330 107.550 ;
        RECT 25.930 106.950 29.880 107.100 ;
        RECT 25.930 106.500 26.330 106.950 ;
        RECT 25.930 106.350 29.880 106.500 ;
        RECT 25.930 105.900 26.330 106.350 ;
        RECT 25.930 105.750 29.880 105.900 ;
        RECT 25.930 105.300 26.330 105.750 ;
        RECT 25.930 105.150 29.880 105.300 ;
        RECT 25.930 104.700 26.330 105.150 ;
        RECT 25.930 104.550 29.880 104.700 ;
        RECT 25.930 104.400 26.330 104.550 ;
        RECT 23.130 104.100 26.330 104.400 ;
        RECT 19.580 103.950 29.880 104.100 ;
        RECT 23.130 103.500 26.330 103.950 ;
        RECT 19.580 103.350 29.880 103.500 ;
        RECT 23.130 102.900 26.330 103.350 ;
        RECT 19.580 102.750 29.880 102.900 ;
        RECT 23.130 102.300 26.330 102.750 ;
        RECT 19.580 102.150 29.880 102.300 ;
        RECT 23.530 101.200 25.930 102.150 ;
        RECT 30.480 101.600 30.630 109.800 ;
        RECT 31.080 101.600 31.230 109.800 ;
        RECT 31.680 101.600 31.830 109.800 ;
        RECT 32.280 101.600 32.430 109.800 ;
        RECT 32.880 101.600 33.030 109.800 ;
        RECT 33.480 101.600 33.630 109.800 ;
        RECT 34.080 101.600 34.230 109.800 ;
        RECT 35.230 110.200 35.380 118.400 ;
        RECT 35.830 110.200 35.980 118.400 ;
        RECT 36.430 110.200 36.580 118.400 ;
        RECT 37.030 110.200 37.180 118.400 ;
        RECT 37.630 110.200 37.780 118.400 ;
        RECT 38.230 110.200 38.380 118.400 ;
        RECT 38.830 110.200 38.980 118.400 ;
        RECT 43.530 117.850 45.940 118.800 ;
        RECT 39.580 117.700 49.880 117.850 ;
        RECT 43.130 117.250 46.330 117.700 ;
        RECT 39.580 117.100 49.880 117.250 ;
        RECT 43.130 116.650 46.330 117.100 ;
        RECT 39.580 116.500 49.880 116.650 ;
        RECT 43.130 116.050 46.330 116.500 ;
        RECT 39.580 115.900 49.880 116.050 ;
        RECT 43.130 115.600 46.330 115.900 ;
        RECT 43.130 115.450 43.530 115.600 ;
        RECT 39.580 115.300 43.530 115.450 ;
        RECT 43.130 114.850 43.530 115.300 ;
        RECT 39.580 114.700 43.530 114.850 ;
        RECT 43.130 114.250 43.530 114.700 ;
        RECT 39.580 114.100 43.530 114.250 ;
        RECT 43.130 113.650 43.530 114.100 ;
        RECT 39.580 113.500 43.530 113.650 ;
        RECT 43.130 113.050 43.530 113.500 ;
        RECT 39.580 112.900 43.530 113.050 ;
        RECT 43.130 112.450 43.530 112.900 ;
        RECT 39.580 112.300 43.530 112.450 ;
        RECT 43.130 111.850 43.530 112.300 ;
        RECT 39.580 111.700 43.530 111.850 ;
        RECT 43.130 111.250 43.530 111.700 ;
        RECT 39.580 111.100 43.530 111.250 ;
        RECT 43.130 110.650 43.530 111.100 ;
        RECT 39.580 110.500 43.530 110.650 ;
        RECT 43.130 110.200 43.530 110.500 ;
        RECT 35.230 109.800 43.530 110.200 ;
        RECT 35.230 101.600 35.380 109.800 ;
        RECT 35.830 101.600 35.980 109.800 ;
        RECT 36.430 101.600 36.580 109.800 ;
        RECT 37.030 101.600 37.180 109.800 ;
        RECT 37.630 101.600 37.780 109.800 ;
        RECT 38.230 101.600 38.380 109.800 ;
        RECT 38.830 101.600 38.980 109.800 ;
        RECT 43.130 109.500 43.530 109.800 ;
        RECT 39.580 109.350 43.530 109.500 ;
        RECT 43.130 108.900 43.530 109.350 ;
        RECT 39.580 108.750 43.530 108.900 ;
        RECT 43.130 108.300 43.530 108.750 ;
        RECT 39.580 108.150 43.530 108.300 ;
        RECT 43.130 107.700 43.530 108.150 ;
        RECT 39.580 107.550 43.530 107.700 ;
        RECT 43.130 107.100 43.530 107.550 ;
        RECT 39.580 106.950 43.530 107.100 ;
        RECT 43.130 106.500 43.530 106.950 ;
        RECT 39.580 106.350 43.530 106.500 ;
        RECT 43.130 105.900 43.530 106.350 ;
        RECT 39.580 105.750 43.530 105.900 ;
        RECT 43.130 105.300 43.530 105.750 ;
        RECT 39.580 105.150 43.530 105.300 ;
        RECT 43.130 104.700 43.530 105.150 ;
        RECT 39.580 104.550 43.530 104.700 ;
        RECT 43.130 104.400 43.530 104.550 ;
        RECT 45.930 115.450 46.330 115.600 ;
        RECT 45.930 115.300 49.880 115.450 ;
        RECT 45.930 114.850 46.330 115.300 ;
        RECT 45.930 114.700 49.880 114.850 ;
        RECT 45.930 114.250 46.330 114.700 ;
        RECT 45.930 114.100 49.880 114.250 ;
        RECT 45.930 113.650 46.330 114.100 ;
        RECT 45.930 113.500 49.880 113.650 ;
        RECT 45.930 113.050 46.330 113.500 ;
        RECT 45.930 112.900 49.880 113.050 ;
        RECT 45.930 112.450 46.330 112.900 ;
        RECT 45.930 112.300 49.880 112.450 ;
        RECT 45.930 111.850 46.330 112.300 ;
        RECT 45.930 111.700 49.880 111.850 ;
        RECT 45.930 111.250 46.330 111.700 ;
        RECT 45.930 111.100 49.880 111.250 ;
        RECT 45.930 110.650 46.330 111.100 ;
        RECT 45.930 110.500 49.880 110.650 ;
        RECT 45.930 110.200 46.330 110.500 ;
        RECT 50.480 110.200 50.630 118.400 ;
        RECT 51.080 110.200 51.230 118.400 ;
        RECT 51.680 110.200 51.830 118.400 ;
        RECT 52.280 110.200 52.430 118.400 ;
        RECT 52.880 110.200 53.030 118.400 ;
        RECT 53.480 110.200 53.630 118.400 ;
        RECT 54.080 110.200 54.230 118.400 ;
        RECT 45.930 109.800 54.230 110.200 ;
        RECT 45.930 109.500 46.330 109.800 ;
        RECT 45.930 109.350 49.880 109.500 ;
        RECT 45.930 108.900 46.330 109.350 ;
        RECT 45.930 108.750 49.880 108.900 ;
        RECT 45.930 108.300 46.330 108.750 ;
        RECT 45.930 108.150 49.880 108.300 ;
        RECT 45.930 107.700 46.330 108.150 ;
        RECT 45.930 107.550 49.880 107.700 ;
        RECT 45.930 107.100 46.330 107.550 ;
        RECT 45.930 106.950 49.880 107.100 ;
        RECT 45.930 106.500 46.330 106.950 ;
        RECT 45.930 106.350 49.880 106.500 ;
        RECT 45.930 105.900 46.330 106.350 ;
        RECT 45.930 105.750 49.880 105.900 ;
        RECT 45.930 105.300 46.330 105.750 ;
        RECT 45.930 105.150 49.880 105.300 ;
        RECT 45.930 104.700 46.330 105.150 ;
        RECT 45.930 104.550 49.880 104.700 ;
        RECT 45.930 104.400 46.330 104.550 ;
        RECT 43.130 104.100 46.330 104.400 ;
        RECT 39.580 103.950 49.880 104.100 ;
        RECT 43.130 103.500 46.330 103.950 ;
        RECT 39.580 103.350 49.880 103.500 ;
        RECT 43.130 102.900 46.330 103.350 ;
        RECT 39.580 102.750 49.880 102.900 ;
        RECT 43.130 102.300 46.330 102.750 ;
        RECT 39.580 102.150 49.880 102.300 ;
        RECT 43.530 101.200 45.930 102.150 ;
        RECT 50.480 101.600 50.630 109.800 ;
        RECT 51.080 101.600 51.230 109.800 ;
        RECT 51.680 101.600 51.830 109.800 ;
        RECT 52.280 101.600 52.430 109.800 ;
        RECT 52.880 101.600 53.030 109.800 ;
        RECT 53.480 101.600 53.630 109.800 ;
        RECT 54.080 101.600 54.230 109.800 ;
        RECT 55.230 110.200 55.380 118.400 ;
        RECT 55.830 110.200 55.980 118.400 ;
        RECT 56.430 110.200 56.580 118.400 ;
        RECT 57.030 110.200 57.180 118.400 ;
        RECT 57.630 110.200 57.780 118.400 ;
        RECT 58.230 110.200 58.380 118.400 ;
        RECT 58.830 110.200 58.980 118.400 ;
        RECT 63.530 117.850 65.940 118.800 ;
        RECT 59.580 117.700 69.880 117.850 ;
        RECT 63.130 117.250 66.330 117.700 ;
        RECT 59.580 117.100 69.880 117.250 ;
        RECT 63.130 116.650 66.330 117.100 ;
        RECT 59.580 116.500 69.880 116.650 ;
        RECT 63.130 116.050 66.330 116.500 ;
        RECT 59.580 115.900 69.880 116.050 ;
        RECT 63.130 115.600 66.330 115.900 ;
        RECT 63.130 115.450 63.530 115.600 ;
        RECT 59.580 115.300 63.530 115.450 ;
        RECT 63.130 114.850 63.530 115.300 ;
        RECT 59.580 114.700 63.530 114.850 ;
        RECT 63.130 114.250 63.530 114.700 ;
        RECT 59.580 114.100 63.530 114.250 ;
        RECT 63.130 113.650 63.530 114.100 ;
        RECT 59.580 113.500 63.530 113.650 ;
        RECT 63.130 113.050 63.530 113.500 ;
        RECT 59.580 112.900 63.530 113.050 ;
        RECT 63.130 112.450 63.530 112.900 ;
        RECT 59.580 112.300 63.530 112.450 ;
        RECT 63.130 111.850 63.530 112.300 ;
        RECT 59.580 111.700 63.530 111.850 ;
        RECT 63.130 111.250 63.530 111.700 ;
        RECT 59.580 111.100 63.530 111.250 ;
        RECT 63.130 110.650 63.530 111.100 ;
        RECT 59.580 110.500 63.530 110.650 ;
        RECT 63.130 110.200 63.530 110.500 ;
        RECT 55.230 109.800 63.530 110.200 ;
        RECT 55.230 101.600 55.380 109.800 ;
        RECT 55.830 101.600 55.980 109.800 ;
        RECT 56.430 101.600 56.580 109.800 ;
        RECT 57.030 101.600 57.180 109.800 ;
        RECT 57.630 101.600 57.780 109.800 ;
        RECT 58.230 101.600 58.380 109.800 ;
        RECT 58.830 101.600 58.980 109.800 ;
        RECT 63.130 109.500 63.530 109.800 ;
        RECT 59.580 109.350 63.530 109.500 ;
        RECT 63.130 108.900 63.530 109.350 ;
        RECT 59.580 108.750 63.530 108.900 ;
        RECT 63.130 108.300 63.530 108.750 ;
        RECT 59.580 108.150 63.530 108.300 ;
        RECT 63.130 107.700 63.530 108.150 ;
        RECT 59.580 107.550 63.530 107.700 ;
        RECT 63.130 107.100 63.530 107.550 ;
        RECT 59.580 106.950 63.530 107.100 ;
        RECT 63.130 106.500 63.530 106.950 ;
        RECT 59.580 106.350 63.530 106.500 ;
        RECT 63.130 105.900 63.530 106.350 ;
        RECT 59.580 105.750 63.530 105.900 ;
        RECT 63.130 105.300 63.530 105.750 ;
        RECT 59.580 105.150 63.530 105.300 ;
        RECT 63.130 104.700 63.530 105.150 ;
        RECT 59.580 104.550 63.530 104.700 ;
        RECT 63.130 104.400 63.530 104.550 ;
        RECT 65.930 115.450 66.330 115.600 ;
        RECT 65.930 115.300 69.880 115.450 ;
        RECT 65.930 114.850 66.330 115.300 ;
        RECT 65.930 114.700 69.880 114.850 ;
        RECT 65.930 114.250 66.330 114.700 ;
        RECT 65.930 114.100 69.880 114.250 ;
        RECT 65.930 113.650 66.330 114.100 ;
        RECT 65.930 113.500 69.880 113.650 ;
        RECT 65.930 113.050 66.330 113.500 ;
        RECT 65.930 112.900 69.880 113.050 ;
        RECT 65.930 112.450 66.330 112.900 ;
        RECT 65.930 112.300 69.880 112.450 ;
        RECT 65.930 111.850 66.330 112.300 ;
        RECT 65.930 111.700 69.880 111.850 ;
        RECT 65.930 111.250 66.330 111.700 ;
        RECT 65.930 111.100 69.880 111.250 ;
        RECT 65.930 110.650 66.330 111.100 ;
        RECT 65.930 110.500 69.880 110.650 ;
        RECT 65.930 110.200 66.330 110.500 ;
        RECT 70.480 110.200 70.630 118.400 ;
        RECT 71.080 110.200 71.230 118.400 ;
        RECT 71.680 110.200 71.830 118.400 ;
        RECT 72.280 110.200 72.430 118.400 ;
        RECT 72.880 110.200 73.030 118.400 ;
        RECT 73.480 110.200 73.630 118.400 ;
        RECT 74.080 110.200 74.230 118.400 ;
        RECT 65.930 109.800 74.230 110.200 ;
        RECT 65.930 109.500 66.330 109.800 ;
        RECT 65.930 109.350 69.880 109.500 ;
        RECT 65.930 108.900 66.330 109.350 ;
        RECT 65.930 108.750 69.880 108.900 ;
        RECT 65.930 108.300 66.330 108.750 ;
        RECT 65.930 108.150 69.880 108.300 ;
        RECT 65.930 107.700 66.330 108.150 ;
        RECT 65.930 107.550 69.880 107.700 ;
        RECT 65.930 107.100 66.330 107.550 ;
        RECT 65.930 106.950 69.880 107.100 ;
        RECT 65.930 106.500 66.330 106.950 ;
        RECT 65.930 106.350 69.880 106.500 ;
        RECT 65.930 105.900 66.330 106.350 ;
        RECT 65.930 105.750 69.880 105.900 ;
        RECT 65.930 105.300 66.330 105.750 ;
        RECT 65.930 105.150 69.880 105.300 ;
        RECT 65.930 104.700 66.330 105.150 ;
        RECT 65.930 104.550 69.880 104.700 ;
        RECT 65.930 104.400 66.330 104.550 ;
        RECT 63.130 104.100 66.330 104.400 ;
        RECT 59.580 103.950 69.880 104.100 ;
        RECT 63.130 103.500 66.330 103.950 ;
        RECT 59.580 103.350 69.880 103.500 ;
        RECT 63.130 102.900 66.330 103.350 ;
        RECT 59.580 102.750 69.880 102.900 ;
        RECT 63.130 102.300 66.330 102.750 ;
        RECT 59.580 102.150 69.880 102.300 ;
        RECT 63.530 101.200 65.930 102.150 ;
        RECT 70.480 101.600 70.630 109.800 ;
        RECT 71.080 101.600 71.230 109.800 ;
        RECT 71.680 101.600 71.830 109.800 ;
        RECT 72.280 101.600 72.430 109.800 ;
        RECT 72.880 101.600 73.030 109.800 ;
        RECT 73.480 101.600 73.630 109.800 ;
        RECT 74.080 101.600 74.230 109.800 ;
        RECT 75.230 110.200 75.380 118.400 ;
        RECT 75.830 110.200 75.980 118.400 ;
        RECT 76.430 110.200 76.580 118.400 ;
        RECT 77.030 110.200 77.180 118.400 ;
        RECT 77.630 110.200 77.780 118.400 ;
        RECT 78.230 110.200 78.380 118.400 ;
        RECT 78.830 110.200 78.980 118.400 ;
        RECT 83.530 117.850 85.940 118.800 ;
        RECT 79.580 117.700 89.880 117.850 ;
        RECT 83.130 117.250 86.330 117.700 ;
        RECT 79.580 117.100 89.880 117.250 ;
        RECT 83.130 116.650 86.330 117.100 ;
        RECT 79.580 116.500 89.880 116.650 ;
        RECT 83.130 116.050 86.330 116.500 ;
        RECT 79.580 115.900 89.880 116.050 ;
        RECT 83.130 115.600 86.330 115.900 ;
        RECT 83.130 115.450 83.530 115.600 ;
        RECT 79.580 115.300 83.530 115.450 ;
        RECT 83.130 114.850 83.530 115.300 ;
        RECT 79.580 114.700 83.530 114.850 ;
        RECT 83.130 114.250 83.530 114.700 ;
        RECT 79.580 114.100 83.530 114.250 ;
        RECT 83.130 113.650 83.530 114.100 ;
        RECT 79.580 113.500 83.530 113.650 ;
        RECT 83.130 113.050 83.530 113.500 ;
        RECT 79.580 112.900 83.530 113.050 ;
        RECT 83.130 112.450 83.530 112.900 ;
        RECT 79.580 112.300 83.530 112.450 ;
        RECT 83.130 111.850 83.530 112.300 ;
        RECT 79.580 111.700 83.530 111.850 ;
        RECT 83.130 111.250 83.530 111.700 ;
        RECT 79.580 111.100 83.530 111.250 ;
        RECT 83.130 110.650 83.530 111.100 ;
        RECT 79.580 110.500 83.530 110.650 ;
        RECT 83.130 110.200 83.530 110.500 ;
        RECT 75.230 109.800 83.530 110.200 ;
        RECT 75.230 101.600 75.380 109.800 ;
        RECT 75.830 101.600 75.980 109.800 ;
        RECT 76.430 101.600 76.580 109.800 ;
        RECT 77.030 101.600 77.180 109.800 ;
        RECT 77.630 101.600 77.780 109.800 ;
        RECT 78.230 101.600 78.380 109.800 ;
        RECT 78.830 101.600 78.980 109.800 ;
        RECT 83.130 109.500 83.530 109.800 ;
        RECT 79.580 109.350 83.530 109.500 ;
        RECT 83.130 108.900 83.530 109.350 ;
        RECT 79.580 108.750 83.530 108.900 ;
        RECT 83.130 108.300 83.530 108.750 ;
        RECT 79.580 108.150 83.530 108.300 ;
        RECT 83.130 107.700 83.530 108.150 ;
        RECT 79.580 107.550 83.530 107.700 ;
        RECT 83.130 107.100 83.530 107.550 ;
        RECT 79.580 106.950 83.530 107.100 ;
        RECT 83.130 106.500 83.530 106.950 ;
        RECT 79.580 106.350 83.530 106.500 ;
        RECT 83.130 105.900 83.530 106.350 ;
        RECT 79.580 105.750 83.530 105.900 ;
        RECT 83.130 105.300 83.530 105.750 ;
        RECT 79.580 105.150 83.530 105.300 ;
        RECT 83.130 104.700 83.530 105.150 ;
        RECT 79.580 104.550 83.530 104.700 ;
        RECT 83.130 104.400 83.530 104.550 ;
        RECT 85.930 115.450 86.330 115.600 ;
        RECT 85.930 115.300 89.880 115.450 ;
        RECT 85.930 114.850 86.330 115.300 ;
        RECT 85.930 114.700 89.880 114.850 ;
        RECT 85.930 114.250 86.330 114.700 ;
        RECT 85.930 114.100 89.880 114.250 ;
        RECT 85.930 113.650 86.330 114.100 ;
        RECT 85.930 113.500 89.880 113.650 ;
        RECT 85.930 113.050 86.330 113.500 ;
        RECT 85.930 112.900 89.880 113.050 ;
        RECT 85.930 112.450 86.330 112.900 ;
        RECT 85.930 112.300 89.880 112.450 ;
        RECT 85.930 111.850 86.330 112.300 ;
        RECT 85.930 111.700 89.880 111.850 ;
        RECT 85.930 111.250 86.330 111.700 ;
        RECT 85.930 111.100 89.880 111.250 ;
        RECT 85.930 110.650 86.330 111.100 ;
        RECT 85.930 110.500 89.880 110.650 ;
        RECT 85.930 110.200 86.330 110.500 ;
        RECT 90.480 110.200 90.630 118.400 ;
        RECT 91.080 110.200 91.230 118.400 ;
        RECT 91.680 110.200 91.830 118.400 ;
        RECT 92.280 110.200 92.430 118.400 ;
        RECT 92.880 110.200 93.030 118.400 ;
        RECT 93.480 110.200 93.630 118.400 ;
        RECT 94.080 110.200 94.230 118.400 ;
        RECT 85.930 109.800 94.230 110.200 ;
        RECT 85.930 109.500 86.330 109.800 ;
        RECT 85.930 109.350 89.880 109.500 ;
        RECT 85.930 108.900 86.330 109.350 ;
        RECT 85.930 108.750 89.880 108.900 ;
        RECT 85.930 108.300 86.330 108.750 ;
        RECT 85.930 108.150 89.880 108.300 ;
        RECT 85.930 107.700 86.330 108.150 ;
        RECT 85.930 107.550 89.880 107.700 ;
        RECT 85.930 107.100 86.330 107.550 ;
        RECT 85.930 106.950 89.880 107.100 ;
        RECT 85.930 106.500 86.330 106.950 ;
        RECT 85.930 106.350 89.880 106.500 ;
        RECT 85.930 105.900 86.330 106.350 ;
        RECT 85.930 105.750 89.880 105.900 ;
        RECT 85.930 105.300 86.330 105.750 ;
        RECT 85.930 105.150 89.880 105.300 ;
        RECT 85.930 104.700 86.330 105.150 ;
        RECT 85.930 104.550 89.880 104.700 ;
        RECT 85.930 104.400 86.330 104.550 ;
        RECT 83.130 104.100 86.330 104.400 ;
        RECT 79.580 103.950 89.880 104.100 ;
        RECT 83.130 103.500 86.330 103.950 ;
        RECT 79.580 103.350 89.880 103.500 ;
        RECT 83.130 102.900 86.330 103.350 ;
        RECT 79.580 102.750 89.880 102.900 ;
        RECT 83.130 102.300 86.330 102.750 ;
        RECT 79.580 102.150 89.880 102.300 ;
        RECT 83.530 101.200 85.930 102.150 ;
        RECT 90.480 101.600 90.630 109.800 ;
        RECT 91.080 101.600 91.230 109.800 ;
        RECT 91.680 101.600 91.830 109.800 ;
        RECT 92.280 101.600 92.430 109.800 ;
        RECT 92.880 101.600 93.030 109.800 ;
        RECT 93.480 101.600 93.630 109.800 ;
        RECT 94.080 101.600 94.230 109.800 ;
        RECT 95.230 110.200 95.380 118.400 ;
        RECT 95.830 110.200 95.980 118.400 ;
        RECT 96.430 110.200 96.580 118.400 ;
        RECT 97.030 110.200 97.180 118.400 ;
        RECT 97.630 110.200 97.780 118.400 ;
        RECT 98.230 110.200 98.380 118.400 ;
        RECT 98.830 110.200 98.980 118.400 ;
        RECT 103.530 117.850 105.940 118.800 ;
        RECT 99.580 117.700 109.880 117.850 ;
        RECT 103.130 117.250 106.330 117.700 ;
        RECT 99.580 117.100 109.880 117.250 ;
        RECT 103.130 116.650 106.330 117.100 ;
        RECT 99.580 116.500 109.880 116.650 ;
        RECT 103.130 116.050 106.330 116.500 ;
        RECT 99.580 115.900 109.880 116.050 ;
        RECT 103.130 115.600 106.330 115.900 ;
        RECT 103.130 115.450 103.530 115.600 ;
        RECT 99.580 115.300 103.530 115.450 ;
        RECT 103.130 114.850 103.530 115.300 ;
        RECT 99.580 114.700 103.530 114.850 ;
        RECT 103.130 114.250 103.530 114.700 ;
        RECT 99.580 114.100 103.530 114.250 ;
        RECT 103.130 113.650 103.530 114.100 ;
        RECT 99.580 113.500 103.530 113.650 ;
        RECT 103.130 113.050 103.530 113.500 ;
        RECT 99.580 112.900 103.530 113.050 ;
        RECT 103.130 112.450 103.530 112.900 ;
        RECT 99.580 112.300 103.530 112.450 ;
        RECT 103.130 111.850 103.530 112.300 ;
        RECT 99.580 111.700 103.530 111.850 ;
        RECT 103.130 111.250 103.530 111.700 ;
        RECT 99.580 111.100 103.530 111.250 ;
        RECT 103.130 110.650 103.530 111.100 ;
        RECT 99.580 110.500 103.530 110.650 ;
        RECT 103.130 110.200 103.530 110.500 ;
        RECT 95.230 109.800 103.530 110.200 ;
        RECT 95.230 101.600 95.380 109.800 ;
        RECT 95.830 101.600 95.980 109.800 ;
        RECT 96.430 101.600 96.580 109.800 ;
        RECT 97.030 101.600 97.180 109.800 ;
        RECT 97.630 101.600 97.780 109.800 ;
        RECT 98.230 101.600 98.380 109.800 ;
        RECT 98.830 101.600 98.980 109.800 ;
        RECT 103.130 109.500 103.530 109.800 ;
        RECT 99.580 109.350 103.530 109.500 ;
        RECT 103.130 108.900 103.530 109.350 ;
        RECT 99.580 108.750 103.530 108.900 ;
        RECT 103.130 108.300 103.530 108.750 ;
        RECT 99.580 108.150 103.530 108.300 ;
        RECT 103.130 107.700 103.530 108.150 ;
        RECT 99.580 107.550 103.530 107.700 ;
        RECT 103.130 107.100 103.530 107.550 ;
        RECT 99.580 106.950 103.530 107.100 ;
        RECT 103.130 106.500 103.530 106.950 ;
        RECT 99.580 106.350 103.530 106.500 ;
        RECT 103.130 105.900 103.530 106.350 ;
        RECT 99.580 105.750 103.530 105.900 ;
        RECT 103.130 105.300 103.530 105.750 ;
        RECT 99.580 105.150 103.530 105.300 ;
        RECT 103.130 104.700 103.530 105.150 ;
        RECT 99.580 104.550 103.530 104.700 ;
        RECT 103.130 104.400 103.530 104.550 ;
        RECT 105.930 115.450 106.330 115.600 ;
        RECT 105.930 115.300 109.880 115.450 ;
        RECT 105.930 114.850 106.330 115.300 ;
        RECT 105.930 114.700 109.880 114.850 ;
        RECT 105.930 114.250 106.330 114.700 ;
        RECT 105.930 114.100 109.880 114.250 ;
        RECT 105.930 113.650 106.330 114.100 ;
        RECT 105.930 113.500 109.880 113.650 ;
        RECT 105.930 113.050 106.330 113.500 ;
        RECT 105.930 112.900 109.880 113.050 ;
        RECT 105.930 112.450 106.330 112.900 ;
        RECT 105.930 112.300 109.880 112.450 ;
        RECT 105.930 111.850 106.330 112.300 ;
        RECT 105.930 111.700 109.880 111.850 ;
        RECT 105.930 111.250 106.330 111.700 ;
        RECT 105.930 111.100 109.880 111.250 ;
        RECT 105.930 110.650 106.330 111.100 ;
        RECT 105.930 110.500 109.880 110.650 ;
        RECT 105.930 110.200 106.330 110.500 ;
        RECT 110.480 110.200 110.630 118.400 ;
        RECT 111.080 110.200 111.230 118.400 ;
        RECT 111.680 110.200 111.830 118.400 ;
        RECT 112.280 110.200 112.430 118.400 ;
        RECT 112.880 110.200 113.030 118.400 ;
        RECT 113.480 110.200 113.630 118.400 ;
        RECT 114.080 110.200 114.230 118.400 ;
        RECT 105.930 109.800 114.230 110.200 ;
        RECT 105.930 109.500 106.330 109.800 ;
        RECT 105.930 109.350 109.880 109.500 ;
        RECT 105.930 108.900 106.330 109.350 ;
        RECT 105.930 108.750 109.880 108.900 ;
        RECT 105.930 108.300 106.330 108.750 ;
        RECT 105.930 108.150 109.880 108.300 ;
        RECT 105.930 107.700 106.330 108.150 ;
        RECT 105.930 107.550 109.880 107.700 ;
        RECT 105.930 107.100 106.330 107.550 ;
        RECT 105.930 106.950 109.880 107.100 ;
        RECT 105.930 106.500 106.330 106.950 ;
        RECT 105.930 106.350 109.880 106.500 ;
        RECT 105.930 105.900 106.330 106.350 ;
        RECT 105.930 105.750 109.880 105.900 ;
        RECT 105.930 105.300 106.330 105.750 ;
        RECT 105.930 105.150 109.880 105.300 ;
        RECT 105.930 104.700 106.330 105.150 ;
        RECT 105.930 104.550 109.880 104.700 ;
        RECT 105.930 104.400 106.330 104.550 ;
        RECT 103.130 104.100 106.330 104.400 ;
        RECT 99.580 103.950 109.880 104.100 ;
        RECT 103.130 103.500 106.330 103.950 ;
        RECT 99.580 103.350 109.880 103.500 ;
        RECT 103.130 102.900 106.330 103.350 ;
        RECT 99.580 102.750 109.880 102.900 ;
        RECT 103.130 102.300 106.330 102.750 ;
        RECT 99.580 102.150 109.880 102.300 ;
        RECT 103.530 101.200 105.930 102.150 ;
        RECT 110.480 101.600 110.630 109.800 ;
        RECT 111.080 101.600 111.230 109.800 ;
        RECT 111.680 101.600 111.830 109.800 ;
        RECT 112.280 101.600 112.430 109.800 ;
        RECT 112.880 101.600 113.030 109.800 ;
        RECT 113.480 101.600 113.630 109.800 ;
        RECT 114.080 101.600 114.230 109.800 ;
        RECT 115.230 110.200 115.380 118.400 ;
        RECT 115.830 110.200 115.980 118.400 ;
        RECT 116.430 110.200 116.580 118.400 ;
        RECT 117.030 110.200 117.180 118.400 ;
        RECT 117.630 110.200 117.780 118.400 ;
        RECT 118.230 110.200 118.380 118.400 ;
        RECT 118.830 110.200 118.980 118.400 ;
        RECT 123.530 117.850 124.730 118.800 ;
        RECT 119.580 117.700 124.730 117.850 ;
        RECT 123.130 117.250 124.730 117.700 ;
        RECT 119.580 117.100 124.730 117.250 ;
        RECT 123.130 116.650 124.730 117.100 ;
        RECT 119.580 116.500 124.730 116.650 ;
        RECT 123.130 116.050 124.730 116.500 ;
        RECT 125.135 116.060 127.135 117.335 ;
        RECT 119.580 115.900 124.730 116.050 ;
        RECT 123.130 115.600 124.730 115.900 ;
        RECT 123.130 115.450 123.530 115.600 ;
        RECT 119.580 115.300 123.530 115.450 ;
        RECT 123.130 114.850 123.530 115.300 ;
        RECT 119.580 114.700 123.530 114.850 ;
        RECT 123.130 114.250 123.530 114.700 ;
        RECT 119.580 114.100 123.530 114.250 ;
        RECT 123.130 113.650 123.530 114.100 ;
        RECT 119.580 113.500 123.530 113.650 ;
        RECT 123.130 113.050 123.530 113.500 ;
        RECT 119.580 112.900 123.530 113.050 ;
        RECT 123.130 112.450 123.530 112.900 ;
        RECT 119.580 112.300 123.530 112.450 ;
        RECT 123.130 111.850 123.530 112.300 ;
        RECT 119.580 111.700 123.530 111.850 ;
        RECT 123.130 111.250 123.530 111.700 ;
        RECT 119.580 111.100 123.530 111.250 ;
        RECT 123.130 110.650 123.530 111.100 ;
        RECT 119.580 110.500 123.530 110.650 ;
        RECT 123.130 110.200 123.530 110.500 ;
        RECT 115.230 109.800 123.530 110.200 ;
        RECT 115.230 101.600 115.380 109.800 ;
        RECT 115.830 101.600 115.980 109.800 ;
        RECT 116.430 101.600 116.580 109.800 ;
        RECT 117.030 101.600 117.180 109.800 ;
        RECT 117.630 101.600 117.780 109.800 ;
        RECT 118.230 101.600 118.380 109.800 ;
        RECT 118.830 101.600 118.980 109.800 ;
        RECT 123.130 109.500 123.530 109.800 ;
        RECT 119.580 109.350 123.530 109.500 ;
        RECT 123.130 108.900 123.530 109.350 ;
        RECT 119.580 108.750 123.530 108.900 ;
        RECT 123.130 108.300 123.530 108.750 ;
        RECT 119.580 108.150 123.530 108.300 ;
        RECT 123.130 107.700 123.530 108.150 ;
        RECT 119.580 107.550 123.530 107.700 ;
        RECT 123.130 107.100 123.530 107.550 ;
        RECT 119.580 106.950 123.530 107.100 ;
        RECT 123.130 106.500 123.530 106.950 ;
        RECT 119.580 106.350 123.530 106.500 ;
        RECT 123.130 105.900 123.530 106.350 ;
        RECT 119.580 105.750 123.530 105.900 ;
        RECT 123.130 105.300 123.530 105.750 ;
        RECT 119.580 105.150 123.530 105.300 ;
        RECT 123.130 104.700 123.530 105.150 ;
        RECT 119.580 104.550 123.530 104.700 ;
        RECT 123.130 104.400 123.530 104.550 ;
        RECT 123.130 104.100 124.730 104.400 ;
        RECT 119.580 103.950 124.730 104.100 ;
        RECT 123.130 103.500 124.730 103.950 ;
        RECT 119.580 103.350 124.730 103.500 ;
        RECT 123.130 102.900 124.730 103.350 ;
        RECT 119.580 102.750 124.730 102.900 ;
        RECT 123.130 102.300 124.730 102.750 ;
        RECT 119.580 102.150 124.730 102.300 ;
        RECT 123.530 101.200 124.730 102.150 ;
        RECT 125.140 101.845 127.140 103.120 ;
        RECT 4.730 98.800 9.130 101.200 ;
        RECT 20.330 98.800 29.130 101.200 ;
        RECT 40.330 98.800 49.130 101.200 ;
        RECT 60.330 98.800 69.130 101.200 ;
        RECT 80.330 98.800 89.130 101.200 ;
        RECT 100.330 98.800 109.130 101.200 ;
        RECT 120.330 98.800 124.730 101.200 ;
        RECT 4.730 97.850 5.940 98.800 ;
        RECT 2.315 96.570 4.320 97.845 ;
        RECT 4.730 97.700 9.880 97.850 ;
        RECT 4.730 97.250 6.330 97.700 ;
        RECT 4.730 97.100 9.880 97.250 ;
        RECT 4.730 96.650 6.330 97.100 ;
        RECT 4.730 96.500 9.880 96.650 ;
        RECT 4.730 96.050 6.330 96.500 ;
        RECT 4.730 95.900 9.880 96.050 ;
        RECT 4.730 95.600 6.330 95.900 ;
        RECT 2.315 93.250 4.315 95.545 ;
        RECT 5.930 95.450 6.330 95.600 ;
        RECT 5.930 95.300 9.880 95.450 ;
        RECT 5.930 94.850 6.330 95.300 ;
        RECT 5.930 94.700 9.880 94.850 ;
        RECT 5.930 94.250 6.330 94.700 ;
        RECT 5.930 94.100 9.880 94.250 ;
        RECT 5.930 93.650 6.330 94.100 ;
        RECT 5.930 93.500 9.880 93.650 ;
        RECT 5.930 93.050 6.330 93.500 ;
        RECT 5.930 92.900 9.880 93.050 ;
        RECT 5.930 92.450 6.330 92.900 ;
        RECT 5.930 92.300 9.880 92.450 ;
        RECT 5.930 91.850 6.330 92.300 ;
        RECT 5.930 91.700 9.880 91.850 ;
        RECT 5.930 91.250 6.330 91.700 ;
        RECT 5.930 91.100 9.880 91.250 ;
        RECT 5.930 90.650 6.330 91.100 ;
        RECT 5.930 90.500 9.880 90.650 ;
        RECT 5.930 90.200 6.330 90.500 ;
        RECT 10.480 90.200 10.630 98.400 ;
        RECT 11.080 90.200 11.230 98.400 ;
        RECT 11.680 90.200 11.830 98.400 ;
        RECT 12.280 90.200 12.430 98.400 ;
        RECT 12.880 90.200 13.030 98.400 ;
        RECT 13.480 90.200 13.630 98.400 ;
        RECT 14.080 90.200 14.230 98.400 ;
        RECT 5.930 89.800 14.230 90.200 ;
        RECT 5.930 89.500 6.330 89.800 ;
        RECT 5.930 89.350 9.880 89.500 ;
        RECT 5.930 88.900 6.330 89.350 ;
        RECT 5.930 88.750 9.880 88.900 ;
        RECT 5.930 88.300 6.330 88.750 ;
        RECT 5.930 88.150 9.880 88.300 ;
        RECT 5.930 87.700 6.330 88.150 ;
        RECT 5.930 87.550 9.880 87.700 ;
        RECT 5.930 87.100 6.330 87.550 ;
        RECT 5.930 86.950 9.880 87.100 ;
        RECT 2.315 84.455 4.315 86.750 ;
        RECT 5.930 86.500 6.330 86.950 ;
        RECT 5.930 86.350 9.880 86.500 ;
        RECT 5.930 85.900 6.330 86.350 ;
        RECT 5.930 85.750 9.880 85.900 ;
        RECT 5.930 85.300 6.330 85.750 ;
        RECT 5.930 85.150 9.880 85.300 ;
        RECT 5.930 84.700 6.330 85.150 ;
        RECT 5.930 84.550 9.880 84.700 ;
        RECT 5.930 84.400 6.330 84.550 ;
        RECT 4.730 84.100 6.330 84.400 ;
        RECT 4.730 83.950 9.880 84.100 ;
        RECT 4.730 83.500 6.330 83.950 ;
        RECT 2.315 82.195 4.320 83.470 ;
        RECT 4.730 83.350 9.880 83.500 ;
        RECT 4.730 82.900 6.330 83.350 ;
        RECT 4.730 82.750 9.880 82.900 ;
        RECT 4.730 82.300 6.330 82.750 ;
        RECT 4.730 82.150 9.880 82.300 ;
        RECT 4.730 81.200 5.930 82.150 ;
        RECT 10.480 81.600 10.630 89.800 ;
        RECT 11.080 81.600 11.230 89.800 ;
        RECT 11.680 81.600 11.830 89.800 ;
        RECT 12.280 81.600 12.430 89.800 ;
        RECT 12.880 81.600 13.030 89.800 ;
        RECT 13.480 81.600 13.630 89.800 ;
        RECT 14.080 81.600 14.230 89.800 ;
        RECT 15.230 90.200 15.380 98.400 ;
        RECT 15.830 90.200 15.980 98.400 ;
        RECT 16.430 90.200 16.580 98.400 ;
        RECT 17.030 90.200 17.180 98.400 ;
        RECT 17.630 90.200 17.780 98.400 ;
        RECT 18.230 90.200 18.380 98.400 ;
        RECT 18.830 90.200 18.980 98.400 ;
        RECT 23.530 97.850 25.940 98.800 ;
        RECT 19.580 97.700 29.880 97.850 ;
        RECT 23.130 97.250 26.330 97.700 ;
        RECT 19.580 97.100 29.880 97.250 ;
        RECT 23.130 96.650 26.330 97.100 ;
        RECT 19.580 96.500 29.880 96.650 ;
        RECT 23.130 96.050 26.330 96.500 ;
        RECT 19.580 95.900 29.880 96.050 ;
        RECT 23.130 95.600 26.330 95.900 ;
        RECT 23.130 95.450 23.530 95.600 ;
        RECT 19.580 95.300 23.530 95.450 ;
        RECT 23.130 94.850 23.530 95.300 ;
        RECT 19.580 94.700 23.530 94.850 ;
        RECT 23.130 94.250 23.530 94.700 ;
        RECT 19.580 94.100 23.530 94.250 ;
        RECT 23.130 93.650 23.530 94.100 ;
        RECT 19.580 93.500 23.530 93.650 ;
        RECT 23.130 93.050 23.530 93.500 ;
        RECT 19.580 92.900 23.530 93.050 ;
        RECT 23.130 92.450 23.530 92.900 ;
        RECT 19.580 92.300 23.530 92.450 ;
        RECT 23.130 91.850 23.530 92.300 ;
        RECT 19.580 91.700 23.530 91.850 ;
        RECT 23.130 91.250 23.530 91.700 ;
        RECT 19.580 91.100 23.530 91.250 ;
        RECT 23.130 90.650 23.530 91.100 ;
        RECT 19.580 90.500 23.530 90.650 ;
        RECT 23.130 90.200 23.530 90.500 ;
        RECT 15.230 89.800 23.530 90.200 ;
        RECT 15.230 81.600 15.380 89.800 ;
        RECT 15.830 81.600 15.980 89.800 ;
        RECT 16.430 81.600 16.580 89.800 ;
        RECT 17.030 81.600 17.180 89.800 ;
        RECT 17.630 81.600 17.780 89.800 ;
        RECT 18.230 81.600 18.380 89.800 ;
        RECT 18.830 81.600 18.980 89.800 ;
        RECT 23.130 89.500 23.530 89.800 ;
        RECT 19.580 89.350 23.530 89.500 ;
        RECT 23.130 88.900 23.530 89.350 ;
        RECT 19.580 88.750 23.530 88.900 ;
        RECT 23.130 88.300 23.530 88.750 ;
        RECT 19.580 88.150 23.530 88.300 ;
        RECT 23.130 87.700 23.530 88.150 ;
        RECT 19.580 87.550 23.530 87.700 ;
        RECT 23.130 87.100 23.530 87.550 ;
        RECT 19.580 86.950 23.530 87.100 ;
        RECT 23.130 86.500 23.530 86.950 ;
        RECT 19.580 86.350 23.530 86.500 ;
        RECT 23.130 85.900 23.530 86.350 ;
        RECT 19.580 85.750 23.530 85.900 ;
        RECT 23.130 85.300 23.530 85.750 ;
        RECT 19.580 85.150 23.530 85.300 ;
        RECT 23.130 84.700 23.530 85.150 ;
        RECT 19.580 84.550 23.530 84.700 ;
        RECT 23.130 84.400 23.530 84.550 ;
        RECT 25.930 95.450 26.330 95.600 ;
        RECT 25.930 95.300 29.880 95.450 ;
        RECT 25.930 94.850 26.330 95.300 ;
        RECT 25.930 94.700 29.880 94.850 ;
        RECT 25.930 94.250 26.330 94.700 ;
        RECT 25.930 94.100 29.880 94.250 ;
        RECT 25.930 93.650 26.330 94.100 ;
        RECT 25.930 93.500 29.880 93.650 ;
        RECT 25.930 93.050 26.330 93.500 ;
        RECT 25.930 92.900 29.880 93.050 ;
        RECT 25.930 92.450 26.330 92.900 ;
        RECT 25.930 92.300 29.880 92.450 ;
        RECT 25.930 91.850 26.330 92.300 ;
        RECT 25.930 91.700 29.880 91.850 ;
        RECT 25.930 91.250 26.330 91.700 ;
        RECT 25.930 91.100 29.880 91.250 ;
        RECT 25.930 90.650 26.330 91.100 ;
        RECT 25.930 90.500 29.880 90.650 ;
        RECT 25.930 90.200 26.330 90.500 ;
        RECT 30.480 90.200 30.630 98.400 ;
        RECT 31.080 90.200 31.230 98.400 ;
        RECT 31.680 90.200 31.830 98.400 ;
        RECT 32.280 90.200 32.430 98.400 ;
        RECT 32.880 90.200 33.030 98.400 ;
        RECT 33.480 90.200 33.630 98.400 ;
        RECT 34.080 90.200 34.230 98.400 ;
        RECT 25.930 89.800 34.230 90.200 ;
        RECT 25.930 89.500 26.330 89.800 ;
        RECT 25.930 89.350 29.880 89.500 ;
        RECT 25.930 88.900 26.330 89.350 ;
        RECT 25.930 88.750 29.880 88.900 ;
        RECT 25.930 88.300 26.330 88.750 ;
        RECT 25.930 88.150 29.880 88.300 ;
        RECT 25.930 87.700 26.330 88.150 ;
        RECT 25.930 87.550 29.880 87.700 ;
        RECT 25.930 87.100 26.330 87.550 ;
        RECT 25.930 86.950 29.880 87.100 ;
        RECT 25.930 86.500 26.330 86.950 ;
        RECT 25.930 86.350 29.880 86.500 ;
        RECT 25.930 85.900 26.330 86.350 ;
        RECT 25.930 85.750 29.880 85.900 ;
        RECT 25.930 85.300 26.330 85.750 ;
        RECT 25.930 85.150 29.880 85.300 ;
        RECT 25.930 84.700 26.330 85.150 ;
        RECT 25.930 84.550 29.880 84.700 ;
        RECT 25.930 84.400 26.330 84.550 ;
        RECT 23.130 84.100 26.330 84.400 ;
        RECT 19.580 83.950 29.880 84.100 ;
        RECT 23.130 83.500 26.330 83.950 ;
        RECT 19.580 83.350 29.880 83.500 ;
        RECT 23.130 82.900 26.330 83.350 ;
        RECT 19.580 82.750 29.880 82.900 ;
        RECT 23.130 82.300 26.330 82.750 ;
        RECT 19.580 82.150 29.880 82.300 ;
        RECT 23.530 81.200 25.930 82.150 ;
        RECT 30.480 81.600 30.630 89.800 ;
        RECT 31.080 81.600 31.230 89.800 ;
        RECT 31.680 81.600 31.830 89.800 ;
        RECT 32.280 81.600 32.430 89.800 ;
        RECT 32.880 81.600 33.030 89.800 ;
        RECT 33.480 81.600 33.630 89.800 ;
        RECT 34.080 81.600 34.230 89.800 ;
        RECT 35.230 90.200 35.380 98.400 ;
        RECT 35.830 90.200 35.980 98.400 ;
        RECT 36.430 90.200 36.580 98.400 ;
        RECT 37.030 90.200 37.180 98.400 ;
        RECT 37.630 90.200 37.780 98.400 ;
        RECT 38.230 90.200 38.380 98.400 ;
        RECT 38.830 90.200 38.980 98.400 ;
        RECT 43.530 97.850 45.940 98.800 ;
        RECT 39.580 97.700 49.880 97.850 ;
        RECT 43.130 97.250 46.330 97.700 ;
        RECT 39.580 97.100 49.880 97.250 ;
        RECT 43.130 96.650 46.330 97.100 ;
        RECT 39.580 96.500 49.880 96.650 ;
        RECT 43.130 96.050 46.330 96.500 ;
        RECT 39.580 95.900 49.880 96.050 ;
        RECT 43.130 95.600 46.330 95.900 ;
        RECT 43.130 95.450 43.530 95.600 ;
        RECT 39.580 95.300 43.530 95.450 ;
        RECT 43.130 94.850 43.530 95.300 ;
        RECT 39.580 94.700 43.530 94.850 ;
        RECT 43.130 94.250 43.530 94.700 ;
        RECT 39.580 94.100 43.530 94.250 ;
        RECT 43.130 93.650 43.530 94.100 ;
        RECT 39.580 93.500 43.530 93.650 ;
        RECT 43.130 93.050 43.530 93.500 ;
        RECT 39.580 92.900 43.530 93.050 ;
        RECT 43.130 92.450 43.530 92.900 ;
        RECT 39.580 92.300 43.530 92.450 ;
        RECT 43.130 91.850 43.530 92.300 ;
        RECT 39.580 91.700 43.530 91.850 ;
        RECT 43.130 91.250 43.530 91.700 ;
        RECT 39.580 91.100 43.530 91.250 ;
        RECT 43.130 90.650 43.530 91.100 ;
        RECT 39.580 90.500 43.530 90.650 ;
        RECT 43.130 90.200 43.530 90.500 ;
        RECT 35.230 89.800 43.530 90.200 ;
        RECT 35.230 81.600 35.380 89.800 ;
        RECT 35.830 81.600 35.980 89.800 ;
        RECT 36.430 81.600 36.580 89.800 ;
        RECT 37.030 81.600 37.180 89.800 ;
        RECT 37.630 81.600 37.780 89.800 ;
        RECT 38.230 81.600 38.380 89.800 ;
        RECT 38.830 81.600 38.980 89.800 ;
        RECT 43.130 89.500 43.530 89.800 ;
        RECT 39.580 89.350 43.530 89.500 ;
        RECT 43.130 88.900 43.530 89.350 ;
        RECT 39.580 88.750 43.530 88.900 ;
        RECT 43.130 88.300 43.530 88.750 ;
        RECT 39.580 88.150 43.530 88.300 ;
        RECT 43.130 87.700 43.530 88.150 ;
        RECT 39.580 87.550 43.530 87.700 ;
        RECT 43.130 87.100 43.530 87.550 ;
        RECT 39.580 86.950 43.530 87.100 ;
        RECT 43.130 86.500 43.530 86.950 ;
        RECT 39.580 86.350 43.530 86.500 ;
        RECT 43.130 85.900 43.530 86.350 ;
        RECT 39.580 85.750 43.530 85.900 ;
        RECT 43.130 85.300 43.530 85.750 ;
        RECT 39.580 85.150 43.530 85.300 ;
        RECT 43.130 84.700 43.530 85.150 ;
        RECT 39.580 84.550 43.530 84.700 ;
        RECT 43.130 84.400 43.530 84.550 ;
        RECT 45.930 95.450 46.330 95.600 ;
        RECT 45.930 95.300 49.880 95.450 ;
        RECT 45.930 94.850 46.330 95.300 ;
        RECT 45.930 94.700 49.880 94.850 ;
        RECT 45.930 94.250 46.330 94.700 ;
        RECT 45.930 94.100 49.880 94.250 ;
        RECT 45.930 93.650 46.330 94.100 ;
        RECT 45.930 93.500 49.880 93.650 ;
        RECT 45.930 93.050 46.330 93.500 ;
        RECT 45.930 92.900 49.880 93.050 ;
        RECT 45.930 92.450 46.330 92.900 ;
        RECT 45.930 92.300 49.880 92.450 ;
        RECT 45.930 91.850 46.330 92.300 ;
        RECT 45.930 91.700 49.880 91.850 ;
        RECT 45.930 91.250 46.330 91.700 ;
        RECT 45.930 91.100 49.880 91.250 ;
        RECT 45.930 90.650 46.330 91.100 ;
        RECT 45.930 90.500 49.880 90.650 ;
        RECT 45.930 90.200 46.330 90.500 ;
        RECT 50.480 90.200 50.630 98.400 ;
        RECT 51.080 90.200 51.230 98.400 ;
        RECT 51.680 90.200 51.830 98.400 ;
        RECT 52.280 90.200 52.430 98.400 ;
        RECT 52.880 90.200 53.030 98.400 ;
        RECT 53.480 90.200 53.630 98.400 ;
        RECT 54.080 90.200 54.230 98.400 ;
        RECT 45.930 89.800 54.230 90.200 ;
        RECT 45.930 89.500 46.330 89.800 ;
        RECT 45.930 89.350 49.880 89.500 ;
        RECT 45.930 88.900 46.330 89.350 ;
        RECT 45.930 88.750 49.880 88.900 ;
        RECT 45.930 88.300 46.330 88.750 ;
        RECT 45.930 88.150 49.880 88.300 ;
        RECT 45.930 87.700 46.330 88.150 ;
        RECT 45.930 87.550 49.880 87.700 ;
        RECT 45.930 87.100 46.330 87.550 ;
        RECT 45.930 86.950 49.880 87.100 ;
        RECT 45.930 86.500 46.330 86.950 ;
        RECT 45.930 86.350 49.880 86.500 ;
        RECT 45.930 85.900 46.330 86.350 ;
        RECT 45.930 85.750 49.880 85.900 ;
        RECT 45.930 85.300 46.330 85.750 ;
        RECT 45.930 85.150 49.880 85.300 ;
        RECT 45.930 84.700 46.330 85.150 ;
        RECT 45.930 84.550 49.880 84.700 ;
        RECT 45.930 84.400 46.330 84.550 ;
        RECT 43.130 84.100 46.330 84.400 ;
        RECT 39.580 83.950 49.880 84.100 ;
        RECT 43.130 83.500 46.330 83.950 ;
        RECT 39.580 83.350 49.880 83.500 ;
        RECT 43.130 82.900 46.330 83.350 ;
        RECT 39.580 82.750 49.880 82.900 ;
        RECT 43.130 82.300 46.330 82.750 ;
        RECT 39.580 82.150 49.880 82.300 ;
        RECT 43.530 81.200 45.930 82.150 ;
        RECT 50.480 81.600 50.630 89.800 ;
        RECT 51.080 81.600 51.230 89.800 ;
        RECT 51.680 81.600 51.830 89.800 ;
        RECT 52.280 81.600 52.430 89.800 ;
        RECT 52.880 81.600 53.030 89.800 ;
        RECT 53.480 81.600 53.630 89.800 ;
        RECT 54.080 81.600 54.230 89.800 ;
        RECT 55.230 90.200 55.380 98.400 ;
        RECT 55.830 90.200 55.980 98.400 ;
        RECT 56.430 90.200 56.580 98.400 ;
        RECT 57.030 90.200 57.180 98.400 ;
        RECT 57.630 90.200 57.780 98.400 ;
        RECT 58.230 90.200 58.380 98.400 ;
        RECT 58.830 90.200 58.980 98.400 ;
        RECT 63.530 97.850 65.940 98.800 ;
        RECT 59.580 97.700 69.880 97.850 ;
        RECT 63.130 97.250 66.330 97.700 ;
        RECT 59.580 97.100 69.880 97.250 ;
        RECT 63.130 96.650 66.330 97.100 ;
        RECT 59.580 96.500 69.880 96.650 ;
        RECT 63.130 96.050 66.330 96.500 ;
        RECT 59.580 95.900 69.880 96.050 ;
        RECT 63.130 95.600 66.330 95.900 ;
        RECT 63.130 95.450 63.530 95.600 ;
        RECT 59.580 95.300 63.530 95.450 ;
        RECT 63.130 94.850 63.530 95.300 ;
        RECT 59.580 94.700 63.530 94.850 ;
        RECT 63.130 94.250 63.530 94.700 ;
        RECT 59.580 94.100 63.530 94.250 ;
        RECT 63.130 93.650 63.530 94.100 ;
        RECT 59.580 93.500 63.530 93.650 ;
        RECT 63.130 93.050 63.530 93.500 ;
        RECT 59.580 92.900 63.530 93.050 ;
        RECT 63.130 92.450 63.530 92.900 ;
        RECT 59.580 92.300 63.530 92.450 ;
        RECT 63.130 91.850 63.530 92.300 ;
        RECT 59.580 91.700 63.530 91.850 ;
        RECT 63.130 91.250 63.530 91.700 ;
        RECT 59.580 91.100 63.530 91.250 ;
        RECT 63.130 90.650 63.530 91.100 ;
        RECT 59.580 90.500 63.530 90.650 ;
        RECT 63.130 90.200 63.530 90.500 ;
        RECT 55.230 89.800 63.530 90.200 ;
        RECT 55.230 81.600 55.380 89.800 ;
        RECT 55.830 81.600 55.980 89.800 ;
        RECT 56.430 81.600 56.580 89.800 ;
        RECT 57.030 81.600 57.180 89.800 ;
        RECT 57.630 81.600 57.780 89.800 ;
        RECT 58.230 81.600 58.380 89.800 ;
        RECT 58.830 81.600 58.980 89.800 ;
        RECT 63.130 89.500 63.530 89.800 ;
        RECT 59.580 89.350 63.530 89.500 ;
        RECT 63.130 88.900 63.530 89.350 ;
        RECT 59.580 88.750 63.530 88.900 ;
        RECT 63.130 88.300 63.530 88.750 ;
        RECT 59.580 88.150 63.530 88.300 ;
        RECT 63.130 87.700 63.530 88.150 ;
        RECT 59.580 87.550 63.530 87.700 ;
        RECT 63.130 87.100 63.530 87.550 ;
        RECT 59.580 86.950 63.530 87.100 ;
        RECT 63.130 86.500 63.530 86.950 ;
        RECT 59.580 86.350 63.530 86.500 ;
        RECT 63.130 85.900 63.530 86.350 ;
        RECT 59.580 85.750 63.530 85.900 ;
        RECT 63.130 85.300 63.530 85.750 ;
        RECT 59.580 85.150 63.530 85.300 ;
        RECT 63.130 84.700 63.530 85.150 ;
        RECT 59.580 84.550 63.530 84.700 ;
        RECT 63.130 84.400 63.530 84.550 ;
        RECT 65.930 95.450 66.330 95.600 ;
        RECT 65.930 95.300 69.880 95.450 ;
        RECT 65.930 94.850 66.330 95.300 ;
        RECT 65.930 94.700 69.880 94.850 ;
        RECT 65.930 94.250 66.330 94.700 ;
        RECT 65.930 94.100 69.880 94.250 ;
        RECT 65.930 93.650 66.330 94.100 ;
        RECT 65.930 93.500 69.880 93.650 ;
        RECT 65.930 93.050 66.330 93.500 ;
        RECT 65.930 92.900 69.880 93.050 ;
        RECT 65.930 92.450 66.330 92.900 ;
        RECT 65.930 92.300 69.880 92.450 ;
        RECT 65.930 91.850 66.330 92.300 ;
        RECT 65.930 91.700 69.880 91.850 ;
        RECT 65.930 91.250 66.330 91.700 ;
        RECT 65.930 91.100 69.880 91.250 ;
        RECT 65.930 90.650 66.330 91.100 ;
        RECT 65.930 90.500 69.880 90.650 ;
        RECT 65.930 90.200 66.330 90.500 ;
        RECT 70.480 90.200 70.630 98.400 ;
        RECT 71.080 90.200 71.230 98.400 ;
        RECT 71.680 90.200 71.830 98.400 ;
        RECT 72.280 90.200 72.430 98.400 ;
        RECT 72.880 90.200 73.030 98.400 ;
        RECT 73.480 90.200 73.630 98.400 ;
        RECT 74.080 90.200 74.230 98.400 ;
        RECT 65.930 89.800 74.230 90.200 ;
        RECT 65.930 89.500 66.330 89.800 ;
        RECT 65.930 89.350 69.880 89.500 ;
        RECT 65.930 88.900 66.330 89.350 ;
        RECT 65.930 88.750 69.880 88.900 ;
        RECT 65.930 88.300 66.330 88.750 ;
        RECT 65.930 88.150 69.880 88.300 ;
        RECT 65.930 87.700 66.330 88.150 ;
        RECT 65.930 87.550 69.880 87.700 ;
        RECT 65.930 87.100 66.330 87.550 ;
        RECT 65.930 86.950 69.880 87.100 ;
        RECT 65.930 86.500 66.330 86.950 ;
        RECT 65.930 86.350 69.880 86.500 ;
        RECT 65.930 85.900 66.330 86.350 ;
        RECT 65.930 85.750 69.880 85.900 ;
        RECT 65.930 85.300 66.330 85.750 ;
        RECT 65.930 85.150 69.880 85.300 ;
        RECT 65.930 84.700 66.330 85.150 ;
        RECT 65.930 84.550 69.880 84.700 ;
        RECT 65.930 84.400 66.330 84.550 ;
        RECT 63.130 84.100 66.330 84.400 ;
        RECT 59.580 83.950 69.880 84.100 ;
        RECT 63.130 83.500 66.330 83.950 ;
        RECT 59.580 83.350 69.880 83.500 ;
        RECT 63.130 82.900 66.330 83.350 ;
        RECT 59.580 82.750 69.880 82.900 ;
        RECT 63.130 82.300 66.330 82.750 ;
        RECT 59.580 82.150 69.880 82.300 ;
        RECT 63.530 81.200 65.930 82.150 ;
        RECT 70.480 81.600 70.630 89.800 ;
        RECT 71.080 81.600 71.230 89.800 ;
        RECT 71.680 81.600 71.830 89.800 ;
        RECT 72.280 81.600 72.430 89.800 ;
        RECT 72.880 81.600 73.030 89.800 ;
        RECT 73.480 81.600 73.630 89.800 ;
        RECT 74.080 81.600 74.230 89.800 ;
        RECT 75.230 90.200 75.380 98.400 ;
        RECT 75.830 90.200 75.980 98.400 ;
        RECT 76.430 90.200 76.580 98.400 ;
        RECT 77.030 90.200 77.180 98.400 ;
        RECT 77.630 90.200 77.780 98.400 ;
        RECT 78.230 90.200 78.380 98.400 ;
        RECT 78.830 90.200 78.980 98.400 ;
        RECT 83.530 97.850 85.940 98.800 ;
        RECT 79.580 97.700 89.880 97.850 ;
        RECT 83.130 97.250 86.330 97.700 ;
        RECT 79.580 97.100 89.880 97.250 ;
        RECT 83.130 96.650 86.330 97.100 ;
        RECT 79.580 96.500 89.880 96.650 ;
        RECT 83.130 96.050 86.330 96.500 ;
        RECT 79.580 95.900 89.880 96.050 ;
        RECT 83.130 95.600 86.330 95.900 ;
        RECT 83.130 95.450 83.530 95.600 ;
        RECT 79.580 95.300 83.530 95.450 ;
        RECT 83.130 94.850 83.530 95.300 ;
        RECT 79.580 94.700 83.530 94.850 ;
        RECT 83.130 94.250 83.530 94.700 ;
        RECT 79.580 94.100 83.530 94.250 ;
        RECT 83.130 93.650 83.530 94.100 ;
        RECT 79.580 93.500 83.530 93.650 ;
        RECT 83.130 93.050 83.530 93.500 ;
        RECT 79.580 92.900 83.530 93.050 ;
        RECT 83.130 92.450 83.530 92.900 ;
        RECT 79.580 92.300 83.530 92.450 ;
        RECT 83.130 91.850 83.530 92.300 ;
        RECT 79.580 91.700 83.530 91.850 ;
        RECT 83.130 91.250 83.530 91.700 ;
        RECT 79.580 91.100 83.530 91.250 ;
        RECT 83.130 90.650 83.530 91.100 ;
        RECT 79.580 90.500 83.530 90.650 ;
        RECT 83.130 90.200 83.530 90.500 ;
        RECT 75.230 89.800 83.530 90.200 ;
        RECT 75.230 81.600 75.380 89.800 ;
        RECT 75.830 81.600 75.980 89.800 ;
        RECT 76.430 81.600 76.580 89.800 ;
        RECT 77.030 81.600 77.180 89.800 ;
        RECT 77.630 81.600 77.780 89.800 ;
        RECT 78.230 81.600 78.380 89.800 ;
        RECT 78.830 81.600 78.980 89.800 ;
        RECT 83.130 89.500 83.530 89.800 ;
        RECT 79.580 89.350 83.530 89.500 ;
        RECT 83.130 88.900 83.530 89.350 ;
        RECT 79.580 88.750 83.530 88.900 ;
        RECT 83.130 88.300 83.530 88.750 ;
        RECT 79.580 88.150 83.530 88.300 ;
        RECT 83.130 87.700 83.530 88.150 ;
        RECT 79.580 87.550 83.530 87.700 ;
        RECT 83.130 87.100 83.530 87.550 ;
        RECT 79.580 86.950 83.530 87.100 ;
        RECT 83.130 86.500 83.530 86.950 ;
        RECT 79.580 86.350 83.530 86.500 ;
        RECT 83.130 85.900 83.530 86.350 ;
        RECT 79.580 85.750 83.530 85.900 ;
        RECT 83.130 85.300 83.530 85.750 ;
        RECT 79.580 85.150 83.530 85.300 ;
        RECT 83.130 84.700 83.530 85.150 ;
        RECT 79.580 84.550 83.530 84.700 ;
        RECT 83.130 84.400 83.530 84.550 ;
        RECT 85.930 95.450 86.330 95.600 ;
        RECT 85.930 95.300 89.880 95.450 ;
        RECT 85.930 94.850 86.330 95.300 ;
        RECT 85.930 94.700 89.880 94.850 ;
        RECT 85.930 94.250 86.330 94.700 ;
        RECT 85.930 94.100 89.880 94.250 ;
        RECT 85.930 93.650 86.330 94.100 ;
        RECT 85.930 93.500 89.880 93.650 ;
        RECT 85.930 93.050 86.330 93.500 ;
        RECT 85.930 92.900 89.880 93.050 ;
        RECT 85.930 92.450 86.330 92.900 ;
        RECT 85.930 92.300 89.880 92.450 ;
        RECT 85.930 91.850 86.330 92.300 ;
        RECT 85.930 91.700 89.880 91.850 ;
        RECT 85.930 91.250 86.330 91.700 ;
        RECT 85.930 91.100 89.880 91.250 ;
        RECT 85.930 90.650 86.330 91.100 ;
        RECT 85.930 90.500 89.880 90.650 ;
        RECT 85.930 90.200 86.330 90.500 ;
        RECT 90.480 90.200 90.630 98.400 ;
        RECT 91.080 90.200 91.230 98.400 ;
        RECT 91.680 90.200 91.830 98.400 ;
        RECT 92.280 90.200 92.430 98.400 ;
        RECT 92.880 90.200 93.030 98.400 ;
        RECT 93.480 90.200 93.630 98.400 ;
        RECT 94.080 90.200 94.230 98.400 ;
        RECT 85.930 89.800 94.230 90.200 ;
        RECT 85.930 89.500 86.330 89.800 ;
        RECT 85.930 89.350 89.880 89.500 ;
        RECT 85.930 88.900 86.330 89.350 ;
        RECT 85.930 88.750 89.880 88.900 ;
        RECT 85.930 88.300 86.330 88.750 ;
        RECT 85.930 88.150 89.880 88.300 ;
        RECT 85.930 87.700 86.330 88.150 ;
        RECT 85.930 87.550 89.880 87.700 ;
        RECT 85.930 87.100 86.330 87.550 ;
        RECT 85.930 86.950 89.880 87.100 ;
        RECT 85.930 86.500 86.330 86.950 ;
        RECT 85.930 86.350 89.880 86.500 ;
        RECT 85.930 85.900 86.330 86.350 ;
        RECT 85.930 85.750 89.880 85.900 ;
        RECT 85.930 85.300 86.330 85.750 ;
        RECT 85.930 85.150 89.880 85.300 ;
        RECT 85.930 84.700 86.330 85.150 ;
        RECT 85.930 84.550 89.880 84.700 ;
        RECT 85.930 84.400 86.330 84.550 ;
        RECT 83.130 84.100 86.330 84.400 ;
        RECT 79.580 83.950 89.880 84.100 ;
        RECT 83.130 83.500 86.330 83.950 ;
        RECT 79.580 83.350 89.880 83.500 ;
        RECT 83.130 82.900 86.330 83.350 ;
        RECT 79.580 82.750 89.880 82.900 ;
        RECT 83.130 82.300 86.330 82.750 ;
        RECT 79.580 82.150 89.880 82.300 ;
        RECT 83.530 81.200 85.930 82.150 ;
        RECT 90.480 81.600 90.630 89.800 ;
        RECT 91.080 81.600 91.230 89.800 ;
        RECT 91.680 81.600 91.830 89.800 ;
        RECT 92.280 81.600 92.430 89.800 ;
        RECT 92.880 81.600 93.030 89.800 ;
        RECT 93.480 81.600 93.630 89.800 ;
        RECT 94.080 81.600 94.230 89.800 ;
        RECT 95.230 90.200 95.380 98.400 ;
        RECT 95.830 90.200 95.980 98.400 ;
        RECT 96.430 90.200 96.580 98.400 ;
        RECT 97.030 90.200 97.180 98.400 ;
        RECT 97.630 90.200 97.780 98.400 ;
        RECT 98.230 90.200 98.380 98.400 ;
        RECT 98.830 90.200 98.980 98.400 ;
        RECT 103.530 97.850 105.940 98.800 ;
        RECT 99.580 97.700 109.880 97.850 ;
        RECT 103.130 97.250 106.330 97.700 ;
        RECT 99.580 97.100 109.880 97.250 ;
        RECT 103.130 96.650 106.330 97.100 ;
        RECT 99.580 96.500 109.880 96.650 ;
        RECT 103.130 96.050 106.330 96.500 ;
        RECT 99.580 95.900 109.880 96.050 ;
        RECT 103.130 95.600 106.330 95.900 ;
        RECT 103.130 95.450 103.530 95.600 ;
        RECT 99.580 95.300 103.530 95.450 ;
        RECT 103.130 94.850 103.530 95.300 ;
        RECT 99.580 94.700 103.530 94.850 ;
        RECT 103.130 94.250 103.530 94.700 ;
        RECT 99.580 94.100 103.530 94.250 ;
        RECT 103.130 93.650 103.530 94.100 ;
        RECT 99.580 93.500 103.530 93.650 ;
        RECT 103.130 93.050 103.530 93.500 ;
        RECT 99.580 92.900 103.530 93.050 ;
        RECT 103.130 92.450 103.530 92.900 ;
        RECT 99.580 92.300 103.530 92.450 ;
        RECT 103.130 91.850 103.530 92.300 ;
        RECT 99.580 91.700 103.530 91.850 ;
        RECT 103.130 91.250 103.530 91.700 ;
        RECT 99.580 91.100 103.530 91.250 ;
        RECT 103.130 90.650 103.530 91.100 ;
        RECT 99.580 90.500 103.530 90.650 ;
        RECT 103.130 90.200 103.530 90.500 ;
        RECT 95.230 89.800 103.530 90.200 ;
        RECT 95.230 81.600 95.380 89.800 ;
        RECT 95.830 81.600 95.980 89.800 ;
        RECT 96.430 81.600 96.580 89.800 ;
        RECT 97.030 81.600 97.180 89.800 ;
        RECT 97.630 81.600 97.780 89.800 ;
        RECT 98.230 81.600 98.380 89.800 ;
        RECT 98.830 81.600 98.980 89.800 ;
        RECT 103.130 89.500 103.530 89.800 ;
        RECT 99.580 89.350 103.530 89.500 ;
        RECT 103.130 88.900 103.530 89.350 ;
        RECT 99.580 88.750 103.530 88.900 ;
        RECT 103.130 88.300 103.530 88.750 ;
        RECT 99.580 88.150 103.530 88.300 ;
        RECT 103.130 87.700 103.530 88.150 ;
        RECT 99.580 87.550 103.530 87.700 ;
        RECT 103.130 87.100 103.530 87.550 ;
        RECT 99.580 86.950 103.530 87.100 ;
        RECT 103.130 86.500 103.530 86.950 ;
        RECT 99.580 86.350 103.530 86.500 ;
        RECT 103.130 85.900 103.530 86.350 ;
        RECT 99.580 85.750 103.530 85.900 ;
        RECT 103.130 85.300 103.530 85.750 ;
        RECT 99.580 85.150 103.530 85.300 ;
        RECT 103.130 84.700 103.530 85.150 ;
        RECT 99.580 84.550 103.530 84.700 ;
        RECT 103.130 84.400 103.530 84.550 ;
        RECT 105.930 95.450 106.330 95.600 ;
        RECT 105.930 95.300 109.880 95.450 ;
        RECT 105.930 94.850 106.330 95.300 ;
        RECT 105.930 94.700 109.880 94.850 ;
        RECT 105.930 94.250 106.330 94.700 ;
        RECT 105.930 94.100 109.880 94.250 ;
        RECT 105.930 93.650 106.330 94.100 ;
        RECT 105.930 93.500 109.880 93.650 ;
        RECT 105.930 93.050 106.330 93.500 ;
        RECT 105.930 92.900 109.880 93.050 ;
        RECT 105.930 92.450 106.330 92.900 ;
        RECT 105.930 92.300 109.880 92.450 ;
        RECT 105.930 91.850 106.330 92.300 ;
        RECT 105.930 91.700 109.880 91.850 ;
        RECT 105.930 91.250 106.330 91.700 ;
        RECT 105.930 91.100 109.880 91.250 ;
        RECT 105.930 90.650 106.330 91.100 ;
        RECT 105.930 90.500 109.880 90.650 ;
        RECT 105.930 90.200 106.330 90.500 ;
        RECT 110.480 90.200 110.630 98.400 ;
        RECT 111.080 90.200 111.230 98.400 ;
        RECT 111.680 90.200 111.830 98.400 ;
        RECT 112.280 90.200 112.430 98.400 ;
        RECT 112.880 90.200 113.030 98.400 ;
        RECT 113.480 90.200 113.630 98.400 ;
        RECT 114.080 90.200 114.230 98.400 ;
        RECT 105.930 89.800 114.230 90.200 ;
        RECT 105.930 89.500 106.330 89.800 ;
        RECT 105.930 89.350 109.880 89.500 ;
        RECT 105.930 88.900 106.330 89.350 ;
        RECT 105.930 88.750 109.880 88.900 ;
        RECT 105.930 88.300 106.330 88.750 ;
        RECT 105.930 88.150 109.880 88.300 ;
        RECT 105.930 87.700 106.330 88.150 ;
        RECT 105.930 87.550 109.880 87.700 ;
        RECT 105.930 87.100 106.330 87.550 ;
        RECT 105.930 86.950 109.880 87.100 ;
        RECT 105.930 86.500 106.330 86.950 ;
        RECT 105.930 86.350 109.880 86.500 ;
        RECT 105.930 85.900 106.330 86.350 ;
        RECT 105.930 85.750 109.880 85.900 ;
        RECT 105.930 85.300 106.330 85.750 ;
        RECT 105.930 85.150 109.880 85.300 ;
        RECT 105.930 84.700 106.330 85.150 ;
        RECT 105.930 84.550 109.880 84.700 ;
        RECT 105.930 84.400 106.330 84.550 ;
        RECT 103.130 84.100 106.330 84.400 ;
        RECT 99.580 83.950 109.880 84.100 ;
        RECT 103.130 83.500 106.330 83.950 ;
        RECT 99.580 83.350 109.880 83.500 ;
        RECT 103.130 82.900 106.330 83.350 ;
        RECT 99.580 82.750 109.880 82.900 ;
        RECT 103.130 82.300 106.330 82.750 ;
        RECT 99.580 82.150 109.880 82.300 ;
        RECT 103.530 81.200 105.930 82.150 ;
        RECT 110.480 81.600 110.630 89.800 ;
        RECT 111.080 81.600 111.230 89.800 ;
        RECT 111.680 81.600 111.830 89.800 ;
        RECT 112.280 81.600 112.430 89.800 ;
        RECT 112.880 81.600 113.030 89.800 ;
        RECT 113.480 81.600 113.630 89.800 ;
        RECT 114.080 81.600 114.230 89.800 ;
        RECT 115.230 90.200 115.380 98.400 ;
        RECT 115.830 90.200 115.980 98.400 ;
        RECT 116.430 90.200 116.580 98.400 ;
        RECT 117.030 90.200 117.180 98.400 ;
        RECT 117.630 90.200 117.780 98.400 ;
        RECT 118.230 90.200 118.380 98.400 ;
        RECT 118.830 90.200 118.980 98.400 ;
        RECT 123.530 97.850 124.730 98.800 ;
        RECT 119.580 97.700 124.730 97.850 ;
        RECT 123.130 97.250 124.730 97.700 ;
        RECT 119.580 97.100 124.730 97.250 ;
        RECT 123.130 96.650 124.730 97.100 ;
        RECT 119.580 96.500 124.730 96.650 ;
        RECT 123.130 96.050 124.730 96.500 ;
        RECT 119.580 95.900 124.730 96.050 ;
        RECT 125.140 95.970 127.140 97.245 ;
        RECT 123.130 95.600 124.730 95.900 ;
        RECT 123.130 95.450 123.530 95.600 ;
        RECT 119.580 95.300 123.530 95.450 ;
        RECT 123.130 94.850 123.530 95.300 ;
        RECT 119.580 94.700 123.530 94.850 ;
        RECT 123.130 94.250 123.530 94.700 ;
        RECT 119.580 94.100 123.530 94.250 ;
        RECT 123.130 93.650 123.530 94.100 ;
        RECT 119.580 93.500 123.530 93.650 ;
        RECT 123.130 93.050 123.530 93.500 ;
        RECT 119.580 92.900 123.530 93.050 ;
        RECT 123.130 92.450 123.530 92.900 ;
        RECT 119.580 92.300 123.530 92.450 ;
        RECT 123.130 91.850 123.530 92.300 ;
        RECT 119.580 91.700 123.530 91.850 ;
        RECT 123.130 91.250 123.530 91.700 ;
        RECT 119.580 91.100 123.530 91.250 ;
        RECT 123.130 90.650 123.530 91.100 ;
        RECT 119.580 90.500 123.530 90.650 ;
        RECT 123.130 90.200 123.530 90.500 ;
        RECT 115.230 89.800 123.530 90.200 ;
        RECT 115.230 81.600 115.380 89.800 ;
        RECT 115.830 81.600 115.980 89.800 ;
        RECT 116.430 81.600 116.580 89.800 ;
        RECT 117.030 81.600 117.180 89.800 ;
        RECT 117.630 81.600 117.780 89.800 ;
        RECT 118.230 81.600 118.380 89.800 ;
        RECT 118.830 81.600 118.980 89.800 ;
        RECT 123.130 89.500 123.530 89.800 ;
        RECT 119.580 89.350 123.530 89.500 ;
        RECT 123.130 88.900 123.530 89.350 ;
        RECT 119.580 88.750 123.530 88.900 ;
        RECT 123.130 88.300 123.530 88.750 ;
        RECT 119.580 88.150 123.530 88.300 ;
        RECT 123.130 87.700 123.530 88.150 ;
        RECT 119.580 87.550 123.530 87.700 ;
        RECT 123.130 87.100 123.530 87.550 ;
        RECT 119.580 86.950 123.530 87.100 ;
        RECT 123.130 86.500 123.530 86.950 ;
        RECT 119.580 86.350 123.530 86.500 ;
        RECT 123.130 85.900 123.530 86.350 ;
        RECT 119.580 85.750 123.530 85.900 ;
        RECT 123.130 85.300 123.530 85.750 ;
        RECT 119.580 85.150 123.530 85.300 ;
        RECT 123.130 84.700 123.530 85.150 ;
        RECT 119.580 84.550 123.530 84.700 ;
        RECT 123.130 84.400 123.530 84.550 ;
        RECT 123.130 84.100 124.730 84.400 ;
        RECT 119.580 83.950 124.730 84.100 ;
        RECT 123.130 83.500 124.730 83.950 ;
        RECT 119.580 83.350 124.730 83.500 ;
        RECT 123.130 82.900 124.730 83.350 ;
        RECT 119.580 82.750 124.730 82.900 ;
        RECT 123.130 82.300 124.730 82.750 ;
        RECT 119.580 82.150 124.730 82.300 ;
        RECT 123.530 81.200 124.730 82.150 ;
        RECT 125.135 81.765 127.135 83.040 ;
        RECT 4.730 78.800 9.130 81.200 ;
        RECT 20.330 78.800 29.130 81.200 ;
        RECT 40.330 78.800 49.130 81.200 ;
        RECT 60.330 78.800 69.130 81.200 ;
        RECT 80.330 78.800 89.130 81.200 ;
        RECT 100.330 78.800 109.130 81.200 ;
        RECT 120.330 78.800 124.730 81.200 ;
        RECT 2.315 76.690 4.320 77.965 ;
        RECT 4.730 77.850 5.940 78.800 ;
        RECT 4.730 77.700 9.880 77.850 ;
        RECT 4.730 77.250 6.330 77.700 ;
        RECT 4.730 77.100 9.880 77.250 ;
        RECT 4.730 76.650 6.330 77.100 ;
        RECT 4.730 76.500 9.880 76.650 ;
        RECT 4.730 76.050 6.330 76.500 ;
        RECT 4.730 75.900 9.880 76.050 ;
        RECT 4.730 75.600 6.330 75.900 ;
        RECT 2.315 73.250 4.315 75.545 ;
        RECT 5.930 75.450 6.330 75.600 ;
        RECT 5.930 75.300 9.880 75.450 ;
        RECT 5.930 74.850 6.330 75.300 ;
        RECT 5.930 74.700 9.880 74.850 ;
        RECT 5.930 74.250 6.330 74.700 ;
        RECT 5.930 74.100 9.880 74.250 ;
        RECT 5.930 73.650 6.330 74.100 ;
        RECT 5.930 73.500 9.880 73.650 ;
        RECT 5.930 73.050 6.330 73.500 ;
        RECT 5.930 72.900 9.880 73.050 ;
        RECT 5.930 72.450 6.330 72.900 ;
        RECT 5.930 72.300 9.880 72.450 ;
        RECT 5.930 71.850 6.330 72.300 ;
        RECT 5.930 71.700 9.880 71.850 ;
        RECT 5.930 71.250 6.330 71.700 ;
        RECT 5.930 71.100 9.880 71.250 ;
        RECT 5.930 70.650 6.330 71.100 ;
        RECT 5.930 70.500 9.880 70.650 ;
        RECT 5.930 70.200 6.330 70.500 ;
        RECT 10.480 70.200 10.630 78.400 ;
        RECT 11.080 70.200 11.230 78.400 ;
        RECT 11.680 70.200 11.830 78.400 ;
        RECT 12.280 70.200 12.430 78.400 ;
        RECT 12.880 70.200 13.030 78.400 ;
        RECT 13.480 70.200 13.630 78.400 ;
        RECT 14.080 70.200 14.230 78.400 ;
        RECT 5.930 69.800 14.230 70.200 ;
        RECT 5.930 69.500 6.330 69.800 ;
        RECT 5.930 69.350 9.880 69.500 ;
        RECT 5.930 68.900 6.330 69.350 ;
        RECT 5.930 68.750 9.880 68.900 ;
        RECT 5.930 68.300 6.330 68.750 ;
        RECT 5.930 68.150 9.880 68.300 ;
        RECT 5.930 67.700 6.330 68.150 ;
        RECT 5.930 67.550 9.880 67.700 ;
        RECT 5.930 67.100 6.330 67.550 ;
        RECT 5.930 66.950 9.880 67.100 ;
        RECT 2.315 64.450 4.315 66.745 ;
        RECT 5.930 66.500 6.330 66.950 ;
        RECT 5.930 66.350 9.880 66.500 ;
        RECT 5.930 65.900 6.330 66.350 ;
        RECT 5.930 65.750 9.880 65.900 ;
        RECT 5.930 65.300 6.330 65.750 ;
        RECT 5.930 65.150 9.880 65.300 ;
        RECT 5.930 64.700 6.330 65.150 ;
        RECT 5.930 64.550 9.880 64.700 ;
        RECT 5.930 64.400 6.330 64.550 ;
        RECT 4.730 64.100 6.330 64.400 ;
        RECT 4.730 63.950 9.880 64.100 ;
        RECT 2.315 62.360 4.325 63.635 ;
        RECT 4.730 63.500 6.330 63.950 ;
        RECT 4.730 63.350 9.880 63.500 ;
        RECT 4.730 62.900 6.330 63.350 ;
        RECT 4.730 62.750 9.880 62.900 ;
        RECT 4.730 62.300 6.330 62.750 ;
        RECT 4.730 62.150 9.880 62.300 ;
        RECT 4.730 61.200 5.930 62.150 ;
        RECT 10.480 61.600 10.630 69.800 ;
        RECT 11.080 61.600 11.230 69.800 ;
        RECT 11.680 61.600 11.830 69.800 ;
        RECT 12.280 61.600 12.430 69.800 ;
        RECT 12.880 61.600 13.030 69.800 ;
        RECT 13.480 61.600 13.630 69.800 ;
        RECT 14.080 61.600 14.230 69.800 ;
        RECT 15.230 70.200 15.380 78.400 ;
        RECT 15.830 70.200 15.980 78.400 ;
        RECT 16.430 70.200 16.580 78.400 ;
        RECT 17.030 70.200 17.180 78.400 ;
        RECT 17.630 70.200 17.780 78.400 ;
        RECT 18.230 70.200 18.380 78.400 ;
        RECT 18.830 70.200 18.980 78.400 ;
        RECT 23.530 77.850 25.940 78.800 ;
        RECT 19.580 77.700 29.880 77.850 ;
        RECT 23.130 77.250 26.330 77.700 ;
        RECT 19.580 77.100 29.880 77.250 ;
        RECT 23.130 76.650 26.330 77.100 ;
        RECT 19.580 76.500 29.880 76.650 ;
        RECT 23.130 76.050 26.330 76.500 ;
        RECT 19.580 75.900 29.880 76.050 ;
        RECT 23.130 75.600 26.330 75.900 ;
        RECT 23.130 75.450 23.530 75.600 ;
        RECT 19.580 75.300 23.530 75.450 ;
        RECT 23.130 74.850 23.530 75.300 ;
        RECT 19.580 74.700 23.530 74.850 ;
        RECT 23.130 74.250 23.530 74.700 ;
        RECT 19.580 74.100 23.530 74.250 ;
        RECT 23.130 73.650 23.530 74.100 ;
        RECT 19.580 73.500 23.530 73.650 ;
        RECT 23.130 73.050 23.530 73.500 ;
        RECT 19.580 72.900 23.530 73.050 ;
        RECT 23.130 72.450 23.530 72.900 ;
        RECT 19.580 72.300 23.530 72.450 ;
        RECT 23.130 71.850 23.530 72.300 ;
        RECT 19.580 71.700 23.530 71.850 ;
        RECT 23.130 71.250 23.530 71.700 ;
        RECT 19.580 71.100 23.530 71.250 ;
        RECT 23.130 70.650 23.530 71.100 ;
        RECT 19.580 70.500 23.530 70.650 ;
        RECT 23.130 70.200 23.530 70.500 ;
        RECT 15.230 69.800 23.530 70.200 ;
        RECT 15.230 61.600 15.380 69.800 ;
        RECT 15.830 61.600 15.980 69.800 ;
        RECT 16.430 61.600 16.580 69.800 ;
        RECT 17.030 61.600 17.180 69.800 ;
        RECT 17.630 61.600 17.780 69.800 ;
        RECT 18.230 61.600 18.380 69.800 ;
        RECT 18.830 61.600 18.980 69.800 ;
        RECT 23.130 69.500 23.530 69.800 ;
        RECT 19.580 69.350 23.530 69.500 ;
        RECT 23.130 68.900 23.530 69.350 ;
        RECT 19.580 68.750 23.530 68.900 ;
        RECT 23.130 68.300 23.530 68.750 ;
        RECT 19.580 68.150 23.530 68.300 ;
        RECT 23.130 67.700 23.530 68.150 ;
        RECT 19.580 67.550 23.530 67.700 ;
        RECT 23.130 67.100 23.530 67.550 ;
        RECT 19.580 66.950 23.530 67.100 ;
        RECT 23.130 66.500 23.530 66.950 ;
        RECT 19.580 66.350 23.530 66.500 ;
        RECT 23.130 65.900 23.530 66.350 ;
        RECT 19.580 65.750 23.530 65.900 ;
        RECT 23.130 65.300 23.530 65.750 ;
        RECT 19.580 65.150 23.530 65.300 ;
        RECT 23.130 64.700 23.530 65.150 ;
        RECT 19.580 64.550 23.530 64.700 ;
        RECT 23.130 64.400 23.530 64.550 ;
        RECT 25.930 75.450 26.330 75.600 ;
        RECT 25.930 75.300 29.880 75.450 ;
        RECT 25.930 74.850 26.330 75.300 ;
        RECT 25.930 74.700 29.880 74.850 ;
        RECT 25.930 74.250 26.330 74.700 ;
        RECT 25.930 74.100 29.880 74.250 ;
        RECT 25.930 73.650 26.330 74.100 ;
        RECT 25.930 73.500 29.880 73.650 ;
        RECT 25.930 73.050 26.330 73.500 ;
        RECT 25.930 72.900 29.880 73.050 ;
        RECT 25.930 72.450 26.330 72.900 ;
        RECT 25.930 72.300 29.880 72.450 ;
        RECT 25.930 71.850 26.330 72.300 ;
        RECT 25.930 71.700 29.880 71.850 ;
        RECT 25.930 71.250 26.330 71.700 ;
        RECT 25.930 71.100 29.880 71.250 ;
        RECT 25.930 70.650 26.330 71.100 ;
        RECT 25.930 70.500 29.880 70.650 ;
        RECT 25.930 70.200 26.330 70.500 ;
        RECT 30.480 70.200 30.630 78.400 ;
        RECT 31.080 70.200 31.230 78.400 ;
        RECT 31.680 70.200 31.830 78.400 ;
        RECT 32.280 70.200 32.430 78.400 ;
        RECT 32.880 70.200 33.030 78.400 ;
        RECT 33.480 70.200 33.630 78.400 ;
        RECT 34.080 70.200 34.230 78.400 ;
        RECT 25.930 69.800 34.230 70.200 ;
        RECT 25.930 69.500 26.330 69.800 ;
        RECT 25.930 69.350 29.880 69.500 ;
        RECT 25.930 68.900 26.330 69.350 ;
        RECT 25.930 68.750 29.880 68.900 ;
        RECT 25.930 68.300 26.330 68.750 ;
        RECT 25.930 68.150 29.880 68.300 ;
        RECT 25.930 67.700 26.330 68.150 ;
        RECT 25.930 67.550 29.880 67.700 ;
        RECT 25.930 67.100 26.330 67.550 ;
        RECT 25.930 66.950 29.880 67.100 ;
        RECT 25.930 66.500 26.330 66.950 ;
        RECT 25.930 66.350 29.880 66.500 ;
        RECT 25.930 65.900 26.330 66.350 ;
        RECT 25.930 65.750 29.880 65.900 ;
        RECT 25.930 65.300 26.330 65.750 ;
        RECT 25.930 65.150 29.880 65.300 ;
        RECT 25.930 64.700 26.330 65.150 ;
        RECT 25.930 64.550 29.880 64.700 ;
        RECT 25.930 64.400 26.330 64.550 ;
        RECT 23.130 64.100 26.330 64.400 ;
        RECT 19.580 63.950 29.880 64.100 ;
        RECT 23.130 63.500 26.330 63.950 ;
        RECT 19.580 63.350 29.880 63.500 ;
        RECT 23.130 62.900 26.330 63.350 ;
        RECT 19.580 62.750 29.880 62.900 ;
        RECT 23.130 62.300 26.330 62.750 ;
        RECT 19.580 62.150 29.880 62.300 ;
        RECT 23.530 61.200 25.930 62.150 ;
        RECT 30.480 61.600 30.630 69.800 ;
        RECT 31.080 61.600 31.230 69.800 ;
        RECT 31.680 61.600 31.830 69.800 ;
        RECT 32.280 61.600 32.430 69.800 ;
        RECT 32.880 61.600 33.030 69.800 ;
        RECT 33.480 61.600 33.630 69.800 ;
        RECT 34.080 61.600 34.230 69.800 ;
        RECT 35.230 70.200 35.380 78.400 ;
        RECT 35.830 70.200 35.980 78.400 ;
        RECT 36.430 70.200 36.580 78.400 ;
        RECT 37.030 70.200 37.180 78.400 ;
        RECT 37.630 70.200 37.780 78.400 ;
        RECT 38.230 70.200 38.380 78.400 ;
        RECT 38.830 70.200 38.980 78.400 ;
        RECT 43.530 77.850 45.940 78.800 ;
        RECT 39.580 77.700 49.880 77.850 ;
        RECT 43.130 77.250 46.330 77.700 ;
        RECT 39.580 77.100 49.880 77.250 ;
        RECT 43.130 76.650 46.330 77.100 ;
        RECT 39.580 76.500 49.880 76.650 ;
        RECT 43.130 76.050 46.330 76.500 ;
        RECT 39.580 75.900 49.880 76.050 ;
        RECT 43.130 75.600 46.330 75.900 ;
        RECT 43.130 75.450 43.530 75.600 ;
        RECT 39.580 75.300 43.530 75.450 ;
        RECT 43.130 74.850 43.530 75.300 ;
        RECT 39.580 74.700 43.530 74.850 ;
        RECT 43.130 74.250 43.530 74.700 ;
        RECT 39.580 74.100 43.530 74.250 ;
        RECT 43.130 73.650 43.530 74.100 ;
        RECT 39.580 73.500 43.530 73.650 ;
        RECT 43.130 73.050 43.530 73.500 ;
        RECT 39.580 72.900 43.530 73.050 ;
        RECT 43.130 72.450 43.530 72.900 ;
        RECT 39.580 72.300 43.530 72.450 ;
        RECT 43.130 71.850 43.530 72.300 ;
        RECT 39.580 71.700 43.530 71.850 ;
        RECT 43.130 71.250 43.530 71.700 ;
        RECT 39.580 71.100 43.530 71.250 ;
        RECT 43.130 70.650 43.530 71.100 ;
        RECT 39.580 70.500 43.530 70.650 ;
        RECT 43.130 70.200 43.530 70.500 ;
        RECT 35.230 69.800 43.530 70.200 ;
        RECT 35.230 61.600 35.380 69.800 ;
        RECT 35.830 61.600 35.980 69.800 ;
        RECT 36.430 61.600 36.580 69.800 ;
        RECT 37.030 61.600 37.180 69.800 ;
        RECT 37.630 61.600 37.780 69.800 ;
        RECT 38.230 61.600 38.380 69.800 ;
        RECT 38.830 61.600 38.980 69.800 ;
        RECT 43.130 69.500 43.530 69.800 ;
        RECT 39.580 69.350 43.530 69.500 ;
        RECT 43.130 68.900 43.530 69.350 ;
        RECT 39.580 68.750 43.530 68.900 ;
        RECT 43.130 68.300 43.530 68.750 ;
        RECT 39.580 68.150 43.530 68.300 ;
        RECT 43.130 67.700 43.530 68.150 ;
        RECT 39.580 67.550 43.530 67.700 ;
        RECT 43.130 67.100 43.530 67.550 ;
        RECT 39.580 66.950 43.530 67.100 ;
        RECT 43.130 66.500 43.530 66.950 ;
        RECT 39.580 66.350 43.530 66.500 ;
        RECT 43.130 65.900 43.530 66.350 ;
        RECT 39.580 65.750 43.530 65.900 ;
        RECT 43.130 65.300 43.530 65.750 ;
        RECT 39.580 65.150 43.530 65.300 ;
        RECT 43.130 64.700 43.530 65.150 ;
        RECT 39.580 64.550 43.530 64.700 ;
        RECT 43.130 64.400 43.530 64.550 ;
        RECT 45.930 75.450 46.330 75.600 ;
        RECT 45.930 75.300 49.880 75.450 ;
        RECT 45.930 74.850 46.330 75.300 ;
        RECT 45.930 74.700 49.880 74.850 ;
        RECT 45.930 74.250 46.330 74.700 ;
        RECT 45.930 74.100 49.880 74.250 ;
        RECT 45.930 73.650 46.330 74.100 ;
        RECT 45.930 73.500 49.880 73.650 ;
        RECT 45.930 73.050 46.330 73.500 ;
        RECT 45.930 72.900 49.880 73.050 ;
        RECT 45.930 72.450 46.330 72.900 ;
        RECT 45.930 72.300 49.880 72.450 ;
        RECT 45.930 71.850 46.330 72.300 ;
        RECT 45.930 71.700 49.880 71.850 ;
        RECT 45.930 71.250 46.330 71.700 ;
        RECT 45.930 71.100 49.880 71.250 ;
        RECT 45.930 70.650 46.330 71.100 ;
        RECT 45.930 70.500 49.880 70.650 ;
        RECT 45.930 70.200 46.330 70.500 ;
        RECT 50.480 70.200 50.630 78.400 ;
        RECT 51.080 70.200 51.230 78.400 ;
        RECT 51.680 70.200 51.830 78.400 ;
        RECT 52.280 70.200 52.430 78.400 ;
        RECT 52.880 70.200 53.030 78.400 ;
        RECT 53.480 70.200 53.630 78.400 ;
        RECT 54.080 70.200 54.230 78.400 ;
        RECT 45.930 69.800 54.230 70.200 ;
        RECT 45.930 69.500 46.330 69.800 ;
        RECT 45.930 69.350 49.880 69.500 ;
        RECT 45.930 68.900 46.330 69.350 ;
        RECT 45.930 68.750 49.880 68.900 ;
        RECT 45.930 68.300 46.330 68.750 ;
        RECT 45.930 68.150 49.880 68.300 ;
        RECT 45.930 67.700 46.330 68.150 ;
        RECT 45.930 67.550 49.880 67.700 ;
        RECT 45.930 67.100 46.330 67.550 ;
        RECT 45.930 66.950 49.880 67.100 ;
        RECT 45.930 66.500 46.330 66.950 ;
        RECT 45.930 66.350 49.880 66.500 ;
        RECT 45.930 65.900 46.330 66.350 ;
        RECT 45.930 65.750 49.880 65.900 ;
        RECT 45.930 65.300 46.330 65.750 ;
        RECT 45.930 65.150 49.880 65.300 ;
        RECT 45.930 64.700 46.330 65.150 ;
        RECT 45.930 64.550 49.880 64.700 ;
        RECT 45.930 64.400 46.330 64.550 ;
        RECT 43.130 64.100 46.330 64.400 ;
        RECT 39.580 63.950 49.880 64.100 ;
        RECT 43.130 63.500 46.330 63.950 ;
        RECT 39.580 63.350 49.880 63.500 ;
        RECT 43.130 62.900 46.330 63.350 ;
        RECT 39.580 62.750 49.880 62.900 ;
        RECT 43.130 62.300 46.330 62.750 ;
        RECT 39.580 62.150 49.880 62.300 ;
        RECT 43.530 61.200 45.930 62.150 ;
        RECT 50.480 61.600 50.630 69.800 ;
        RECT 51.080 61.600 51.230 69.800 ;
        RECT 51.680 61.600 51.830 69.800 ;
        RECT 52.280 61.600 52.430 69.800 ;
        RECT 52.880 61.600 53.030 69.800 ;
        RECT 53.480 61.600 53.630 69.800 ;
        RECT 54.080 61.600 54.230 69.800 ;
        RECT 55.230 70.200 55.380 78.400 ;
        RECT 55.830 70.200 55.980 78.400 ;
        RECT 56.430 70.200 56.580 78.400 ;
        RECT 57.030 70.200 57.180 78.400 ;
        RECT 57.630 70.200 57.780 78.400 ;
        RECT 58.230 70.200 58.380 78.400 ;
        RECT 58.830 70.200 58.980 78.400 ;
        RECT 63.530 77.850 65.940 78.800 ;
        RECT 59.580 77.700 69.880 77.850 ;
        RECT 63.130 77.250 66.330 77.700 ;
        RECT 59.580 77.100 69.880 77.250 ;
        RECT 63.130 76.650 66.330 77.100 ;
        RECT 59.580 76.500 69.880 76.650 ;
        RECT 63.130 76.050 66.330 76.500 ;
        RECT 59.580 75.900 69.880 76.050 ;
        RECT 63.130 75.600 66.330 75.900 ;
        RECT 63.130 75.450 63.530 75.600 ;
        RECT 59.580 75.300 63.530 75.450 ;
        RECT 63.130 74.850 63.530 75.300 ;
        RECT 59.580 74.700 63.530 74.850 ;
        RECT 63.130 74.250 63.530 74.700 ;
        RECT 59.580 74.100 63.530 74.250 ;
        RECT 63.130 73.650 63.530 74.100 ;
        RECT 59.580 73.500 63.530 73.650 ;
        RECT 63.130 73.050 63.530 73.500 ;
        RECT 59.580 72.900 63.530 73.050 ;
        RECT 63.130 72.450 63.530 72.900 ;
        RECT 59.580 72.300 63.530 72.450 ;
        RECT 63.130 71.850 63.530 72.300 ;
        RECT 59.580 71.700 63.530 71.850 ;
        RECT 63.130 71.250 63.530 71.700 ;
        RECT 59.580 71.100 63.530 71.250 ;
        RECT 63.130 70.650 63.530 71.100 ;
        RECT 59.580 70.500 63.530 70.650 ;
        RECT 63.130 70.200 63.530 70.500 ;
        RECT 55.230 69.800 63.530 70.200 ;
        RECT 55.230 61.600 55.380 69.800 ;
        RECT 55.830 61.600 55.980 69.800 ;
        RECT 56.430 61.600 56.580 69.800 ;
        RECT 57.030 61.600 57.180 69.800 ;
        RECT 57.630 61.600 57.780 69.800 ;
        RECT 58.230 61.600 58.380 69.800 ;
        RECT 58.830 61.600 58.980 69.800 ;
        RECT 63.130 69.500 63.530 69.800 ;
        RECT 59.580 69.350 63.530 69.500 ;
        RECT 63.130 68.900 63.530 69.350 ;
        RECT 59.580 68.750 63.530 68.900 ;
        RECT 63.130 68.300 63.530 68.750 ;
        RECT 59.580 68.150 63.530 68.300 ;
        RECT 63.130 67.700 63.530 68.150 ;
        RECT 59.580 67.550 63.530 67.700 ;
        RECT 63.130 67.100 63.530 67.550 ;
        RECT 59.580 66.950 63.530 67.100 ;
        RECT 63.130 66.500 63.530 66.950 ;
        RECT 59.580 66.350 63.530 66.500 ;
        RECT 63.130 65.900 63.530 66.350 ;
        RECT 59.580 65.750 63.530 65.900 ;
        RECT 63.130 65.300 63.530 65.750 ;
        RECT 59.580 65.150 63.530 65.300 ;
        RECT 63.130 64.700 63.530 65.150 ;
        RECT 59.580 64.550 63.530 64.700 ;
        RECT 63.130 64.400 63.530 64.550 ;
        RECT 65.930 75.450 66.330 75.600 ;
        RECT 65.930 75.300 69.880 75.450 ;
        RECT 65.930 74.850 66.330 75.300 ;
        RECT 65.930 74.700 69.880 74.850 ;
        RECT 65.930 74.250 66.330 74.700 ;
        RECT 65.930 74.100 69.880 74.250 ;
        RECT 65.930 73.650 66.330 74.100 ;
        RECT 65.930 73.500 69.880 73.650 ;
        RECT 65.930 73.050 66.330 73.500 ;
        RECT 65.930 72.900 69.880 73.050 ;
        RECT 65.930 72.450 66.330 72.900 ;
        RECT 65.930 72.300 69.880 72.450 ;
        RECT 65.930 71.850 66.330 72.300 ;
        RECT 65.930 71.700 69.880 71.850 ;
        RECT 65.930 71.250 66.330 71.700 ;
        RECT 65.930 71.100 69.880 71.250 ;
        RECT 65.930 70.650 66.330 71.100 ;
        RECT 65.930 70.500 69.880 70.650 ;
        RECT 65.930 70.200 66.330 70.500 ;
        RECT 70.480 70.200 70.630 78.400 ;
        RECT 71.080 70.200 71.230 78.400 ;
        RECT 71.680 70.200 71.830 78.400 ;
        RECT 72.280 70.200 72.430 78.400 ;
        RECT 72.880 70.200 73.030 78.400 ;
        RECT 73.480 70.200 73.630 78.400 ;
        RECT 74.080 70.200 74.230 78.400 ;
        RECT 65.930 69.800 74.230 70.200 ;
        RECT 65.930 69.500 66.330 69.800 ;
        RECT 65.930 69.350 69.880 69.500 ;
        RECT 65.930 68.900 66.330 69.350 ;
        RECT 65.930 68.750 69.880 68.900 ;
        RECT 65.930 68.300 66.330 68.750 ;
        RECT 65.930 68.150 69.880 68.300 ;
        RECT 65.930 67.700 66.330 68.150 ;
        RECT 65.930 67.550 69.880 67.700 ;
        RECT 65.930 67.100 66.330 67.550 ;
        RECT 65.930 66.950 69.880 67.100 ;
        RECT 65.930 66.500 66.330 66.950 ;
        RECT 65.930 66.350 69.880 66.500 ;
        RECT 65.930 65.900 66.330 66.350 ;
        RECT 65.930 65.750 69.880 65.900 ;
        RECT 65.930 65.300 66.330 65.750 ;
        RECT 65.930 65.150 69.880 65.300 ;
        RECT 65.930 64.700 66.330 65.150 ;
        RECT 65.930 64.550 69.880 64.700 ;
        RECT 65.930 64.400 66.330 64.550 ;
        RECT 63.130 64.100 66.330 64.400 ;
        RECT 59.580 63.950 69.880 64.100 ;
        RECT 63.130 63.500 66.330 63.950 ;
        RECT 59.580 63.350 69.880 63.500 ;
        RECT 63.130 62.900 66.330 63.350 ;
        RECT 59.580 62.750 69.880 62.900 ;
        RECT 63.130 62.300 66.330 62.750 ;
        RECT 59.580 62.150 69.880 62.300 ;
        RECT 63.530 61.200 65.930 62.150 ;
        RECT 70.480 61.600 70.630 69.800 ;
        RECT 71.080 61.600 71.230 69.800 ;
        RECT 71.680 61.600 71.830 69.800 ;
        RECT 72.280 61.600 72.430 69.800 ;
        RECT 72.880 61.600 73.030 69.800 ;
        RECT 73.480 61.600 73.630 69.800 ;
        RECT 74.080 61.600 74.230 69.800 ;
        RECT 75.230 70.200 75.380 78.400 ;
        RECT 75.830 70.200 75.980 78.400 ;
        RECT 76.430 70.200 76.580 78.400 ;
        RECT 77.030 70.200 77.180 78.400 ;
        RECT 77.630 70.200 77.780 78.400 ;
        RECT 78.230 70.200 78.380 78.400 ;
        RECT 78.830 70.200 78.980 78.400 ;
        RECT 83.530 77.850 85.940 78.800 ;
        RECT 79.580 77.700 89.880 77.850 ;
        RECT 83.130 77.250 86.330 77.700 ;
        RECT 79.580 77.100 89.880 77.250 ;
        RECT 83.130 76.650 86.330 77.100 ;
        RECT 79.580 76.500 89.880 76.650 ;
        RECT 83.130 76.050 86.330 76.500 ;
        RECT 79.580 75.900 89.880 76.050 ;
        RECT 83.130 75.600 86.330 75.900 ;
        RECT 83.130 75.450 83.530 75.600 ;
        RECT 79.580 75.300 83.530 75.450 ;
        RECT 83.130 74.850 83.530 75.300 ;
        RECT 79.580 74.700 83.530 74.850 ;
        RECT 83.130 74.250 83.530 74.700 ;
        RECT 79.580 74.100 83.530 74.250 ;
        RECT 83.130 73.650 83.530 74.100 ;
        RECT 79.580 73.500 83.530 73.650 ;
        RECT 83.130 73.050 83.530 73.500 ;
        RECT 79.580 72.900 83.530 73.050 ;
        RECT 83.130 72.450 83.530 72.900 ;
        RECT 79.580 72.300 83.530 72.450 ;
        RECT 83.130 71.850 83.530 72.300 ;
        RECT 79.580 71.700 83.530 71.850 ;
        RECT 83.130 71.250 83.530 71.700 ;
        RECT 79.580 71.100 83.530 71.250 ;
        RECT 83.130 70.650 83.530 71.100 ;
        RECT 79.580 70.500 83.530 70.650 ;
        RECT 83.130 70.200 83.530 70.500 ;
        RECT 75.230 69.800 83.530 70.200 ;
        RECT 75.230 61.600 75.380 69.800 ;
        RECT 75.830 61.600 75.980 69.800 ;
        RECT 76.430 61.600 76.580 69.800 ;
        RECT 77.030 61.600 77.180 69.800 ;
        RECT 77.630 61.600 77.780 69.800 ;
        RECT 78.230 61.600 78.380 69.800 ;
        RECT 78.830 61.600 78.980 69.800 ;
        RECT 83.130 69.500 83.530 69.800 ;
        RECT 79.580 69.350 83.530 69.500 ;
        RECT 83.130 68.900 83.530 69.350 ;
        RECT 79.580 68.750 83.530 68.900 ;
        RECT 83.130 68.300 83.530 68.750 ;
        RECT 79.580 68.150 83.530 68.300 ;
        RECT 83.130 67.700 83.530 68.150 ;
        RECT 79.580 67.550 83.530 67.700 ;
        RECT 83.130 67.100 83.530 67.550 ;
        RECT 79.580 66.950 83.530 67.100 ;
        RECT 83.130 66.500 83.530 66.950 ;
        RECT 79.580 66.350 83.530 66.500 ;
        RECT 83.130 65.900 83.530 66.350 ;
        RECT 79.580 65.750 83.530 65.900 ;
        RECT 83.130 65.300 83.530 65.750 ;
        RECT 79.580 65.150 83.530 65.300 ;
        RECT 83.130 64.700 83.530 65.150 ;
        RECT 79.580 64.550 83.530 64.700 ;
        RECT 83.130 64.400 83.530 64.550 ;
        RECT 85.930 75.450 86.330 75.600 ;
        RECT 85.930 75.300 89.880 75.450 ;
        RECT 85.930 74.850 86.330 75.300 ;
        RECT 85.930 74.700 89.880 74.850 ;
        RECT 85.930 74.250 86.330 74.700 ;
        RECT 85.930 74.100 89.880 74.250 ;
        RECT 85.930 73.650 86.330 74.100 ;
        RECT 85.930 73.500 89.880 73.650 ;
        RECT 85.930 73.050 86.330 73.500 ;
        RECT 85.930 72.900 89.880 73.050 ;
        RECT 85.930 72.450 86.330 72.900 ;
        RECT 85.930 72.300 89.880 72.450 ;
        RECT 85.930 71.850 86.330 72.300 ;
        RECT 85.930 71.700 89.880 71.850 ;
        RECT 85.930 71.250 86.330 71.700 ;
        RECT 85.930 71.100 89.880 71.250 ;
        RECT 85.930 70.650 86.330 71.100 ;
        RECT 85.930 70.500 89.880 70.650 ;
        RECT 85.930 70.200 86.330 70.500 ;
        RECT 90.480 70.200 90.630 78.400 ;
        RECT 91.080 70.200 91.230 78.400 ;
        RECT 91.680 70.200 91.830 78.400 ;
        RECT 92.280 70.200 92.430 78.400 ;
        RECT 92.880 70.200 93.030 78.400 ;
        RECT 93.480 70.200 93.630 78.400 ;
        RECT 94.080 70.200 94.230 78.400 ;
        RECT 85.930 69.800 94.230 70.200 ;
        RECT 85.930 69.500 86.330 69.800 ;
        RECT 85.930 69.350 89.880 69.500 ;
        RECT 85.930 68.900 86.330 69.350 ;
        RECT 85.930 68.750 89.880 68.900 ;
        RECT 85.930 68.300 86.330 68.750 ;
        RECT 85.930 68.150 89.880 68.300 ;
        RECT 85.930 67.700 86.330 68.150 ;
        RECT 85.930 67.550 89.880 67.700 ;
        RECT 85.930 67.100 86.330 67.550 ;
        RECT 85.930 66.950 89.880 67.100 ;
        RECT 85.930 66.500 86.330 66.950 ;
        RECT 85.930 66.350 89.880 66.500 ;
        RECT 85.930 65.900 86.330 66.350 ;
        RECT 85.930 65.750 89.880 65.900 ;
        RECT 85.930 65.300 86.330 65.750 ;
        RECT 85.930 65.150 89.880 65.300 ;
        RECT 85.930 64.700 86.330 65.150 ;
        RECT 85.930 64.550 89.880 64.700 ;
        RECT 85.930 64.400 86.330 64.550 ;
        RECT 83.130 64.100 86.330 64.400 ;
        RECT 79.580 63.950 89.880 64.100 ;
        RECT 83.130 63.500 86.330 63.950 ;
        RECT 79.580 63.350 89.880 63.500 ;
        RECT 83.130 62.900 86.330 63.350 ;
        RECT 79.580 62.750 89.880 62.900 ;
        RECT 83.130 62.300 86.330 62.750 ;
        RECT 79.580 62.150 89.880 62.300 ;
        RECT 83.530 61.200 85.930 62.150 ;
        RECT 90.480 61.600 90.630 69.800 ;
        RECT 91.080 61.600 91.230 69.800 ;
        RECT 91.680 61.600 91.830 69.800 ;
        RECT 92.280 61.600 92.430 69.800 ;
        RECT 92.880 61.600 93.030 69.800 ;
        RECT 93.480 61.600 93.630 69.800 ;
        RECT 94.080 61.600 94.230 69.800 ;
        RECT 95.230 70.200 95.380 78.400 ;
        RECT 95.830 70.200 95.980 78.400 ;
        RECT 96.430 70.200 96.580 78.400 ;
        RECT 97.030 70.200 97.180 78.400 ;
        RECT 97.630 70.200 97.780 78.400 ;
        RECT 98.230 70.200 98.380 78.400 ;
        RECT 98.830 70.200 98.980 78.400 ;
        RECT 103.530 77.850 105.940 78.800 ;
        RECT 99.580 77.700 109.880 77.850 ;
        RECT 103.130 77.250 106.330 77.700 ;
        RECT 99.580 77.100 109.880 77.250 ;
        RECT 103.130 76.650 106.330 77.100 ;
        RECT 99.580 76.500 109.880 76.650 ;
        RECT 103.130 76.050 106.330 76.500 ;
        RECT 99.580 75.900 109.880 76.050 ;
        RECT 103.130 75.600 106.330 75.900 ;
        RECT 103.130 75.450 103.530 75.600 ;
        RECT 99.580 75.300 103.530 75.450 ;
        RECT 103.130 74.850 103.530 75.300 ;
        RECT 99.580 74.700 103.530 74.850 ;
        RECT 103.130 74.250 103.530 74.700 ;
        RECT 99.580 74.100 103.530 74.250 ;
        RECT 103.130 73.650 103.530 74.100 ;
        RECT 99.580 73.500 103.530 73.650 ;
        RECT 103.130 73.050 103.530 73.500 ;
        RECT 99.580 72.900 103.530 73.050 ;
        RECT 103.130 72.450 103.530 72.900 ;
        RECT 99.580 72.300 103.530 72.450 ;
        RECT 103.130 71.850 103.530 72.300 ;
        RECT 99.580 71.700 103.530 71.850 ;
        RECT 103.130 71.250 103.530 71.700 ;
        RECT 99.580 71.100 103.530 71.250 ;
        RECT 103.130 70.650 103.530 71.100 ;
        RECT 99.580 70.500 103.530 70.650 ;
        RECT 103.130 70.200 103.530 70.500 ;
        RECT 95.230 69.800 103.530 70.200 ;
        RECT 95.230 61.600 95.380 69.800 ;
        RECT 95.830 61.600 95.980 69.800 ;
        RECT 96.430 61.600 96.580 69.800 ;
        RECT 97.030 61.600 97.180 69.800 ;
        RECT 97.630 61.600 97.780 69.800 ;
        RECT 98.230 61.600 98.380 69.800 ;
        RECT 98.830 61.600 98.980 69.800 ;
        RECT 103.130 69.500 103.530 69.800 ;
        RECT 99.580 69.350 103.530 69.500 ;
        RECT 103.130 68.900 103.530 69.350 ;
        RECT 99.580 68.750 103.530 68.900 ;
        RECT 103.130 68.300 103.530 68.750 ;
        RECT 99.580 68.150 103.530 68.300 ;
        RECT 103.130 67.700 103.530 68.150 ;
        RECT 99.580 67.550 103.530 67.700 ;
        RECT 103.130 67.100 103.530 67.550 ;
        RECT 99.580 66.950 103.530 67.100 ;
        RECT 103.130 66.500 103.530 66.950 ;
        RECT 99.580 66.350 103.530 66.500 ;
        RECT 103.130 65.900 103.530 66.350 ;
        RECT 99.580 65.750 103.530 65.900 ;
        RECT 103.130 65.300 103.530 65.750 ;
        RECT 99.580 65.150 103.530 65.300 ;
        RECT 103.130 64.700 103.530 65.150 ;
        RECT 99.580 64.550 103.530 64.700 ;
        RECT 103.130 64.400 103.530 64.550 ;
        RECT 105.930 75.450 106.330 75.600 ;
        RECT 105.930 75.300 109.880 75.450 ;
        RECT 105.930 74.850 106.330 75.300 ;
        RECT 105.930 74.700 109.880 74.850 ;
        RECT 105.930 74.250 106.330 74.700 ;
        RECT 105.930 74.100 109.880 74.250 ;
        RECT 105.930 73.650 106.330 74.100 ;
        RECT 105.930 73.500 109.880 73.650 ;
        RECT 105.930 73.050 106.330 73.500 ;
        RECT 105.930 72.900 109.880 73.050 ;
        RECT 105.930 72.450 106.330 72.900 ;
        RECT 105.930 72.300 109.880 72.450 ;
        RECT 105.930 71.850 106.330 72.300 ;
        RECT 105.930 71.700 109.880 71.850 ;
        RECT 105.930 71.250 106.330 71.700 ;
        RECT 105.930 71.100 109.880 71.250 ;
        RECT 105.930 70.650 106.330 71.100 ;
        RECT 105.930 70.500 109.880 70.650 ;
        RECT 105.930 70.200 106.330 70.500 ;
        RECT 110.480 70.200 110.630 78.400 ;
        RECT 111.080 70.200 111.230 78.400 ;
        RECT 111.680 70.200 111.830 78.400 ;
        RECT 112.280 70.200 112.430 78.400 ;
        RECT 112.880 70.200 113.030 78.400 ;
        RECT 113.480 70.200 113.630 78.400 ;
        RECT 114.080 70.200 114.230 78.400 ;
        RECT 105.930 69.800 114.230 70.200 ;
        RECT 105.930 69.500 106.330 69.800 ;
        RECT 105.930 69.350 109.880 69.500 ;
        RECT 105.930 68.900 106.330 69.350 ;
        RECT 105.930 68.750 109.880 68.900 ;
        RECT 105.930 68.300 106.330 68.750 ;
        RECT 105.930 68.150 109.880 68.300 ;
        RECT 105.930 67.700 106.330 68.150 ;
        RECT 105.930 67.550 109.880 67.700 ;
        RECT 105.930 67.100 106.330 67.550 ;
        RECT 105.930 66.950 109.880 67.100 ;
        RECT 105.930 66.500 106.330 66.950 ;
        RECT 105.930 66.350 109.880 66.500 ;
        RECT 105.930 65.900 106.330 66.350 ;
        RECT 105.930 65.750 109.880 65.900 ;
        RECT 105.930 65.300 106.330 65.750 ;
        RECT 105.930 65.150 109.880 65.300 ;
        RECT 105.930 64.700 106.330 65.150 ;
        RECT 105.930 64.550 109.880 64.700 ;
        RECT 105.930 64.400 106.330 64.550 ;
        RECT 103.130 64.100 106.330 64.400 ;
        RECT 99.580 63.950 109.880 64.100 ;
        RECT 103.130 63.500 106.330 63.950 ;
        RECT 99.580 63.350 109.880 63.500 ;
        RECT 103.130 62.900 106.330 63.350 ;
        RECT 99.580 62.750 109.880 62.900 ;
        RECT 103.130 62.300 106.330 62.750 ;
        RECT 99.580 62.150 109.880 62.300 ;
        RECT 103.530 61.200 105.930 62.150 ;
        RECT 110.480 61.600 110.630 69.800 ;
        RECT 111.080 61.600 111.230 69.800 ;
        RECT 111.680 61.600 111.830 69.800 ;
        RECT 112.280 61.600 112.430 69.800 ;
        RECT 112.880 61.600 113.030 69.800 ;
        RECT 113.480 61.600 113.630 69.800 ;
        RECT 114.080 61.600 114.230 69.800 ;
        RECT 115.230 70.200 115.380 78.400 ;
        RECT 115.830 70.200 115.980 78.400 ;
        RECT 116.430 70.200 116.580 78.400 ;
        RECT 117.030 70.200 117.180 78.400 ;
        RECT 117.630 70.200 117.780 78.400 ;
        RECT 118.230 70.200 118.380 78.400 ;
        RECT 118.830 70.200 118.980 78.400 ;
        RECT 123.530 77.850 124.730 78.800 ;
        RECT 119.580 77.700 124.730 77.850 ;
        RECT 123.130 77.250 124.730 77.700 ;
        RECT 119.580 77.100 124.730 77.250 ;
        RECT 123.130 76.650 124.730 77.100 ;
        RECT 119.580 76.500 124.730 76.650 ;
        RECT 123.130 76.050 124.730 76.500 ;
        RECT 119.580 75.900 124.730 76.050 ;
        RECT 125.135 75.910 127.135 77.185 ;
        RECT 123.130 75.600 124.730 75.900 ;
        RECT 123.130 75.450 123.530 75.600 ;
        RECT 119.580 75.300 123.530 75.450 ;
        RECT 123.130 74.850 123.530 75.300 ;
        RECT 119.580 74.700 123.530 74.850 ;
        RECT 123.130 74.250 123.530 74.700 ;
        RECT 119.580 74.100 123.530 74.250 ;
        RECT 123.130 73.650 123.530 74.100 ;
        RECT 119.580 73.500 123.530 73.650 ;
        RECT 123.130 73.050 123.530 73.500 ;
        RECT 119.580 72.900 123.530 73.050 ;
        RECT 123.130 72.450 123.530 72.900 ;
        RECT 119.580 72.300 123.530 72.450 ;
        RECT 123.130 71.850 123.530 72.300 ;
        RECT 119.580 71.700 123.530 71.850 ;
        RECT 123.130 71.250 123.530 71.700 ;
        RECT 119.580 71.100 123.530 71.250 ;
        RECT 123.130 70.650 123.530 71.100 ;
        RECT 119.580 70.500 123.530 70.650 ;
        RECT 123.130 70.200 123.530 70.500 ;
        RECT 115.230 69.800 123.530 70.200 ;
        RECT 115.230 61.600 115.380 69.800 ;
        RECT 115.830 61.600 115.980 69.800 ;
        RECT 116.430 61.600 116.580 69.800 ;
        RECT 117.030 61.600 117.180 69.800 ;
        RECT 117.630 61.600 117.780 69.800 ;
        RECT 118.230 61.600 118.380 69.800 ;
        RECT 118.830 61.600 118.980 69.800 ;
        RECT 123.130 69.500 123.530 69.800 ;
        RECT 119.580 69.350 123.530 69.500 ;
        RECT 123.130 68.900 123.530 69.350 ;
        RECT 119.580 68.750 123.530 68.900 ;
        RECT 123.130 68.300 123.530 68.750 ;
        RECT 119.580 68.150 123.530 68.300 ;
        RECT 123.130 67.700 123.530 68.150 ;
        RECT 119.580 67.550 123.530 67.700 ;
        RECT 123.130 67.100 123.530 67.550 ;
        RECT 119.580 66.950 123.530 67.100 ;
        RECT 123.130 66.500 123.530 66.950 ;
        RECT 119.580 66.350 123.530 66.500 ;
        RECT 123.130 65.900 123.530 66.350 ;
        RECT 119.580 65.750 123.530 65.900 ;
        RECT 123.130 65.300 123.530 65.750 ;
        RECT 119.580 65.150 123.530 65.300 ;
        RECT 123.130 64.700 123.530 65.150 ;
        RECT 119.580 64.550 123.530 64.700 ;
        RECT 123.130 64.400 123.530 64.550 ;
        RECT 123.130 64.100 124.730 64.400 ;
        RECT 119.580 63.950 124.730 64.100 ;
        RECT 123.130 63.500 124.730 63.950 ;
        RECT 119.580 63.350 124.730 63.500 ;
        RECT 123.130 62.900 124.730 63.350 ;
        RECT 119.580 62.750 124.730 62.900 ;
        RECT 123.130 62.300 124.730 62.750 ;
        RECT 119.580 62.150 124.730 62.300 ;
        RECT 123.530 61.200 124.730 62.150 ;
        RECT 125.135 62.105 127.135 63.380 ;
        RECT 4.730 58.800 9.130 61.200 ;
        RECT 20.330 58.800 29.130 61.200 ;
        RECT 40.330 58.800 49.130 61.200 ;
        RECT 60.330 58.800 69.130 61.200 ;
        RECT 80.330 58.800 89.130 61.200 ;
        RECT 100.330 58.800 109.130 61.200 ;
        RECT 120.330 58.800 124.730 61.200 ;
        RECT 4.730 57.850 5.940 58.800 ;
        RECT 4.730 57.700 9.880 57.850 ;
        RECT 2.315 56.280 4.330 57.555 ;
        RECT 4.730 57.250 6.330 57.700 ;
        RECT 4.730 57.100 9.880 57.250 ;
        RECT 4.730 56.650 6.330 57.100 ;
        RECT 4.730 56.500 9.880 56.650 ;
        RECT 4.730 56.050 6.330 56.500 ;
        RECT 4.730 55.900 9.880 56.050 ;
        RECT 4.730 55.600 6.330 55.900 ;
        RECT 2.315 53.250 4.315 55.545 ;
        RECT 5.930 55.450 6.330 55.600 ;
        RECT 5.930 55.300 9.880 55.450 ;
        RECT 5.930 54.850 6.330 55.300 ;
        RECT 5.930 54.700 9.880 54.850 ;
        RECT 5.930 54.250 6.330 54.700 ;
        RECT 5.930 54.100 9.880 54.250 ;
        RECT 5.930 53.650 6.330 54.100 ;
        RECT 5.930 53.500 9.880 53.650 ;
        RECT 5.930 53.050 6.330 53.500 ;
        RECT 5.930 52.900 9.880 53.050 ;
        RECT 5.930 52.450 6.330 52.900 ;
        RECT 5.930 52.300 9.880 52.450 ;
        RECT 5.930 51.850 6.330 52.300 ;
        RECT 5.930 51.700 9.880 51.850 ;
        RECT 5.930 51.250 6.330 51.700 ;
        RECT 5.930 51.100 9.880 51.250 ;
        RECT 5.930 50.650 6.330 51.100 ;
        RECT 5.930 50.500 9.880 50.650 ;
        RECT 5.930 50.200 6.330 50.500 ;
        RECT 10.480 50.200 10.630 58.400 ;
        RECT 11.080 50.200 11.230 58.400 ;
        RECT 11.680 50.200 11.830 58.400 ;
        RECT 12.280 50.200 12.430 58.400 ;
        RECT 12.880 50.200 13.030 58.400 ;
        RECT 13.480 50.200 13.630 58.400 ;
        RECT 14.080 50.200 14.230 58.400 ;
        RECT 5.930 49.800 14.230 50.200 ;
        RECT 5.930 49.500 6.330 49.800 ;
        RECT 5.930 49.350 9.880 49.500 ;
        RECT 5.930 48.900 6.330 49.350 ;
        RECT 5.930 48.750 9.880 48.900 ;
        RECT 5.930 48.300 6.330 48.750 ;
        RECT 5.930 48.150 9.880 48.300 ;
        RECT 5.930 47.700 6.330 48.150 ;
        RECT 5.930 47.550 9.880 47.700 ;
        RECT 5.930 47.100 6.330 47.550 ;
        RECT 5.930 46.950 9.880 47.100 ;
        RECT 2.315 44.450 4.315 46.745 ;
        RECT 5.930 46.500 6.330 46.950 ;
        RECT 5.930 46.350 9.880 46.500 ;
        RECT 5.930 45.900 6.330 46.350 ;
        RECT 5.930 45.750 9.880 45.900 ;
        RECT 5.930 45.300 6.330 45.750 ;
        RECT 5.930 45.150 9.880 45.300 ;
        RECT 5.930 44.700 6.330 45.150 ;
        RECT 5.930 44.550 9.880 44.700 ;
        RECT 5.930 44.400 6.330 44.550 ;
        RECT 4.730 44.100 6.330 44.400 ;
        RECT 4.730 43.950 9.880 44.100 ;
        RECT 4.730 43.500 6.330 43.950 ;
        RECT 4.730 43.350 9.880 43.500 ;
        RECT 2.315 41.955 4.320 43.230 ;
        RECT 4.730 42.900 6.330 43.350 ;
        RECT 4.730 42.750 9.880 42.900 ;
        RECT 4.730 42.300 6.330 42.750 ;
        RECT 4.730 42.150 9.880 42.300 ;
        RECT 4.730 41.200 5.930 42.150 ;
        RECT 10.480 41.600 10.630 49.800 ;
        RECT 11.080 41.600 11.230 49.800 ;
        RECT 11.680 41.600 11.830 49.800 ;
        RECT 12.280 41.600 12.430 49.800 ;
        RECT 12.880 41.600 13.030 49.800 ;
        RECT 13.480 41.600 13.630 49.800 ;
        RECT 14.080 41.600 14.230 49.800 ;
        RECT 15.230 50.200 15.380 58.400 ;
        RECT 15.830 50.200 15.980 58.400 ;
        RECT 16.430 50.200 16.580 58.400 ;
        RECT 17.030 50.200 17.180 58.400 ;
        RECT 17.630 50.200 17.780 58.400 ;
        RECT 18.230 50.200 18.380 58.400 ;
        RECT 18.830 50.200 18.980 58.400 ;
        RECT 23.530 57.850 25.940 58.800 ;
        RECT 19.580 57.700 29.880 57.850 ;
        RECT 23.130 57.250 26.330 57.700 ;
        RECT 19.580 57.100 29.880 57.250 ;
        RECT 23.130 56.650 26.330 57.100 ;
        RECT 19.580 56.500 29.880 56.650 ;
        RECT 23.130 56.050 26.330 56.500 ;
        RECT 19.580 55.900 29.880 56.050 ;
        RECT 23.130 55.600 26.330 55.900 ;
        RECT 23.130 55.450 23.530 55.600 ;
        RECT 19.580 55.300 23.530 55.450 ;
        RECT 23.130 54.850 23.530 55.300 ;
        RECT 19.580 54.700 23.530 54.850 ;
        RECT 23.130 54.250 23.530 54.700 ;
        RECT 19.580 54.100 23.530 54.250 ;
        RECT 23.130 53.650 23.530 54.100 ;
        RECT 19.580 53.500 23.530 53.650 ;
        RECT 23.130 53.050 23.530 53.500 ;
        RECT 19.580 52.900 23.530 53.050 ;
        RECT 23.130 52.450 23.530 52.900 ;
        RECT 19.580 52.300 23.530 52.450 ;
        RECT 23.130 51.850 23.530 52.300 ;
        RECT 19.580 51.700 23.530 51.850 ;
        RECT 23.130 51.250 23.530 51.700 ;
        RECT 19.580 51.100 23.530 51.250 ;
        RECT 23.130 50.650 23.530 51.100 ;
        RECT 19.580 50.500 23.530 50.650 ;
        RECT 23.130 50.200 23.530 50.500 ;
        RECT 15.230 49.800 23.530 50.200 ;
        RECT 15.230 41.600 15.380 49.800 ;
        RECT 15.830 41.600 15.980 49.800 ;
        RECT 16.430 41.600 16.580 49.800 ;
        RECT 17.030 41.600 17.180 49.800 ;
        RECT 17.630 41.600 17.780 49.800 ;
        RECT 18.230 41.600 18.380 49.800 ;
        RECT 18.830 41.600 18.980 49.800 ;
        RECT 23.130 49.500 23.530 49.800 ;
        RECT 19.580 49.350 23.530 49.500 ;
        RECT 23.130 48.900 23.530 49.350 ;
        RECT 19.580 48.750 23.530 48.900 ;
        RECT 23.130 48.300 23.530 48.750 ;
        RECT 19.580 48.150 23.530 48.300 ;
        RECT 23.130 47.700 23.530 48.150 ;
        RECT 19.580 47.550 23.530 47.700 ;
        RECT 23.130 47.100 23.530 47.550 ;
        RECT 19.580 46.950 23.530 47.100 ;
        RECT 23.130 46.500 23.530 46.950 ;
        RECT 19.580 46.350 23.530 46.500 ;
        RECT 23.130 45.900 23.530 46.350 ;
        RECT 19.580 45.750 23.530 45.900 ;
        RECT 23.130 45.300 23.530 45.750 ;
        RECT 19.580 45.150 23.530 45.300 ;
        RECT 23.130 44.700 23.530 45.150 ;
        RECT 19.580 44.550 23.530 44.700 ;
        RECT 23.130 44.400 23.530 44.550 ;
        RECT 25.930 55.450 26.330 55.600 ;
        RECT 25.930 55.300 29.880 55.450 ;
        RECT 25.930 54.850 26.330 55.300 ;
        RECT 25.930 54.700 29.880 54.850 ;
        RECT 25.930 54.250 26.330 54.700 ;
        RECT 25.930 54.100 29.880 54.250 ;
        RECT 25.930 53.650 26.330 54.100 ;
        RECT 25.930 53.500 29.880 53.650 ;
        RECT 25.930 53.050 26.330 53.500 ;
        RECT 25.930 52.900 29.880 53.050 ;
        RECT 25.930 52.450 26.330 52.900 ;
        RECT 25.930 52.300 29.880 52.450 ;
        RECT 25.930 51.850 26.330 52.300 ;
        RECT 25.930 51.700 29.880 51.850 ;
        RECT 25.930 51.250 26.330 51.700 ;
        RECT 25.930 51.100 29.880 51.250 ;
        RECT 25.930 50.650 26.330 51.100 ;
        RECT 25.930 50.500 29.880 50.650 ;
        RECT 25.930 50.200 26.330 50.500 ;
        RECT 30.480 50.200 30.630 58.400 ;
        RECT 31.080 50.200 31.230 58.400 ;
        RECT 31.680 50.200 31.830 58.400 ;
        RECT 32.280 50.200 32.430 58.400 ;
        RECT 32.880 50.200 33.030 58.400 ;
        RECT 33.480 50.200 33.630 58.400 ;
        RECT 34.080 50.200 34.230 58.400 ;
        RECT 25.930 49.800 34.230 50.200 ;
        RECT 25.930 49.500 26.330 49.800 ;
        RECT 25.930 49.350 29.880 49.500 ;
        RECT 25.930 48.900 26.330 49.350 ;
        RECT 25.930 48.750 29.880 48.900 ;
        RECT 25.930 48.300 26.330 48.750 ;
        RECT 25.930 48.150 29.880 48.300 ;
        RECT 25.930 47.700 26.330 48.150 ;
        RECT 25.930 47.550 29.880 47.700 ;
        RECT 25.930 47.100 26.330 47.550 ;
        RECT 25.930 46.950 29.880 47.100 ;
        RECT 25.930 46.500 26.330 46.950 ;
        RECT 25.930 46.350 29.880 46.500 ;
        RECT 25.930 45.900 26.330 46.350 ;
        RECT 25.930 45.750 29.880 45.900 ;
        RECT 25.930 45.300 26.330 45.750 ;
        RECT 25.930 45.150 29.880 45.300 ;
        RECT 25.930 44.700 26.330 45.150 ;
        RECT 25.930 44.550 29.880 44.700 ;
        RECT 25.930 44.400 26.330 44.550 ;
        RECT 23.130 44.100 26.330 44.400 ;
        RECT 19.580 43.950 29.880 44.100 ;
        RECT 23.130 43.500 26.330 43.950 ;
        RECT 19.580 43.350 29.880 43.500 ;
        RECT 23.130 42.900 26.330 43.350 ;
        RECT 19.580 42.750 29.880 42.900 ;
        RECT 23.130 42.300 26.330 42.750 ;
        RECT 19.580 42.150 29.880 42.300 ;
        RECT 23.530 41.200 25.930 42.150 ;
        RECT 30.480 41.600 30.630 49.800 ;
        RECT 31.080 41.600 31.230 49.800 ;
        RECT 31.680 41.600 31.830 49.800 ;
        RECT 32.280 41.600 32.430 49.800 ;
        RECT 32.880 41.600 33.030 49.800 ;
        RECT 33.480 41.600 33.630 49.800 ;
        RECT 34.080 41.600 34.230 49.800 ;
        RECT 35.230 50.200 35.380 58.400 ;
        RECT 35.830 50.200 35.980 58.400 ;
        RECT 36.430 50.200 36.580 58.400 ;
        RECT 37.030 50.200 37.180 58.400 ;
        RECT 37.630 50.200 37.780 58.400 ;
        RECT 38.230 50.200 38.380 58.400 ;
        RECT 38.830 50.200 38.980 58.400 ;
        RECT 43.530 57.850 45.940 58.800 ;
        RECT 39.580 57.700 49.880 57.850 ;
        RECT 43.130 57.250 46.330 57.700 ;
        RECT 39.580 57.100 49.880 57.250 ;
        RECT 43.130 56.650 46.330 57.100 ;
        RECT 39.580 56.500 49.880 56.650 ;
        RECT 43.130 56.050 46.330 56.500 ;
        RECT 39.580 55.900 49.880 56.050 ;
        RECT 43.130 55.600 46.330 55.900 ;
        RECT 43.130 55.450 43.530 55.600 ;
        RECT 39.580 55.300 43.530 55.450 ;
        RECT 43.130 54.850 43.530 55.300 ;
        RECT 39.580 54.700 43.530 54.850 ;
        RECT 43.130 54.250 43.530 54.700 ;
        RECT 39.580 54.100 43.530 54.250 ;
        RECT 43.130 53.650 43.530 54.100 ;
        RECT 39.580 53.500 43.530 53.650 ;
        RECT 43.130 53.050 43.530 53.500 ;
        RECT 39.580 52.900 43.530 53.050 ;
        RECT 43.130 52.450 43.530 52.900 ;
        RECT 39.580 52.300 43.530 52.450 ;
        RECT 43.130 51.850 43.530 52.300 ;
        RECT 39.580 51.700 43.530 51.850 ;
        RECT 43.130 51.250 43.530 51.700 ;
        RECT 39.580 51.100 43.530 51.250 ;
        RECT 43.130 50.650 43.530 51.100 ;
        RECT 39.580 50.500 43.530 50.650 ;
        RECT 43.130 50.200 43.530 50.500 ;
        RECT 35.230 49.800 43.530 50.200 ;
        RECT 35.230 41.600 35.380 49.800 ;
        RECT 35.830 41.600 35.980 49.800 ;
        RECT 36.430 41.600 36.580 49.800 ;
        RECT 37.030 41.600 37.180 49.800 ;
        RECT 37.630 41.600 37.780 49.800 ;
        RECT 38.230 41.600 38.380 49.800 ;
        RECT 38.830 41.600 38.980 49.800 ;
        RECT 43.130 49.500 43.530 49.800 ;
        RECT 39.580 49.350 43.530 49.500 ;
        RECT 43.130 48.900 43.530 49.350 ;
        RECT 39.580 48.750 43.530 48.900 ;
        RECT 43.130 48.300 43.530 48.750 ;
        RECT 39.580 48.150 43.530 48.300 ;
        RECT 43.130 47.700 43.530 48.150 ;
        RECT 39.580 47.550 43.530 47.700 ;
        RECT 43.130 47.100 43.530 47.550 ;
        RECT 39.580 46.950 43.530 47.100 ;
        RECT 43.130 46.500 43.530 46.950 ;
        RECT 39.580 46.350 43.530 46.500 ;
        RECT 43.130 45.900 43.530 46.350 ;
        RECT 39.580 45.750 43.530 45.900 ;
        RECT 43.130 45.300 43.530 45.750 ;
        RECT 39.580 45.150 43.530 45.300 ;
        RECT 43.130 44.700 43.530 45.150 ;
        RECT 39.580 44.550 43.530 44.700 ;
        RECT 43.130 44.400 43.530 44.550 ;
        RECT 45.930 55.450 46.330 55.600 ;
        RECT 45.930 55.300 49.880 55.450 ;
        RECT 45.930 54.850 46.330 55.300 ;
        RECT 45.930 54.700 49.880 54.850 ;
        RECT 45.930 54.250 46.330 54.700 ;
        RECT 45.930 54.100 49.880 54.250 ;
        RECT 45.930 53.650 46.330 54.100 ;
        RECT 45.930 53.500 49.880 53.650 ;
        RECT 45.930 53.050 46.330 53.500 ;
        RECT 45.930 52.900 49.880 53.050 ;
        RECT 45.930 52.450 46.330 52.900 ;
        RECT 45.930 52.300 49.880 52.450 ;
        RECT 45.930 51.850 46.330 52.300 ;
        RECT 45.930 51.700 49.880 51.850 ;
        RECT 45.930 51.250 46.330 51.700 ;
        RECT 45.930 51.100 49.880 51.250 ;
        RECT 45.930 50.650 46.330 51.100 ;
        RECT 45.930 50.500 49.880 50.650 ;
        RECT 45.930 50.200 46.330 50.500 ;
        RECT 50.480 50.200 50.630 58.400 ;
        RECT 51.080 50.200 51.230 58.400 ;
        RECT 51.680 50.200 51.830 58.400 ;
        RECT 52.280 50.200 52.430 58.400 ;
        RECT 52.880 50.200 53.030 58.400 ;
        RECT 53.480 50.200 53.630 58.400 ;
        RECT 54.080 50.200 54.230 58.400 ;
        RECT 45.930 49.800 54.230 50.200 ;
        RECT 45.930 49.500 46.330 49.800 ;
        RECT 45.930 49.350 49.880 49.500 ;
        RECT 45.930 48.900 46.330 49.350 ;
        RECT 45.930 48.750 49.880 48.900 ;
        RECT 45.930 48.300 46.330 48.750 ;
        RECT 45.930 48.150 49.880 48.300 ;
        RECT 45.930 47.700 46.330 48.150 ;
        RECT 45.930 47.550 49.880 47.700 ;
        RECT 45.930 47.100 46.330 47.550 ;
        RECT 45.930 46.950 49.880 47.100 ;
        RECT 45.930 46.500 46.330 46.950 ;
        RECT 45.930 46.350 49.880 46.500 ;
        RECT 45.930 45.900 46.330 46.350 ;
        RECT 45.930 45.750 49.880 45.900 ;
        RECT 45.930 45.300 46.330 45.750 ;
        RECT 45.930 45.150 49.880 45.300 ;
        RECT 45.930 44.700 46.330 45.150 ;
        RECT 45.930 44.550 49.880 44.700 ;
        RECT 45.930 44.400 46.330 44.550 ;
        RECT 43.130 44.100 46.330 44.400 ;
        RECT 39.580 43.950 49.880 44.100 ;
        RECT 43.130 43.500 46.330 43.950 ;
        RECT 39.580 43.350 49.880 43.500 ;
        RECT 43.130 42.900 46.330 43.350 ;
        RECT 39.580 42.750 49.880 42.900 ;
        RECT 43.130 42.300 46.330 42.750 ;
        RECT 39.580 42.150 49.880 42.300 ;
        RECT 43.530 41.200 45.930 42.150 ;
        RECT 50.480 41.600 50.630 49.800 ;
        RECT 51.080 41.600 51.230 49.800 ;
        RECT 51.680 41.600 51.830 49.800 ;
        RECT 52.280 41.600 52.430 49.800 ;
        RECT 52.880 41.600 53.030 49.800 ;
        RECT 53.480 41.600 53.630 49.800 ;
        RECT 54.080 41.600 54.230 49.800 ;
        RECT 55.230 50.200 55.380 58.400 ;
        RECT 55.830 50.200 55.980 58.400 ;
        RECT 56.430 50.200 56.580 58.400 ;
        RECT 57.030 50.200 57.180 58.400 ;
        RECT 57.630 50.200 57.780 58.400 ;
        RECT 58.230 50.200 58.380 58.400 ;
        RECT 58.830 50.200 58.980 58.400 ;
        RECT 63.530 57.850 65.940 58.800 ;
        RECT 59.580 57.700 69.880 57.850 ;
        RECT 63.130 57.250 66.330 57.700 ;
        RECT 59.580 57.100 69.880 57.250 ;
        RECT 63.130 56.650 66.330 57.100 ;
        RECT 59.580 56.500 69.880 56.650 ;
        RECT 63.130 56.050 66.330 56.500 ;
        RECT 59.580 55.900 69.880 56.050 ;
        RECT 63.130 55.600 66.330 55.900 ;
        RECT 63.130 55.450 63.530 55.600 ;
        RECT 59.580 55.300 63.530 55.450 ;
        RECT 63.130 54.850 63.530 55.300 ;
        RECT 59.580 54.700 63.530 54.850 ;
        RECT 63.130 54.250 63.530 54.700 ;
        RECT 59.580 54.100 63.530 54.250 ;
        RECT 63.130 53.650 63.530 54.100 ;
        RECT 59.580 53.500 63.530 53.650 ;
        RECT 63.130 53.050 63.530 53.500 ;
        RECT 59.580 52.900 63.530 53.050 ;
        RECT 63.130 52.450 63.530 52.900 ;
        RECT 59.580 52.300 63.530 52.450 ;
        RECT 63.130 51.850 63.530 52.300 ;
        RECT 59.580 51.700 63.530 51.850 ;
        RECT 63.130 51.250 63.530 51.700 ;
        RECT 59.580 51.100 63.530 51.250 ;
        RECT 63.130 50.650 63.530 51.100 ;
        RECT 59.580 50.500 63.530 50.650 ;
        RECT 63.130 50.200 63.530 50.500 ;
        RECT 55.230 49.800 63.530 50.200 ;
        RECT 55.230 41.600 55.380 49.800 ;
        RECT 55.830 41.600 55.980 49.800 ;
        RECT 56.430 41.600 56.580 49.800 ;
        RECT 57.030 41.600 57.180 49.800 ;
        RECT 57.630 41.600 57.780 49.800 ;
        RECT 58.230 41.600 58.380 49.800 ;
        RECT 58.830 41.600 58.980 49.800 ;
        RECT 63.130 49.500 63.530 49.800 ;
        RECT 59.580 49.350 63.530 49.500 ;
        RECT 63.130 48.900 63.530 49.350 ;
        RECT 59.580 48.750 63.530 48.900 ;
        RECT 63.130 48.300 63.530 48.750 ;
        RECT 59.580 48.150 63.530 48.300 ;
        RECT 63.130 47.700 63.530 48.150 ;
        RECT 59.580 47.550 63.530 47.700 ;
        RECT 63.130 47.100 63.530 47.550 ;
        RECT 59.580 46.950 63.530 47.100 ;
        RECT 63.130 46.500 63.530 46.950 ;
        RECT 59.580 46.350 63.530 46.500 ;
        RECT 63.130 45.900 63.530 46.350 ;
        RECT 59.580 45.750 63.530 45.900 ;
        RECT 63.130 45.300 63.530 45.750 ;
        RECT 59.580 45.150 63.530 45.300 ;
        RECT 63.130 44.700 63.530 45.150 ;
        RECT 59.580 44.550 63.530 44.700 ;
        RECT 63.130 44.400 63.530 44.550 ;
        RECT 65.930 55.450 66.330 55.600 ;
        RECT 65.930 55.300 69.880 55.450 ;
        RECT 65.930 54.850 66.330 55.300 ;
        RECT 65.930 54.700 69.880 54.850 ;
        RECT 65.930 54.250 66.330 54.700 ;
        RECT 65.930 54.100 69.880 54.250 ;
        RECT 65.930 53.650 66.330 54.100 ;
        RECT 65.930 53.500 69.880 53.650 ;
        RECT 65.930 53.050 66.330 53.500 ;
        RECT 65.930 52.900 69.880 53.050 ;
        RECT 65.930 52.450 66.330 52.900 ;
        RECT 65.930 52.300 69.880 52.450 ;
        RECT 65.930 51.850 66.330 52.300 ;
        RECT 65.930 51.700 69.880 51.850 ;
        RECT 65.930 51.250 66.330 51.700 ;
        RECT 65.930 51.100 69.880 51.250 ;
        RECT 65.930 50.650 66.330 51.100 ;
        RECT 65.930 50.500 69.880 50.650 ;
        RECT 65.930 50.200 66.330 50.500 ;
        RECT 70.480 50.200 70.630 58.400 ;
        RECT 71.080 50.200 71.230 58.400 ;
        RECT 71.680 50.200 71.830 58.400 ;
        RECT 72.280 50.200 72.430 58.400 ;
        RECT 72.880 50.200 73.030 58.400 ;
        RECT 73.480 50.200 73.630 58.400 ;
        RECT 74.080 50.200 74.230 58.400 ;
        RECT 65.930 49.800 74.230 50.200 ;
        RECT 65.930 49.500 66.330 49.800 ;
        RECT 65.930 49.350 69.880 49.500 ;
        RECT 65.930 48.900 66.330 49.350 ;
        RECT 65.930 48.750 69.880 48.900 ;
        RECT 65.930 48.300 66.330 48.750 ;
        RECT 65.930 48.150 69.880 48.300 ;
        RECT 65.930 47.700 66.330 48.150 ;
        RECT 65.930 47.550 69.880 47.700 ;
        RECT 65.930 47.100 66.330 47.550 ;
        RECT 65.930 46.950 69.880 47.100 ;
        RECT 65.930 46.500 66.330 46.950 ;
        RECT 65.930 46.350 69.880 46.500 ;
        RECT 65.930 45.900 66.330 46.350 ;
        RECT 65.930 45.750 69.880 45.900 ;
        RECT 65.930 45.300 66.330 45.750 ;
        RECT 65.930 45.150 69.880 45.300 ;
        RECT 65.930 44.700 66.330 45.150 ;
        RECT 65.930 44.550 69.880 44.700 ;
        RECT 65.930 44.400 66.330 44.550 ;
        RECT 63.130 44.100 66.330 44.400 ;
        RECT 59.580 43.950 69.880 44.100 ;
        RECT 63.130 43.500 66.330 43.950 ;
        RECT 59.580 43.350 69.880 43.500 ;
        RECT 63.130 42.900 66.330 43.350 ;
        RECT 59.580 42.750 69.880 42.900 ;
        RECT 63.130 42.300 66.330 42.750 ;
        RECT 59.580 42.150 69.880 42.300 ;
        RECT 63.530 41.200 65.930 42.150 ;
        RECT 70.480 41.600 70.630 49.800 ;
        RECT 71.080 41.600 71.230 49.800 ;
        RECT 71.680 41.600 71.830 49.800 ;
        RECT 72.280 41.600 72.430 49.800 ;
        RECT 72.880 41.600 73.030 49.800 ;
        RECT 73.480 41.600 73.630 49.800 ;
        RECT 74.080 41.600 74.230 49.800 ;
        RECT 75.230 50.200 75.380 58.400 ;
        RECT 75.830 50.200 75.980 58.400 ;
        RECT 76.430 50.200 76.580 58.400 ;
        RECT 77.030 50.200 77.180 58.400 ;
        RECT 77.630 50.200 77.780 58.400 ;
        RECT 78.230 50.200 78.380 58.400 ;
        RECT 78.830 50.200 78.980 58.400 ;
        RECT 83.530 57.850 85.940 58.800 ;
        RECT 79.580 57.700 89.880 57.850 ;
        RECT 83.130 57.250 86.330 57.700 ;
        RECT 79.580 57.100 89.880 57.250 ;
        RECT 83.130 56.650 86.330 57.100 ;
        RECT 79.580 56.500 89.880 56.650 ;
        RECT 83.130 56.050 86.330 56.500 ;
        RECT 79.580 55.900 89.880 56.050 ;
        RECT 83.130 55.600 86.330 55.900 ;
        RECT 83.130 55.450 83.530 55.600 ;
        RECT 79.580 55.300 83.530 55.450 ;
        RECT 83.130 54.850 83.530 55.300 ;
        RECT 79.580 54.700 83.530 54.850 ;
        RECT 83.130 54.250 83.530 54.700 ;
        RECT 79.580 54.100 83.530 54.250 ;
        RECT 83.130 53.650 83.530 54.100 ;
        RECT 79.580 53.500 83.530 53.650 ;
        RECT 83.130 53.050 83.530 53.500 ;
        RECT 79.580 52.900 83.530 53.050 ;
        RECT 83.130 52.450 83.530 52.900 ;
        RECT 79.580 52.300 83.530 52.450 ;
        RECT 83.130 51.850 83.530 52.300 ;
        RECT 79.580 51.700 83.530 51.850 ;
        RECT 83.130 51.250 83.530 51.700 ;
        RECT 79.580 51.100 83.530 51.250 ;
        RECT 83.130 50.650 83.530 51.100 ;
        RECT 79.580 50.500 83.530 50.650 ;
        RECT 83.130 50.200 83.530 50.500 ;
        RECT 75.230 49.800 83.530 50.200 ;
        RECT 75.230 41.600 75.380 49.800 ;
        RECT 75.830 41.600 75.980 49.800 ;
        RECT 76.430 41.600 76.580 49.800 ;
        RECT 77.030 41.600 77.180 49.800 ;
        RECT 77.630 41.600 77.780 49.800 ;
        RECT 78.230 41.600 78.380 49.800 ;
        RECT 78.830 41.600 78.980 49.800 ;
        RECT 83.130 49.500 83.530 49.800 ;
        RECT 79.580 49.350 83.530 49.500 ;
        RECT 83.130 48.900 83.530 49.350 ;
        RECT 79.580 48.750 83.530 48.900 ;
        RECT 83.130 48.300 83.530 48.750 ;
        RECT 79.580 48.150 83.530 48.300 ;
        RECT 83.130 47.700 83.530 48.150 ;
        RECT 79.580 47.550 83.530 47.700 ;
        RECT 83.130 47.100 83.530 47.550 ;
        RECT 79.580 46.950 83.530 47.100 ;
        RECT 83.130 46.500 83.530 46.950 ;
        RECT 79.580 46.350 83.530 46.500 ;
        RECT 83.130 45.900 83.530 46.350 ;
        RECT 79.580 45.750 83.530 45.900 ;
        RECT 83.130 45.300 83.530 45.750 ;
        RECT 79.580 45.150 83.530 45.300 ;
        RECT 83.130 44.700 83.530 45.150 ;
        RECT 79.580 44.550 83.530 44.700 ;
        RECT 83.130 44.400 83.530 44.550 ;
        RECT 85.930 55.450 86.330 55.600 ;
        RECT 85.930 55.300 89.880 55.450 ;
        RECT 85.930 54.850 86.330 55.300 ;
        RECT 85.930 54.700 89.880 54.850 ;
        RECT 85.930 54.250 86.330 54.700 ;
        RECT 85.930 54.100 89.880 54.250 ;
        RECT 85.930 53.650 86.330 54.100 ;
        RECT 85.930 53.500 89.880 53.650 ;
        RECT 85.930 53.050 86.330 53.500 ;
        RECT 85.930 52.900 89.880 53.050 ;
        RECT 85.930 52.450 86.330 52.900 ;
        RECT 85.930 52.300 89.880 52.450 ;
        RECT 85.930 51.850 86.330 52.300 ;
        RECT 85.930 51.700 89.880 51.850 ;
        RECT 85.930 51.250 86.330 51.700 ;
        RECT 85.930 51.100 89.880 51.250 ;
        RECT 85.930 50.650 86.330 51.100 ;
        RECT 85.930 50.500 89.880 50.650 ;
        RECT 85.930 50.200 86.330 50.500 ;
        RECT 90.480 50.200 90.630 58.400 ;
        RECT 91.080 50.200 91.230 58.400 ;
        RECT 91.680 50.200 91.830 58.400 ;
        RECT 92.280 50.200 92.430 58.400 ;
        RECT 92.880 50.200 93.030 58.400 ;
        RECT 93.480 50.200 93.630 58.400 ;
        RECT 94.080 50.200 94.230 58.400 ;
        RECT 85.930 49.800 94.230 50.200 ;
        RECT 85.930 49.500 86.330 49.800 ;
        RECT 85.930 49.350 89.880 49.500 ;
        RECT 85.930 48.900 86.330 49.350 ;
        RECT 85.930 48.750 89.880 48.900 ;
        RECT 85.930 48.300 86.330 48.750 ;
        RECT 85.930 48.150 89.880 48.300 ;
        RECT 85.930 47.700 86.330 48.150 ;
        RECT 85.930 47.550 89.880 47.700 ;
        RECT 85.930 47.100 86.330 47.550 ;
        RECT 85.930 46.950 89.880 47.100 ;
        RECT 85.930 46.500 86.330 46.950 ;
        RECT 85.930 46.350 89.880 46.500 ;
        RECT 85.930 45.900 86.330 46.350 ;
        RECT 85.930 45.750 89.880 45.900 ;
        RECT 85.930 45.300 86.330 45.750 ;
        RECT 85.930 45.150 89.880 45.300 ;
        RECT 85.930 44.700 86.330 45.150 ;
        RECT 85.930 44.550 89.880 44.700 ;
        RECT 85.930 44.400 86.330 44.550 ;
        RECT 83.130 44.100 86.330 44.400 ;
        RECT 79.580 43.950 89.880 44.100 ;
        RECT 83.130 43.500 86.330 43.950 ;
        RECT 79.580 43.350 89.880 43.500 ;
        RECT 83.130 42.900 86.330 43.350 ;
        RECT 79.580 42.750 89.880 42.900 ;
        RECT 83.130 42.300 86.330 42.750 ;
        RECT 79.580 42.150 89.880 42.300 ;
        RECT 83.530 41.200 85.930 42.150 ;
        RECT 90.480 41.600 90.630 49.800 ;
        RECT 91.080 41.600 91.230 49.800 ;
        RECT 91.680 41.600 91.830 49.800 ;
        RECT 92.280 41.600 92.430 49.800 ;
        RECT 92.880 41.600 93.030 49.800 ;
        RECT 93.480 41.600 93.630 49.800 ;
        RECT 94.080 41.600 94.230 49.800 ;
        RECT 95.230 50.200 95.380 58.400 ;
        RECT 95.830 50.200 95.980 58.400 ;
        RECT 96.430 50.200 96.580 58.400 ;
        RECT 97.030 50.200 97.180 58.400 ;
        RECT 97.630 50.200 97.780 58.400 ;
        RECT 98.230 50.200 98.380 58.400 ;
        RECT 98.830 50.200 98.980 58.400 ;
        RECT 103.530 57.850 105.940 58.800 ;
        RECT 99.580 57.700 109.880 57.850 ;
        RECT 103.130 57.250 106.330 57.700 ;
        RECT 99.580 57.100 109.880 57.250 ;
        RECT 103.130 56.650 106.330 57.100 ;
        RECT 99.580 56.500 109.880 56.650 ;
        RECT 103.130 56.050 106.330 56.500 ;
        RECT 99.580 55.900 109.880 56.050 ;
        RECT 103.130 55.600 106.330 55.900 ;
        RECT 103.130 55.450 103.530 55.600 ;
        RECT 99.580 55.300 103.530 55.450 ;
        RECT 103.130 54.850 103.530 55.300 ;
        RECT 99.580 54.700 103.530 54.850 ;
        RECT 103.130 54.250 103.530 54.700 ;
        RECT 99.580 54.100 103.530 54.250 ;
        RECT 103.130 53.650 103.530 54.100 ;
        RECT 99.580 53.500 103.530 53.650 ;
        RECT 103.130 53.050 103.530 53.500 ;
        RECT 99.580 52.900 103.530 53.050 ;
        RECT 103.130 52.450 103.530 52.900 ;
        RECT 99.580 52.300 103.530 52.450 ;
        RECT 103.130 51.850 103.530 52.300 ;
        RECT 99.580 51.700 103.530 51.850 ;
        RECT 103.130 51.250 103.530 51.700 ;
        RECT 99.580 51.100 103.530 51.250 ;
        RECT 103.130 50.650 103.530 51.100 ;
        RECT 99.580 50.500 103.530 50.650 ;
        RECT 103.130 50.200 103.530 50.500 ;
        RECT 95.230 49.800 103.530 50.200 ;
        RECT 95.230 41.600 95.380 49.800 ;
        RECT 95.830 41.600 95.980 49.800 ;
        RECT 96.430 41.600 96.580 49.800 ;
        RECT 97.030 41.600 97.180 49.800 ;
        RECT 97.630 41.600 97.780 49.800 ;
        RECT 98.230 41.600 98.380 49.800 ;
        RECT 98.830 41.600 98.980 49.800 ;
        RECT 103.130 49.500 103.530 49.800 ;
        RECT 99.580 49.350 103.530 49.500 ;
        RECT 103.130 48.900 103.530 49.350 ;
        RECT 99.580 48.750 103.530 48.900 ;
        RECT 103.130 48.300 103.530 48.750 ;
        RECT 99.580 48.150 103.530 48.300 ;
        RECT 103.130 47.700 103.530 48.150 ;
        RECT 99.580 47.550 103.530 47.700 ;
        RECT 103.130 47.100 103.530 47.550 ;
        RECT 99.580 46.950 103.530 47.100 ;
        RECT 103.130 46.500 103.530 46.950 ;
        RECT 99.580 46.350 103.530 46.500 ;
        RECT 103.130 45.900 103.530 46.350 ;
        RECT 99.580 45.750 103.530 45.900 ;
        RECT 103.130 45.300 103.530 45.750 ;
        RECT 99.580 45.150 103.530 45.300 ;
        RECT 103.130 44.700 103.530 45.150 ;
        RECT 99.580 44.550 103.530 44.700 ;
        RECT 103.130 44.400 103.530 44.550 ;
        RECT 105.930 55.450 106.330 55.600 ;
        RECT 105.930 55.300 109.880 55.450 ;
        RECT 105.930 54.850 106.330 55.300 ;
        RECT 105.930 54.700 109.880 54.850 ;
        RECT 105.930 54.250 106.330 54.700 ;
        RECT 105.930 54.100 109.880 54.250 ;
        RECT 105.930 53.650 106.330 54.100 ;
        RECT 105.930 53.500 109.880 53.650 ;
        RECT 105.930 53.050 106.330 53.500 ;
        RECT 105.930 52.900 109.880 53.050 ;
        RECT 105.930 52.450 106.330 52.900 ;
        RECT 105.930 52.300 109.880 52.450 ;
        RECT 105.930 51.850 106.330 52.300 ;
        RECT 105.930 51.700 109.880 51.850 ;
        RECT 105.930 51.250 106.330 51.700 ;
        RECT 105.930 51.100 109.880 51.250 ;
        RECT 105.930 50.650 106.330 51.100 ;
        RECT 105.930 50.500 109.880 50.650 ;
        RECT 105.930 50.200 106.330 50.500 ;
        RECT 110.480 50.200 110.630 58.400 ;
        RECT 111.080 50.200 111.230 58.400 ;
        RECT 111.680 50.200 111.830 58.400 ;
        RECT 112.280 50.200 112.430 58.400 ;
        RECT 112.880 50.200 113.030 58.400 ;
        RECT 113.480 50.200 113.630 58.400 ;
        RECT 114.080 50.200 114.230 58.400 ;
        RECT 105.930 49.800 114.230 50.200 ;
        RECT 105.930 49.500 106.330 49.800 ;
        RECT 105.930 49.350 109.880 49.500 ;
        RECT 105.930 48.900 106.330 49.350 ;
        RECT 105.930 48.750 109.880 48.900 ;
        RECT 105.930 48.300 106.330 48.750 ;
        RECT 105.930 48.150 109.880 48.300 ;
        RECT 105.930 47.700 106.330 48.150 ;
        RECT 105.930 47.550 109.880 47.700 ;
        RECT 105.930 47.100 106.330 47.550 ;
        RECT 105.930 46.950 109.880 47.100 ;
        RECT 105.930 46.500 106.330 46.950 ;
        RECT 105.930 46.350 109.880 46.500 ;
        RECT 105.930 45.900 106.330 46.350 ;
        RECT 105.930 45.750 109.880 45.900 ;
        RECT 105.930 45.300 106.330 45.750 ;
        RECT 105.930 45.150 109.880 45.300 ;
        RECT 105.930 44.700 106.330 45.150 ;
        RECT 105.930 44.550 109.880 44.700 ;
        RECT 105.930 44.400 106.330 44.550 ;
        RECT 103.130 44.100 106.330 44.400 ;
        RECT 99.580 43.950 109.880 44.100 ;
        RECT 103.130 43.500 106.330 43.950 ;
        RECT 99.580 43.350 109.880 43.500 ;
        RECT 103.130 42.900 106.330 43.350 ;
        RECT 99.580 42.750 109.880 42.900 ;
        RECT 103.130 42.300 106.330 42.750 ;
        RECT 99.580 42.150 109.880 42.300 ;
        RECT 103.530 41.200 105.930 42.150 ;
        RECT 110.480 41.600 110.630 49.800 ;
        RECT 111.080 41.600 111.230 49.800 ;
        RECT 111.680 41.600 111.830 49.800 ;
        RECT 112.280 41.600 112.430 49.800 ;
        RECT 112.880 41.600 113.030 49.800 ;
        RECT 113.480 41.600 113.630 49.800 ;
        RECT 114.080 41.600 114.230 49.800 ;
        RECT 115.230 50.200 115.380 58.400 ;
        RECT 115.830 50.200 115.980 58.400 ;
        RECT 116.430 50.200 116.580 58.400 ;
        RECT 117.030 50.200 117.180 58.400 ;
        RECT 117.630 50.200 117.780 58.400 ;
        RECT 118.230 50.200 118.380 58.400 ;
        RECT 118.830 50.200 118.980 58.400 ;
        RECT 123.530 57.850 124.730 58.800 ;
        RECT 119.580 57.700 124.730 57.850 ;
        RECT 123.130 57.250 124.730 57.700 ;
        RECT 119.580 57.100 124.730 57.250 ;
        RECT 123.130 56.650 124.730 57.100 ;
        RECT 119.580 56.500 124.730 56.650 ;
        RECT 123.130 56.050 124.730 56.500 ;
        RECT 119.580 55.900 124.730 56.050 ;
        RECT 125.135 56.035 127.135 57.310 ;
        RECT 123.130 55.600 124.730 55.900 ;
        RECT 123.130 55.450 123.530 55.600 ;
        RECT 119.580 55.300 123.530 55.450 ;
        RECT 123.130 54.850 123.530 55.300 ;
        RECT 119.580 54.700 123.530 54.850 ;
        RECT 123.130 54.250 123.530 54.700 ;
        RECT 119.580 54.100 123.530 54.250 ;
        RECT 123.130 53.650 123.530 54.100 ;
        RECT 119.580 53.500 123.530 53.650 ;
        RECT 123.130 53.050 123.530 53.500 ;
        RECT 119.580 52.900 123.530 53.050 ;
        RECT 123.130 52.450 123.530 52.900 ;
        RECT 119.580 52.300 123.530 52.450 ;
        RECT 123.130 51.850 123.530 52.300 ;
        RECT 119.580 51.700 123.530 51.850 ;
        RECT 123.130 51.250 123.530 51.700 ;
        RECT 119.580 51.100 123.530 51.250 ;
        RECT 123.130 50.650 123.530 51.100 ;
        RECT 119.580 50.500 123.530 50.650 ;
        RECT 123.130 50.200 123.530 50.500 ;
        RECT 115.230 49.800 123.530 50.200 ;
        RECT 115.230 41.600 115.380 49.800 ;
        RECT 115.830 41.600 115.980 49.800 ;
        RECT 116.430 41.600 116.580 49.800 ;
        RECT 117.030 41.600 117.180 49.800 ;
        RECT 117.630 41.600 117.780 49.800 ;
        RECT 118.230 41.600 118.380 49.800 ;
        RECT 118.830 41.600 118.980 49.800 ;
        RECT 123.130 49.500 123.530 49.800 ;
        RECT 119.580 49.350 123.530 49.500 ;
        RECT 123.130 48.900 123.530 49.350 ;
        RECT 119.580 48.750 123.530 48.900 ;
        RECT 123.130 48.300 123.530 48.750 ;
        RECT 119.580 48.150 123.530 48.300 ;
        RECT 123.130 47.700 123.530 48.150 ;
        RECT 119.580 47.550 123.530 47.700 ;
        RECT 123.130 47.100 123.530 47.550 ;
        RECT 119.580 46.950 123.530 47.100 ;
        RECT 123.130 46.500 123.530 46.950 ;
        RECT 119.580 46.350 123.530 46.500 ;
        RECT 123.130 45.900 123.530 46.350 ;
        RECT 119.580 45.750 123.530 45.900 ;
        RECT 123.130 45.300 123.530 45.750 ;
        RECT 119.580 45.150 123.530 45.300 ;
        RECT 123.130 44.700 123.530 45.150 ;
        RECT 119.580 44.550 123.530 44.700 ;
        RECT 123.130 44.400 123.530 44.550 ;
        RECT 123.130 44.100 124.730 44.400 ;
        RECT 119.580 43.950 124.730 44.100 ;
        RECT 123.130 43.500 124.730 43.950 ;
        RECT 119.580 43.350 124.730 43.500 ;
        RECT 123.130 42.900 124.730 43.350 ;
        RECT 119.580 42.750 124.730 42.900 ;
        RECT 123.130 42.300 124.730 42.750 ;
        RECT 119.580 42.150 124.730 42.300 ;
        RECT 123.530 41.200 124.730 42.150 ;
        RECT 125.140 41.820 127.140 43.095 ;
        RECT 4.730 38.800 9.130 41.200 ;
        RECT 20.330 38.800 29.130 41.200 ;
        RECT 40.330 38.800 49.130 41.200 ;
        RECT 60.330 38.800 69.130 41.200 ;
        RECT 80.330 38.800 89.130 41.200 ;
        RECT 100.330 38.800 109.130 41.200 ;
        RECT 120.330 38.800 124.730 41.200 ;
        RECT 4.730 37.850 5.940 38.800 ;
        RECT 4.730 37.700 9.880 37.850 ;
        RECT 2.315 36.345 4.320 37.620 ;
        RECT 4.730 37.250 6.330 37.700 ;
        RECT 4.730 37.100 9.880 37.250 ;
        RECT 4.730 36.650 6.330 37.100 ;
        RECT 4.730 36.500 9.880 36.650 ;
        RECT 4.730 36.050 6.330 36.500 ;
        RECT 4.730 35.900 9.880 36.050 ;
        RECT 4.730 35.600 6.330 35.900 ;
        RECT 2.315 33.255 4.315 35.550 ;
        RECT 5.930 35.450 6.330 35.600 ;
        RECT 5.930 35.300 9.880 35.450 ;
        RECT 5.930 34.850 6.330 35.300 ;
        RECT 5.930 34.700 9.880 34.850 ;
        RECT 5.930 34.250 6.330 34.700 ;
        RECT 5.930 34.100 9.880 34.250 ;
        RECT 5.930 33.650 6.330 34.100 ;
        RECT 5.930 33.500 9.880 33.650 ;
        RECT 5.930 33.050 6.330 33.500 ;
        RECT 5.930 32.900 9.880 33.050 ;
        RECT 5.930 32.450 6.330 32.900 ;
        RECT 5.930 32.300 9.880 32.450 ;
        RECT 5.930 31.850 6.330 32.300 ;
        RECT 5.930 31.700 9.880 31.850 ;
        RECT 5.930 31.250 6.330 31.700 ;
        RECT 5.930 31.100 9.880 31.250 ;
        RECT 5.930 30.650 6.330 31.100 ;
        RECT 5.930 30.500 9.880 30.650 ;
        RECT 5.930 30.200 6.330 30.500 ;
        RECT 10.480 30.200 10.630 38.400 ;
        RECT 11.080 30.200 11.230 38.400 ;
        RECT 11.680 30.200 11.830 38.400 ;
        RECT 12.280 30.200 12.430 38.400 ;
        RECT 12.880 30.200 13.030 38.400 ;
        RECT 13.480 30.200 13.630 38.400 ;
        RECT 14.080 30.200 14.230 38.400 ;
        RECT 5.930 29.800 14.230 30.200 ;
        RECT 5.930 29.500 6.330 29.800 ;
        RECT 5.930 29.350 9.880 29.500 ;
        RECT 5.930 28.900 6.330 29.350 ;
        RECT 5.930 28.750 9.880 28.900 ;
        RECT 5.930 28.300 6.330 28.750 ;
        RECT 5.930 28.150 9.880 28.300 ;
        RECT 5.930 27.700 6.330 28.150 ;
        RECT 5.930 27.550 9.880 27.700 ;
        RECT 5.930 27.100 6.330 27.550 ;
        RECT 5.930 26.950 9.880 27.100 ;
        RECT 2.315 24.445 4.315 26.740 ;
        RECT 5.930 26.500 6.330 26.950 ;
        RECT 5.930 26.350 9.880 26.500 ;
        RECT 5.930 25.900 6.330 26.350 ;
        RECT 5.930 25.750 9.880 25.900 ;
        RECT 5.930 25.300 6.330 25.750 ;
        RECT 5.930 25.150 9.880 25.300 ;
        RECT 5.930 24.700 6.330 25.150 ;
        RECT 5.930 24.550 9.880 24.700 ;
        RECT 5.930 24.400 6.330 24.550 ;
        RECT 4.730 24.100 6.330 24.400 ;
        RECT 4.730 23.950 9.880 24.100 ;
        RECT 4.730 23.500 6.330 23.950 ;
        RECT 4.730 23.350 9.880 23.500 ;
        RECT 2.315 22.045 4.315 23.320 ;
        RECT 4.730 22.900 6.330 23.350 ;
        RECT 4.730 22.750 9.880 22.900 ;
        RECT 4.730 22.300 6.330 22.750 ;
        RECT 4.730 22.150 9.880 22.300 ;
        RECT 4.730 21.200 5.930 22.150 ;
        RECT 10.480 21.600 10.630 29.800 ;
        RECT 11.080 21.600 11.230 29.800 ;
        RECT 11.680 21.600 11.830 29.800 ;
        RECT 12.280 21.600 12.430 29.800 ;
        RECT 12.880 21.600 13.030 29.800 ;
        RECT 13.480 21.600 13.630 29.800 ;
        RECT 14.080 21.600 14.230 29.800 ;
        RECT 15.230 30.200 15.380 38.400 ;
        RECT 15.830 30.200 15.980 38.400 ;
        RECT 16.430 30.200 16.580 38.400 ;
        RECT 17.030 30.200 17.180 38.400 ;
        RECT 17.630 30.200 17.780 38.400 ;
        RECT 18.230 30.200 18.380 38.400 ;
        RECT 18.830 30.200 18.980 38.400 ;
        RECT 23.530 37.850 25.940 38.800 ;
        RECT 19.580 37.700 29.880 37.850 ;
        RECT 23.130 37.250 26.330 37.700 ;
        RECT 19.580 37.100 29.880 37.250 ;
        RECT 23.130 36.650 26.330 37.100 ;
        RECT 19.580 36.500 29.880 36.650 ;
        RECT 23.130 36.050 26.330 36.500 ;
        RECT 19.580 35.900 29.880 36.050 ;
        RECT 23.130 35.600 26.330 35.900 ;
        RECT 23.130 35.450 23.530 35.600 ;
        RECT 19.580 35.300 23.530 35.450 ;
        RECT 23.130 34.850 23.530 35.300 ;
        RECT 19.580 34.700 23.530 34.850 ;
        RECT 23.130 34.250 23.530 34.700 ;
        RECT 19.580 34.100 23.530 34.250 ;
        RECT 23.130 33.650 23.530 34.100 ;
        RECT 19.580 33.500 23.530 33.650 ;
        RECT 23.130 33.050 23.530 33.500 ;
        RECT 19.580 32.900 23.530 33.050 ;
        RECT 23.130 32.450 23.530 32.900 ;
        RECT 19.580 32.300 23.530 32.450 ;
        RECT 23.130 31.850 23.530 32.300 ;
        RECT 19.580 31.700 23.530 31.850 ;
        RECT 23.130 31.250 23.530 31.700 ;
        RECT 19.580 31.100 23.530 31.250 ;
        RECT 23.130 30.650 23.530 31.100 ;
        RECT 19.580 30.500 23.530 30.650 ;
        RECT 23.130 30.200 23.530 30.500 ;
        RECT 15.230 29.800 23.530 30.200 ;
        RECT 15.230 21.600 15.380 29.800 ;
        RECT 15.830 21.600 15.980 29.800 ;
        RECT 16.430 21.600 16.580 29.800 ;
        RECT 17.030 21.600 17.180 29.800 ;
        RECT 17.630 21.600 17.780 29.800 ;
        RECT 18.230 21.600 18.380 29.800 ;
        RECT 18.830 21.600 18.980 29.800 ;
        RECT 23.130 29.500 23.530 29.800 ;
        RECT 19.580 29.350 23.530 29.500 ;
        RECT 23.130 28.900 23.530 29.350 ;
        RECT 19.580 28.750 23.530 28.900 ;
        RECT 23.130 28.300 23.530 28.750 ;
        RECT 19.580 28.150 23.530 28.300 ;
        RECT 23.130 27.700 23.530 28.150 ;
        RECT 19.580 27.550 23.530 27.700 ;
        RECT 23.130 27.100 23.530 27.550 ;
        RECT 19.580 26.950 23.530 27.100 ;
        RECT 23.130 26.500 23.530 26.950 ;
        RECT 19.580 26.350 23.530 26.500 ;
        RECT 23.130 25.900 23.530 26.350 ;
        RECT 19.580 25.750 23.530 25.900 ;
        RECT 23.130 25.300 23.530 25.750 ;
        RECT 19.580 25.150 23.530 25.300 ;
        RECT 23.130 24.700 23.530 25.150 ;
        RECT 19.580 24.550 23.530 24.700 ;
        RECT 23.130 24.400 23.530 24.550 ;
        RECT 25.930 35.450 26.330 35.600 ;
        RECT 25.930 35.300 29.880 35.450 ;
        RECT 25.930 34.850 26.330 35.300 ;
        RECT 25.930 34.700 29.880 34.850 ;
        RECT 25.930 34.250 26.330 34.700 ;
        RECT 25.930 34.100 29.880 34.250 ;
        RECT 25.930 33.650 26.330 34.100 ;
        RECT 25.930 33.500 29.880 33.650 ;
        RECT 25.930 33.050 26.330 33.500 ;
        RECT 25.930 32.900 29.880 33.050 ;
        RECT 25.930 32.450 26.330 32.900 ;
        RECT 25.930 32.300 29.880 32.450 ;
        RECT 25.930 31.850 26.330 32.300 ;
        RECT 25.930 31.700 29.880 31.850 ;
        RECT 25.930 31.250 26.330 31.700 ;
        RECT 25.930 31.100 29.880 31.250 ;
        RECT 25.930 30.650 26.330 31.100 ;
        RECT 25.930 30.500 29.880 30.650 ;
        RECT 25.930 30.200 26.330 30.500 ;
        RECT 30.480 30.200 30.630 38.400 ;
        RECT 31.080 30.200 31.230 38.400 ;
        RECT 31.680 30.200 31.830 38.400 ;
        RECT 32.280 30.200 32.430 38.400 ;
        RECT 32.880 30.200 33.030 38.400 ;
        RECT 33.480 30.200 33.630 38.400 ;
        RECT 34.080 30.200 34.230 38.400 ;
        RECT 25.930 29.800 34.230 30.200 ;
        RECT 25.930 29.500 26.330 29.800 ;
        RECT 25.930 29.350 29.880 29.500 ;
        RECT 25.930 28.900 26.330 29.350 ;
        RECT 25.930 28.750 29.880 28.900 ;
        RECT 25.930 28.300 26.330 28.750 ;
        RECT 25.930 28.150 29.880 28.300 ;
        RECT 25.930 27.700 26.330 28.150 ;
        RECT 25.930 27.550 29.880 27.700 ;
        RECT 25.930 27.100 26.330 27.550 ;
        RECT 25.930 26.950 29.880 27.100 ;
        RECT 25.930 26.500 26.330 26.950 ;
        RECT 25.930 26.350 29.880 26.500 ;
        RECT 25.930 25.900 26.330 26.350 ;
        RECT 25.930 25.750 29.880 25.900 ;
        RECT 25.930 25.300 26.330 25.750 ;
        RECT 25.930 25.150 29.880 25.300 ;
        RECT 25.930 24.700 26.330 25.150 ;
        RECT 25.930 24.550 29.880 24.700 ;
        RECT 25.930 24.400 26.330 24.550 ;
        RECT 23.130 24.100 26.330 24.400 ;
        RECT 19.580 23.950 29.880 24.100 ;
        RECT 23.130 23.500 26.330 23.950 ;
        RECT 19.580 23.350 29.880 23.500 ;
        RECT 23.130 22.900 26.330 23.350 ;
        RECT 19.580 22.750 29.880 22.900 ;
        RECT 23.130 22.300 26.330 22.750 ;
        RECT 19.580 22.150 29.880 22.300 ;
        RECT 23.530 21.200 25.930 22.150 ;
        RECT 30.480 21.600 30.630 29.800 ;
        RECT 31.080 21.600 31.230 29.800 ;
        RECT 31.680 21.600 31.830 29.800 ;
        RECT 32.280 21.600 32.430 29.800 ;
        RECT 32.880 21.600 33.030 29.800 ;
        RECT 33.480 21.600 33.630 29.800 ;
        RECT 34.080 21.600 34.230 29.800 ;
        RECT 35.230 30.200 35.380 38.400 ;
        RECT 35.830 30.200 35.980 38.400 ;
        RECT 36.430 30.200 36.580 38.400 ;
        RECT 37.030 30.200 37.180 38.400 ;
        RECT 37.630 30.200 37.780 38.400 ;
        RECT 38.230 30.200 38.380 38.400 ;
        RECT 38.830 30.200 38.980 38.400 ;
        RECT 43.530 37.850 45.940 38.800 ;
        RECT 39.580 37.700 49.880 37.850 ;
        RECT 43.130 37.250 46.330 37.700 ;
        RECT 39.580 37.100 49.880 37.250 ;
        RECT 43.130 36.650 46.330 37.100 ;
        RECT 39.580 36.500 49.880 36.650 ;
        RECT 43.130 36.050 46.330 36.500 ;
        RECT 39.580 35.900 49.880 36.050 ;
        RECT 43.130 35.600 46.330 35.900 ;
        RECT 43.130 35.450 43.530 35.600 ;
        RECT 39.580 35.300 43.530 35.450 ;
        RECT 43.130 34.850 43.530 35.300 ;
        RECT 39.580 34.700 43.530 34.850 ;
        RECT 43.130 34.250 43.530 34.700 ;
        RECT 39.580 34.100 43.530 34.250 ;
        RECT 43.130 33.650 43.530 34.100 ;
        RECT 39.580 33.500 43.530 33.650 ;
        RECT 43.130 33.050 43.530 33.500 ;
        RECT 39.580 32.900 43.530 33.050 ;
        RECT 43.130 32.450 43.530 32.900 ;
        RECT 39.580 32.300 43.530 32.450 ;
        RECT 43.130 31.850 43.530 32.300 ;
        RECT 39.580 31.700 43.530 31.850 ;
        RECT 43.130 31.250 43.530 31.700 ;
        RECT 39.580 31.100 43.530 31.250 ;
        RECT 43.130 30.650 43.530 31.100 ;
        RECT 39.580 30.500 43.530 30.650 ;
        RECT 43.130 30.200 43.530 30.500 ;
        RECT 35.230 29.800 43.530 30.200 ;
        RECT 35.230 21.600 35.380 29.800 ;
        RECT 35.830 21.600 35.980 29.800 ;
        RECT 36.430 21.600 36.580 29.800 ;
        RECT 37.030 21.600 37.180 29.800 ;
        RECT 37.630 21.600 37.780 29.800 ;
        RECT 38.230 21.600 38.380 29.800 ;
        RECT 38.830 21.600 38.980 29.800 ;
        RECT 43.130 29.500 43.530 29.800 ;
        RECT 39.580 29.350 43.530 29.500 ;
        RECT 43.130 28.900 43.530 29.350 ;
        RECT 39.580 28.750 43.530 28.900 ;
        RECT 43.130 28.300 43.530 28.750 ;
        RECT 39.580 28.150 43.530 28.300 ;
        RECT 43.130 27.700 43.530 28.150 ;
        RECT 39.580 27.550 43.530 27.700 ;
        RECT 43.130 27.100 43.530 27.550 ;
        RECT 39.580 26.950 43.530 27.100 ;
        RECT 43.130 26.500 43.530 26.950 ;
        RECT 39.580 26.350 43.530 26.500 ;
        RECT 43.130 25.900 43.530 26.350 ;
        RECT 39.580 25.750 43.530 25.900 ;
        RECT 43.130 25.300 43.530 25.750 ;
        RECT 39.580 25.150 43.530 25.300 ;
        RECT 43.130 24.700 43.530 25.150 ;
        RECT 39.580 24.550 43.530 24.700 ;
        RECT 43.130 24.400 43.530 24.550 ;
        RECT 45.930 35.450 46.330 35.600 ;
        RECT 45.930 35.300 49.880 35.450 ;
        RECT 45.930 34.850 46.330 35.300 ;
        RECT 45.930 34.700 49.880 34.850 ;
        RECT 45.930 34.250 46.330 34.700 ;
        RECT 45.930 34.100 49.880 34.250 ;
        RECT 45.930 33.650 46.330 34.100 ;
        RECT 45.930 33.500 49.880 33.650 ;
        RECT 45.930 33.050 46.330 33.500 ;
        RECT 45.930 32.900 49.880 33.050 ;
        RECT 45.930 32.450 46.330 32.900 ;
        RECT 45.930 32.300 49.880 32.450 ;
        RECT 45.930 31.850 46.330 32.300 ;
        RECT 45.930 31.700 49.880 31.850 ;
        RECT 45.930 31.250 46.330 31.700 ;
        RECT 45.930 31.100 49.880 31.250 ;
        RECT 45.930 30.650 46.330 31.100 ;
        RECT 45.930 30.500 49.880 30.650 ;
        RECT 45.930 30.200 46.330 30.500 ;
        RECT 50.480 30.200 50.630 38.400 ;
        RECT 51.080 30.200 51.230 38.400 ;
        RECT 51.680 30.200 51.830 38.400 ;
        RECT 52.280 30.200 52.430 38.400 ;
        RECT 52.880 30.200 53.030 38.400 ;
        RECT 53.480 30.200 53.630 38.400 ;
        RECT 54.080 30.200 54.230 38.400 ;
        RECT 45.930 29.800 54.230 30.200 ;
        RECT 45.930 29.500 46.330 29.800 ;
        RECT 45.930 29.350 49.880 29.500 ;
        RECT 45.930 28.900 46.330 29.350 ;
        RECT 45.930 28.750 49.880 28.900 ;
        RECT 45.930 28.300 46.330 28.750 ;
        RECT 45.930 28.150 49.880 28.300 ;
        RECT 45.930 27.700 46.330 28.150 ;
        RECT 45.930 27.550 49.880 27.700 ;
        RECT 45.930 27.100 46.330 27.550 ;
        RECT 45.930 26.950 49.880 27.100 ;
        RECT 45.930 26.500 46.330 26.950 ;
        RECT 45.930 26.350 49.880 26.500 ;
        RECT 45.930 25.900 46.330 26.350 ;
        RECT 45.930 25.750 49.880 25.900 ;
        RECT 45.930 25.300 46.330 25.750 ;
        RECT 45.930 25.150 49.880 25.300 ;
        RECT 45.930 24.700 46.330 25.150 ;
        RECT 45.930 24.550 49.880 24.700 ;
        RECT 45.930 24.400 46.330 24.550 ;
        RECT 43.130 24.100 46.330 24.400 ;
        RECT 39.580 23.950 49.880 24.100 ;
        RECT 43.130 23.500 46.330 23.950 ;
        RECT 39.580 23.350 49.880 23.500 ;
        RECT 43.130 22.900 46.330 23.350 ;
        RECT 39.580 22.750 49.880 22.900 ;
        RECT 43.130 22.300 46.330 22.750 ;
        RECT 39.580 22.150 49.880 22.300 ;
        RECT 43.530 21.200 45.930 22.150 ;
        RECT 50.480 21.600 50.630 29.800 ;
        RECT 51.080 21.600 51.230 29.800 ;
        RECT 51.680 21.600 51.830 29.800 ;
        RECT 52.280 21.600 52.430 29.800 ;
        RECT 52.880 21.600 53.030 29.800 ;
        RECT 53.480 21.600 53.630 29.800 ;
        RECT 54.080 21.600 54.230 29.800 ;
        RECT 55.230 30.200 55.380 38.400 ;
        RECT 55.830 30.200 55.980 38.400 ;
        RECT 56.430 30.200 56.580 38.400 ;
        RECT 57.030 30.200 57.180 38.400 ;
        RECT 57.630 30.200 57.780 38.400 ;
        RECT 58.230 30.200 58.380 38.400 ;
        RECT 58.830 30.200 58.980 38.400 ;
        RECT 63.530 37.850 65.940 38.800 ;
        RECT 59.580 37.700 69.880 37.850 ;
        RECT 63.130 37.250 66.330 37.700 ;
        RECT 59.580 37.100 69.880 37.250 ;
        RECT 63.130 36.650 66.330 37.100 ;
        RECT 59.580 36.500 69.880 36.650 ;
        RECT 63.130 36.050 66.330 36.500 ;
        RECT 59.580 35.900 69.880 36.050 ;
        RECT 63.130 35.600 66.330 35.900 ;
        RECT 63.130 35.450 63.530 35.600 ;
        RECT 59.580 35.300 63.530 35.450 ;
        RECT 63.130 34.850 63.530 35.300 ;
        RECT 59.580 34.700 63.530 34.850 ;
        RECT 63.130 34.250 63.530 34.700 ;
        RECT 59.580 34.100 63.530 34.250 ;
        RECT 63.130 33.650 63.530 34.100 ;
        RECT 59.580 33.500 63.530 33.650 ;
        RECT 63.130 33.050 63.530 33.500 ;
        RECT 59.580 32.900 63.530 33.050 ;
        RECT 63.130 32.450 63.530 32.900 ;
        RECT 59.580 32.300 63.530 32.450 ;
        RECT 63.130 31.850 63.530 32.300 ;
        RECT 59.580 31.700 63.530 31.850 ;
        RECT 63.130 31.250 63.530 31.700 ;
        RECT 59.580 31.100 63.530 31.250 ;
        RECT 63.130 30.650 63.530 31.100 ;
        RECT 59.580 30.500 63.530 30.650 ;
        RECT 63.130 30.200 63.530 30.500 ;
        RECT 55.230 29.800 63.530 30.200 ;
        RECT 55.230 21.600 55.380 29.800 ;
        RECT 55.830 21.600 55.980 29.800 ;
        RECT 56.430 21.600 56.580 29.800 ;
        RECT 57.030 21.600 57.180 29.800 ;
        RECT 57.630 21.600 57.780 29.800 ;
        RECT 58.230 21.600 58.380 29.800 ;
        RECT 58.830 21.600 58.980 29.800 ;
        RECT 63.130 29.500 63.530 29.800 ;
        RECT 59.580 29.350 63.530 29.500 ;
        RECT 63.130 28.900 63.530 29.350 ;
        RECT 59.580 28.750 63.530 28.900 ;
        RECT 63.130 28.300 63.530 28.750 ;
        RECT 59.580 28.150 63.530 28.300 ;
        RECT 63.130 27.700 63.530 28.150 ;
        RECT 59.580 27.550 63.530 27.700 ;
        RECT 63.130 27.100 63.530 27.550 ;
        RECT 59.580 26.950 63.530 27.100 ;
        RECT 63.130 26.500 63.530 26.950 ;
        RECT 59.580 26.350 63.530 26.500 ;
        RECT 63.130 25.900 63.530 26.350 ;
        RECT 59.580 25.750 63.530 25.900 ;
        RECT 63.130 25.300 63.530 25.750 ;
        RECT 59.580 25.150 63.530 25.300 ;
        RECT 63.130 24.700 63.530 25.150 ;
        RECT 59.580 24.550 63.530 24.700 ;
        RECT 63.130 24.400 63.530 24.550 ;
        RECT 65.930 35.450 66.330 35.600 ;
        RECT 65.930 35.300 69.880 35.450 ;
        RECT 65.930 34.850 66.330 35.300 ;
        RECT 65.930 34.700 69.880 34.850 ;
        RECT 65.930 34.250 66.330 34.700 ;
        RECT 65.930 34.100 69.880 34.250 ;
        RECT 65.930 33.650 66.330 34.100 ;
        RECT 65.930 33.500 69.880 33.650 ;
        RECT 65.930 33.050 66.330 33.500 ;
        RECT 65.930 32.900 69.880 33.050 ;
        RECT 65.930 32.450 66.330 32.900 ;
        RECT 65.930 32.300 69.880 32.450 ;
        RECT 65.930 31.850 66.330 32.300 ;
        RECT 65.930 31.700 69.880 31.850 ;
        RECT 65.930 31.250 66.330 31.700 ;
        RECT 65.930 31.100 69.880 31.250 ;
        RECT 65.930 30.650 66.330 31.100 ;
        RECT 65.930 30.500 69.880 30.650 ;
        RECT 65.930 30.200 66.330 30.500 ;
        RECT 70.480 30.200 70.630 38.400 ;
        RECT 71.080 30.200 71.230 38.400 ;
        RECT 71.680 30.200 71.830 38.400 ;
        RECT 72.280 30.200 72.430 38.400 ;
        RECT 72.880 30.200 73.030 38.400 ;
        RECT 73.480 30.200 73.630 38.400 ;
        RECT 74.080 30.200 74.230 38.400 ;
        RECT 65.930 29.800 74.230 30.200 ;
        RECT 65.930 29.500 66.330 29.800 ;
        RECT 65.930 29.350 69.880 29.500 ;
        RECT 65.930 28.900 66.330 29.350 ;
        RECT 65.930 28.750 69.880 28.900 ;
        RECT 65.930 28.300 66.330 28.750 ;
        RECT 65.930 28.150 69.880 28.300 ;
        RECT 65.930 27.700 66.330 28.150 ;
        RECT 65.930 27.550 69.880 27.700 ;
        RECT 65.930 27.100 66.330 27.550 ;
        RECT 65.930 26.950 69.880 27.100 ;
        RECT 65.930 26.500 66.330 26.950 ;
        RECT 65.930 26.350 69.880 26.500 ;
        RECT 65.930 25.900 66.330 26.350 ;
        RECT 65.930 25.750 69.880 25.900 ;
        RECT 65.930 25.300 66.330 25.750 ;
        RECT 65.930 25.150 69.880 25.300 ;
        RECT 65.930 24.700 66.330 25.150 ;
        RECT 65.930 24.550 69.880 24.700 ;
        RECT 65.930 24.400 66.330 24.550 ;
        RECT 63.130 24.100 66.330 24.400 ;
        RECT 59.580 23.950 69.880 24.100 ;
        RECT 63.130 23.500 66.330 23.950 ;
        RECT 59.580 23.350 69.880 23.500 ;
        RECT 63.130 22.900 66.330 23.350 ;
        RECT 59.580 22.750 69.880 22.900 ;
        RECT 63.130 22.300 66.330 22.750 ;
        RECT 59.580 22.150 69.880 22.300 ;
        RECT 63.530 21.200 65.930 22.150 ;
        RECT 70.480 21.600 70.630 29.800 ;
        RECT 71.080 21.600 71.230 29.800 ;
        RECT 71.680 21.600 71.830 29.800 ;
        RECT 72.280 21.600 72.430 29.800 ;
        RECT 72.880 21.600 73.030 29.800 ;
        RECT 73.480 21.600 73.630 29.800 ;
        RECT 74.080 21.600 74.230 29.800 ;
        RECT 75.230 30.200 75.380 38.400 ;
        RECT 75.830 30.200 75.980 38.400 ;
        RECT 76.430 30.200 76.580 38.400 ;
        RECT 77.030 30.200 77.180 38.400 ;
        RECT 77.630 30.200 77.780 38.400 ;
        RECT 78.230 30.200 78.380 38.400 ;
        RECT 78.830 30.200 78.980 38.400 ;
        RECT 83.530 37.850 85.940 38.800 ;
        RECT 79.580 37.700 89.880 37.850 ;
        RECT 83.130 37.250 86.330 37.700 ;
        RECT 79.580 37.100 89.880 37.250 ;
        RECT 83.130 36.650 86.330 37.100 ;
        RECT 79.580 36.500 89.880 36.650 ;
        RECT 83.130 36.050 86.330 36.500 ;
        RECT 79.580 35.900 89.880 36.050 ;
        RECT 83.130 35.600 86.330 35.900 ;
        RECT 83.130 35.450 83.530 35.600 ;
        RECT 79.580 35.300 83.530 35.450 ;
        RECT 83.130 34.850 83.530 35.300 ;
        RECT 79.580 34.700 83.530 34.850 ;
        RECT 83.130 34.250 83.530 34.700 ;
        RECT 79.580 34.100 83.530 34.250 ;
        RECT 83.130 33.650 83.530 34.100 ;
        RECT 79.580 33.500 83.530 33.650 ;
        RECT 83.130 33.050 83.530 33.500 ;
        RECT 79.580 32.900 83.530 33.050 ;
        RECT 83.130 32.450 83.530 32.900 ;
        RECT 79.580 32.300 83.530 32.450 ;
        RECT 83.130 31.850 83.530 32.300 ;
        RECT 79.580 31.700 83.530 31.850 ;
        RECT 83.130 31.250 83.530 31.700 ;
        RECT 79.580 31.100 83.530 31.250 ;
        RECT 83.130 30.650 83.530 31.100 ;
        RECT 79.580 30.500 83.530 30.650 ;
        RECT 83.130 30.200 83.530 30.500 ;
        RECT 75.230 29.800 83.530 30.200 ;
        RECT 75.230 21.600 75.380 29.800 ;
        RECT 75.830 21.600 75.980 29.800 ;
        RECT 76.430 21.600 76.580 29.800 ;
        RECT 77.030 21.600 77.180 29.800 ;
        RECT 77.630 21.600 77.780 29.800 ;
        RECT 78.230 21.600 78.380 29.800 ;
        RECT 78.830 21.600 78.980 29.800 ;
        RECT 83.130 29.500 83.530 29.800 ;
        RECT 79.580 29.350 83.530 29.500 ;
        RECT 83.130 28.900 83.530 29.350 ;
        RECT 79.580 28.750 83.530 28.900 ;
        RECT 83.130 28.300 83.530 28.750 ;
        RECT 79.580 28.150 83.530 28.300 ;
        RECT 83.130 27.700 83.530 28.150 ;
        RECT 79.580 27.550 83.530 27.700 ;
        RECT 83.130 27.100 83.530 27.550 ;
        RECT 79.580 26.950 83.530 27.100 ;
        RECT 83.130 26.500 83.530 26.950 ;
        RECT 79.580 26.350 83.530 26.500 ;
        RECT 83.130 25.900 83.530 26.350 ;
        RECT 79.580 25.750 83.530 25.900 ;
        RECT 83.130 25.300 83.530 25.750 ;
        RECT 79.580 25.150 83.530 25.300 ;
        RECT 83.130 24.700 83.530 25.150 ;
        RECT 79.580 24.550 83.530 24.700 ;
        RECT 83.130 24.400 83.530 24.550 ;
        RECT 85.930 35.450 86.330 35.600 ;
        RECT 85.930 35.300 89.880 35.450 ;
        RECT 85.930 34.850 86.330 35.300 ;
        RECT 85.930 34.700 89.880 34.850 ;
        RECT 85.930 34.250 86.330 34.700 ;
        RECT 85.930 34.100 89.880 34.250 ;
        RECT 85.930 33.650 86.330 34.100 ;
        RECT 85.930 33.500 89.880 33.650 ;
        RECT 85.930 33.050 86.330 33.500 ;
        RECT 85.930 32.900 89.880 33.050 ;
        RECT 85.930 32.450 86.330 32.900 ;
        RECT 85.930 32.300 89.880 32.450 ;
        RECT 85.930 31.850 86.330 32.300 ;
        RECT 85.930 31.700 89.880 31.850 ;
        RECT 85.930 31.250 86.330 31.700 ;
        RECT 85.930 31.100 89.880 31.250 ;
        RECT 85.930 30.650 86.330 31.100 ;
        RECT 85.930 30.500 89.880 30.650 ;
        RECT 85.930 30.200 86.330 30.500 ;
        RECT 90.480 30.200 90.630 38.400 ;
        RECT 91.080 30.200 91.230 38.400 ;
        RECT 91.680 30.200 91.830 38.400 ;
        RECT 92.280 30.200 92.430 38.400 ;
        RECT 92.880 30.200 93.030 38.400 ;
        RECT 93.480 30.200 93.630 38.400 ;
        RECT 94.080 30.200 94.230 38.400 ;
        RECT 85.930 29.800 94.230 30.200 ;
        RECT 85.930 29.500 86.330 29.800 ;
        RECT 85.930 29.350 89.880 29.500 ;
        RECT 85.930 28.900 86.330 29.350 ;
        RECT 85.930 28.750 89.880 28.900 ;
        RECT 85.930 28.300 86.330 28.750 ;
        RECT 85.930 28.150 89.880 28.300 ;
        RECT 85.930 27.700 86.330 28.150 ;
        RECT 85.930 27.550 89.880 27.700 ;
        RECT 85.930 27.100 86.330 27.550 ;
        RECT 85.930 26.950 89.880 27.100 ;
        RECT 85.930 26.500 86.330 26.950 ;
        RECT 85.930 26.350 89.880 26.500 ;
        RECT 85.930 25.900 86.330 26.350 ;
        RECT 85.930 25.750 89.880 25.900 ;
        RECT 85.930 25.300 86.330 25.750 ;
        RECT 85.930 25.150 89.880 25.300 ;
        RECT 85.930 24.700 86.330 25.150 ;
        RECT 85.930 24.550 89.880 24.700 ;
        RECT 85.930 24.400 86.330 24.550 ;
        RECT 83.130 24.100 86.330 24.400 ;
        RECT 79.580 23.950 89.880 24.100 ;
        RECT 83.130 23.500 86.330 23.950 ;
        RECT 79.580 23.350 89.880 23.500 ;
        RECT 83.130 22.900 86.330 23.350 ;
        RECT 79.580 22.750 89.880 22.900 ;
        RECT 83.130 22.300 86.330 22.750 ;
        RECT 79.580 22.150 89.880 22.300 ;
        RECT 83.530 21.200 85.930 22.150 ;
        RECT 90.480 21.600 90.630 29.800 ;
        RECT 91.080 21.600 91.230 29.800 ;
        RECT 91.680 21.600 91.830 29.800 ;
        RECT 92.280 21.600 92.430 29.800 ;
        RECT 92.880 21.600 93.030 29.800 ;
        RECT 93.480 21.600 93.630 29.800 ;
        RECT 94.080 21.600 94.230 29.800 ;
        RECT 95.230 30.200 95.380 38.400 ;
        RECT 95.830 30.200 95.980 38.400 ;
        RECT 96.430 30.200 96.580 38.400 ;
        RECT 97.030 30.200 97.180 38.400 ;
        RECT 97.630 30.200 97.780 38.400 ;
        RECT 98.230 30.200 98.380 38.400 ;
        RECT 98.830 30.200 98.980 38.400 ;
        RECT 103.530 37.850 105.940 38.800 ;
        RECT 99.580 37.700 109.880 37.850 ;
        RECT 103.130 37.250 106.330 37.700 ;
        RECT 99.580 37.100 109.880 37.250 ;
        RECT 103.130 36.650 106.330 37.100 ;
        RECT 99.580 36.500 109.880 36.650 ;
        RECT 103.130 36.050 106.330 36.500 ;
        RECT 99.580 35.900 109.880 36.050 ;
        RECT 103.130 35.600 106.330 35.900 ;
        RECT 103.130 35.450 103.530 35.600 ;
        RECT 99.580 35.300 103.530 35.450 ;
        RECT 103.130 34.850 103.530 35.300 ;
        RECT 99.580 34.700 103.530 34.850 ;
        RECT 103.130 34.250 103.530 34.700 ;
        RECT 99.580 34.100 103.530 34.250 ;
        RECT 103.130 33.650 103.530 34.100 ;
        RECT 99.580 33.500 103.530 33.650 ;
        RECT 103.130 33.050 103.530 33.500 ;
        RECT 99.580 32.900 103.530 33.050 ;
        RECT 103.130 32.450 103.530 32.900 ;
        RECT 99.580 32.300 103.530 32.450 ;
        RECT 103.130 31.850 103.530 32.300 ;
        RECT 99.580 31.700 103.530 31.850 ;
        RECT 103.130 31.250 103.530 31.700 ;
        RECT 99.580 31.100 103.530 31.250 ;
        RECT 103.130 30.650 103.530 31.100 ;
        RECT 99.580 30.500 103.530 30.650 ;
        RECT 103.130 30.200 103.530 30.500 ;
        RECT 95.230 29.800 103.530 30.200 ;
        RECT 95.230 21.600 95.380 29.800 ;
        RECT 95.830 21.600 95.980 29.800 ;
        RECT 96.430 21.600 96.580 29.800 ;
        RECT 97.030 21.600 97.180 29.800 ;
        RECT 97.630 21.600 97.780 29.800 ;
        RECT 98.230 21.600 98.380 29.800 ;
        RECT 98.830 21.600 98.980 29.800 ;
        RECT 103.130 29.500 103.530 29.800 ;
        RECT 99.580 29.350 103.530 29.500 ;
        RECT 103.130 28.900 103.530 29.350 ;
        RECT 99.580 28.750 103.530 28.900 ;
        RECT 103.130 28.300 103.530 28.750 ;
        RECT 99.580 28.150 103.530 28.300 ;
        RECT 103.130 27.700 103.530 28.150 ;
        RECT 99.580 27.550 103.530 27.700 ;
        RECT 103.130 27.100 103.530 27.550 ;
        RECT 99.580 26.950 103.530 27.100 ;
        RECT 103.130 26.500 103.530 26.950 ;
        RECT 99.580 26.350 103.530 26.500 ;
        RECT 103.130 25.900 103.530 26.350 ;
        RECT 99.580 25.750 103.530 25.900 ;
        RECT 103.130 25.300 103.530 25.750 ;
        RECT 99.580 25.150 103.530 25.300 ;
        RECT 103.130 24.700 103.530 25.150 ;
        RECT 99.580 24.550 103.530 24.700 ;
        RECT 103.130 24.400 103.530 24.550 ;
        RECT 105.930 35.450 106.330 35.600 ;
        RECT 105.930 35.300 109.880 35.450 ;
        RECT 105.930 34.850 106.330 35.300 ;
        RECT 105.930 34.700 109.880 34.850 ;
        RECT 105.930 34.250 106.330 34.700 ;
        RECT 105.930 34.100 109.880 34.250 ;
        RECT 105.930 33.650 106.330 34.100 ;
        RECT 105.930 33.500 109.880 33.650 ;
        RECT 105.930 33.050 106.330 33.500 ;
        RECT 105.930 32.900 109.880 33.050 ;
        RECT 105.930 32.450 106.330 32.900 ;
        RECT 105.930 32.300 109.880 32.450 ;
        RECT 105.930 31.850 106.330 32.300 ;
        RECT 105.930 31.700 109.880 31.850 ;
        RECT 105.930 31.250 106.330 31.700 ;
        RECT 105.930 31.100 109.880 31.250 ;
        RECT 105.930 30.650 106.330 31.100 ;
        RECT 105.930 30.500 109.880 30.650 ;
        RECT 105.930 30.200 106.330 30.500 ;
        RECT 110.480 30.200 110.630 38.400 ;
        RECT 111.080 30.200 111.230 38.400 ;
        RECT 111.680 30.200 111.830 38.400 ;
        RECT 112.280 30.200 112.430 38.400 ;
        RECT 112.880 30.200 113.030 38.400 ;
        RECT 113.480 30.200 113.630 38.400 ;
        RECT 114.080 30.200 114.230 38.400 ;
        RECT 105.930 29.800 114.230 30.200 ;
        RECT 105.930 29.500 106.330 29.800 ;
        RECT 105.930 29.350 109.880 29.500 ;
        RECT 105.930 28.900 106.330 29.350 ;
        RECT 105.930 28.750 109.880 28.900 ;
        RECT 105.930 28.300 106.330 28.750 ;
        RECT 105.930 28.150 109.880 28.300 ;
        RECT 105.930 27.700 106.330 28.150 ;
        RECT 105.930 27.550 109.880 27.700 ;
        RECT 105.930 27.100 106.330 27.550 ;
        RECT 105.930 26.950 109.880 27.100 ;
        RECT 105.930 26.500 106.330 26.950 ;
        RECT 105.930 26.350 109.880 26.500 ;
        RECT 105.930 25.900 106.330 26.350 ;
        RECT 105.930 25.750 109.880 25.900 ;
        RECT 105.930 25.300 106.330 25.750 ;
        RECT 105.930 25.150 109.880 25.300 ;
        RECT 105.930 24.700 106.330 25.150 ;
        RECT 105.930 24.550 109.880 24.700 ;
        RECT 105.930 24.400 106.330 24.550 ;
        RECT 103.130 24.100 106.330 24.400 ;
        RECT 99.580 23.950 109.880 24.100 ;
        RECT 103.130 23.500 106.330 23.950 ;
        RECT 99.580 23.350 109.880 23.500 ;
        RECT 103.130 22.900 106.330 23.350 ;
        RECT 99.580 22.750 109.880 22.900 ;
        RECT 103.130 22.300 106.330 22.750 ;
        RECT 99.580 22.150 109.880 22.300 ;
        RECT 103.530 21.200 105.930 22.150 ;
        RECT 110.480 21.600 110.630 29.800 ;
        RECT 111.080 21.600 111.230 29.800 ;
        RECT 111.680 21.600 111.830 29.800 ;
        RECT 112.280 21.600 112.430 29.800 ;
        RECT 112.880 21.600 113.030 29.800 ;
        RECT 113.480 21.600 113.630 29.800 ;
        RECT 114.080 21.600 114.230 29.800 ;
        RECT 115.230 30.200 115.380 38.400 ;
        RECT 115.830 30.200 115.980 38.400 ;
        RECT 116.430 30.200 116.580 38.400 ;
        RECT 117.030 30.200 117.180 38.400 ;
        RECT 117.630 30.200 117.780 38.400 ;
        RECT 118.230 30.200 118.380 38.400 ;
        RECT 118.830 30.200 118.980 38.400 ;
        RECT 123.530 37.850 124.730 38.800 ;
        RECT 119.580 37.700 124.730 37.850 ;
        RECT 123.130 37.250 124.730 37.700 ;
        RECT 119.580 37.100 124.730 37.250 ;
        RECT 123.130 36.650 124.730 37.100 ;
        RECT 119.580 36.500 124.730 36.650 ;
        RECT 123.130 36.050 124.730 36.500 ;
        RECT 119.580 35.900 124.730 36.050 ;
        RECT 125.135 36.035 127.135 37.310 ;
        RECT 123.130 35.600 124.730 35.900 ;
        RECT 123.130 35.450 123.530 35.600 ;
        RECT 119.580 35.300 123.530 35.450 ;
        RECT 123.130 34.850 123.530 35.300 ;
        RECT 119.580 34.700 123.530 34.850 ;
        RECT 123.130 34.250 123.530 34.700 ;
        RECT 119.580 34.100 123.530 34.250 ;
        RECT 123.130 33.650 123.530 34.100 ;
        RECT 119.580 33.500 123.530 33.650 ;
        RECT 123.130 33.050 123.530 33.500 ;
        RECT 119.580 32.900 123.530 33.050 ;
        RECT 123.130 32.450 123.530 32.900 ;
        RECT 119.580 32.300 123.530 32.450 ;
        RECT 123.130 31.850 123.530 32.300 ;
        RECT 119.580 31.700 123.530 31.850 ;
        RECT 123.130 31.250 123.530 31.700 ;
        RECT 119.580 31.100 123.530 31.250 ;
        RECT 123.130 30.650 123.530 31.100 ;
        RECT 119.580 30.500 123.530 30.650 ;
        RECT 123.130 30.200 123.530 30.500 ;
        RECT 115.230 29.800 123.530 30.200 ;
        RECT 115.230 21.600 115.380 29.800 ;
        RECT 115.830 21.600 115.980 29.800 ;
        RECT 116.430 21.600 116.580 29.800 ;
        RECT 117.030 21.600 117.180 29.800 ;
        RECT 117.630 21.600 117.780 29.800 ;
        RECT 118.230 21.600 118.380 29.800 ;
        RECT 118.830 21.600 118.980 29.800 ;
        RECT 123.130 29.500 123.530 29.800 ;
        RECT 119.580 29.350 123.530 29.500 ;
        RECT 123.130 28.900 123.530 29.350 ;
        RECT 119.580 28.750 123.530 28.900 ;
        RECT 123.130 28.300 123.530 28.750 ;
        RECT 119.580 28.150 123.530 28.300 ;
        RECT 123.130 27.700 123.530 28.150 ;
        RECT 119.580 27.550 123.530 27.700 ;
        RECT 123.130 27.100 123.530 27.550 ;
        RECT 119.580 26.950 123.530 27.100 ;
        RECT 123.130 26.500 123.530 26.950 ;
        RECT 119.580 26.350 123.530 26.500 ;
        RECT 123.130 25.900 123.530 26.350 ;
        RECT 119.580 25.750 123.530 25.900 ;
        RECT 123.130 25.300 123.530 25.750 ;
        RECT 119.580 25.150 123.530 25.300 ;
        RECT 123.130 24.700 123.530 25.150 ;
        RECT 119.580 24.550 123.530 24.700 ;
        RECT 123.130 24.400 123.530 24.550 ;
        RECT 123.130 24.100 124.730 24.400 ;
        RECT 119.580 23.950 124.730 24.100 ;
        RECT 123.130 23.500 124.730 23.950 ;
        RECT 119.580 23.350 124.730 23.500 ;
        RECT 123.130 22.900 124.730 23.350 ;
        RECT 119.580 22.750 124.730 22.900 ;
        RECT 123.130 22.300 124.730 22.750 ;
        RECT 119.580 22.150 124.730 22.300 ;
        RECT 123.530 21.200 124.730 22.150 ;
        RECT 125.140 21.820 127.140 23.095 ;
        RECT 4.730 18.800 9.130 21.200 ;
        RECT 20.330 18.800 29.130 21.200 ;
        RECT 40.330 18.800 49.130 21.200 ;
        RECT 60.330 18.800 69.130 21.200 ;
        RECT 80.330 18.800 89.130 21.200 ;
        RECT 100.330 18.800 109.130 21.200 ;
        RECT 120.330 18.800 124.730 21.200 ;
        RECT 4.730 17.850 5.940 18.800 ;
        RECT 2.315 16.490 4.315 17.765 ;
        RECT 4.730 17.700 9.880 17.850 ;
        RECT 4.730 17.250 6.330 17.700 ;
        RECT 4.730 17.100 9.880 17.250 ;
        RECT 4.730 16.650 6.330 17.100 ;
        RECT 4.730 16.500 9.880 16.650 ;
        RECT 4.730 16.050 6.330 16.500 ;
        RECT 4.730 15.900 9.880 16.050 ;
        RECT 4.730 15.600 6.330 15.900 ;
        RECT 2.315 13.255 4.315 15.550 ;
        RECT 5.930 15.450 6.330 15.600 ;
        RECT 5.930 15.300 9.880 15.450 ;
        RECT 5.930 14.850 6.330 15.300 ;
        RECT 5.930 14.700 9.880 14.850 ;
        RECT 5.930 14.250 6.330 14.700 ;
        RECT 5.930 14.100 9.880 14.250 ;
        RECT 5.930 13.650 6.330 14.100 ;
        RECT 5.930 13.500 9.880 13.650 ;
        RECT 5.930 13.050 6.330 13.500 ;
        RECT 5.930 12.900 9.880 13.050 ;
        RECT 5.930 12.450 6.330 12.900 ;
        RECT 5.930 12.300 9.880 12.450 ;
        RECT 5.930 11.850 6.330 12.300 ;
        RECT 5.930 11.700 9.880 11.850 ;
        RECT 5.930 11.250 6.330 11.700 ;
        RECT 5.930 11.100 9.880 11.250 ;
        RECT 5.930 10.650 6.330 11.100 ;
        RECT 5.930 10.500 9.880 10.650 ;
        RECT 5.930 10.200 6.330 10.500 ;
        RECT 10.480 10.200 10.630 18.400 ;
        RECT 11.080 10.200 11.230 18.400 ;
        RECT 11.680 10.200 11.830 18.400 ;
        RECT 12.280 10.200 12.430 18.400 ;
        RECT 12.880 10.200 13.030 18.400 ;
        RECT 13.480 10.200 13.630 18.400 ;
        RECT 14.080 10.200 14.230 18.400 ;
        RECT 5.930 9.800 14.230 10.200 ;
        RECT 5.930 9.500 6.330 9.800 ;
        RECT 5.930 9.350 9.880 9.500 ;
        RECT 5.930 8.900 6.330 9.350 ;
        RECT 5.930 8.750 9.880 8.900 ;
        RECT 5.930 8.300 6.330 8.750 ;
        RECT 5.930 8.150 9.880 8.300 ;
        RECT 5.930 7.700 6.330 8.150 ;
        RECT 5.930 7.550 9.880 7.700 ;
        RECT 5.930 7.100 6.330 7.550 ;
        RECT 5.930 6.950 9.880 7.100 ;
        RECT 2.315 4.450 4.315 6.745 ;
        RECT 5.930 6.500 6.330 6.950 ;
        RECT 5.930 6.350 9.880 6.500 ;
        RECT 5.930 5.900 6.330 6.350 ;
        RECT 5.930 5.750 9.880 5.900 ;
        RECT 5.930 5.300 6.330 5.750 ;
        RECT 5.930 5.150 9.880 5.300 ;
        RECT 5.930 4.700 6.330 5.150 ;
        RECT 5.930 4.550 9.880 4.700 ;
        RECT 5.930 4.400 6.330 4.550 ;
        RECT 4.730 4.100 6.330 4.400 ;
        RECT 4.730 3.950 9.880 4.100 ;
        RECT 2.315 2.375 4.325 3.650 ;
        RECT 4.730 3.500 6.330 3.950 ;
        RECT 4.730 3.350 9.880 3.500 ;
        RECT 4.730 2.900 6.330 3.350 ;
        RECT 4.730 2.750 9.880 2.900 ;
        RECT 4.730 2.300 6.330 2.750 ;
        RECT 4.730 2.150 9.880 2.300 ;
        RECT 4.730 1.200 5.930 2.150 ;
        RECT 10.480 1.600 10.630 9.800 ;
        RECT 11.080 1.600 11.230 9.800 ;
        RECT 11.680 1.600 11.830 9.800 ;
        RECT 12.280 1.600 12.430 9.800 ;
        RECT 12.880 1.600 13.030 9.800 ;
        RECT 13.480 1.600 13.630 9.800 ;
        RECT 14.080 1.600 14.230 9.800 ;
        RECT 15.230 10.200 15.380 18.400 ;
        RECT 15.830 10.200 15.980 18.400 ;
        RECT 16.430 10.200 16.580 18.400 ;
        RECT 17.030 10.200 17.180 18.400 ;
        RECT 17.630 10.200 17.780 18.400 ;
        RECT 18.230 10.200 18.380 18.400 ;
        RECT 18.830 10.200 18.980 18.400 ;
        RECT 23.530 17.850 25.940 18.800 ;
        RECT 19.580 17.700 29.880 17.850 ;
        RECT 23.130 17.250 26.330 17.700 ;
        RECT 19.580 17.100 29.880 17.250 ;
        RECT 23.130 16.650 26.330 17.100 ;
        RECT 19.580 16.500 29.880 16.650 ;
        RECT 23.130 16.050 26.330 16.500 ;
        RECT 19.580 15.900 29.880 16.050 ;
        RECT 23.130 15.600 26.330 15.900 ;
        RECT 23.130 15.450 23.530 15.600 ;
        RECT 19.580 15.300 23.530 15.450 ;
        RECT 23.130 14.850 23.530 15.300 ;
        RECT 19.580 14.700 23.530 14.850 ;
        RECT 23.130 14.250 23.530 14.700 ;
        RECT 19.580 14.100 23.530 14.250 ;
        RECT 23.130 13.650 23.530 14.100 ;
        RECT 19.580 13.500 23.530 13.650 ;
        RECT 23.130 13.050 23.530 13.500 ;
        RECT 19.580 12.900 23.530 13.050 ;
        RECT 23.130 12.450 23.530 12.900 ;
        RECT 19.580 12.300 23.530 12.450 ;
        RECT 23.130 11.850 23.530 12.300 ;
        RECT 19.580 11.700 23.530 11.850 ;
        RECT 23.130 11.250 23.530 11.700 ;
        RECT 19.580 11.100 23.530 11.250 ;
        RECT 23.130 10.650 23.530 11.100 ;
        RECT 19.580 10.500 23.530 10.650 ;
        RECT 23.130 10.200 23.530 10.500 ;
        RECT 15.230 9.800 23.530 10.200 ;
        RECT 15.230 1.600 15.380 9.800 ;
        RECT 15.830 1.600 15.980 9.800 ;
        RECT 16.430 1.600 16.580 9.800 ;
        RECT 17.030 1.600 17.180 9.800 ;
        RECT 17.630 1.600 17.780 9.800 ;
        RECT 18.230 1.600 18.380 9.800 ;
        RECT 18.830 1.600 18.980 9.800 ;
        RECT 23.130 9.500 23.530 9.800 ;
        RECT 19.580 9.350 23.530 9.500 ;
        RECT 23.130 8.900 23.530 9.350 ;
        RECT 19.580 8.750 23.530 8.900 ;
        RECT 23.130 8.300 23.530 8.750 ;
        RECT 19.580 8.150 23.530 8.300 ;
        RECT 23.130 7.700 23.530 8.150 ;
        RECT 19.580 7.550 23.530 7.700 ;
        RECT 23.130 7.100 23.530 7.550 ;
        RECT 19.580 6.950 23.530 7.100 ;
        RECT 23.130 6.500 23.530 6.950 ;
        RECT 19.580 6.350 23.530 6.500 ;
        RECT 23.130 5.900 23.530 6.350 ;
        RECT 19.580 5.750 23.530 5.900 ;
        RECT 23.130 5.300 23.530 5.750 ;
        RECT 19.580 5.150 23.530 5.300 ;
        RECT 23.130 4.700 23.530 5.150 ;
        RECT 19.580 4.550 23.530 4.700 ;
        RECT 23.130 4.400 23.530 4.550 ;
        RECT 25.930 15.450 26.330 15.600 ;
        RECT 25.930 15.300 29.880 15.450 ;
        RECT 25.930 14.850 26.330 15.300 ;
        RECT 25.930 14.700 29.880 14.850 ;
        RECT 25.930 14.250 26.330 14.700 ;
        RECT 25.930 14.100 29.880 14.250 ;
        RECT 25.930 13.650 26.330 14.100 ;
        RECT 25.930 13.500 29.880 13.650 ;
        RECT 25.930 13.050 26.330 13.500 ;
        RECT 25.930 12.900 29.880 13.050 ;
        RECT 25.930 12.450 26.330 12.900 ;
        RECT 25.930 12.300 29.880 12.450 ;
        RECT 25.930 11.850 26.330 12.300 ;
        RECT 25.930 11.700 29.880 11.850 ;
        RECT 25.930 11.250 26.330 11.700 ;
        RECT 25.930 11.100 29.880 11.250 ;
        RECT 25.930 10.650 26.330 11.100 ;
        RECT 25.930 10.500 29.880 10.650 ;
        RECT 25.930 10.200 26.330 10.500 ;
        RECT 30.480 10.200 30.630 18.400 ;
        RECT 31.080 10.200 31.230 18.400 ;
        RECT 31.680 10.200 31.830 18.400 ;
        RECT 32.280 10.200 32.430 18.400 ;
        RECT 32.880 10.200 33.030 18.400 ;
        RECT 33.480 10.200 33.630 18.400 ;
        RECT 34.080 10.200 34.230 18.400 ;
        RECT 25.930 9.800 34.230 10.200 ;
        RECT 25.930 9.500 26.330 9.800 ;
        RECT 25.930 9.350 29.880 9.500 ;
        RECT 25.930 8.900 26.330 9.350 ;
        RECT 25.930 8.750 29.880 8.900 ;
        RECT 25.930 8.300 26.330 8.750 ;
        RECT 25.930 8.150 29.880 8.300 ;
        RECT 25.930 7.700 26.330 8.150 ;
        RECT 25.930 7.550 29.880 7.700 ;
        RECT 25.930 7.100 26.330 7.550 ;
        RECT 25.930 6.950 29.880 7.100 ;
        RECT 25.930 6.500 26.330 6.950 ;
        RECT 25.930 6.350 29.880 6.500 ;
        RECT 25.930 5.900 26.330 6.350 ;
        RECT 25.930 5.750 29.880 5.900 ;
        RECT 25.930 5.300 26.330 5.750 ;
        RECT 25.930 5.150 29.880 5.300 ;
        RECT 25.930 4.700 26.330 5.150 ;
        RECT 25.930 4.550 29.880 4.700 ;
        RECT 25.930 4.400 26.330 4.550 ;
        RECT 23.130 4.100 26.330 4.400 ;
        RECT 19.580 3.950 29.880 4.100 ;
        RECT 23.130 3.500 26.330 3.950 ;
        RECT 19.580 3.350 29.880 3.500 ;
        RECT 23.130 2.900 26.330 3.350 ;
        RECT 19.580 2.750 29.880 2.900 ;
        RECT 23.130 2.300 26.330 2.750 ;
        RECT 19.580 2.150 29.880 2.300 ;
        RECT 23.530 1.200 25.930 2.150 ;
        RECT 30.480 1.600 30.630 9.800 ;
        RECT 31.080 1.600 31.230 9.800 ;
        RECT 31.680 1.600 31.830 9.800 ;
        RECT 32.280 1.600 32.430 9.800 ;
        RECT 32.880 1.600 33.030 9.800 ;
        RECT 33.480 1.600 33.630 9.800 ;
        RECT 34.080 1.600 34.230 9.800 ;
        RECT 35.230 10.200 35.380 18.400 ;
        RECT 35.830 10.200 35.980 18.400 ;
        RECT 36.430 10.200 36.580 18.400 ;
        RECT 37.030 10.200 37.180 18.400 ;
        RECT 37.630 10.200 37.780 18.400 ;
        RECT 38.230 10.200 38.380 18.400 ;
        RECT 38.830 10.200 38.980 18.400 ;
        RECT 43.530 17.850 45.940 18.800 ;
        RECT 39.580 17.700 49.880 17.850 ;
        RECT 43.130 17.250 46.330 17.700 ;
        RECT 39.580 17.100 49.880 17.250 ;
        RECT 43.130 16.650 46.330 17.100 ;
        RECT 39.580 16.500 49.880 16.650 ;
        RECT 43.130 16.050 46.330 16.500 ;
        RECT 39.580 15.900 49.880 16.050 ;
        RECT 43.130 15.600 46.330 15.900 ;
        RECT 43.130 15.450 43.530 15.600 ;
        RECT 39.580 15.300 43.530 15.450 ;
        RECT 43.130 14.850 43.530 15.300 ;
        RECT 39.580 14.700 43.530 14.850 ;
        RECT 43.130 14.250 43.530 14.700 ;
        RECT 39.580 14.100 43.530 14.250 ;
        RECT 43.130 13.650 43.530 14.100 ;
        RECT 39.580 13.500 43.530 13.650 ;
        RECT 43.130 13.050 43.530 13.500 ;
        RECT 39.580 12.900 43.530 13.050 ;
        RECT 43.130 12.450 43.530 12.900 ;
        RECT 39.580 12.300 43.530 12.450 ;
        RECT 43.130 11.850 43.530 12.300 ;
        RECT 39.580 11.700 43.530 11.850 ;
        RECT 43.130 11.250 43.530 11.700 ;
        RECT 39.580 11.100 43.530 11.250 ;
        RECT 43.130 10.650 43.530 11.100 ;
        RECT 39.580 10.500 43.530 10.650 ;
        RECT 43.130 10.200 43.530 10.500 ;
        RECT 35.230 9.800 43.530 10.200 ;
        RECT 35.230 1.600 35.380 9.800 ;
        RECT 35.830 1.600 35.980 9.800 ;
        RECT 36.430 1.600 36.580 9.800 ;
        RECT 37.030 1.600 37.180 9.800 ;
        RECT 37.630 1.600 37.780 9.800 ;
        RECT 38.230 1.600 38.380 9.800 ;
        RECT 38.830 1.600 38.980 9.800 ;
        RECT 43.130 9.500 43.530 9.800 ;
        RECT 39.580 9.350 43.530 9.500 ;
        RECT 43.130 8.900 43.530 9.350 ;
        RECT 39.580 8.750 43.530 8.900 ;
        RECT 43.130 8.300 43.530 8.750 ;
        RECT 39.580 8.150 43.530 8.300 ;
        RECT 43.130 7.700 43.530 8.150 ;
        RECT 39.580 7.550 43.530 7.700 ;
        RECT 43.130 7.100 43.530 7.550 ;
        RECT 39.580 6.950 43.530 7.100 ;
        RECT 43.130 6.500 43.530 6.950 ;
        RECT 39.580 6.350 43.530 6.500 ;
        RECT 43.130 5.900 43.530 6.350 ;
        RECT 39.580 5.750 43.530 5.900 ;
        RECT 43.130 5.300 43.530 5.750 ;
        RECT 39.580 5.150 43.530 5.300 ;
        RECT 43.130 4.700 43.530 5.150 ;
        RECT 39.580 4.550 43.530 4.700 ;
        RECT 43.130 4.400 43.530 4.550 ;
        RECT 45.930 15.450 46.330 15.600 ;
        RECT 45.930 15.300 49.880 15.450 ;
        RECT 45.930 14.850 46.330 15.300 ;
        RECT 45.930 14.700 49.880 14.850 ;
        RECT 45.930 14.250 46.330 14.700 ;
        RECT 45.930 14.100 49.880 14.250 ;
        RECT 45.930 13.650 46.330 14.100 ;
        RECT 45.930 13.500 49.880 13.650 ;
        RECT 45.930 13.050 46.330 13.500 ;
        RECT 45.930 12.900 49.880 13.050 ;
        RECT 45.930 12.450 46.330 12.900 ;
        RECT 45.930 12.300 49.880 12.450 ;
        RECT 45.930 11.850 46.330 12.300 ;
        RECT 45.930 11.700 49.880 11.850 ;
        RECT 45.930 11.250 46.330 11.700 ;
        RECT 45.930 11.100 49.880 11.250 ;
        RECT 45.930 10.650 46.330 11.100 ;
        RECT 45.930 10.500 49.880 10.650 ;
        RECT 45.930 10.200 46.330 10.500 ;
        RECT 50.480 10.200 50.630 18.400 ;
        RECT 51.080 10.200 51.230 18.400 ;
        RECT 51.680 10.200 51.830 18.400 ;
        RECT 52.280 10.200 52.430 18.400 ;
        RECT 52.880 10.200 53.030 18.400 ;
        RECT 53.480 10.200 53.630 18.400 ;
        RECT 54.080 10.200 54.230 18.400 ;
        RECT 45.930 9.800 54.230 10.200 ;
        RECT 45.930 9.500 46.330 9.800 ;
        RECT 45.930 9.350 49.880 9.500 ;
        RECT 45.930 8.900 46.330 9.350 ;
        RECT 45.930 8.750 49.880 8.900 ;
        RECT 45.930 8.300 46.330 8.750 ;
        RECT 45.930 8.150 49.880 8.300 ;
        RECT 45.930 7.700 46.330 8.150 ;
        RECT 45.930 7.550 49.880 7.700 ;
        RECT 45.930 7.100 46.330 7.550 ;
        RECT 45.930 6.950 49.880 7.100 ;
        RECT 45.930 6.500 46.330 6.950 ;
        RECT 45.930 6.350 49.880 6.500 ;
        RECT 45.930 5.900 46.330 6.350 ;
        RECT 45.930 5.750 49.880 5.900 ;
        RECT 45.930 5.300 46.330 5.750 ;
        RECT 45.930 5.150 49.880 5.300 ;
        RECT 45.930 4.700 46.330 5.150 ;
        RECT 45.930 4.550 49.880 4.700 ;
        RECT 45.930 4.400 46.330 4.550 ;
        RECT 43.130 4.100 46.330 4.400 ;
        RECT 39.580 3.950 49.880 4.100 ;
        RECT 43.130 3.500 46.330 3.950 ;
        RECT 39.580 3.350 49.880 3.500 ;
        RECT 43.130 2.900 46.330 3.350 ;
        RECT 39.580 2.750 49.880 2.900 ;
        RECT 43.130 2.300 46.330 2.750 ;
        RECT 39.580 2.150 49.880 2.300 ;
        RECT 43.530 1.200 45.930 2.150 ;
        RECT 50.480 1.600 50.630 9.800 ;
        RECT 51.080 1.600 51.230 9.800 ;
        RECT 51.680 1.600 51.830 9.800 ;
        RECT 52.280 1.600 52.430 9.800 ;
        RECT 52.880 1.600 53.030 9.800 ;
        RECT 53.480 1.600 53.630 9.800 ;
        RECT 54.080 1.600 54.230 9.800 ;
        RECT 55.230 10.200 55.380 18.400 ;
        RECT 55.830 10.200 55.980 18.400 ;
        RECT 56.430 10.200 56.580 18.400 ;
        RECT 57.030 10.200 57.180 18.400 ;
        RECT 57.630 10.200 57.780 18.400 ;
        RECT 58.230 10.200 58.380 18.400 ;
        RECT 58.830 10.200 58.980 18.400 ;
        RECT 63.530 17.850 65.940 18.800 ;
        RECT 59.580 17.700 69.880 17.850 ;
        RECT 63.130 17.250 66.330 17.700 ;
        RECT 59.580 17.100 69.880 17.250 ;
        RECT 63.130 16.650 66.330 17.100 ;
        RECT 59.580 16.500 69.880 16.650 ;
        RECT 63.130 16.050 66.330 16.500 ;
        RECT 59.580 15.900 69.880 16.050 ;
        RECT 63.130 15.600 66.330 15.900 ;
        RECT 63.130 15.450 63.530 15.600 ;
        RECT 59.580 15.300 63.530 15.450 ;
        RECT 63.130 14.850 63.530 15.300 ;
        RECT 59.580 14.700 63.530 14.850 ;
        RECT 63.130 14.250 63.530 14.700 ;
        RECT 59.580 14.100 63.530 14.250 ;
        RECT 63.130 13.650 63.530 14.100 ;
        RECT 59.580 13.500 63.530 13.650 ;
        RECT 63.130 13.050 63.530 13.500 ;
        RECT 59.580 12.900 63.530 13.050 ;
        RECT 63.130 12.450 63.530 12.900 ;
        RECT 59.580 12.300 63.530 12.450 ;
        RECT 63.130 11.850 63.530 12.300 ;
        RECT 59.580 11.700 63.530 11.850 ;
        RECT 63.130 11.250 63.530 11.700 ;
        RECT 59.580 11.100 63.530 11.250 ;
        RECT 63.130 10.650 63.530 11.100 ;
        RECT 59.580 10.500 63.530 10.650 ;
        RECT 63.130 10.200 63.530 10.500 ;
        RECT 55.230 9.800 63.530 10.200 ;
        RECT 55.230 1.600 55.380 9.800 ;
        RECT 55.830 1.600 55.980 9.800 ;
        RECT 56.430 1.600 56.580 9.800 ;
        RECT 57.030 1.600 57.180 9.800 ;
        RECT 57.630 1.600 57.780 9.800 ;
        RECT 58.230 1.600 58.380 9.800 ;
        RECT 58.830 1.600 58.980 9.800 ;
        RECT 63.130 9.500 63.530 9.800 ;
        RECT 59.580 9.350 63.530 9.500 ;
        RECT 63.130 8.900 63.530 9.350 ;
        RECT 59.580 8.750 63.530 8.900 ;
        RECT 63.130 8.300 63.530 8.750 ;
        RECT 59.580 8.150 63.530 8.300 ;
        RECT 63.130 7.700 63.530 8.150 ;
        RECT 59.580 7.550 63.530 7.700 ;
        RECT 63.130 7.100 63.530 7.550 ;
        RECT 59.580 6.950 63.530 7.100 ;
        RECT 63.130 6.500 63.530 6.950 ;
        RECT 59.580 6.350 63.530 6.500 ;
        RECT 63.130 5.900 63.530 6.350 ;
        RECT 59.580 5.750 63.530 5.900 ;
        RECT 63.130 5.300 63.530 5.750 ;
        RECT 59.580 5.150 63.530 5.300 ;
        RECT 63.130 4.700 63.530 5.150 ;
        RECT 59.580 4.550 63.530 4.700 ;
        RECT 63.130 4.400 63.530 4.550 ;
        RECT 65.930 15.450 66.330 15.600 ;
        RECT 65.930 15.300 69.880 15.450 ;
        RECT 65.930 14.850 66.330 15.300 ;
        RECT 65.930 14.700 69.880 14.850 ;
        RECT 65.930 14.250 66.330 14.700 ;
        RECT 65.930 14.100 69.880 14.250 ;
        RECT 65.930 13.650 66.330 14.100 ;
        RECT 65.930 13.500 69.880 13.650 ;
        RECT 65.930 13.050 66.330 13.500 ;
        RECT 65.930 12.900 69.880 13.050 ;
        RECT 65.930 12.450 66.330 12.900 ;
        RECT 65.930 12.300 69.880 12.450 ;
        RECT 65.930 11.850 66.330 12.300 ;
        RECT 65.930 11.700 69.880 11.850 ;
        RECT 65.930 11.250 66.330 11.700 ;
        RECT 65.930 11.100 69.880 11.250 ;
        RECT 65.930 10.650 66.330 11.100 ;
        RECT 65.930 10.500 69.880 10.650 ;
        RECT 65.930 10.200 66.330 10.500 ;
        RECT 70.480 10.200 70.630 18.400 ;
        RECT 71.080 10.200 71.230 18.400 ;
        RECT 71.680 10.200 71.830 18.400 ;
        RECT 72.280 10.200 72.430 18.400 ;
        RECT 72.880 10.200 73.030 18.400 ;
        RECT 73.480 10.200 73.630 18.400 ;
        RECT 74.080 10.200 74.230 18.400 ;
        RECT 65.930 9.800 74.230 10.200 ;
        RECT 65.930 9.500 66.330 9.800 ;
        RECT 65.930 9.350 69.880 9.500 ;
        RECT 65.930 8.900 66.330 9.350 ;
        RECT 65.930 8.750 69.880 8.900 ;
        RECT 65.930 8.300 66.330 8.750 ;
        RECT 65.930 8.150 69.880 8.300 ;
        RECT 65.930 7.700 66.330 8.150 ;
        RECT 65.930 7.550 69.880 7.700 ;
        RECT 65.930 7.100 66.330 7.550 ;
        RECT 65.930 6.950 69.880 7.100 ;
        RECT 65.930 6.500 66.330 6.950 ;
        RECT 65.930 6.350 69.880 6.500 ;
        RECT 65.930 5.900 66.330 6.350 ;
        RECT 65.930 5.750 69.880 5.900 ;
        RECT 65.930 5.300 66.330 5.750 ;
        RECT 65.930 5.150 69.880 5.300 ;
        RECT 65.930 4.700 66.330 5.150 ;
        RECT 65.930 4.550 69.880 4.700 ;
        RECT 65.930 4.400 66.330 4.550 ;
        RECT 63.130 4.100 66.330 4.400 ;
        RECT 59.580 3.950 69.880 4.100 ;
        RECT 63.130 3.500 66.330 3.950 ;
        RECT 59.580 3.350 69.880 3.500 ;
        RECT 63.130 2.900 66.330 3.350 ;
        RECT 59.580 2.750 69.880 2.900 ;
        RECT 63.130 2.300 66.330 2.750 ;
        RECT 59.580 2.150 69.880 2.300 ;
        RECT 63.530 1.200 65.930 2.150 ;
        RECT 70.480 1.600 70.630 9.800 ;
        RECT 71.080 1.600 71.230 9.800 ;
        RECT 71.680 1.600 71.830 9.800 ;
        RECT 72.280 1.600 72.430 9.800 ;
        RECT 72.880 1.600 73.030 9.800 ;
        RECT 73.480 1.600 73.630 9.800 ;
        RECT 74.080 1.600 74.230 9.800 ;
        RECT 75.230 10.200 75.380 18.400 ;
        RECT 75.830 10.200 75.980 18.400 ;
        RECT 76.430 10.200 76.580 18.400 ;
        RECT 77.030 10.200 77.180 18.400 ;
        RECT 77.630 10.200 77.780 18.400 ;
        RECT 78.230 10.200 78.380 18.400 ;
        RECT 78.830 10.200 78.980 18.400 ;
        RECT 83.530 17.850 85.940 18.800 ;
        RECT 79.580 17.700 89.880 17.850 ;
        RECT 83.130 17.250 86.330 17.700 ;
        RECT 79.580 17.100 89.880 17.250 ;
        RECT 83.130 16.650 86.330 17.100 ;
        RECT 79.580 16.500 89.880 16.650 ;
        RECT 83.130 16.050 86.330 16.500 ;
        RECT 79.580 15.900 89.880 16.050 ;
        RECT 83.130 15.600 86.330 15.900 ;
        RECT 83.130 15.450 83.530 15.600 ;
        RECT 79.580 15.300 83.530 15.450 ;
        RECT 83.130 14.850 83.530 15.300 ;
        RECT 79.580 14.700 83.530 14.850 ;
        RECT 83.130 14.250 83.530 14.700 ;
        RECT 79.580 14.100 83.530 14.250 ;
        RECT 83.130 13.650 83.530 14.100 ;
        RECT 79.580 13.500 83.530 13.650 ;
        RECT 83.130 13.050 83.530 13.500 ;
        RECT 79.580 12.900 83.530 13.050 ;
        RECT 83.130 12.450 83.530 12.900 ;
        RECT 79.580 12.300 83.530 12.450 ;
        RECT 83.130 11.850 83.530 12.300 ;
        RECT 79.580 11.700 83.530 11.850 ;
        RECT 83.130 11.250 83.530 11.700 ;
        RECT 79.580 11.100 83.530 11.250 ;
        RECT 83.130 10.650 83.530 11.100 ;
        RECT 79.580 10.500 83.530 10.650 ;
        RECT 83.130 10.200 83.530 10.500 ;
        RECT 75.230 9.800 83.530 10.200 ;
        RECT 75.230 1.600 75.380 9.800 ;
        RECT 75.830 1.600 75.980 9.800 ;
        RECT 76.430 1.600 76.580 9.800 ;
        RECT 77.030 1.600 77.180 9.800 ;
        RECT 77.630 1.600 77.780 9.800 ;
        RECT 78.230 1.600 78.380 9.800 ;
        RECT 78.830 1.600 78.980 9.800 ;
        RECT 83.130 9.500 83.530 9.800 ;
        RECT 79.580 9.350 83.530 9.500 ;
        RECT 83.130 8.900 83.530 9.350 ;
        RECT 79.580 8.750 83.530 8.900 ;
        RECT 83.130 8.300 83.530 8.750 ;
        RECT 79.580 8.150 83.530 8.300 ;
        RECT 83.130 7.700 83.530 8.150 ;
        RECT 79.580 7.550 83.530 7.700 ;
        RECT 83.130 7.100 83.530 7.550 ;
        RECT 79.580 6.950 83.530 7.100 ;
        RECT 83.130 6.500 83.530 6.950 ;
        RECT 79.580 6.350 83.530 6.500 ;
        RECT 83.130 5.900 83.530 6.350 ;
        RECT 79.580 5.750 83.530 5.900 ;
        RECT 83.130 5.300 83.530 5.750 ;
        RECT 79.580 5.150 83.530 5.300 ;
        RECT 83.130 4.700 83.530 5.150 ;
        RECT 79.580 4.550 83.530 4.700 ;
        RECT 83.130 4.400 83.530 4.550 ;
        RECT 85.930 15.450 86.330 15.600 ;
        RECT 85.930 15.300 89.880 15.450 ;
        RECT 85.930 14.850 86.330 15.300 ;
        RECT 85.930 14.700 89.880 14.850 ;
        RECT 85.930 14.250 86.330 14.700 ;
        RECT 85.930 14.100 89.880 14.250 ;
        RECT 85.930 13.650 86.330 14.100 ;
        RECT 85.930 13.500 89.880 13.650 ;
        RECT 85.930 13.050 86.330 13.500 ;
        RECT 85.930 12.900 89.880 13.050 ;
        RECT 85.930 12.450 86.330 12.900 ;
        RECT 85.930 12.300 89.880 12.450 ;
        RECT 85.930 11.850 86.330 12.300 ;
        RECT 85.930 11.700 89.880 11.850 ;
        RECT 85.930 11.250 86.330 11.700 ;
        RECT 85.930 11.100 89.880 11.250 ;
        RECT 85.930 10.650 86.330 11.100 ;
        RECT 85.930 10.500 89.880 10.650 ;
        RECT 85.930 10.200 86.330 10.500 ;
        RECT 90.480 10.200 90.630 18.400 ;
        RECT 91.080 10.200 91.230 18.400 ;
        RECT 91.680 10.200 91.830 18.400 ;
        RECT 92.280 10.200 92.430 18.400 ;
        RECT 92.880 10.200 93.030 18.400 ;
        RECT 93.480 10.200 93.630 18.400 ;
        RECT 94.080 10.200 94.230 18.400 ;
        RECT 85.930 9.800 94.230 10.200 ;
        RECT 85.930 9.500 86.330 9.800 ;
        RECT 85.930 9.350 89.880 9.500 ;
        RECT 85.930 8.900 86.330 9.350 ;
        RECT 85.930 8.750 89.880 8.900 ;
        RECT 85.930 8.300 86.330 8.750 ;
        RECT 85.930 8.150 89.880 8.300 ;
        RECT 85.930 7.700 86.330 8.150 ;
        RECT 85.930 7.550 89.880 7.700 ;
        RECT 85.930 7.100 86.330 7.550 ;
        RECT 85.930 6.950 89.880 7.100 ;
        RECT 85.930 6.500 86.330 6.950 ;
        RECT 85.930 6.350 89.880 6.500 ;
        RECT 85.930 5.900 86.330 6.350 ;
        RECT 85.930 5.750 89.880 5.900 ;
        RECT 85.930 5.300 86.330 5.750 ;
        RECT 85.930 5.150 89.880 5.300 ;
        RECT 85.930 4.700 86.330 5.150 ;
        RECT 85.930 4.550 89.880 4.700 ;
        RECT 85.930 4.400 86.330 4.550 ;
        RECT 83.130 4.100 86.330 4.400 ;
        RECT 79.580 3.950 89.880 4.100 ;
        RECT 83.130 3.500 86.330 3.950 ;
        RECT 79.580 3.350 89.880 3.500 ;
        RECT 83.130 2.900 86.330 3.350 ;
        RECT 79.580 2.750 89.880 2.900 ;
        RECT 83.130 2.300 86.330 2.750 ;
        RECT 79.580 2.150 89.880 2.300 ;
        RECT 83.530 1.200 85.930 2.150 ;
        RECT 90.480 1.600 90.630 9.800 ;
        RECT 91.080 1.600 91.230 9.800 ;
        RECT 91.680 1.600 91.830 9.800 ;
        RECT 92.280 1.600 92.430 9.800 ;
        RECT 92.880 1.600 93.030 9.800 ;
        RECT 93.480 1.600 93.630 9.800 ;
        RECT 94.080 1.600 94.230 9.800 ;
        RECT 95.230 10.200 95.380 18.400 ;
        RECT 95.830 10.200 95.980 18.400 ;
        RECT 96.430 10.200 96.580 18.400 ;
        RECT 97.030 10.200 97.180 18.400 ;
        RECT 97.630 10.200 97.780 18.400 ;
        RECT 98.230 10.200 98.380 18.400 ;
        RECT 98.830 10.200 98.980 18.400 ;
        RECT 103.530 17.850 105.940 18.800 ;
        RECT 99.580 17.700 109.880 17.850 ;
        RECT 103.130 17.250 106.330 17.700 ;
        RECT 99.580 17.100 109.880 17.250 ;
        RECT 103.130 16.650 106.330 17.100 ;
        RECT 99.580 16.500 109.880 16.650 ;
        RECT 103.130 16.050 106.330 16.500 ;
        RECT 99.580 15.900 109.880 16.050 ;
        RECT 103.130 15.600 106.330 15.900 ;
        RECT 103.130 15.450 103.530 15.600 ;
        RECT 99.580 15.300 103.530 15.450 ;
        RECT 103.130 14.850 103.530 15.300 ;
        RECT 99.580 14.700 103.530 14.850 ;
        RECT 103.130 14.250 103.530 14.700 ;
        RECT 99.580 14.100 103.530 14.250 ;
        RECT 103.130 13.650 103.530 14.100 ;
        RECT 99.580 13.500 103.530 13.650 ;
        RECT 103.130 13.050 103.530 13.500 ;
        RECT 99.580 12.900 103.530 13.050 ;
        RECT 103.130 12.450 103.530 12.900 ;
        RECT 99.580 12.300 103.530 12.450 ;
        RECT 103.130 11.850 103.530 12.300 ;
        RECT 99.580 11.700 103.530 11.850 ;
        RECT 103.130 11.250 103.530 11.700 ;
        RECT 99.580 11.100 103.530 11.250 ;
        RECT 103.130 10.650 103.530 11.100 ;
        RECT 99.580 10.500 103.530 10.650 ;
        RECT 103.130 10.200 103.530 10.500 ;
        RECT 95.230 9.800 103.530 10.200 ;
        RECT 95.230 1.600 95.380 9.800 ;
        RECT 95.830 1.600 95.980 9.800 ;
        RECT 96.430 1.600 96.580 9.800 ;
        RECT 97.030 1.600 97.180 9.800 ;
        RECT 97.630 1.600 97.780 9.800 ;
        RECT 98.230 1.600 98.380 9.800 ;
        RECT 98.830 1.600 98.980 9.800 ;
        RECT 103.130 9.500 103.530 9.800 ;
        RECT 99.580 9.350 103.530 9.500 ;
        RECT 103.130 8.900 103.530 9.350 ;
        RECT 99.580 8.750 103.530 8.900 ;
        RECT 103.130 8.300 103.530 8.750 ;
        RECT 99.580 8.150 103.530 8.300 ;
        RECT 103.130 7.700 103.530 8.150 ;
        RECT 99.580 7.550 103.530 7.700 ;
        RECT 103.130 7.100 103.530 7.550 ;
        RECT 99.580 6.950 103.530 7.100 ;
        RECT 103.130 6.500 103.530 6.950 ;
        RECT 99.580 6.350 103.530 6.500 ;
        RECT 103.130 5.900 103.530 6.350 ;
        RECT 99.580 5.750 103.530 5.900 ;
        RECT 103.130 5.300 103.530 5.750 ;
        RECT 99.580 5.150 103.530 5.300 ;
        RECT 103.130 4.700 103.530 5.150 ;
        RECT 99.580 4.550 103.530 4.700 ;
        RECT 103.130 4.400 103.530 4.550 ;
        RECT 105.930 15.450 106.330 15.600 ;
        RECT 105.930 15.300 109.880 15.450 ;
        RECT 105.930 14.850 106.330 15.300 ;
        RECT 105.930 14.700 109.880 14.850 ;
        RECT 105.930 14.250 106.330 14.700 ;
        RECT 105.930 14.100 109.880 14.250 ;
        RECT 105.930 13.650 106.330 14.100 ;
        RECT 105.930 13.500 109.880 13.650 ;
        RECT 105.930 13.050 106.330 13.500 ;
        RECT 105.930 12.900 109.880 13.050 ;
        RECT 105.930 12.450 106.330 12.900 ;
        RECT 105.930 12.300 109.880 12.450 ;
        RECT 105.930 11.850 106.330 12.300 ;
        RECT 105.930 11.700 109.880 11.850 ;
        RECT 105.930 11.250 106.330 11.700 ;
        RECT 105.930 11.100 109.880 11.250 ;
        RECT 105.930 10.650 106.330 11.100 ;
        RECT 105.930 10.500 109.880 10.650 ;
        RECT 105.930 10.200 106.330 10.500 ;
        RECT 110.480 10.200 110.630 18.400 ;
        RECT 111.080 10.200 111.230 18.400 ;
        RECT 111.680 10.200 111.830 18.400 ;
        RECT 112.280 10.200 112.430 18.400 ;
        RECT 112.880 10.200 113.030 18.400 ;
        RECT 113.480 10.200 113.630 18.400 ;
        RECT 114.080 10.200 114.230 18.400 ;
        RECT 105.930 9.800 114.230 10.200 ;
        RECT 105.930 9.500 106.330 9.800 ;
        RECT 105.930 9.350 109.880 9.500 ;
        RECT 105.930 8.900 106.330 9.350 ;
        RECT 105.930 8.750 109.880 8.900 ;
        RECT 105.930 8.300 106.330 8.750 ;
        RECT 105.930 8.150 109.880 8.300 ;
        RECT 105.930 7.700 106.330 8.150 ;
        RECT 105.930 7.550 109.880 7.700 ;
        RECT 105.930 7.100 106.330 7.550 ;
        RECT 105.930 6.950 109.880 7.100 ;
        RECT 105.930 6.500 106.330 6.950 ;
        RECT 105.930 6.350 109.880 6.500 ;
        RECT 105.930 5.900 106.330 6.350 ;
        RECT 105.930 5.750 109.880 5.900 ;
        RECT 105.930 5.300 106.330 5.750 ;
        RECT 105.930 5.150 109.880 5.300 ;
        RECT 105.930 4.700 106.330 5.150 ;
        RECT 105.930 4.550 109.880 4.700 ;
        RECT 105.930 4.400 106.330 4.550 ;
        RECT 103.130 4.100 106.330 4.400 ;
        RECT 99.580 3.950 109.880 4.100 ;
        RECT 103.130 3.500 106.330 3.950 ;
        RECT 99.580 3.350 109.880 3.500 ;
        RECT 103.130 2.900 106.330 3.350 ;
        RECT 99.580 2.750 109.880 2.900 ;
        RECT 103.130 2.300 106.330 2.750 ;
        RECT 99.580 2.150 109.880 2.300 ;
        RECT 103.530 1.200 105.930 2.150 ;
        RECT 110.480 1.600 110.630 9.800 ;
        RECT 111.080 1.600 111.230 9.800 ;
        RECT 111.680 1.600 111.830 9.800 ;
        RECT 112.280 1.600 112.430 9.800 ;
        RECT 112.880 1.600 113.030 9.800 ;
        RECT 113.480 1.600 113.630 9.800 ;
        RECT 114.080 1.600 114.230 9.800 ;
        RECT 115.230 10.200 115.380 18.400 ;
        RECT 115.830 10.200 115.980 18.400 ;
        RECT 116.430 10.200 116.580 18.400 ;
        RECT 117.030 10.200 117.180 18.400 ;
        RECT 117.630 10.200 117.780 18.400 ;
        RECT 118.230 10.200 118.380 18.400 ;
        RECT 118.830 10.200 118.980 18.400 ;
        RECT 123.530 17.850 124.730 18.800 ;
        RECT 119.580 17.700 124.730 17.850 ;
        RECT 123.130 17.250 124.730 17.700 ;
        RECT 119.580 17.100 124.730 17.250 ;
        RECT 123.130 16.650 124.730 17.100 ;
        RECT 119.580 16.500 124.730 16.650 ;
        RECT 123.130 16.050 124.730 16.500 ;
        RECT 119.580 15.900 124.730 16.050 ;
        RECT 125.135 16.035 127.135 17.310 ;
        RECT 123.130 15.600 124.730 15.900 ;
        RECT 123.130 15.450 123.530 15.600 ;
        RECT 119.580 15.300 123.530 15.450 ;
        RECT 123.130 14.850 123.530 15.300 ;
        RECT 119.580 14.700 123.530 14.850 ;
        RECT 123.130 14.250 123.530 14.700 ;
        RECT 119.580 14.100 123.530 14.250 ;
        RECT 123.130 13.650 123.530 14.100 ;
        RECT 119.580 13.500 123.530 13.650 ;
        RECT 123.130 13.050 123.530 13.500 ;
        RECT 119.580 12.900 123.530 13.050 ;
        RECT 123.130 12.450 123.530 12.900 ;
        RECT 119.580 12.300 123.530 12.450 ;
        RECT 123.130 11.850 123.530 12.300 ;
        RECT 119.580 11.700 123.530 11.850 ;
        RECT 123.130 11.250 123.530 11.700 ;
        RECT 119.580 11.100 123.530 11.250 ;
        RECT 123.130 10.650 123.530 11.100 ;
        RECT 119.580 10.500 123.530 10.650 ;
        RECT 123.130 10.200 123.530 10.500 ;
        RECT 115.230 9.800 123.530 10.200 ;
        RECT 115.230 1.600 115.380 9.800 ;
        RECT 115.830 1.600 115.980 9.800 ;
        RECT 116.430 1.600 116.580 9.800 ;
        RECT 117.030 1.600 117.180 9.800 ;
        RECT 117.630 1.600 117.780 9.800 ;
        RECT 118.230 1.600 118.380 9.800 ;
        RECT 118.830 1.600 118.980 9.800 ;
        RECT 123.130 9.500 123.530 9.800 ;
        RECT 119.580 9.350 123.530 9.500 ;
        RECT 123.130 8.900 123.530 9.350 ;
        RECT 119.580 8.750 123.530 8.900 ;
        RECT 123.130 8.300 123.530 8.750 ;
        RECT 119.580 8.150 123.530 8.300 ;
        RECT 123.130 7.700 123.530 8.150 ;
        RECT 119.580 7.550 123.530 7.700 ;
        RECT 123.130 7.100 123.530 7.550 ;
        RECT 119.580 6.950 123.530 7.100 ;
        RECT 123.130 6.500 123.530 6.950 ;
        RECT 119.580 6.350 123.530 6.500 ;
        RECT 123.130 5.900 123.530 6.350 ;
        RECT 119.580 5.750 123.530 5.900 ;
        RECT 123.130 5.300 123.530 5.750 ;
        RECT 119.580 5.150 123.530 5.300 ;
        RECT 123.130 4.700 123.530 5.150 ;
        RECT 119.580 4.550 123.530 4.700 ;
        RECT 123.130 4.400 123.530 4.550 ;
        RECT 123.130 4.100 124.730 4.400 ;
        RECT 119.580 3.950 124.730 4.100 ;
        RECT 123.130 3.500 124.730 3.950 ;
        RECT 119.580 3.350 124.730 3.500 ;
        RECT 123.130 2.900 124.730 3.350 ;
        RECT 119.580 2.750 124.730 2.900 ;
        RECT 123.130 2.300 124.730 2.750 ;
        RECT 119.580 2.150 124.730 2.300 ;
        RECT 123.530 1.200 124.730 2.150 ;
        RECT 125.140 1.820 127.140 3.095 ;
        RECT 4.730 0.000 9.130 1.200 ;
        RECT 20.330 0.000 29.130 1.200 ;
        RECT 40.330 0.000 49.130 1.200 ;
        RECT 60.330 0.000 69.130 1.200 ;
        RECT 80.330 0.000 89.130 1.200 ;
        RECT 100.330 0.000 109.130 1.200 ;
        RECT 120.330 0.000 124.730 1.200 ;
      LAYER via2 ;
        RECT 2.515 336.880 2.875 337.260 ;
        RECT 3.145 336.880 3.505 337.260 ;
        RECT 3.745 336.880 4.105 337.260 ;
        RECT 2.515 336.290 2.875 336.670 ;
        RECT 3.145 336.290 3.505 336.670 ;
        RECT 3.745 336.290 4.105 336.670 ;
        RECT 2.520 334.920 2.880 335.300 ;
        RECT 3.130 334.920 3.490 335.300 ;
        RECT 3.760 334.920 4.120 335.300 ;
        RECT 2.520 334.185 2.880 334.565 ;
        RECT 3.130 334.185 3.490 334.565 ;
        RECT 3.760 334.185 4.120 334.565 ;
        RECT 2.520 333.500 2.880 333.880 ;
        RECT 3.130 333.500 3.490 333.880 ;
        RECT 3.760 333.500 4.120 333.880 ;
        RECT 2.520 326.120 2.880 326.500 ;
        RECT 3.130 326.120 3.490 326.500 ;
        RECT 3.760 326.120 4.120 326.500 ;
        RECT 2.520 325.385 2.880 325.765 ;
        RECT 3.130 325.385 3.490 325.765 ;
        RECT 3.760 325.385 4.120 325.765 ;
        RECT 2.520 324.700 2.880 325.080 ;
        RECT 3.130 324.700 3.490 325.080 ;
        RECT 3.760 324.700 4.120 325.080 ;
        RECT 2.515 323.515 2.875 323.895 ;
        RECT 3.145 323.515 3.505 323.895 ;
        RECT 3.745 323.515 4.105 323.895 ;
        RECT 2.515 322.925 2.875 323.305 ;
        RECT 3.145 322.925 3.505 323.305 ;
        RECT 3.745 322.925 4.105 323.305 ;
        RECT 125.340 337.080 125.700 337.460 ;
        RECT 125.970 337.080 126.330 337.460 ;
        RECT 126.570 337.080 126.930 337.460 ;
        RECT 125.340 336.490 125.700 336.870 ;
        RECT 125.970 336.490 126.330 336.870 ;
        RECT 126.570 336.490 126.930 336.870 ;
        RECT 125.340 323.095 125.700 323.475 ;
        RECT 125.970 323.095 126.330 323.475 ;
        RECT 126.570 323.095 126.930 323.475 ;
        RECT 125.340 322.505 125.700 322.885 ;
        RECT 125.970 322.505 126.330 322.885 ;
        RECT 126.570 322.505 126.930 322.885 ;
        RECT 2.515 316.870 2.875 317.250 ;
        RECT 3.145 316.870 3.505 317.250 ;
        RECT 3.745 316.870 4.105 317.250 ;
        RECT 2.515 316.280 2.875 316.660 ;
        RECT 3.145 316.280 3.505 316.660 ;
        RECT 3.745 316.280 4.105 316.660 ;
        RECT 2.520 314.920 2.880 315.300 ;
        RECT 3.130 314.920 3.490 315.300 ;
        RECT 3.760 314.920 4.120 315.300 ;
        RECT 2.520 314.185 2.880 314.565 ;
        RECT 3.130 314.185 3.490 314.565 ;
        RECT 3.760 314.185 4.120 314.565 ;
        RECT 2.520 313.500 2.880 313.880 ;
        RECT 3.130 313.500 3.490 313.880 ;
        RECT 3.760 313.500 4.120 313.880 ;
        RECT 2.520 306.125 2.880 306.505 ;
        RECT 3.130 306.125 3.490 306.505 ;
        RECT 3.760 306.125 4.120 306.505 ;
        RECT 2.520 305.390 2.880 305.770 ;
        RECT 3.130 305.390 3.490 305.770 ;
        RECT 3.760 305.390 4.120 305.770 ;
        RECT 2.520 304.705 2.880 305.085 ;
        RECT 3.130 304.705 3.490 305.085 ;
        RECT 3.760 304.705 4.120 305.085 ;
        RECT 2.515 303.170 2.875 303.550 ;
        RECT 3.145 303.170 3.505 303.550 ;
        RECT 3.745 303.170 4.105 303.550 ;
        RECT 2.515 302.580 2.875 302.960 ;
        RECT 3.145 302.580 3.505 302.960 ;
        RECT 3.745 302.580 4.105 302.960 ;
        RECT 125.340 317.080 125.700 317.460 ;
        RECT 125.970 317.080 126.330 317.460 ;
        RECT 126.570 317.080 126.930 317.460 ;
        RECT 125.340 316.490 125.700 316.870 ;
        RECT 125.970 316.490 126.330 316.870 ;
        RECT 126.570 316.490 126.930 316.870 ;
        RECT 125.340 303.095 125.700 303.475 ;
        RECT 125.970 303.095 126.330 303.475 ;
        RECT 126.570 303.095 126.930 303.475 ;
        RECT 125.340 302.505 125.700 302.885 ;
        RECT 125.970 302.505 126.330 302.885 ;
        RECT 126.570 302.505 126.930 302.885 ;
        RECT 2.515 297.280 2.875 297.660 ;
        RECT 3.145 297.280 3.505 297.660 ;
        RECT 3.745 297.280 4.105 297.660 ;
        RECT 2.515 296.690 2.875 297.070 ;
        RECT 3.145 296.690 3.505 297.070 ;
        RECT 3.745 296.690 4.105 297.070 ;
        RECT 2.520 294.920 2.880 295.300 ;
        RECT 3.130 294.920 3.490 295.300 ;
        RECT 3.760 294.920 4.120 295.300 ;
        RECT 2.520 294.185 2.880 294.565 ;
        RECT 3.130 294.185 3.490 294.565 ;
        RECT 3.760 294.185 4.120 294.565 ;
        RECT 2.520 293.500 2.880 293.880 ;
        RECT 3.130 293.500 3.490 293.880 ;
        RECT 3.760 293.500 4.120 293.880 ;
        RECT 2.520 286.125 2.880 286.505 ;
        RECT 3.130 286.125 3.490 286.505 ;
        RECT 3.760 286.125 4.120 286.505 ;
        RECT 2.520 285.390 2.880 285.770 ;
        RECT 3.130 285.390 3.490 285.770 ;
        RECT 3.760 285.390 4.120 285.770 ;
        RECT 2.520 284.705 2.880 285.085 ;
        RECT 3.130 284.705 3.490 285.085 ;
        RECT 3.760 284.705 4.120 285.085 ;
        RECT 2.515 283.040 2.875 283.420 ;
        RECT 3.145 283.040 3.505 283.420 ;
        RECT 3.745 283.040 4.105 283.420 ;
        RECT 2.515 282.450 2.875 282.830 ;
        RECT 3.145 282.450 3.505 282.830 ;
        RECT 3.745 282.450 4.105 282.830 ;
        RECT 125.340 297.080 125.700 297.460 ;
        RECT 125.970 297.080 126.330 297.460 ;
        RECT 126.570 297.080 126.930 297.460 ;
        RECT 125.340 296.490 125.700 296.870 ;
        RECT 125.970 296.490 126.330 296.870 ;
        RECT 126.570 296.490 126.930 296.870 ;
        RECT 125.340 283.095 125.700 283.475 ;
        RECT 125.970 283.095 126.330 283.475 ;
        RECT 126.570 283.095 126.930 283.475 ;
        RECT 125.340 282.505 125.700 282.885 ;
        RECT 125.970 282.505 126.330 282.885 ;
        RECT 126.570 282.505 126.930 282.885 ;
        RECT 2.515 277.025 2.875 277.405 ;
        RECT 3.145 277.025 3.505 277.405 ;
        RECT 3.745 277.025 4.105 277.405 ;
        RECT 2.515 276.435 2.875 276.815 ;
        RECT 3.145 276.435 3.505 276.815 ;
        RECT 3.745 276.435 4.105 276.815 ;
        RECT 2.520 274.920 2.880 275.300 ;
        RECT 3.130 274.920 3.490 275.300 ;
        RECT 3.760 274.920 4.120 275.300 ;
        RECT 2.520 274.185 2.880 274.565 ;
        RECT 3.130 274.185 3.490 274.565 ;
        RECT 3.760 274.185 4.120 274.565 ;
        RECT 2.520 273.500 2.880 273.880 ;
        RECT 3.130 273.500 3.490 273.880 ;
        RECT 3.760 273.500 4.120 273.880 ;
        RECT 2.520 266.115 2.880 266.495 ;
        RECT 3.130 266.115 3.490 266.495 ;
        RECT 3.760 266.115 4.120 266.495 ;
        RECT 2.520 265.380 2.880 265.760 ;
        RECT 3.130 265.380 3.490 265.760 ;
        RECT 3.760 265.380 4.120 265.760 ;
        RECT 2.520 264.695 2.880 265.075 ;
        RECT 3.130 264.695 3.490 265.075 ;
        RECT 3.760 264.695 4.120 265.075 ;
        RECT 2.515 263.140 2.875 263.520 ;
        RECT 3.145 263.140 3.505 263.520 ;
        RECT 3.745 263.140 4.105 263.520 ;
        RECT 2.515 262.550 2.875 262.930 ;
        RECT 3.145 262.550 3.505 262.930 ;
        RECT 3.745 262.550 4.105 262.930 ;
        RECT 125.340 277.350 125.700 277.730 ;
        RECT 125.970 277.350 126.330 277.730 ;
        RECT 126.570 277.350 126.930 277.730 ;
        RECT 125.340 276.760 125.700 277.140 ;
        RECT 125.970 276.760 126.330 277.140 ;
        RECT 126.570 276.760 126.930 277.140 ;
        RECT 125.340 262.770 125.700 263.150 ;
        RECT 125.970 262.770 126.330 263.150 ;
        RECT 126.570 262.770 126.930 263.150 ;
        RECT 125.340 262.180 125.700 262.560 ;
        RECT 125.970 262.180 126.330 262.560 ;
        RECT 126.570 262.180 126.930 262.560 ;
        RECT 2.515 257.105 2.875 257.485 ;
        RECT 3.145 257.105 3.505 257.485 ;
        RECT 3.745 257.105 4.105 257.485 ;
        RECT 2.515 256.515 2.875 256.895 ;
        RECT 3.145 256.515 3.505 256.895 ;
        RECT 3.745 256.515 4.105 256.895 ;
        RECT 2.520 254.920 2.880 255.300 ;
        RECT 3.130 254.920 3.490 255.300 ;
        RECT 3.760 254.920 4.120 255.300 ;
        RECT 2.520 254.185 2.880 254.565 ;
        RECT 3.130 254.185 3.490 254.565 ;
        RECT 3.760 254.185 4.120 254.565 ;
        RECT 2.520 253.500 2.880 253.880 ;
        RECT 3.130 253.500 3.490 253.880 ;
        RECT 3.760 253.500 4.120 253.880 ;
        RECT 2.520 246.125 2.880 246.505 ;
        RECT 3.130 246.125 3.490 246.505 ;
        RECT 3.760 246.125 4.120 246.505 ;
        RECT 2.520 245.390 2.880 245.770 ;
        RECT 3.130 245.390 3.490 245.770 ;
        RECT 3.760 245.390 4.120 245.770 ;
        RECT 2.520 244.705 2.880 245.085 ;
        RECT 3.130 244.705 3.490 245.085 ;
        RECT 3.760 244.705 4.120 245.085 ;
        RECT 2.515 243.275 2.875 243.655 ;
        RECT 3.145 243.275 3.505 243.655 ;
        RECT 3.745 243.275 4.105 243.655 ;
        RECT 2.515 242.685 2.875 243.065 ;
        RECT 3.145 242.685 3.505 243.065 ;
        RECT 3.745 242.685 4.105 243.065 ;
        RECT 125.340 256.855 125.700 257.235 ;
        RECT 125.970 256.855 126.330 257.235 ;
        RECT 126.570 256.855 126.930 257.235 ;
        RECT 125.340 256.265 125.700 256.645 ;
        RECT 125.970 256.265 126.330 256.645 ;
        RECT 126.570 256.265 126.930 256.645 ;
        RECT 125.340 242.495 125.700 242.875 ;
        RECT 125.970 242.495 126.330 242.875 ;
        RECT 126.570 242.495 126.930 242.875 ;
        RECT 125.340 241.905 125.700 242.285 ;
        RECT 125.970 241.905 126.330 242.285 ;
        RECT 126.570 241.905 126.930 242.285 ;
        RECT 2.515 237.340 2.875 237.720 ;
        RECT 3.145 237.340 3.505 237.720 ;
        RECT 3.745 237.340 4.105 237.720 ;
        RECT 2.515 236.750 2.875 237.130 ;
        RECT 3.145 236.750 3.505 237.130 ;
        RECT 3.745 236.750 4.105 237.130 ;
        RECT 2.520 234.920 2.880 235.300 ;
        RECT 3.130 234.920 3.490 235.300 ;
        RECT 3.760 234.920 4.120 235.300 ;
        RECT 2.520 234.185 2.880 234.565 ;
        RECT 3.130 234.185 3.490 234.565 ;
        RECT 3.760 234.185 4.120 234.565 ;
        RECT 2.520 233.500 2.880 233.880 ;
        RECT 3.130 233.500 3.490 233.880 ;
        RECT 3.760 233.500 4.120 233.880 ;
        RECT 2.520 226.125 2.880 226.505 ;
        RECT 3.130 226.125 3.490 226.505 ;
        RECT 3.760 226.125 4.120 226.505 ;
        RECT 2.520 225.390 2.880 225.770 ;
        RECT 3.130 225.390 3.490 225.770 ;
        RECT 3.760 225.390 4.120 225.770 ;
        RECT 2.520 224.705 2.880 225.085 ;
        RECT 3.130 224.705 3.490 225.085 ;
        RECT 3.760 224.705 4.120 225.085 ;
        RECT 2.515 223.230 2.875 223.610 ;
        RECT 3.145 223.230 3.505 223.610 ;
        RECT 3.745 223.230 4.105 223.610 ;
        RECT 2.515 222.640 2.875 223.020 ;
        RECT 3.145 222.640 3.505 223.020 ;
        RECT 3.745 222.640 4.105 223.020 ;
        RECT 125.340 236.820 125.700 237.200 ;
        RECT 125.970 236.820 126.330 237.200 ;
        RECT 126.570 236.820 126.930 237.200 ;
        RECT 125.340 236.230 125.700 236.610 ;
        RECT 125.970 236.230 126.330 236.610 ;
        RECT 126.570 236.230 126.930 236.610 ;
        RECT 125.340 223.025 125.700 223.405 ;
        RECT 125.970 223.025 126.330 223.405 ;
        RECT 126.570 223.025 126.930 223.405 ;
        RECT 125.340 222.435 125.700 222.815 ;
        RECT 125.970 222.435 126.330 222.815 ;
        RECT 126.570 222.435 126.930 222.815 ;
        RECT 2.515 217.465 2.875 217.845 ;
        RECT 3.145 217.465 3.505 217.845 ;
        RECT 3.745 217.465 4.105 217.845 ;
        RECT 2.515 216.875 2.875 217.255 ;
        RECT 3.145 216.875 3.505 217.255 ;
        RECT 3.745 216.875 4.105 217.255 ;
        RECT 2.520 214.920 2.880 215.300 ;
        RECT 3.130 214.920 3.490 215.300 ;
        RECT 3.760 214.920 4.120 215.300 ;
        RECT 2.520 214.185 2.880 214.565 ;
        RECT 3.130 214.185 3.490 214.565 ;
        RECT 3.760 214.185 4.120 214.565 ;
        RECT 2.520 213.500 2.880 213.880 ;
        RECT 3.130 213.500 3.490 213.880 ;
        RECT 3.760 213.500 4.120 213.880 ;
        RECT 2.520 206.120 2.880 206.500 ;
        RECT 3.130 206.120 3.490 206.500 ;
        RECT 3.760 206.120 4.120 206.500 ;
        RECT 2.520 205.385 2.880 205.765 ;
        RECT 3.130 205.385 3.490 205.765 ;
        RECT 3.760 205.385 4.120 205.765 ;
        RECT 2.520 204.700 2.880 205.080 ;
        RECT 3.130 204.700 3.490 205.080 ;
        RECT 3.760 204.700 4.120 205.080 ;
        RECT 2.515 202.165 2.875 202.545 ;
        RECT 3.145 202.165 3.505 202.545 ;
        RECT 3.745 202.165 4.105 202.545 ;
        RECT 2.515 201.575 2.875 201.955 ;
        RECT 3.145 201.575 3.505 201.955 ;
        RECT 3.745 201.575 4.105 201.955 ;
        RECT 125.340 217.260 125.700 217.640 ;
        RECT 125.970 217.260 126.330 217.640 ;
        RECT 126.570 217.260 126.930 217.640 ;
        RECT 125.340 216.670 125.700 217.050 ;
        RECT 125.970 216.670 126.330 217.050 ;
        RECT 126.570 216.670 126.930 217.050 ;
        RECT 125.340 201.680 125.700 202.060 ;
        RECT 125.970 201.680 126.330 202.060 ;
        RECT 126.570 201.680 126.930 202.060 ;
        RECT 125.340 201.090 125.700 201.470 ;
        RECT 125.970 201.090 126.330 201.470 ;
        RECT 126.570 201.090 126.930 201.470 ;
        RECT 2.395 175.260 2.805 175.650 ;
        RECT 2.965 175.260 3.375 175.650 ;
        RECT 3.535 175.260 3.945 175.650 ;
        RECT 2.395 169.820 2.805 170.210 ;
        RECT 2.965 169.820 3.375 170.210 ;
        RECT 3.535 169.820 3.945 170.210 ;
        RECT 2.395 164.380 2.805 164.770 ;
        RECT 2.965 164.380 3.375 164.770 ;
        RECT 3.535 164.380 3.945 164.770 ;
        RECT 125.305 174.460 125.705 174.860 ;
        RECT 125.930 174.460 126.330 174.860 ;
        RECT 126.555 174.460 126.955 174.860 ;
        RECT 125.300 173.860 125.700 174.260 ;
        RECT 125.925 173.860 126.325 174.260 ;
        RECT 126.550 173.860 126.950 174.260 ;
        RECT 125.345 171.580 125.705 171.960 ;
        RECT 125.955 171.580 126.315 171.960 ;
        RECT 126.585 171.580 126.945 171.960 ;
        RECT 125.345 170.845 125.705 171.225 ;
        RECT 125.955 170.845 126.315 171.225 ;
        RECT 126.585 170.845 126.945 171.225 ;
        RECT 125.345 170.160 125.705 170.540 ;
        RECT 125.955 170.160 126.315 170.540 ;
        RECT 126.585 170.160 126.945 170.540 ;
        RECT 125.345 162.780 125.705 163.160 ;
        RECT 125.955 162.780 126.315 163.160 ;
        RECT 126.585 162.780 126.945 163.160 ;
        RECT 125.345 162.045 125.705 162.425 ;
        RECT 125.955 162.045 126.315 162.425 ;
        RECT 126.585 162.045 126.945 162.425 ;
        RECT 125.345 161.360 125.705 161.740 ;
        RECT 125.955 161.360 126.315 161.740 ;
        RECT 126.585 161.360 126.945 161.740 ;
        RECT 125.300 159.185 125.700 159.585 ;
        RECT 125.925 159.185 126.325 159.585 ;
        RECT 126.550 159.185 126.950 159.585 ;
        RECT 125.295 158.585 125.695 158.985 ;
        RECT 125.920 158.585 126.320 158.985 ;
        RECT 126.545 158.585 126.945 158.985 ;
        RECT 2.515 141.130 2.875 141.510 ;
        RECT 3.145 141.130 3.505 141.510 ;
        RECT 3.745 141.130 4.105 141.510 ;
        RECT 2.515 140.540 2.875 140.920 ;
        RECT 3.145 140.540 3.505 140.920 ;
        RECT 3.745 140.540 4.105 140.920 ;
        RECT 125.340 141.130 125.700 141.510 ;
        RECT 125.970 141.130 126.330 141.510 ;
        RECT 126.570 141.130 126.930 141.510 ;
        RECT 125.340 140.540 125.700 140.920 ;
        RECT 125.970 140.540 126.330 140.920 ;
        RECT 126.570 140.540 126.930 140.920 ;
        RECT 2.515 137.220 2.875 137.600 ;
        RECT 3.145 137.220 3.505 137.600 ;
        RECT 3.745 137.220 4.105 137.600 ;
        RECT 2.515 136.630 2.875 137.010 ;
        RECT 3.145 136.630 3.505 137.010 ;
        RECT 3.745 136.630 4.105 137.010 ;
        RECT 2.520 134.925 2.880 135.305 ;
        RECT 3.130 134.925 3.490 135.305 ;
        RECT 3.760 134.925 4.120 135.305 ;
        RECT 2.520 134.190 2.880 134.570 ;
        RECT 3.130 134.190 3.490 134.570 ;
        RECT 3.760 134.190 4.120 134.570 ;
        RECT 2.520 133.505 2.880 133.885 ;
        RECT 3.130 133.505 3.490 133.885 ;
        RECT 3.760 133.505 4.120 133.885 ;
        RECT 2.520 126.090 2.880 126.470 ;
        RECT 3.130 126.090 3.490 126.470 ;
        RECT 3.760 126.090 4.120 126.470 ;
        RECT 2.520 125.355 2.880 125.735 ;
        RECT 3.130 125.355 3.490 125.735 ;
        RECT 3.760 125.355 4.120 125.735 ;
        RECT 2.520 124.670 2.880 125.050 ;
        RECT 3.130 124.670 3.490 125.050 ;
        RECT 3.760 124.670 4.120 125.050 ;
        RECT 2.515 122.660 2.875 123.040 ;
        RECT 3.145 122.660 3.505 123.040 ;
        RECT 3.745 122.660 4.105 123.040 ;
        RECT 2.515 122.070 2.875 122.450 ;
        RECT 3.145 122.070 3.505 122.450 ;
        RECT 3.745 122.070 4.105 122.450 ;
        RECT 125.340 137.220 125.700 137.600 ;
        RECT 125.970 137.220 126.330 137.600 ;
        RECT 126.570 137.220 126.930 137.600 ;
        RECT 125.340 136.630 125.700 137.010 ;
        RECT 125.970 136.630 126.330 137.010 ;
        RECT 126.570 136.630 126.930 137.010 ;
        RECT 125.340 122.415 125.700 122.795 ;
        RECT 125.970 122.415 126.330 122.795 ;
        RECT 126.570 122.415 126.930 122.795 ;
        RECT 125.340 121.825 125.700 122.205 ;
        RECT 125.970 121.825 126.330 122.205 ;
        RECT 126.570 121.825 126.930 122.205 ;
        RECT 2.515 117.640 2.875 118.020 ;
        RECT 3.145 117.640 3.505 118.020 ;
        RECT 3.745 117.640 4.105 118.020 ;
        RECT 2.515 117.050 2.875 117.430 ;
        RECT 3.145 117.050 3.505 117.430 ;
        RECT 3.745 117.050 4.105 117.430 ;
        RECT 2.520 114.920 2.880 115.300 ;
        RECT 3.130 114.920 3.490 115.300 ;
        RECT 3.760 114.920 4.120 115.300 ;
        RECT 2.520 114.185 2.880 114.565 ;
        RECT 3.130 114.185 3.490 114.565 ;
        RECT 3.760 114.185 4.120 114.565 ;
        RECT 2.520 113.500 2.880 113.880 ;
        RECT 3.130 113.500 3.490 113.880 ;
        RECT 3.760 113.500 4.120 113.880 ;
        RECT 2.520 106.120 2.880 106.500 ;
        RECT 3.130 106.120 3.490 106.500 ;
        RECT 3.760 106.120 4.120 106.500 ;
        RECT 2.520 105.385 2.880 105.765 ;
        RECT 3.130 105.385 3.490 105.765 ;
        RECT 3.760 105.385 4.120 105.765 ;
        RECT 2.520 104.700 2.880 105.080 ;
        RECT 3.130 104.700 3.490 105.080 ;
        RECT 3.760 104.700 4.120 105.080 ;
        RECT 2.515 102.750 2.875 103.130 ;
        RECT 3.145 102.750 3.505 103.130 ;
        RECT 3.745 102.750 4.105 103.130 ;
        RECT 2.515 102.160 2.875 102.540 ;
        RECT 3.145 102.160 3.505 102.540 ;
        RECT 3.745 102.160 4.105 102.540 ;
        RECT 125.340 116.830 125.700 117.210 ;
        RECT 125.970 116.830 126.330 117.210 ;
        RECT 126.570 116.830 126.930 117.210 ;
        RECT 125.340 116.240 125.700 116.620 ;
        RECT 125.970 116.240 126.330 116.620 ;
        RECT 126.570 116.240 126.930 116.620 ;
        RECT 125.340 102.615 125.700 102.995 ;
        RECT 125.970 102.615 126.330 102.995 ;
        RECT 126.570 102.615 126.930 102.995 ;
        RECT 125.340 102.025 125.700 102.405 ;
        RECT 125.970 102.025 126.330 102.405 ;
        RECT 126.570 102.025 126.930 102.405 ;
        RECT 2.515 97.340 2.875 97.720 ;
        RECT 3.145 97.340 3.505 97.720 ;
        RECT 3.745 97.340 4.105 97.720 ;
        RECT 2.515 96.750 2.875 97.130 ;
        RECT 3.145 96.750 3.505 97.130 ;
        RECT 3.745 96.750 4.105 97.130 ;
        RECT 2.520 94.920 2.880 95.300 ;
        RECT 3.130 94.920 3.490 95.300 ;
        RECT 3.760 94.920 4.120 95.300 ;
        RECT 2.520 94.185 2.880 94.565 ;
        RECT 3.130 94.185 3.490 94.565 ;
        RECT 3.760 94.185 4.120 94.565 ;
        RECT 2.520 93.500 2.880 93.880 ;
        RECT 3.130 93.500 3.490 93.880 ;
        RECT 3.760 93.500 4.120 93.880 ;
        RECT 2.520 86.125 2.880 86.505 ;
        RECT 3.130 86.125 3.490 86.505 ;
        RECT 3.760 86.125 4.120 86.505 ;
        RECT 2.520 85.390 2.880 85.770 ;
        RECT 3.130 85.390 3.490 85.770 ;
        RECT 3.760 85.390 4.120 85.770 ;
        RECT 2.520 84.705 2.880 85.085 ;
        RECT 3.130 84.705 3.490 85.085 ;
        RECT 3.760 84.705 4.120 85.085 ;
        RECT 2.515 82.965 2.875 83.345 ;
        RECT 3.145 82.965 3.505 83.345 ;
        RECT 3.745 82.965 4.105 83.345 ;
        RECT 2.515 82.375 2.875 82.755 ;
        RECT 3.145 82.375 3.505 82.755 ;
        RECT 3.745 82.375 4.105 82.755 ;
        RECT 125.340 96.740 125.700 97.120 ;
        RECT 125.970 96.740 126.330 97.120 ;
        RECT 126.570 96.740 126.930 97.120 ;
        RECT 125.340 96.150 125.700 96.530 ;
        RECT 125.970 96.150 126.330 96.530 ;
        RECT 126.570 96.150 126.930 96.530 ;
        RECT 125.340 82.535 125.700 82.915 ;
        RECT 125.970 82.535 126.330 82.915 ;
        RECT 126.570 82.535 126.930 82.915 ;
        RECT 125.340 81.945 125.700 82.325 ;
        RECT 125.970 81.945 126.330 82.325 ;
        RECT 126.570 81.945 126.930 82.325 ;
        RECT 2.515 77.460 2.875 77.840 ;
        RECT 3.145 77.460 3.505 77.840 ;
        RECT 3.745 77.460 4.105 77.840 ;
        RECT 2.515 76.870 2.875 77.250 ;
        RECT 3.145 76.870 3.505 77.250 ;
        RECT 3.745 76.870 4.105 77.250 ;
        RECT 2.520 74.920 2.880 75.300 ;
        RECT 3.130 74.920 3.490 75.300 ;
        RECT 3.760 74.920 4.120 75.300 ;
        RECT 2.520 74.185 2.880 74.565 ;
        RECT 3.130 74.185 3.490 74.565 ;
        RECT 3.760 74.185 4.120 74.565 ;
        RECT 2.520 73.500 2.880 73.880 ;
        RECT 3.130 73.500 3.490 73.880 ;
        RECT 3.760 73.500 4.120 73.880 ;
        RECT 2.520 66.120 2.880 66.500 ;
        RECT 3.130 66.120 3.490 66.500 ;
        RECT 3.760 66.120 4.120 66.500 ;
        RECT 2.520 65.385 2.880 65.765 ;
        RECT 3.130 65.385 3.490 65.765 ;
        RECT 3.760 65.385 4.120 65.765 ;
        RECT 2.520 64.700 2.880 65.080 ;
        RECT 3.130 64.700 3.490 65.080 ;
        RECT 3.760 64.700 4.120 65.080 ;
        RECT 2.515 63.130 2.875 63.510 ;
        RECT 3.145 63.130 3.505 63.510 ;
        RECT 3.745 63.130 4.105 63.510 ;
        RECT 2.515 62.540 2.875 62.920 ;
        RECT 3.145 62.540 3.505 62.920 ;
        RECT 3.745 62.540 4.105 62.920 ;
        RECT 125.340 76.680 125.700 77.060 ;
        RECT 125.970 76.680 126.330 77.060 ;
        RECT 126.570 76.680 126.930 77.060 ;
        RECT 125.340 76.090 125.700 76.470 ;
        RECT 125.970 76.090 126.330 76.470 ;
        RECT 126.570 76.090 126.930 76.470 ;
        RECT 125.340 62.875 125.700 63.255 ;
        RECT 125.970 62.875 126.330 63.255 ;
        RECT 126.570 62.875 126.930 63.255 ;
        RECT 125.340 62.285 125.700 62.665 ;
        RECT 125.970 62.285 126.330 62.665 ;
        RECT 126.570 62.285 126.930 62.665 ;
        RECT 2.515 57.050 2.875 57.430 ;
        RECT 3.145 57.050 3.505 57.430 ;
        RECT 3.745 57.050 4.105 57.430 ;
        RECT 2.515 56.460 2.875 56.840 ;
        RECT 3.145 56.460 3.505 56.840 ;
        RECT 3.745 56.460 4.105 56.840 ;
        RECT 2.520 54.920 2.880 55.300 ;
        RECT 3.130 54.920 3.490 55.300 ;
        RECT 3.760 54.920 4.120 55.300 ;
        RECT 2.520 54.185 2.880 54.565 ;
        RECT 3.130 54.185 3.490 54.565 ;
        RECT 3.760 54.185 4.120 54.565 ;
        RECT 2.520 53.500 2.880 53.880 ;
        RECT 3.130 53.500 3.490 53.880 ;
        RECT 3.760 53.500 4.120 53.880 ;
        RECT 2.520 46.120 2.880 46.500 ;
        RECT 3.130 46.120 3.490 46.500 ;
        RECT 3.760 46.120 4.120 46.500 ;
        RECT 2.520 45.385 2.880 45.765 ;
        RECT 3.130 45.385 3.490 45.765 ;
        RECT 3.760 45.385 4.120 45.765 ;
        RECT 2.520 44.700 2.880 45.080 ;
        RECT 3.130 44.700 3.490 45.080 ;
        RECT 3.760 44.700 4.120 45.080 ;
        RECT 2.515 42.725 2.875 43.105 ;
        RECT 3.145 42.725 3.505 43.105 ;
        RECT 3.745 42.725 4.105 43.105 ;
        RECT 2.515 42.135 2.875 42.515 ;
        RECT 3.145 42.135 3.505 42.515 ;
        RECT 3.745 42.135 4.105 42.515 ;
        RECT 125.340 56.805 125.700 57.185 ;
        RECT 125.970 56.805 126.330 57.185 ;
        RECT 126.570 56.805 126.930 57.185 ;
        RECT 125.340 56.215 125.700 56.595 ;
        RECT 125.970 56.215 126.330 56.595 ;
        RECT 126.570 56.215 126.930 56.595 ;
        RECT 125.340 42.590 125.700 42.970 ;
        RECT 125.970 42.590 126.330 42.970 ;
        RECT 126.570 42.590 126.930 42.970 ;
        RECT 125.340 42.000 125.700 42.380 ;
        RECT 125.970 42.000 126.330 42.380 ;
        RECT 126.570 42.000 126.930 42.380 ;
        RECT 2.515 37.115 2.875 37.495 ;
        RECT 3.145 37.115 3.505 37.495 ;
        RECT 3.745 37.115 4.105 37.495 ;
        RECT 2.515 36.525 2.875 36.905 ;
        RECT 3.145 36.525 3.505 36.905 ;
        RECT 3.745 36.525 4.105 36.905 ;
        RECT 2.520 34.925 2.880 35.305 ;
        RECT 3.130 34.925 3.490 35.305 ;
        RECT 3.760 34.925 4.120 35.305 ;
        RECT 2.520 34.190 2.880 34.570 ;
        RECT 3.130 34.190 3.490 34.570 ;
        RECT 3.760 34.190 4.120 34.570 ;
        RECT 2.520 33.505 2.880 33.885 ;
        RECT 3.130 33.505 3.490 33.885 ;
        RECT 3.760 33.505 4.120 33.885 ;
        RECT 2.520 26.115 2.880 26.495 ;
        RECT 3.130 26.115 3.490 26.495 ;
        RECT 3.760 26.115 4.120 26.495 ;
        RECT 2.520 25.380 2.880 25.760 ;
        RECT 3.130 25.380 3.490 25.760 ;
        RECT 3.760 25.380 4.120 25.760 ;
        RECT 2.520 24.695 2.880 25.075 ;
        RECT 3.130 24.695 3.490 25.075 ;
        RECT 3.760 24.695 4.120 25.075 ;
        RECT 2.515 22.815 2.875 23.195 ;
        RECT 3.145 22.815 3.505 23.195 ;
        RECT 3.745 22.815 4.105 23.195 ;
        RECT 2.515 22.225 2.875 22.605 ;
        RECT 3.145 22.225 3.505 22.605 ;
        RECT 3.745 22.225 4.105 22.605 ;
        RECT 125.340 36.805 125.700 37.185 ;
        RECT 125.970 36.805 126.330 37.185 ;
        RECT 126.570 36.805 126.930 37.185 ;
        RECT 125.340 36.215 125.700 36.595 ;
        RECT 125.970 36.215 126.330 36.595 ;
        RECT 126.570 36.215 126.930 36.595 ;
        RECT 125.340 22.590 125.700 22.970 ;
        RECT 125.970 22.590 126.330 22.970 ;
        RECT 126.570 22.590 126.930 22.970 ;
        RECT 125.340 22.000 125.700 22.380 ;
        RECT 125.970 22.000 126.330 22.380 ;
        RECT 126.570 22.000 126.930 22.380 ;
        RECT 2.515 17.260 2.875 17.640 ;
        RECT 3.145 17.260 3.505 17.640 ;
        RECT 3.745 17.260 4.105 17.640 ;
        RECT 2.515 16.670 2.875 17.050 ;
        RECT 3.145 16.670 3.505 17.050 ;
        RECT 3.745 16.670 4.105 17.050 ;
        RECT 2.520 14.925 2.880 15.305 ;
        RECT 3.130 14.925 3.490 15.305 ;
        RECT 3.760 14.925 4.120 15.305 ;
        RECT 2.520 14.190 2.880 14.570 ;
        RECT 3.130 14.190 3.490 14.570 ;
        RECT 3.760 14.190 4.120 14.570 ;
        RECT 2.520 13.505 2.880 13.885 ;
        RECT 3.130 13.505 3.490 13.885 ;
        RECT 3.760 13.505 4.120 13.885 ;
        RECT 2.520 6.120 2.880 6.500 ;
        RECT 3.130 6.120 3.490 6.500 ;
        RECT 3.760 6.120 4.120 6.500 ;
        RECT 2.520 5.385 2.880 5.765 ;
        RECT 3.130 5.385 3.490 5.765 ;
        RECT 3.760 5.385 4.120 5.765 ;
        RECT 2.520 4.700 2.880 5.080 ;
        RECT 3.130 4.700 3.490 5.080 ;
        RECT 3.760 4.700 4.120 5.080 ;
        RECT 2.515 3.145 2.875 3.525 ;
        RECT 3.145 3.145 3.505 3.525 ;
        RECT 3.745 3.145 4.105 3.525 ;
        RECT 2.515 2.555 2.875 2.935 ;
        RECT 3.145 2.555 3.505 2.935 ;
        RECT 3.745 2.555 4.105 2.935 ;
        RECT 125.340 16.805 125.700 17.185 ;
        RECT 125.970 16.805 126.330 17.185 ;
        RECT 126.570 16.805 126.930 17.185 ;
        RECT 125.340 16.215 125.700 16.595 ;
        RECT 125.970 16.215 126.330 16.595 ;
        RECT 126.570 16.215 126.930 16.595 ;
        RECT 125.340 2.590 125.700 2.970 ;
        RECT 125.970 2.590 126.330 2.970 ;
        RECT 126.570 2.590 126.930 2.970 ;
        RECT 125.340 2.000 125.700 2.380 ;
        RECT 125.970 2.000 126.330 2.380 ;
        RECT 126.570 2.000 126.930 2.380 ;
      LAYER met3 ;
        RECT 2.315 336.110 4.320 337.385 ;
        RECT 125.130 336.310 127.130 337.585 ;
        RECT 2.315 333.250 4.315 335.545 ;
        RECT 2.315 324.450 4.315 326.745 ;
        RECT 2.315 322.745 4.320 324.020 ;
        RECT 125.140 322.325 127.140 323.600 ;
        RECT 2.315 316.100 4.320 317.375 ;
        RECT 125.130 316.310 127.130 317.585 ;
        RECT 2.315 313.250 4.315 315.545 ;
        RECT 2.315 304.455 4.315 306.750 ;
        RECT 2.315 302.400 4.320 303.675 ;
        RECT 125.140 302.325 127.140 303.600 ;
        RECT 2.315 296.510 4.320 297.785 ;
        RECT 125.130 296.310 127.130 297.585 ;
        RECT 2.320 295.340 4.320 295.545 ;
        RECT 2.315 293.250 4.320 295.340 ;
        RECT 2.315 284.455 4.315 286.750 ;
        RECT 2.315 282.270 4.330 283.545 ;
        RECT 125.140 282.325 127.140 283.600 ;
        RECT 2.315 276.255 4.320 277.530 ;
        RECT 125.135 276.580 127.135 277.855 ;
        RECT 2.320 275.340 4.320 275.545 ;
        RECT 2.315 273.250 4.320 275.340 ;
        RECT 2.315 264.445 4.315 266.740 ;
        RECT 2.315 262.370 4.320 263.645 ;
        RECT 125.140 262.000 127.140 263.275 ;
        RECT 2.315 256.335 4.330 257.610 ;
        RECT 125.135 256.085 127.135 257.360 ;
        RECT 2.315 253.250 4.315 255.545 ;
        RECT 2.315 244.455 4.315 246.750 ;
        RECT 2.315 242.505 4.320 243.780 ;
        RECT 125.140 241.725 127.140 243.000 ;
        RECT 2.315 236.570 4.320 237.845 ;
        RECT 125.140 236.050 127.140 237.325 ;
        RECT 2.315 233.250 4.315 235.545 ;
        RECT 2.315 224.455 4.315 226.750 ;
        RECT 2.315 222.460 4.320 223.735 ;
        RECT 125.140 222.255 127.140 223.530 ;
        RECT 2.315 216.695 4.320 217.970 ;
        RECT 125.140 216.490 127.140 217.765 ;
        RECT 2.315 213.250 4.315 215.545 ;
        RECT 2.315 204.455 4.315 206.750 ;
        RECT 2.315 204.450 4.180 204.455 ;
        RECT 2.315 201.395 4.315 202.670 ;
        RECT 125.140 200.910 127.140 202.185 ;
        RECT 2.315 175.215 4.025 175.695 ;
        RECT 42.635 175.410 47.035 176.660 ;
        RECT 58.235 175.410 67.035 176.660 ;
        RECT 78.235 175.410 87.035 176.660 ;
        RECT 98.235 175.410 107.035 176.660 ;
        RECT 118.235 175.410 122.635 176.660 ;
        RECT 42.635 172.260 122.635 175.410 ;
        RECT 125.140 173.715 127.140 174.990 ;
        RECT 2.315 169.775 4.025 170.255 ;
        RECT 2.315 164.335 4.025 164.815 ;
        RECT 43.885 161.060 61.385 172.260 ;
        RECT 63.885 161.060 81.385 172.260 ;
        RECT 83.885 161.060 101.385 172.260 ;
        RECT 103.885 161.060 121.385 172.260 ;
        RECT 125.140 169.915 127.140 172.210 ;
        RECT 125.140 169.910 127.005 169.915 ;
        RECT 125.140 161.115 127.140 163.410 ;
        RECT 125.140 161.110 127.005 161.115 ;
        RECT 42.635 157.910 122.635 161.060 ;
        RECT 125.135 158.440 127.135 159.715 ;
        RECT 42.635 156.660 47.035 157.910 ;
        RECT 58.235 156.660 67.035 157.910 ;
        RECT 78.235 156.660 87.035 157.910 ;
        RECT 98.235 156.660 107.035 157.910 ;
        RECT 118.235 156.660 122.635 157.910 ;
        RECT 2.315 140.360 4.330 141.800 ;
        RECT 125.125 140.360 127.140 141.800 ;
        RECT 4.730 138.750 9.130 140.000 ;
        RECT 20.330 138.750 29.130 140.000 ;
        RECT 40.330 138.750 49.130 140.000 ;
        RECT 60.330 138.750 69.130 140.000 ;
        RECT 80.330 138.750 89.130 140.000 ;
        RECT 100.330 138.750 109.130 140.000 ;
        RECT 120.330 138.750 124.730 140.000 ;
        RECT 2.315 136.450 4.315 137.725 ;
        RECT 4.730 135.600 124.730 138.750 ;
        RECT 125.140 136.450 127.140 137.725 ;
        RECT 2.315 133.255 4.315 135.555 ;
        RECT 2.315 124.425 4.315 126.745 ;
        RECT 2.315 124.420 4.310 124.425 ;
        RECT 5.980 124.400 23.480 135.600 ;
        RECT 25.980 124.400 43.480 135.600 ;
        RECT 45.980 124.400 63.480 135.600 ;
        RECT 65.980 124.400 83.480 135.600 ;
        RECT 85.980 124.400 103.480 135.600 ;
        RECT 105.980 124.400 123.480 135.600 ;
        RECT 2.315 121.890 4.315 123.165 ;
        RECT 4.730 121.250 124.730 124.400 ;
        RECT 125.140 121.645 127.140 122.920 ;
        RECT 4.730 118.750 9.130 121.250 ;
        RECT 20.330 118.750 29.130 121.250 ;
        RECT 40.330 118.750 49.130 121.250 ;
        RECT 60.330 118.750 69.130 121.250 ;
        RECT 80.330 118.750 89.130 121.250 ;
        RECT 100.330 118.750 109.130 121.250 ;
        RECT 120.330 118.750 124.730 121.250 ;
        RECT 2.315 116.870 4.315 118.145 ;
        RECT 4.730 115.600 124.730 118.750 ;
        RECT 125.135 116.060 127.135 117.335 ;
        RECT 2.315 113.250 4.315 115.545 ;
        RECT 2.315 104.450 4.315 106.745 ;
        RECT 5.980 104.400 23.480 115.600 ;
        RECT 25.980 104.400 43.480 115.600 ;
        RECT 45.980 104.400 63.480 115.600 ;
        RECT 65.980 104.400 83.480 115.600 ;
        RECT 85.980 104.400 103.480 115.600 ;
        RECT 105.980 104.400 123.480 115.600 ;
        RECT 2.315 101.980 4.320 103.255 ;
        RECT 4.730 101.250 124.730 104.400 ;
        RECT 125.140 101.845 127.140 103.120 ;
        RECT 4.730 98.750 9.130 101.250 ;
        RECT 20.330 98.750 29.130 101.250 ;
        RECT 40.330 98.750 49.130 101.250 ;
        RECT 60.330 98.750 69.130 101.250 ;
        RECT 80.330 98.750 89.130 101.250 ;
        RECT 100.330 98.750 109.130 101.250 ;
        RECT 120.330 98.750 124.730 101.250 ;
        RECT 2.315 96.570 4.320 97.845 ;
        RECT 4.730 95.600 124.730 98.750 ;
        RECT 125.140 95.970 127.140 97.245 ;
        RECT 2.315 93.250 4.315 95.545 ;
        RECT 2.315 84.455 4.315 86.750 ;
        RECT 5.980 84.400 23.480 95.600 ;
        RECT 25.980 84.400 43.480 95.600 ;
        RECT 45.980 84.400 63.480 95.600 ;
        RECT 65.980 84.400 83.480 95.600 ;
        RECT 85.980 84.400 103.480 95.600 ;
        RECT 105.980 84.400 123.480 95.600 ;
        RECT 2.315 82.195 4.320 83.470 ;
        RECT 4.730 81.250 124.730 84.400 ;
        RECT 125.135 81.765 127.135 83.040 ;
        RECT 4.730 78.750 9.130 81.250 ;
        RECT 20.330 78.750 29.130 81.250 ;
        RECT 40.330 78.750 49.130 81.250 ;
        RECT 60.330 78.750 69.130 81.250 ;
        RECT 80.330 78.750 89.130 81.250 ;
        RECT 100.330 78.750 109.130 81.250 ;
        RECT 120.330 78.750 124.730 81.250 ;
        RECT 2.315 76.690 4.320 77.965 ;
        RECT 4.730 75.600 124.730 78.750 ;
        RECT 125.135 75.910 127.135 77.185 ;
        RECT 2.315 73.250 4.315 75.545 ;
        RECT 2.315 64.450 4.315 66.745 ;
        RECT 5.980 64.400 23.480 75.600 ;
        RECT 25.980 64.400 43.480 75.600 ;
        RECT 45.980 64.400 63.480 75.600 ;
        RECT 65.980 64.400 83.480 75.600 ;
        RECT 85.980 64.400 103.480 75.600 ;
        RECT 105.980 64.400 123.480 75.600 ;
        RECT 2.315 62.360 4.325 63.635 ;
        RECT 4.730 61.250 124.730 64.400 ;
        RECT 125.135 62.105 127.135 63.380 ;
        RECT 4.730 58.750 9.130 61.250 ;
        RECT 20.330 58.750 29.130 61.250 ;
        RECT 40.330 58.750 49.130 61.250 ;
        RECT 60.330 58.750 69.130 61.250 ;
        RECT 80.330 58.750 89.130 61.250 ;
        RECT 100.330 58.750 109.130 61.250 ;
        RECT 120.330 58.750 124.730 61.250 ;
        RECT 2.315 56.280 4.330 57.555 ;
        RECT 4.730 55.600 124.730 58.750 ;
        RECT 125.135 56.035 127.135 57.310 ;
        RECT 2.315 53.250 4.315 55.545 ;
        RECT 2.315 44.450 4.315 46.745 ;
        RECT 5.980 44.400 23.480 55.600 ;
        RECT 25.980 44.400 43.480 55.600 ;
        RECT 45.980 44.400 63.480 55.600 ;
        RECT 65.980 44.400 83.480 55.600 ;
        RECT 85.980 44.400 103.480 55.600 ;
        RECT 105.980 44.400 123.480 55.600 ;
        RECT 2.315 41.955 4.320 43.230 ;
        RECT 4.730 41.250 124.730 44.400 ;
        RECT 125.140 41.820 127.140 43.095 ;
        RECT 4.730 38.750 9.130 41.250 ;
        RECT 20.330 38.750 29.130 41.250 ;
        RECT 40.330 38.750 49.130 41.250 ;
        RECT 60.330 38.750 69.130 41.250 ;
        RECT 80.330 38.750 89.130 41.250 ;
        RECT 100.330 38.750 109.130 41.250 ;
        RECT 120.330 38.750 124.730 41.250 ;
        RECT 2.315 36.345 4.320 37.620 ;
        RECT 4.730 35.600 124.730 38.750 ;
        RECT 125.135 36.035 127.135 37.310 ;
        RECT 2.315 33.255 4.315 35.550 ;
        RECT 2.315 24.445 4.315 26.740 ;
        RECT 5.980 24.400 23.480 35.600 ;
        RECT 25.980 24.400 43.480 35.600 ;
        RECT 45.980 24.400 63.480 35.600 ;
        RECT 65.980 24.400 83.480 35.600 ;
        RECT 85.980 24.400 103.480 35.600 ;
        RECT 105.980 24.400 123.480 35.600 ;
        RECT 2.315 22.045 4.315 23.320 ;
        RECT 4.730 21.250 124.730 24.400 ;
        RECT 125.140 21.820 127.140 23.095 ;
        RECT 4.730 18.750 9.130 21.250 ;
        RECT 20.330 18.750 29.130 21.250 ;
        RECT 40.330 18.750 49.130 21.250 ;
        RECT 60.330 18.750 69.130 21.250 ;
        RECT 80.330 18.750 89.130 21.250 ;
        RECT 100.330 18.750 109.130 21.250 ;
        RECT 120.330 18.750 124.730 21.250 ;
        RECT 2.315 16.490 4.315 17.765 ;
        RECT 4.730 15.600 124.730 18.750 ;
        RECT 125.135 16.035 127.135 17.310 ;
        RECT 2.315 13.255 4.315 15.550 ;
        RECT 2.315 4.450 4.315 6.745 ;
        RECT 5.980 4.400 23.480 15.600 ;
        RECT 25.980 4.400 43.480 15.600 ;
        RECT 45.980 4.400 63.480 15.600 ;
        RECT 65.980 4.400 83.480 15.600 ;
        RECT 85.980 4.400 103.480 15.600 ;
        RECT 105.980 4.400 123.480 15.600 ;
        RECT 2.315 2.375 4.325 3.650 ;
        RECT 4.730 1.250 124.730 4.400 ;
        RECT 125.140 1.820 127.140 3.095 ;
        RECT 4.730 0.000 9.130 1.250 ;
        RECT 20.330 0.000 29.130 1.250 ;
        RECT 40.330 0.000 49.130 1.250 ;
        RECT 60.330 0.000 69.130 1.250 ;
        RECT 80.330 0.000 89.130 1.250 ;
        RECT 100.330 0.000 109.130 1.250 ;
        RECT 120.330 0.000 124.730 1.250 ;
      LAYER via3 ;
        RECT 2.515 336.880 2.875 337.260 ;
        RECT 3.145 336.880 3.505 337.260 ;
        RECT 3.745 336.880 4.105 337.260 ;
        RECT 2.515 336.290 2.875 336.670 ;
        RECT 3.145 336.290 3.505 336.670 ;
        RECT 3.745 336.290 4.105 336.670 ;
        RECT 125.340 337.080 125.700 337.460 ;
        RECT 125.970 337.080 126.330 337.460 ;
        RECT 126.570 337.080 126.930 337.460 ;
        RECT 125.340 336.490 125.700 336.870 ;
        RECT 125.970 336.490 126.330 336.870 ;
        RECT 126.570 336.490 126.930 336.870 ;
        RECT 2.520 334.920 2.880 335.300 ;
        RECT 3.130 334.920 3.490 335.300 ;
        RECT 3.760 334.920 4.120 335.300 ;
        RECT 2.520 334.185 2.880 334.565 ;
        RECT 3.130 334.185 3.490 334.565 ;
        RECT 3.760 334.185 4.120 334.565 ;
        RECT 2.520 333.500 2.880 333.880 ;
        RECT 3.130 333.500 3.490 333.880 ;
        RECT 3.760 333.500 4.120 333.880 ;
        RECT 2.520 326.120 2.880 326.500 ;
        RECT 3.130 326.120 3.490 326.500 ;
        RECT 3.760 326.120 4.120 326.500 ;
        RECT 2.520 325.385 2.880 325.765 ;
        RECT 3.130 325.385 3.490 325.765 ;
        RECT 3.760 325.385 4.120 325.765 ;
        RECT 2.520 324.700 2.880 325.080 ;
        RECT 3.130 324.700 3.490 325.080 ;
        RECT 3.760 324.700 4.120 325.080 ;
        RECT 2.515 323.515 2.875 323.895 ;
        RECT 3.145 323.515 3.505 323.895 ;
        RECT 3.745 323.515 4.105 323.895 ;
        RECT 2.515 322.925 2.875 323.305 ;
        RECT 3.145 322.925 3.505 323.305 ;
        RECT 3.745 322.925 4.105 323.305 ;
        RECT 125.340 323.095 125.700 323.475 ;
        RECT 125.970 323.095 126.330 323.475 ;
        RECT 126.570 323.095 126.930 323.475 ;
        RECT 125.340 322.505 125.700 322.885 ;
        RECT 125.970 322.505 126.330 322.885 ;
        RECT 126.570 322.505 126.930 322.885 ;
        RECT 2.515 316.870 2.875 317.250 ;
        RECT 3.145 316.870 3.505 317.250 ;
        RECT 3.745 316.870 4.105 317.250 ;
        RECT 2.515 316.280 2.875 316.660 ;
        RECT 3.145 316.280 3.505 316.660 ;
        RECT 3.745 316.280 4.105 316.660 ;
        RECT 125.340 317.080 125.700 317.460 ;
        RECT 125.970 317.080 126.330 317.460 ;
        RECT 126.570 317.080 126.930 317.460 ;
        RECT 125.340 316.490 125.700 316.870 ;
        RECT 125.970 316.490 126.330 316.870 ;
        RECT 126.570 316.490 126.930 316.870 ;
        RECT 2.520 314.920 2.880 315.300 ;
        RECT 3.130 314.920 3.490 315.300 ;
        RECT 3.760 314.920 4.120 315.300 ;
        RECT 2.520 314.185 2.880 314.565 ;
        RECT 3.130 314.185 3.490 314.565 ;
        RECT 3.760 314.185 4.120 314.565 ;
        RECT 2.520 313.500 2.880 313.880 ;
        RECT 3.130 313.500 3.490 313.880 ;
        RECT 3.760 313.500 4.120 313.880 ;
        RECT 2.520 306.125 2.880 306.505 ;
        RECT 3.130 306.125 3.490 306.505 ;
        RECT 3.760 306.125 4.120 306.505 ;
        RECT 2.520 305.390 2.880 305.770 ;
        RECT 3.130 305.390 3.490 305.770 ;
        RECT 3.760 305.390 4.120 305.770 ;
        RECT 2.520 304.705 2.880 305.085 ;
        RECT 3.130 304.705 3.490 305.085 ;
        RECT 3.760 304.705 4.120 305.085 ;
        RECT 2.515 303.170 2.875 303.550 ;
        RECT 3.145 303.170 3.505 303.550 ;
        RECT 3.745 303.170 4.105 303.550 ;
        RECT 2.515 302.580 2.875 302.960 ;
        RECT 3.145 302.580 3.505 302.960 ;
        RECT 3.745 302.580 4.105 302.960 ;
        RECT 125.340 303.095 125.700 303.475 ;
        RECT 125.970 303.095 126.330 303.475 ;
        RECT 126.570 303.095 126.930 303.475 ;
        RECT 125.340 302.505 125.700 302.885 ;
        RECT 125.970 302.505 126.330 302.885 ;
        RECT 126.570 302.505 126.930 302.885 ;
        RECT 2.515 297.280 2.875 297.660 ;
        RECT 3.145 297.280 3.505 297.660 ;
        RECT 3.745 297.280 4.105 297.660 ;
        RECT 2.515 296.690 2.875 297.070 ;
        RECT 3.145 296.690 3.505 297.070 ;
        RECT 3.745 296.690 4.105 297.070 ;
        RECT 125.340 297.080 125.700 297.460 ;
        RECT 125.970 297.080 126.330 297.460 ;
        RECT 126.570 297.080 126.930 297.460 ;
        RECT 125.340 296.490 125.700 296.870 ;
        RECT 125.970 296.490 126.330 296.870 ;
        RECT 126.570 296.490 126.930 296.870 ;
        RECT 2.520 294.920 2.880 295.300 ;
        RECT 3.130 294.920 3.490 295.300 ;
        RECT 3.760 294.920 4.120 295.300 ;
        RECT 2.520 294.185 2.880 294.565 ;
        RECT 3.130 294.185 3.490 294.565 ;
        RECT 3.760 294.185 4.120 294.565 ;
        RECT 2.520 293.500 2.880 293.880 ;
        RECT 3.130 293.500 3.490 293.880 ;
        RECT 3.760 293.500 4.120 293.880 ;
        RECT 2.520 286.125 2.880 286.505 ;
        RECT 3.130 286.125 3.490 286.505 ;
        RECT 3.760 286.125 4.120 286.505 ;
        RECT 2.520 285.390 2.880 285.770 ;
        RECT 3.130 285.390 3.490 285.770 ;
        RECT 3.760 285.390 4.120 285.770 ;
        RECT 2.520 284.705 2.880 285.085 ;
        RECT 3.130 284.705 3.490 285.085 ;
        RECT 3.760 284.705 4.120 285.085 ;
        RECT 2.515 283.040 2.875 283.420 ;
        RECT 3.145 283.040 3.505 283.420 ;
        RECT 3.745 283.040 4.105 283.420 ;
        RECT 2.515 282.450 2.875 282.830 ;
        RECT 3.145 282.450 3.505 282.830 ;
        RECT 3.745 282.450 4.105 282.830 ;
        RECT 125.340 283.095 125.700 283.475 ;
        RECT 125.970 283.095 126.330 283.475 ;
        RECT 126.570 283.095 126.930 283.475 ;
        RECT 125.340 282.505 125.700 282.885 ;
        RECT 125.970 282.505 126.330 282.885 ;
        RECT 126.570 282.505 126.930 282.885 ;
        RECT 2.515 277.025 2.875 277.405 ;
        RECT 3.145 277.025 3.505 277.405 ;
        RECT 3.745 277.025 4.105 277.405 ;
        RECT 2.515 276.435 2.875 276.815 ;
        RECT 3.145 276.435 3.505 276.815 ;
        RECT 3.745 276.435 4.105 276.815 ;
        RECT 125.340 277.350 125.700 277.730 ;
        RECT 125.970 277.350 126.330 277.730 ;
        RECT 126.570 277.350 126.930 277.730 ;
        RECT 125.340 276.760 125.700 277.140 ;
        RECT 125.970 276.760 126.330 277.140 ;
        RECT 126.570 276.760 126.930 277.140 ;
        RECT 2.520 274.920 2.880 275.300 ;
        RECT 3.130 274.920 3.490 275.300 ;
        RECT 3.760 274.920 4.120 275.300 ;
        RECT 2.520 274.185 2.880 274.565 ;
        RECT 3.130 274.185 3.490 274.565 ;
        RECT 3.760 274.185 4.120 274.565 ;
        RECT 2.520 273.500 2.880 273.880 ;
        RECT 3.130 273.500 3.490 273.880 ;
        RECT 3.760 273.500 4.120 273.880 ;
        RECT 2.520 266.115 2.880 266.495 ;
        RECT 3.130 266.115 3.490 266.495 ;
        RECT 3.760 266.115 4.120 266.495 ;
        RECT 2.520 265.380 2.880 265.760 ;
        RECT 3.130 265.380 3.490 265.760 ;
        RECT 3.760 265.380 4.120 265.760 ;
        RECT 2.520 264.695 2.880 265.075 ;
        RECT 3.130 264.695 3.490 265.075 ;
        RECT 3.760 264.695 4.120 265.075 ;
        RECT 2.515 263.140 2.875 263.520 ;
        RECT 3.145 263.140 3.505 263.520 ;
        RECT 3.745 263.140 4.105 263.520 ;
        RECT 2.515 262.550 2.875 262.930 ;
        RECT 3.145 262.550 3.505 262.930 ;
        RECT 3.745 262.550 4.105 262.930 ;
        RECT 125.340 262.770 125.700 263.150 ;
        RECT 125.970 262.770 126.330 263.150 ;
        RECT 126.570 262.770 126.930 263.150 ;
        RECT 125.340 262.180 125.700 262.560 ;
        RECT 125.970 262.180 126.330 262.560 ;
        RECT 126.570 262.180 126.930 262.560 ;
        RECT 2.515 257.105 2.875 257.485 ;
        RECT 3.145 257.105 3.505 257.485 ;
        RECT 3.745 257.105 4.105 257.485 ;
        RECT 2.515 256.515 2.875 256.895 ;
        RECT 3.145 256.515 3.505 256.895 ;
        RECT 3.745 256.515 4.105 256.895 ;
        RECT 125.340 256.855 125.700 257.235 ;
        RECT 125.970 256.855 126.330 257.235 ;
        RECT 126.570 256.855 126.930 257.235 ;
        RECT 125.340 256.265 125.700 256.645 ;
        RECT 125.970 256.265 126.330 256.645 ;
        RECT 126.570 256.265 126.930 256.645 ;
        RECT 2.520 254.920 2.880 255.300 ;
        RECT 3.130 254.920 3.490 255.300 ;
        RECT 3.760 254.920 4.120 255.300 ;
        RECT 2.520 254.185 2.880 254.565 ;
        RECT 3.130 254.185 3.490 254.565 ;
        RECT 3.760 254.185 4.120 254.565 ;
        RECT 2.520 253.500 2.880 253.880 ;
        RECT 3.130 253.500 3.490 253.880 ;
        RECT 3.760 253.500 4.120 253.880 ;
        RECT 2.520 246.125 2.880 246.505 ;
        RECT 3.130 246.125 3.490 246.505 ;
        RECT 3.760 246.125 4.120 246.505 ;
        RECT 2.520 245.390 2.880 245.770 ;
        RECT 3.130 245.390 3.490 245.770 ;
        RECT 3.760 245.390 4.120 245.770 ;
        RECT 2.520 244.705 2.880 245.085 ;
        RECT 3.130 244.705 3.490 245.085 ;
        RECT 3.760 244.705 4.120 245.085 ;
        RECT 2.515 243.275 2.875 243.655 ;
        RECT 3.145 243.275 3.505 243.655 ;
        RECT 3.745 243.275 4.105 243.655 ;
        RECT 2.515 242.685 2.875 243.065 ;
        RECT 3.145 242.685 3.505 243.065 ;
        RECT 3.745 242.685 4.105 243.065 ;
        RECT 125.340 242.495 125.700 242.875 ;
        RECT 125.970 242.495 126.330 242.875 ;
        RECT 126.570 242.495 126.930 242.875 ;
        RECT 125.340 241.905 125.700 242.285 ;
        RECT 125.970 241.905 126.330 242.285 ;
        RECT 126.570 241.905 126.930 242.285 ;
        RECT 2.515 237.340 2.875 237.720 ;
        RECT 3.145 237.340 3.505 237.720 ;
        RECT 3.745 237.340 4.105 237.720 ;
        RECT 2.515 236.750 2.875 237.130 ;
        RECT 3.145 236.750 3.505 237.130 ;
        RECT 3.745 236.750 4.105 237.130 ;
        RECT 125.340 236.820 125.700 237.200 ;
        RECT 125.970 236.820 126.330 237.200 ;
        RECT 126.570 236.820 126.930 237.200 ;
        RECT 125.340 236.230 125.700 236.610 ;
        RECT 125.970 236.230 126.330 236.610 ;
        RECT 126.570 236.230 126.930 236.610 ;
        RECT 2.520 234.920 2.880 235.300 ;
        RECT 3.130 234.920 3.490 235.300 ;
        RECT 3.760 234.920 4.120 235.300 ;
        RECT 2.520 234.185 2.880 234.565 ;
        RECT 3.130 234.185 3.490 234.565 ;
        RECT 3.760 234.185 4.120 234.565 ;
        RECT 2.520 233.500 2.880 233.880 ;
        RECT 3.130 233.500 3.490 233.880 ;
        RECT 3.760 233.500 4.120 233.880 ;
        RECT 2.520 226.125 2.880 226.505 ;
        RECT 3.130 226.125 3.490 226.505 ;
        RECT 3.760 226.125 4.120 226.505 ;
        RECT 2.520 225.390 2.880 225.770 ;
        RECT 3.130 225.390 3.490 225.770 ;
        RECT 3.760 225.390 4.120 225.770 ;
        RECT 2.520 224.705 2.880 225.085 ;
        RECT 3.130 224.705 3.490 225.085 ;
        RECT 3.760 224.705 4.120 225.085 ;
        RECT 2.515 223.230 2.875 223.610 ;
        RECT 3.145 223.230 3.505 223.610 ;
        RECT 3.745 223.230 4.105 223.610 ;
        RECT 2.515 222.640 2.875 223.020 ;
        RECT 3.145 222.640 3.505 223.020 ;
        RECT 3.745 222.640 4.105 223.020 ;
        RECT 125.340 223.025 125.700 223.405 ;
        RECT 125.970 223.025 126.330 223.405 ;
        RECT 126.570 223.025 126.930 223.405 ;
        RECT 125.340 222.435 125.700 222.815 ;
        RECT 125.970 222.435 126.330 222.815 ;
        RECT 126.570 222.435 126.930 222.815 ;
        RECT 2.515 217.465 2.875 217.845 ;
        RECT 3.145 217.465 3.505 217.845 ;
        RECT 3.745 217.465 4.105 217.845 ;
        RECT 2.515 216.875 2.875 217.255 ;
        RECT 3.145 216.875 3.505 217.255 ;
        RECT 3.745 216.875 4.105 217.255 ;
        RECT 125.340 217.260 125.700 217.640 ;
        RECT 125.970 217.260 126.330 217.640 ;
        RECT 126.570 217.260 126.930 217.640 ;
        RECT 125.340 216.670 125.700 217.050 ;
        RECT 125.970 216.670 126.330 217.050 ;
        RECT 126.570 216.670 126.930 217.050 ;
        RECT 2.520 214.920 2.880 215.300 ;
        RECT 3.130 214.920 3.490 215.300 ;
        RECT 3.760 214.920 4.120 215.300 ;
        RECT 2.520 214.185 2.880 214.565 ;
        RECT 3.130 214.185 3.490 214.565 ;
        RECT 3.760 214.185 4.120 214.565 ;
        RECT 2.520 213.500 2.880 213.880 ;
        RECT 3.130 213.500 3.490 213.880 ;
        RECT 3.760 213.500 4.120 213.880 ;
        RECT 2.520 206.120 2.880 206.500 ;
        RECT 3.130 206.120 3.490 206.500 ;
        RECT 3.760 206.120 4.120 206.500 ;
        RECT 2.520 205.385 2.880 205.765 ;
        RECT 3.130 205.385 3.490 205.765 ;
        RECT 3.760 205.385 4.120 205.765 ;
        RECT 2.520 204.700 2.880 205.080 ;
        RECT 3.130 204.700 3.490 205.080 ;
        RECT 3.760 204.700 4.120 205.080 ;
        RECT 2.515 202.165 2.875 202.545 ;
        RECT 3.145 202.165 3.505 202.545 ;
        RECT 3.745 202.165 4.105 202.545 ;
        RECT 2.515 201.575 2.875 201.955 ;
        RECT 3.145 201.575 3.505 201.955 ;
        RECT 3.745 201.575 4.105 201.955 ;
        RECT 125.340 201.680 125.700 202.060 ;
        RECT 125.970 201.680 126.330 202.060 ;
        RECT 126.570 201.680 126.930 202.060 ;
        RECT 125.340 201.090 125.700 201.470 ;
        RECT 125.970 201.090 126.330 201.470 ;
        RECT 126.570 201.090 126.930 201.470 ;
        RECT 42.735 175.710 43.585 176.560 ;
        RECT 43.685 175.710 44.535 176.560 ;
        RECT 45.135 175.710 45.985 176.560 ;
        RECT 46.085 175.710 46.935 176.560 ;
        RECT 2.390 175.255 2.810 175.655 ;
        RECT 2.960 175.255 3.380 175.655 ;
        RECT 3.530 175.255 3.950 175.655 ;
        RECT 42.735 174.760 43.585 175.610 ;
        RECT 58.335 175.710 59.185 176.560 ;
        RECT 59.285 175.710 60.135 176.560 ;
        RECT 60.735 175.710 61.585 176.560 ;
        RECT 61.685 175.710 62.535 176.560 ;
        RECT 62.735 175.710 63.585 176.560 ;
        RECT 63.685 175.710 64.535 176.560 ;
        RECT 65.135 175.710 65.985 176.560 ;
        RECT 66.085 175.710 66.935 176.560 ;
        RECT 61.685 174.760 62.535 175.610 ;
        RECT 62.735 174.760 63.585 175.610 ;
        RECT 78.335 175.710 79.185 176.560 ;
        RECT 79.285 175.710 80.135 176.560 ;
        RECT 80.735 175.710 81.585 176.560 ;
        RECT 81.685 175.710 82.535 176.560 ;
        RECT 82.735 175.710 83.585 176.560 ;
        RECT 83.685 175.710 84.535 176.560 ;
        RECT 85.135 175.710 85.985 176.560 ;
        RECT 86.085 175.710 86.935 176.560 ;
        RECT 81.685 174.760 82.535 175.610 ;
        RECT 82.735 174.760 83.585 175.610 ;
        RECT 98.335 175.710 99.185 176.560 ;
        RECT 99.285 175.710 100.135 176.560 ;
        RECT 100.735 175.710 101.585 176.560 ;
        RECT 101.685 175.710 102.535 176.560 ;
        RECT 102.735 175.710 103.585 176.560 ;
        RECT 103.685 175.710 104.535 176.560 ;
        RECT 105.135 175.710 105.985 176.560 ;
        RECT 106.085 175.710 106.935 176.560 ;
        RECT 101.685 174.760 102.535 175.610 ;
        RECT 102.735 174.760 103.585 175.610 ;
        RECT 118.335 175.710 119.185 176.560 ;
        RECT 119.285 175.710 120.135 176.560 ;
        RECT 120.735 175.710 121.585 176.560 ;
        RECT 121.685 175.710 122.535 176.560 ;
        RECT 121.685 174.760 122.535 175.610 ;
        RECT 42.735 173.310 43.585 174.160 ;
        RECT 61.685 173.310 62.535 174.160 ;
        RECT 62.735 173.310 63.585 174.160 ;
        RECT 81.685 173.310 82.535 174.160 ;
        RECT 82.735 173.310 83.585 174.160 ;
        RECT 101.685 173.310 102.535 174.160 ;
        RECT 102.735 173.310 103.585 174.160 ;
        RECT 121.685 173.310 122.535 174.160 ;
        RECT 125.305 174.460 125.705 174.860 ;
        RECT 125.930 174.460 126.330 174.860 ;
        RECT 126.555 174.460 126.955 174.860 ;
        RECT 125.300 173.860 125.700 174.260 ;
        RECT 125.925 173.860 126.325 174.260 ;
        RECT 126.550 173.860 126.950 174.260 ;
        RECT 42.735 172.360 43.585 173.210 ;
        RECT 61.685 172.360 62.535 173.210 ;
        RECT 62.735 172.360 63.585 173.210 ;
        RECT 81.685 172.360 82.535 173.210 ;
        RECT 82.735 172.360 83.585 173.210 ;
        RECT 101.685 172.360 102.535 173.210 ;
        RECT 102.735 172.360 103.585 173.210 ;
        RECT 121.685 172.360 122.535 173.210 ;
        RECT 2.390 169.815 2.810 170.215 ;
        RECT 2.960 169.815 3.380 170.215 ;
        RECT 3.530 169.815 3.950 170.215 ;
        RECT 2.390 164.375 2.810 164.775 ;
        RECT 2.960 164.375 3.380 164.775 ;
        RECT 3.530 164.375 3.950 164.775 ;
        RECT 125.345 171.580 125.705 171.960 ;
        RECT 125.955 171.580 126.315 171.960 ;
        RECT 126.585 171.580 126.945 171.960 ;
        RECT 125.345 170.845 125.705 171.225 ;
        RECT 125.955 170.845 126.315 171.225 ;
        RECT 126.585 170.845 126.945 171.225 ;
        RECT 125.345 170.160 125.705 170.540 ;
        RECT 125.955 170.160 126.315 170.540 ;
        RECT 126.585 170.160 126.945 170.540 ;
        RECT 125.345 162.780 125.705 163.160 ;
        RECT 125.955 162.780 126.315 163.160 ;
        RECT 126.585 162.780 126.945 163.160 ;
        RECT 125.345 162.045 125.705 162.425 ;
        RECT 125.955 162.045 126.315 162.425 ;
        RECT 126.585 162.045 126.945 162.425 ;
        RECT 125.345 161.360 125.705 161.740 ;
        RECT 125.955 161.360 126.315 161.740 ;
        RECT 126.585 161.360 126.945 161.740 ;
        RECT 42.735 160.110 43.585 160.960 ;
        RECT 61.685 160.110 62.535 160.960 ;
        RECT 62.735 160.110 63.585 160.960 ;
        RECT 81.685 160.110 82.535 160.960 ;
        RECT 82.735 160.110 83.585 160.960 ;
        RECT 101.685 160.110 102.535 160.960 ;
        RECT 102.735 160.110 103.585 160.960 ;
        RECT 121.685 160.110 122.535 160.960 ;
        RECT 42.735 159.160 43.585 160.010 ;
        RECT 61.685 159.160 62.535 160.010 ;
        RECT 62.735 159.160 63.585 160.010 ;
        RECT 81.685 159.160 82.535 160.010 ;
        RECT 82.735 159.160 83.585 160.010 ;
        RECT 101.685 159.160 102.535 160.010 ;
        RECT 102.735 159.160 103.585 160.010 ;
        RECT 121.685 159.160 122.535 160.010 ;
        RECT 42.735 157.710 43.585 158.560 ;
        RECT 42.735 156.760 43.585 157.610 ;
        RECT 43.685 156.760 44.535 157.610 ;
        RECT 45.135 156.760 45.985 157.610 ;
        RECT 46.085 156.760 46.935 157.610 ;
        RECT 61.685 157.710 62.535 158.560 ;
        RECT 62.735 157.710 63.585 158.560 ;
        RECT 58.335 156.760 59.185 157.610 ;
        RECT 59.285 156.760 60.135 157.610 ;
        RECT 60.735 156.760 61.585 157.610 ;
        RECT 61.685 156.760 62.535 157.610 ;
        RECT 62.735 156.760 63.585 157.610 ;
        RECT 63.685 156.760 64.535 157.610 ;
        RECT 65.135 156.760 65.985 157.610 ;
        RECT 66.085 156.760 66.935 157.610 ;
        RECT 81.685 157.710 82.535 158.560 ;
        RECT 82.735 157.710 83.585 158.560 ;
        RECT 78.335 156.760 79.185 157.610 ;
        RECT 79.285 156.760 80.135 157.610 ;
        RECT 80.735 156.760 81.585 157.610 ;
        RECT 81.685 156.760 82.535 157.610 ;
        RECT 82.735 156.760 83.585 157.610 ;
        RECT 83.685 156.760 84.535 157.610 ;
        RECT 85.135 156.760 85.985 157.610 ;
        RECT 86.085 156.760 86.935 157.610 ;
        RECT 101.685 157.710 102.535 158.560 ;
        RECT 102.735 157.710 103.585 158.560 ;
        RECT 98.335 156.760 99.185 157.610 ;
        RECT 99.285 156.760 100.135 157.610 ;
        RECT 100.735 156.760 101.585 157.610 ;
        RECT 101.685 156.760 102.535 157.610 ;
        RECT 102.735 156.760 103.585 157.610 ;
        RECT 103.685 156.760 104.535 157.610 ;
        RECT 105.135 156.760 105.985 157.610 ;
        RECT 106.085 156.760 106.935 157.610 ;
        RECT 121.685 157.710 122.535 158.560 ;
        RECT 125.300 159.185 125.700 159.585 ;
        RECT 125.925 159.185 126.325 159.585 ;
        RECT 126.550 159.185 126.950 159.585 ;
        RECT 125.295 158.585 125.695 158.985 ;
        RECT 125.920 158.585 126.320 158.985 ;
        RECT 126.545 158.585 126.945 158.985 ;
        RECT 118.335 156.760 119.185 157.610 ;
        RECT 119.285 156.760 120.135 157.610 ;
        RECT 120.735 156.760 121.585 157.610 ;
        RECT 121.685 156.760 122.535 157.610 ;
        RECT 2.515 141.130 2.875 141.510 ;
        RECT 3.145 141.130 3.505 141.510 ;
        RECT 3.745 141.130 4.105 141.510 ;
        RECT 2.515 140.540 2.875 140.920 ;
        RECT 3.145 140.540 3.505 140.920 ;
        RECT 3.745 140.540 4.105 140.920 ;
        RECT 125.340 141.130 125.700 141.510 ;
        RECT 125.970 141.130 126.330 141.510 ;
        RECT 126.570 141.130 126.930 141.510 ;
        RECT 125.340 140.540 125.700 140.920 ;
        RECT 125.970 140.540 126.330 140.920 ;
        RECT 126.570 140.540 126.930 140.920 ;
        RECT 4.830 139.050 5.680 139.900 ;
        RECT 5.780 139.050 6.630 139.900 ;
        RECT 7.230 139.050 8.080 139.900 ;
        RECT 8.180 139.050 9.030 139.900 ;
        RECT 4.830 138.100 5.680 138.950 ;
        RECT 20.430 139.050 21.280 139.900 ;
        RECT 21.380 139.050 22.230 139.900 ;
        RECT 22.830 139.050 23.680 139.900 ;
        RECT 23.780 139.050 24.630 139.900 ;
        RECT 24.830 139.050 25.680 139.900 ;
        RECT 25.780 139.050 26.630 139.900 ;
        RECT 27.230 139.050 28.080 139.900 ;
        RECT 28.180 139.050 29.030 139.900 ;
        RECT 23.780 138.100 24.630 138.950 ;
        RECT 24.830 138.100 25.680 138.950 ;
        RECT 40.430 139.050 41.280 139.900 ;
        RECT 41.380 139.050 42.230 139.900 ;
        RECT 42.830 139.050 43.680 139.900 ;
        RECT 43.780 139.050 44.630 139.900 ;
        RECT 44.830 139.050 45.680 139.900 ;
        RECT 45.780 139.050 46.630 139.900 ;
        RECT 47.230 139.050 48.080 139.900 ;
        RECT 48.180 139.050 49.030 139.900 ;
        RECT 43.780 138.100 44.630 138.950 ;
        RECT 44.830 138.100 45.680 138.950 ;
        RECT 60.430 139.050 61.280 139.900 ;
        RECT 61.380 139.050 62.230 139.900 ;
        RECT 62.830 139.050 63.680 139.900 ;
        RECT 63.780 139.050 64.630 139.900 ;
        RECT 64.830 139.050 65.680 139.900 ;
        RECT 65.780 139.050 66.630 139.900 ;
        RECT 67.230 139.050 68.080 139.900 ;
        RECT 68.180 139.050 69.030 139.900 ;
        RECT 63.780 138.100 64.630 138.950 ;
        RECT 64.830 138.100 65.680 138.950 ;
        RECT 80.430 139.050 81.280 139.900 ;
        RECT 81.380 139.050 82.230 139.900 ;
        RECT 82.830 139.050 83.680 139.900 ;
        RECT 83.780 139.050 84.630 139.900 ;
        RECT 84.830 139.050 85.680 139.900 ;
        RECT 85.780 139.050 86.630 139.900 ;
        RECT 87.230 139.050 88.080 139.900 ;
        RECT 88.180 139.050 89.030 139.900 ;
        RECT 83.780 138.100 84.630 138.950 ;
        RECT 84.830 138.100 85.680 138.950 ;
        RECT 100.430 139.050 101.280 139.900 ;
        RECT 101.380 139.050 102.230 139.900 ;
        RECT 102.830 139.050 103.680 139.900 ;
        RECT 103.780 139.050 104.630 139.900 ;
        RECT 104.830 139.050 105.680 139.900 ;
        RECT 105.780 139.050 106.630 139.900 ;
        RECT 107.230 139.050 108.080 139.900 ;
        RECT 108.180 139.050 109.030 139.900 ;
        RECT 103.780 138.100 104.630 138.950 ;
        RECT 104.830 138.100 105.680 138.950 ;
        RECT 120.430 139.050 121.280 139.900 ;
        RECT 121.380 139.050 122.230 139.900 ;
        RECT 122.830 139.050 123.680 139.900 ;
        RECT 123.780 139.050 124.630 139.900 ;
        RECT 123.780 138.100 124.630 138.950 ;
        RECT 2.515 137.220 2.875 137.600 ;
        RECT 3.145 137.220 3.505 137.600 ;
        RECT 3.745 137.220 4.105 137.600 ;
        RECT 2.515 136.630 2.875 137.010 ;
        RECT 3.145 136.630 3.505 137.010 ;
        RECT 3.745 136.630 4.105 137.010 ;
        RECT 4.830 136.650 5.680 137.500 ;
        RECT 23.780 136.650 24.630 137.500 ;
        RECT 24.830 136.650 25.680 137.500 ;
        RECT 43.780 136.650 44.630 137.500 ;
        RECT 44.830 136.650 45.680 137.500 ;
        RECT 63.780 136.650 64.630 137.500 ;
        RECT 64.830 136.650 65.680 137.500 ;
        RECT 83.780 136.650 84.630 137.500 ;
        RECT 84.830 136.650 85.680 137.500 ;
        RECT 103.780 136.650 104.630 137.500 ;
        RECT 104.830 136.650 105.680 137.500 ;
        RECT 123.780 136.650 124.630 137.500 ;
        RECT 4.830 135.700 5.680 136.550 ;
        RECT 23.780 135.700 24.630 136.550 ;
        RECT 24.830 135.700 25.680 136.550 ;
        RECT 43.780 135.700 44.630 136.550 ;
        RECT 44.830 135.700 45.680 136.550 ;
        RECT 63.780 135.700 64.630 136.550 ;
        RECT 64.830 135.700 65.680 136.550 ;
        RECT 83.780 135.700 84.630 136.550 ;
        RECT 84.830 135.700 85.680 136.550 ;
        RECT 103.780 135.700 104.630 136.550 ;
        RECT 104.830 135.700 105.680 136.550 ;
        RECT 123.780 135.700 124.630 136.550 ;
        RECT 125.340 137.220 125.700 137.600 ;
        RECT 125.970 137.220 126.330 137.600 ;
        RECT 126.570 137.220 126.930 137.600 ;
        RECT 125.340 136.630 125.700 137.010 ;
        RECT 125.970 136.630 126.330 137.010 ;
        RECT 126.570 136.630 126.930 137.010 ;
        RECT 2.520 134.925 2.880 135.305 ;
        RECT 3.130 134.925 3.490 135.305 ;
        RECT 3.760 134.925 4.120 135.305 ;
        RECT 2.520 134.190 2.880 134.570 ;
        RECT 3.130 134.190 3.490 134.570 ;
        RECT 3.760 134.190 4.120 134.570 ;
        RECT 2.520 133.505 2.880 133.885 ;
        RECT 3.130 133.505 3.490 133.885 ;
        RECT 3.760 133.505 4.120 133.885 ;
        RECT 2.520 126.090 2.880 126.470 ;
        RECT 3.130 126.090 3.490 126.470 ;
        RECT 3.760 126.090 4.120 126.470 ;
        RECT 2.520 125.355 2.880 125.735 ;
        RECT 3.130 125.355 3.490 125.735 ;
        RECT 3.760 125.355 4.120 125.735 ;
        RECT 2.520 124.670 2.880 125.050 ;
        RECT 3.130 124.670 3.490 125.050 ;
        RECT 3.760 124.670 4.120 125.050 ;
        RECT 4.830 123.450 5.680 124.300 ;
        RECT 23.780 123.450 24.630 124.300 ;
        RECT 24.830 123.450 25.680 124.300 ;
        RECT 43.780 123.450 44.630 124.300 ;
        RECT 44.830 123.450 45.680 124.300 ;
        RECT 63.780 123.450 64.630 124.300 ;
        RECT 64.830 123.450 65.680 124.300 ;
        RECT 83.780 123.450 84.630 124.300 ;
        RECT 84.830 123.450 85.680 124.300 ;
        RECT 103.780 123.450 104.630 124.300 ;
        RECT 104.830 123.450 105.680 124.300 ;
        RECT 123.780 123.450 124.630 124.300 ;
        RECT 2.515 122.660 2.875 123.040 ;
        RECT 3.145 122.660 3.505 123.040 ;
        RECT 3.745 122.660 4.105 123.040 ;
        RECT 2.515 122.070 2.875 122.450 ;
        RECT 3.145 122.070 3.505 122.450 ;
        RECT 3.745 122.070 4.105 122.450 ;
        RECT 4.830 122.500 5.680 123.350 ;
        RECT 23.780 122.500 24.630 123.350 ;
        RECT 24.830 122.500 25.680 123.350 ;
        RECT 43.780 122.500 44.630 123.350 ;
        RECT 44.830 122.500 45.680 123.350 ;
        RECT 63.780 122.500 64.630 123.350 ;
        RECT 64.830 122.500 65.680 123.350 ;
        RECT 83.780 122.500 84.630 123.350 ;
        RECT 84.830 122.500 85.680 123.350 ;
        RECT 103.780 122.500 104.630 123.350 ;
        RECT 104.830 122.500 105.680 123.350 ;
        RECT 123.780 122.500 124.630 123.350 ;
        RECT 4.830 121.050 5.680 121.900 ;
        RECT 4.830 120.100 5.680 120.950 ;
        RECT 5.780 120.100 6.630 120.950 ;
        RECT 7.230 120.100 8.080 120.950 ;
        RECT 8.180 120.100 9.030 120.950 ;
        RECT 4.830 119.050 5.680 119.900 ;
        RECT 5.780 119.050 6.630 119.900 ;
        RECT 7.230 119.050 8.080 119.900 ;
        RECT 8.180 119.050 9.030 119.900 ;
        RECT 2.515 117.640 2.875 118.020 ;
        RECT 3.145 117.640 3.505 118.020 ;
        RECT 3.745 117.640 4.105 118.020 ;
        RECT 2.515 117.050 2.875 117.430 ;
        RECT 3.145 117.050 3.505 117.430 ;
        RECT 3.745 117.050 4.105 117.430 ;
        RECT 4.830 118.100 5.680 118.950 ;
        RECT 23.780 121.050 24.630 121.900 ;
        RECT 24.830 121.050 25.680 121.900 ;
        RECT 20.430 120.100 21.280 120.950 ;
        RECT 21.380 120.100 22.230 120.950 ;
        RECT 22.830 120.100 23.680 120.950 ;
        RECT 23.780 120.100 24.630 120.950 ;
        RECT 24.830 120.100 25.680 120.950 ;
        RECT 25.780 120.100 26.630 120.950 ;
        RECT 27.230 120.100 28.080 120.950 ;
        RECT 28.180 120.100 29.030 120.950 ;
        RECT 20.430 119.050 21.280 119.900 ;
        RECT 21.380 119.050 22.230 119.900 ;
        RECT 22.830 119.050 23.680 119.900 ;
        RECT 23.780 119.050 24.630 119.900 ;
        RECT 24.830 119.050 25.680 119.900 ;
        RECT 25.780 119.050 26.630 119.900 ;
        RECT 27.230 119.050 28.080 119.900 ;
        RECT 28.180 119.050 29.030 119.900 ;
        RECT 23.780 118.100 24.630 118.950 ;
        RECT 24.830 118.100 25.680 118.950 ;
        RECT 43.780 121.050 44.630 121.900 ;
        RECT 44.830 121.050 45.680 121.900 ;
        RECT 40.430 120.100 41.280 120.950 ;
        RECT 41.380 120.100 42.230 120.950 ;
        RECT 42.830 120.100 43.680 120.950 ;
        RECT 43.780 120.100 44.630 120.950 ;
        RECT 44.830 120.100 45.680 120.950 ;
        RECT 45.780 120.100 46.630 120.950 ;
        RECT 47.230 120.100 48.080 120.950 ;
        RECT 48.180 120.100 49.030 120.950 ;
        RECT 40.430 119.050 41.280 119.900 ;
        RECT 41.380 119.050 42.230 119.900 ;
        RECT 42.830 119.050 43.680 119.900 ;
        RECT 43.780 119.050 44.630 119.900 ;
        RECT 44.830 119.050 45.680 119.900 ;
        RECT 45.780 119.050 46.630 119.900 ;
        RECT 47.230 119.050 48.080 119.900 ;
        RECT 48.180 119.050 49.030 119.900 ;
        RECT 43.780 118.100 44.630 118.950 ;
        RECT 44.830 118.100 45.680 118.950 ;
        RECT 63.780 121.050 64.630 121.900 ;
        RECT 64.830 121.050 65.680 121.900 ;
        RECT 60.430 120.100 61.280 120.950 ;
        RECT 61.380 120.100 62.230 120.950 ;
        RECT 62.830 120.100 63.680 120.950 ;
        RECT 63.780 120.100 64.630 120.950 ;
        RECT 64.830 120.100 65.680 120.950 ;
        RECT 65.780 120.100 66.630 120.950 ;
        RECT 67.230 120.100 68.080 120.950 ;
        RECT 68.180 120.100 69.030 120.950 ;
        RECT 60.430 119.050 61.280 119.900 ;
        RECT 61.380 119.050 62.230 119.900 ;
        RECT 62.830 119.050 63.680 119.900 ;
        RECT 63.780 119.050 64.630 119.900 ;
        RECT 64.830 119.050 65.680 119.900 ;
        RECT 65.780 119.050 66.630 119.900 ;
        RECT 67.230 119.050 68.080 119.900 ;
        RECT 68.180 119.050 69.030 119.900 ;
        RECT 63.780 118.100 64.630 118.950 ;
        RECT 64.830 118.100 65.680 118.950 ;
        RECT 83.780 121.050 84.630 121.900 ;
        RECT 84.830 121.050 85.680 121.900 ;
        RECT 80.430 120.100 81.280 120.950 ;
        RECT 81.380 120.100 82.230 120.950 ;
        RECT 82.830 120.100 83.680 120.950 ;
        RECT 83.780 120.100 84.630 120.950 ;
        RECT 84.830 120.100 85.680 120.950 ;
        RECT 85.780 120.100 86.630 120.950 ;
        RECT 87.230 120.100 88.080 120.950 ;
        RECT 88.180 120.100 89.030 120.950 ;
        RECT 80.430 119.050 81.280 119.900 ;
        RECT 81.380 119.050 82.230 119.900 ;
        RECT 82.830 119.050 83.680 119.900 ;
        RECT 83.780 119.050 84.630 119.900 ;
        RECT 84.830 119.050 85.680 119.900 ;
        RECT 85.780 119.050 86.630 119.900 ;
        RECT 87.230 119.050 88.080 119.900 ;
        RECT 88.180 119.050 89.030 119.900 ;
        RECT 83.780 118.100 84.630 118.950 ;
        RECT 84.830 118.100 85.680 118.950 ;
        RECT 103.780 121.050 104.630 121.900 ;
        RECT 104.830 121.050 105.680 121.900 ;
        RECT 100.430 120.100 101.280 120.950 ;
        RECT 101.380 120.100 102.230 120.950 ;
        RECT 102.830 120.100 103.680 120.950 ;
        RECT 103.780 120.100 104.630 120.950 ;
        RECT 104.830 120.100 105.680 120.950 ;
        RECT 105.780 120.100 106.630 120.950 ;
        RECT 107.230 120.100 108.080 120.950 ;
        RECT 108.180 120.100 109.030 120.950 ;
        RECT 100.430 119.050 101.280 119.900 ;
        RECT 101.380 119.050 102.230 119.900 ;
        RECT 102.830 119.050 103.680 119.900 ;
        RECT 103.780 119.050 104.630 119.900 ;
        RECT 104.830 119.050 105.680 119.900 ;
        RECT 105.780 119.050 106.630 119.900 ;
        RECT 107.230 119.050 108.080 119.900 ;
        RECT 108.180 119.050 109.030 119.900 ;
        RECT 103.780 118.100 104.630 118.950 ;
        RECT 104.830 118.100 105.680 118.950 ;
        RECT 123.780 121.050 124.630 121.900 ;
        RECT 125.340 122.415 125.700 122.795 ;
        RECT 125.970 122.415 126.330 122.795 ;
        RECT 126.570 122.415 126.930 122.795 ;
        RECT 125.340 121.825 125.700 122.205 ;
        RECT 125.970 121.825 126.330 122.205 ;
        RECT 126.570 121.825 126.930 122.205 ;
        RECT 120.430 120.100 121.280 120.950 ;
        RECT 121.380 120.100 122.230 120.950 ;
        RECT 122.830 120.100 123.680 120.950 ;
        RECT 123.780 120.100 124.630 120.950 ;
        RECT 120.430 119.050 121.280 119.900 ;
        RECT 121.380 119.050 122.230 119.900 ;
        RECT 122.830 119.050 123.680 119.900 ;
        RECT 123.780 119.050 124.630 119.900 ;
        RECT 123.780 118.100 124.630 118.950 ;
        RECT 4.830 116.650 5.680 117.500 ;
        RECT 23.780 116.650 24.630 117.500 ;
        RECT 24.830 116.650 25.680 117.500 ;
        RECT 43.780 116.650 44.630 117.500 ;
        RECT 44.830 116.650 45.680 117.500 ;
        RECT 63.780 116.650 64.630 117.500 ;
        RECT 64.830 116.650 65.680 117.500 ;
        RECT 83.780 116.650 84.630 117.500 ;
        RECT 84.830 116.650 85.680 117.500 ;
        RECT 103.780 116.650 104.630 117.500 ;
        RECT 104.830 116.650 105.680 117.500 ;
        RECT 123.780 116.650 124.630 117.500 ;
        RECT 4.830 115.700 5.680 116.550 ;
        RECT 23.780 115.700 24.630 116.550 ;
        RECT 24.830 115.700 25.680 116.550 ;
        RECT 43.780 115.700 44.630 116.550 ;
        RECT 44.830 115.700 45.680 116.550 ;
        RECT 63.780 115.700 64.630 116.550 ;
        RECT 64.830 115.700 65.680 116.550 ;
        RECT 83.780 115.700 84.630 116.550 ;
        RECT 84.830 115.700 85.680 116.550 ;
        RECT 103.780 115.700 104.630 116.550 ;
        RECT 104.830 115.700 105.680 116.550 ;
        RECT 123.780 115.700 124.630 116.550 ;
        RECT 125.340 116.830 125.700 117.210 ;
        RECT 125.970 116.830 126.330 117.210 ;
        RECT 126.570 116.830 126.930 117.210 ;
        RECT 125.340 116.240 125.700 116.620 ;
        RECT 125.970 116.240 126.330 116.620 ;
        RECT 126.570 116.240 126.930 116.620 ;
        RECT 2.520 114.920 2.880 115.300 ;
        RECT 3.130 114.920 3.490 115.300 ;
        RECT 3.760 114.920 4.120 115.300 ;
        RECT 2.520 114.185 2.880 114.565 ;
        RECT 3.130 114.185 3.490 114.565 ;
        RECT 3.760 114.185 4.120 114.565 ;
        RECT 2.520 113.500 2.880 113.880 ;
        RECT 3.130 113.500 3.490 113.880 ;
        RECT 3.760 113.500 4.120 113.880 ;
        RECT 2.520 106.120 2.880 106.500 ;
        RECT 3.130 106.120 3.490 106.500 ;
        RECT 3.760 106.120 4.120 106.500 ;
        RECT 2.520 105.385 2.880 105.765 ;
        RECT 3.130 105.385 3.490 105.765 ;
        RECT 3.760 105.385 4.120 105.765 ;
        RECT 2.520 104.700 2.880 105.080 ;
        RECT 3.130 104.700 3.490 105.080 ;
        RECT 3.760 104.700 4.120 105.080 ;
        RECT 4.830 103.450 5.680 104.300 ;
        RECT 23.780 103.450 24.630 104.300 ;
        RECT 24.830 103.450 25.680 104.300 ;
        RECT 43.780 103.450 44.630 104.300 ;
        RECT 44.830 103.450 45.680 104.300 ;
        RECT 63.780 103.450 64.630 104.300 ;
        RECT 64.830 103.450 65.680 104.300 ;
        RECT 83.780 103.450 84.630 104.300 ;
        RECT 84.830 103.450 85.680 104.300 ;
        RECT 103.780 103.450 104.630 104.300 ;
        RECT 104.830 103.450 105.680 104.300 ;
        RECT 123.780 103.450 124.630 104.300 ;
        RECT 2.515 102.750 2.875 103.130 ;
        RECT 3.145 102.750 3.505 103.130 ;
        RECT 3.745 102.750 4.105 103.130 ;
        RECT 2.515 102.160 2.875 102.540 ;
        RECT 3.145 102.160 3.505 102.540 ;
        RECT 3.745 102.160 4.105 102.540 ;
        RECT 4.830 102.500 5.680 103.350 ;
        RECT 23.780 102.500 24.630 103.350 ;
        RECT 24.830 102.500 25.680 103.350 ;
        RECT 43.780 102.500 44.630 103.350 ;
        RECT 44.830 102.500 45.680 103.350 ;
        RECT 63.780 102.500 64.630 103.350 ;
        RECT 64.830 102.500 65.680 103.350 ;
        RECT 83.780 102.500 84.630 103.350 ;
        RECT 84.830 102.500 85.680 103.350 ;
        RECT 103.780 102.500 104.630 103.350 ;
        RECT 104.830 102.500 105.680 103.350 ;
        RECT 123.780 102.500 124.630 103.350 ;
        RECT 4.830 101.050 5.680 101.900 ;
        RECT 4.830 100.100 5.680 100.950 ;
        RECT 5.780 100.100 6.630 100.950 ;
        RECT 7.230 100.100 8.080 100.950 ;
        RECT 8.180 100.100 9.030 100.950 ;
        RECT 4.830 99.050 5.680 99.900 ;
        RECT 5.780 99.050 6.630 99.900 ;
        RECT 7.230 99.050 8.080 99.900 ;
        RECT 8.180 99.050 9.030 99.900 ;
        RECT 4.830 98.100 5.680 98.950 ;
        RECT 23.780 101.050 24.630 101.900 ;
        RECT 24.830 101.050 25.680 101.900 ;
        RECT 20.430 100.100 21.280 100.950 ;
        RECT 21.380 100.100 22.230 100.950 ;
        RECT 22.830 100.100 23.680 100.950 ;
        RECT 23.780 100.100 24.630 100.950 ;
        RECT 24.830 100.100 25.680 100.950 ;
        RECT 25.780 100.100 26.630 100.950 ;
        RECT 27.230 100.100 28.080 100.950 ;
        RECT 28.180 100.100 29.030 100.950 ;
        RECT 20.430 99.050 21.280 99.900 ;
        RECT 21.380 99.050 22.230 99.900 ;
        RECT 22.830 99.050 23.680 99.900 ;
        RECT 23.780 99.050 24.630 99.900 ;
        RECT 24.830 99.050 25.680 99.900 ;
        RECT 25.780 99.050 26.630 99.900 ;
        RECT 27.230 99.050 28.080 99.900 ;
        RECT 28.180 99.050 29.030 99.900 ;
        RECT 23.780 98.100 24.630 98.950 ;
        RECT 24.830 98.100 25.680 98.950 ;
        RECT 43.780 101.050 44.630 101.900 ;
        RECT 44.830 101.050 45.680 101.900 ;
        RECT 40.430 100.100 41.280 100.950 ;
        RECT 41.380 100.100 42.230 100.950 ;
        RECT 42.830 100.100 43.680 100.950 ;
        RECT 43.780 100.100 44.630 100.950 ;
        RECT 44.830 100.100 45.680 100.950 ;
        RECT 45.780 100.100 46.630 100.950 ;
        RECT 47.230 100.100 48.080 100.950 ;
        RECT 48.180 100.100 49.030 100.950 ;
        RECT 40.430 99.050 41.280 99.900 ;
        RECT 41.380 99.050 42.230 99.900 ;
        RECT 42.830 99.050 43.680 99.900 ;
        RECT 43.780 99.050 44.630 99.900 ;
        RECT 44.830 99.050 45.680 99.900 ;
        RECT 45.780 99.050 46.630 99.900 ;
        RECT 47.230 99.050 48.080 99.900 ;
        RECT 48.180 99.050 49.030 99.900 ;
        RECT 43.780 98.100 44.630 98.950 ;
        RECT 44.830 98.100 45.680 98.950 ;
        RECT 63.780 101.050 64.630 101.900 ;
        RECT 64.830 101.050 65.680 101.900 ;
        RECT 60.430 100.100 61.280 100.950 ;
        RECT 61.380 100.100 62.230 100.950 ;
        RECT 62.830 100.100 63.680 100.950 ;
        RECT 63.780 100.100 64.630 100.950 ;
        RECT 64.830 100.100 65.680 100.950 ;
        RECT 65.780 100.100 66.630 100.950 ;
        RECT 67.230 100.100 68.080 100.950 ;
        RECT 68.180 100.100 69.030 100.950 ;
        RECT 60.430 99.050 61.280 99.900 ;
        RECT 61.380 99.050 62.230 99.900 ;
        RECT 62.830 99.050 63.680 99.900 ;
        RECT 63.780 99.050 64.630 99.900 ;
        RECT 64.830 99.050 65.680 99.900 ;
        RECT 65.780 99.050 66.630 99.900 ;
        RECT 67.230 99.050 68.080 99.900 ;
        RECT 68.180 99.050 69.030 99.900 ;
        RECT 63.780 98.100 64.630 98.950 ;
        RECT 64.830 98.100 65.680 98.950 ;
        RECT 83.780 101.050 84.630 101.900 ;
        RECT 84.830 101.050 85.680 101.900 ;
        RECT 80.430 100.100 81.280 100.950 ;
        RECT 81.380 100.100 82.230 100.950 ;
        RECT 82.830 100.100 83.680 100.950 ;
        RECT 83.780 100.100 84.630 100.950 ;
        RECT 84.830 100.100 85.680 100.950 ;
        RECT 85.780 100.100 86.630 100.950 ;
        RECT 87.230 100.100 88.080 100.950 ;
        RECT 88.180 100.100 89.030 100.950 ;
        RECT 80.430 99.050 81.280 99.900 ;
        RECT 81.380 99.050 82.230 99.900 ;
        RECT 82.830 99.050 83.680 99.900 ;
        RECT 83.780 99.050 84.630 99.900 ;
        RECT 84.830 99.050 85.680 99.900 ;
        RECT 85.780 99.050 86.630 99.900 ;
        RECT 87.230 99.050 88.080 99.900 ;
        RECT 88.180 99.050 89.030 99.900 ;
        RECT 83.780 98.100 84.630 98.950 ;
        RECT 84.830 98.100 85.680 98.950 ;
        RECT 103.780 101.050 104.630 101.900 ;
        RECT 104.830 101.050 105.680 101.900 ;
        RECT 100.430 100.100 101.280 100.950 ;
        RECT 101.380 100.100 102.230 100.950 ;
        RECT 102.830 100.100 103.680 100.950 ;
        RECT 103.780 100.100 104.630 100.950 ;
        RECT 104.830 100.100 105.680 100.950 ;
        RECT 105.780 100.100 106.630 100.950 ;
        RECT 107.230 100.100 108.080 100.950 ;
        RECT 108.180 100.100 109.030 100.950 ;
        RECT 100.430 99.050 101.280 99.900 ;
        RECT 101.380 99.050 102.230 99.900 ;
        RECT 102.830 99.050 103.680 99.900 ;
        RECT 103.780 99.050 104.630 99.900 ;
        RECT 104.830 99.050 105.680 99.900 ;
        RECT 105.780 99.050 106.630 99.900 ;
        RECT 107.230 99.050 108.080 99.900 ;
        RECT 108.180 99.050 109.030 99.900 ;
        RECT 103.780 98.100 104.630 98.950 ;
        RECT 104.830 98.100 105.680 98.950 ;
        RECT 123.780 101.050 124.630 101.900 ;
        RECT 125.340 102.615 125.700 102.995 ;
        RECT 125.970 102.615 126.330 102.995 ;
        RECT 126.570 102.615 126.930 102.995 ;
        RECT 125.340 102.025 125.700 102.405 ;
        RECT 125.970 102.025 126.330 102.405 ;
        RECT 126.570 102.025 126.930 102.405 ;
        RECT 120.430 100.100 121.280 100.950 ;
        RECT 121.380 100.100 122.230 100.950 ;
        RECT 122.830 100.100 123.680 100.950 ;
        RECT 123.780 100.100 124.630 100.950 ;
        RECT 120.430 99.050 121.280 99.900 ;
        RECT 121.380 99.050 122.230 99.900 ;
        RECT 122.830 99.050 123.680 99.900 ;
        RECT 123.780 99.050 124.630 99.900 ;
        RECT 123.780 98.100 124.630 98.950 ;
        RECT 2.515 97.340 2.875 97.720 ;
        RECT 3.145 97.340 3.505 97.720 ;
        RECT 3.745 97.340 4.105 97.720 ;
        RECT 2.515 96.750 2.875 97.130 ;
        RECT 3.145 96.750 3.505 97.130 ;
        RECT 3.745 96.750 4.105 97.130 ;
        RECT 4.830 96.650 5.680 97.500 ;
        RECT 23.780 96.650 24.630 97.500 ;
        RECT 24.830 96.650 25.680 97.500 ;
        RECT 43.780 96.650 44.630 97.500 ;
        RECT 44.830 96.650 45.680 97.500 ;
        RECT 63.780 96.650 64.630 97.500 ;
        RECT 64.830 96.650 65.680 97.500 ;
        RECT 83.780 96.650 84.630 97.500 ;
        RECT 84.830 96.650 85.680 97.500 ;
        RECT 103.780 96.650 104.630 97.500 ;
        RECT 104.830 96.650 105.680 97.500 ;
        RECT 123.780 96.650 124.630 97.500 ;
        RECT 4.830 95.700 5.680 96.550 ;
        RECT 23.780 95.700 24.630 96.550 ;
        RECT 24.830 95.700 25.680 96.550 ;
        RECT 43.780 95.700 44.630 96.550 ;
        RECT 44.830 95.700 45.680 96.550 ;
        RECT 63.780 95.700 64.630 96.550 ;
        RECT 64.830 95.700 65.680 96.550 ;
        RECT 83.780 95.700 84.630 96.550 ;
        RECT 84.830 95.700 85.680 96.550 ;
        RECT 103.780 95.700 104.630 96.550 ;
        RECT 104.830 95.700 105.680 96.550 ;
        RECT 123.780 95.700 124.630 96.550 ;
        RECT 125.340 96.740 125.700 97.120 ;
        RECT 125.970 96.740 126.330 97.120 ;
        RECT 126.570 96.740 126.930 97.120 ;
        RECT 125.340 96.150 125.700 96.530 ;
        RECT 125.970 96.150 126.330 96.530 ;
        RECT 126.570 96.150 126.930 96.530 ;
        RECT 2.520 94.920 2.880 95.300 ;
        RECT 3.130 94.920 3.490 95.300 ;
        RECT 3.760 94.920 4.120 95.300 ;
        RECT 2.520 94.185 2.880 94.565 ;
        RECT 3.130 94.185 3.490 94.565 ;
        RECT 3.760 94.185 4.120 94.565 ;
        RECT 2.520 93.500 2.880 93.880 ;
        RECT 3.130 93.500 3.490 93.880 ;
        RECT 3.760 93.500 4.120 93.880 ;
        RECT 2.520 86.125 2.880 86.505 ;
        RECT 3.130 86.125 3.490 86.505 ;
        RECT 3.760 86.125 4.120 86.505 ;
        RECT 2.520 85.390 2.880 85.770 ;
        RECT 3.130 85.390 3.490 85.770 ;
        RECT 3.760 85.390 4.120 85.770 ;
        RECT 2.520 84.705 2.880 85.085 ;
        RECT 3.130 84.705 3.490 85.085 ;
        RECT 3.760 84.705 4.120 85.085 ;
        RECT 2.515 82.965 2.875 83.345 ;
        RECT 3.145 82.965 3.505 83.345 ;
        RECT 3.745 82.965 4.105 83.345 ;
        RECT 2.515 82.375 2.875 82.755 ;
        RECT 3.145 82.375 3.505 82.755 ;
        RECT 3.745 82.375 4.105 82.755 ;
        RECT 4.830 83.450 5.680 84.300 ;
        RECT 23.780 83.450 24.630 84.300 ;
        RECT 24.830 83.450 25.680 84.300 ;
        RECT 43.780 83.450 44.630 84.300 ;
        RECT 44.830 83.450 45.680 84.300 ;
        RECT 63.780 83.450 64.630 84.300 ;
        RECT 64.830 83.450 65.680 84.300 ;
        RECT 83.780 83.450 84.630 84.300 ;
        RECT 84.830 83.450 85.680 84.300 ;
        RECT 103.780 83.450 104.630 84.300 ;
        RECT 104.830 83.450 105.680 84.300 ;
        RECT 123.780 83.450 124.630 84.300 ;
        RECT 4.830 82.500 5.680 83.350 ;
        RECT 23.780 82.500 24.630 83.350 ;
        RECT 24.830 82.500 25.680 83.350 ;
        RECT 43.780 82.500 44.630 83.350 ;
        RECT 44.830 82.500 45.680 83.350 ;
        RECT 63.780 82.500 64.630 83.350 ;
        RECT 64.830 82.500 65.680 83.350 ;
        RECT 83.780 82.500 84.630 83.350 ;
        RECT 84.830 82.500 85.680 83.350 ;
        RECT 103.780 82.500 104.630 83.350 ;
        RECT 104.830 82.500 105.680 83.350 ;
        RECT 123.780 82.500 124.630 83.350 ;
        RECT 4.830 81.050 5.680 81.900 ;
        RECT 4.830 80.100 5.680 80.950 ;
        RECT 5.780 80.100 6.630 80.950 ;
        RECT 7.230 80.100 8.080 80.950 ;
        RECT 8.180 80.100 9.030 80.950 ;
        RECT 4.830 79.050 5.680 79.900 ;
        RECT 5.780 79.050 6.630 79.900 ;
        RECT 7.230 79.050 8.080 79.900 ;
        RECT 8.180 79.050 9.030 79.900 ;
        RECT 4.830 78.100 5.680 78.950 ;
        RECT 23.780 81.050 24.630 81.900 ;
        RECT 24.830 81.050 25.680 81.900 ;
        RECT 20.430 80.100 21.280 80.950 ;
        RECT 21.380 80.100 22.230 80.950 ;
        RECT 22.830 80.100 23.680 80.950 ;
        RECT 23.780 80.100 24.630 80.950 ;
        RECT 24.830 80.100 25.680 80.950 ;
        RECT 25.780 80.100 26.630 80.950 ;
        RECT 27.230 80.100 28.080 80.950 ;
        RECT 28.180 80.100 29.030 80.950 ;
        RECT 20.430 79.050 21.280 79.900 ;
        RECT 21.380 79.050 22.230 79.900 ;
        RECT 22.830 79.050 23.680 79.900 ;
        RECT 23.780 79.050 24.630 79.900 ;
        RECT 24.830 79.050 25.680 79.900 ;
        RECT 25.780 79.050 26.630 79.900 ;
        RECT 27.230 79.050 28.080 79.900 ;
        RECT 28.180 79.050 29.030 79.900 ;
        RECT 23.780 78.100 24.630 78.950 ;
        RECT 24.830 78.100 25.680 78.950 ;
        RECT 43.780 81.050 44.630 81.900 ;
        RECT 44.830 81.050 45.680 81.900 ;
        RECT 40.430 80.100 41.280 80.950 ;
        RECT 41.380 80.100 42.230 80.950 ;
        RECT 42.830 80.100 43.680 80.950 ;
        RECT 43.780 80.100 44.630 80.950 ;
        RECT 44.830 80.100 45.680 80.950 ;
        RECT 45.780 80.100 46.630 80.950 ;
        RECT 47.230 80.100 48.080 80.950 ;
        RECT 48.180 80.100 49.030 80.950 ;
        RECT 40.430 79.050 41.280 79.900 ;
        RECT 41.380 79.050 42.230 79.900 ;
        RECT 42.830 79.050 43.680 79.900 ;
        RECT 43.780 79.050 44.630 79.900 ;
        RECT 44.830 79.050 45.680 79.900 ;
        RECT 45.780 79.050 46.630 79.900 ;
        RECT 47.230 79.050 48.080 79.900 ;
        RECT 48.180 79.050 49.030 79.900 ;
        RECT 43.780 78.100 44.630 78.950 ;
        RECT 44.830 78.100 45.680 78.950 ;
        RECT 63.780 81.050 64.630 81.900 ;
        RECT 64.830 81.050 65.680 81.900 ;
        RECT 60.430 80.100 61.280 80.950 ;
        RECT 61.380 80.100 62.230 80.950 ;
        RECT 62.830 80.100 63.680 80.950 ;
        RECT 63.780 80.100 64.630 80.950 ;
        RECT 64.830 80.100 65.680 80.950 ;
        RECT 65.780 80.100 66.630 80.950 ;
        RECT 67.230 80.100 68.080 80.950 ;
        RECT 68.180 80.100 69.030 80.950 ;
        RECT 60.430 79.050 61.280 79.900 ;
        RECT 61.380 79.050 62.230 79.900 ;
        RECT 62.830 79.050 63.680 79.900 ;
        RECT 63.780 79.050 64.630 79.900 ;
        RECT 64.830 79.050 65.680 79.900 ;
        RECT 65.780 79.050 66.630 79.900 ;
        RECT 67.230 79.050 68.080 79.900 ;
        RECT 68.180 79.050 69.030 79.900 ;
        RECT 63.780 78.100 64.630 78.950 ;
        RECT 64.830 78.100 65.680 78.950 ;
        RECT 83.780 81.050 84.630 81.900 ;
        RECT 84.830 81.050 85.680 81.900 ;
        RECT 80.430 80.100 81.280 80.950 ;
        RECT 81.380 80.100 82.230 80.950 ;
        RECT 82.830 80.100 83.680 80.950 ;
        RECT 83.780 80.100 84.630 80.950 ;
        RECT 84.830 80.100 85.680 80.950 ;
        RECT 85.780 80.100 86.630 80.950 ;
        RECT 87.230 80.100 88.080 80.950 ;
        RECT 88.180 80.100 89.030 80.950 ;
        RECT 80.430 79.050 81.280 79.900 ;
        RECT 81.380 79.050 82.230 79.900 ;
        RECT 82.830 79.050 83.680 79.900 ;
        RECT 83.780 79.050 84.630 79.900 ;
        RECT 84.830 79.050 85.680 79.900 ;
        RECT 85.780 79.050 86.630 79.900 ;
        RECT 87.230 79.050 88.080 79.900 ;
        RECT 88.180 79.050 89.030 79.900 ;
        RECT 83.780 78.100 84.630 78.950 ;
        RECT 84.830 78.100 85.680 78.950 ;
        RECT 103.780 81.050 104.630 81.900 ;
        RECT 104.830 81.050 105.680 81.900 ;
        RECT 100.430 80.100 101.280 80.950 ;
        RECT 101.380 80.100 102.230 80.950 ;
        RECT 102.830 80.100 103.680 80.950 ;
        RECT 103.780 80.100 104.630 80.950 ;
        RECT 104.830 80.100 105.680 80.950 ;
        RECT 105.780 80.100 106.630 80.950 ;
        RECT 107.230 80.100 108.080 80.950 ;
        RECT 108.180 80.100 109.030 80.950 ;
        RECT 100.430 79.050 101.280 79.900 ;
        RECT 101.380 79.050 102.230 79.900 ;
        RECT 102.830 79.050 103.680 79.900 ;
        RECT 103.780 79.050 104.630 79.900 ;
        RECT 104.830 79.050 105.680 79.900 ;
        RECT 105.780 79.050 106.630 79.900 ;
        RECT 107.230 79.050 108.080 79.900 ;
        RECT 108.180 79.050 109.030 79.900 ;
        RECT 103.780 78.100 104.630 78.950 ;
        RECT 104.830 78.100 105.680 78.950 ;
        RECT 123.780 81.050 124.630 81.900 ;
        RECT 125.340 82.535 125.700 82.915 ;
        RECT 125.970 82.535 126.330 82.915 ;
        RECT 126.570 82.535 126.930 82.915 ;
        RECT 125.340 81.945 125.700 82.325 ;
        RECT 125.970 81.945 126.330 82.325 ;
        RECT 126.570 81.945 126.930 82.325 ;
        RECT 120.430 80.100 121.280 80.950 ;
        RECT 121.380 80.100 122.230 80.950 ;
        RECT 122.830 80.100 123.680 80.950 ;
        RECT 123.780 80.100 124.630 80.950 ;
        RECT 120.430 79.050 121.280 79.900 ;
        RECT 121.380 79.050 122.230 79.900 ;
        RECT 122.830 79.050 123.680 79.900 ;
        RECT 123.780 79.050 124.630 79.900 ;
        RECT 123.780 78.100 124.630 78.950 ;
        RECT 2.515 77.460 2.875 77.840 ;
        RECT 3.145 77.460 3.505 77.840 ;
        RECT 3.745 77.460 4.105 77.840 ;
        RECT 2.515 76.870 2.875 77.250 ;
        RECT 3.145 76.870 3.505 77.250 ;
        RECT 3.745 76.870 4.105 77.250 ;
        RECT 4.830 76.650 5.680 77.500 ;
        RECT 23.780 76.650 24.630 77.500 ;
        RECT 24.830 76.650 25.680 77.500 ;
        RECT 43.780 76.650 44.630 77.500 ;
        RECT 44.830 76.650 45.680 77.500 ;
        RECT 63.780 76.650 64.630 77.500 ;
        RECT 64.830 76.650 65.680 77.500 ;
        RECT 83.780 76.650 84.630 77.500 ;
        RECT 84.830 76.650 85.680 77.500 ;
        RECT 103.780 76.650 104.630 77.500 ;
        RECT 104.830 76.650 105.680 77.500 ;
        RECT 123.780 76.650 124.630 77.500 ;
        RECT 4.830 75.700 5.680 76.550 ;
        RECT 23.780 75.700 24.630 76.550 ;
        RECT 24.830 75.700 25.680 76.550 ;
        RECT 43.780 75.700 44.630 76.550 ;
        RECT 44.830 75.700 45.680 76.550 ;
        RECT 63.780 75.700 64.630 76.550 ;
        RECT 64.830 75.700 65.680 76.550 ;
        RECT 83.780 75.700 84.630 76.550 ;
        RECT 84.830 75.700 85.680 76.550 ;
        RECT 103.780 75.700 104.630 76.550 ;
        RECT 104.830 75.700 105.680 76.550 ;
        RECT 123.780 75.700 124.630 76.550 ;
        RECT 125.340 76.680 125.700 77.060 ;
        RECT 125.970 76.680 126.330 77.060 ;
        RECT 126.570 76.680 126.930 77.060 ;
        RECT 125.340 76.090 125.700 76.470 ;
        RECT 125.970 76.090 126.330 76.470 ;
        RECT 126.570 76.090 126.930 76.470 ;
        RECT 2.520 74.920 2.880 75.300 ;
        RECT 3.130 74.920 3.490 75.300 ;
        RECT 3.760 74.920 4.120 75.300 ;
        RECT 2.520 74.185 2.880 74.565 ;
        RECT 3.130 74.185 3.490 74.565 ;
        RECT 3.760 74.185 4.120 74.565 ;
        RECT 2.520 73.500 2.880 73.880 ;
        RECT 3.130 73.500 3.490 73.880 ;
        RECT 3.760 73.500 4.120 73.880 ;
        RECT 2.520 66.120 2.880 66.500 ;
        RECT 3.130 66.120 3.490 66.500 ;
        RECT 3.760 66.120 4.120 66.500 ;
        RECT 2.520 65.385 2.880 65.765 ;
        RECT 3.130 65.385 3.490 65.765 ;
        RECT 3.760 65.385 4.120 65.765 ;
        RECT 2.520 64.700 2.880 65.080 ;
        RECT 3.130 64.700 3.490 65.080 ;
        RECT 3.760 64.700 4.120 65.080 ;
        RECT 2.515 63.130 2.875 63.510 ;
        RECT 3.145 63.130 3.505 63.510 ;
        RECT 3.745 63.130 4.105 63.510 ;
        RECT 2.515 62.540 2.875 62.920 ;
        RECT 3.145 62.540 3.505 62.920 ;
        RECT 3.745 62.540 4.105 62.920 ;
        RECT 4.830 63.450 5.680 64.300 ;
        RECT 23.780 63.450 24.630 64.300 ;
        RECT 24.830 63.450 25.680 64.300 ;
        RECT 43.780 63.450 44.630 64.300 ;
        RECT 44.830 63.450 45.680 64.300 ;
        RECT 63.780 63.450 64.630 64.300 ;
        RECT 64.830 63.450 65.680 64.300 ;
        RECT 83.780 63.450 84.630 64.300 ;
        RECT 84.830 63.450 85.680 64.300 ;
        RECT 103.780 63.450 104.630 64.300 ;
        RECT 104.830 63.450 105.680 64.300 ;
        RECT 123.780 63.450 124.630 64.300 ;
        RECT 4.830 62.500 5.680 63.350 ;
        RECT 23.780 62.500 24.630 63.350 ;
        RECT 24.830 62.500 25.680 63.350 ;
        RECT 43.780 62.500 44.630 63.350 ;
        RECT 44.830 62.500 45.680 63.350 ;
        RECT 63.780 62.500 64.630 63.350 ;
        RECT 64.830 62.500 65.680 63.350 ;
        RECT 83.780 62.500 84.630 63.350 ;
        RECT 84.830 62.500 85.680 63.350 ;
        RECT 103.780 62.500 104.630 63.350 ;
        RECT 104.830 62.500 105.680 63.350 ;
        RECT 123.780 62.500 124.630 63.350 ;
        RECT 125.340 62.875 125.700 63.255 ;
        RECT 125.970 62.875 126.330 63.255 ;
        RECT 126.570 62.875 126.930 63.255 ;
        RECT 125.340 62.285 125.700 62.665 ;
        RECT 125.970 62.285 126.330 62.665 ;
        RECT 126.570 62.285 126.930 62.665 ;
        RECT 4.830 61.050 5.680 61.900 ;
        RECT 4.830 60.100 5.680 60.950 ;
        RECT 5.780 60.100 6.630 60.950 ;
        RECT 7.230 60.100 8.080 60.950 ;
        RECT 8.180 60.100 9.030 60.950 ;
        RECT 4.830 59.050 5.680 59.900 ;
        RECT 5.780 59.050 6.630 59.900 ;
        RECT 7.230 59.050 8.080 59.900 ;
        RECT 8.180 59.050 9.030 59.900 ;
        RECT 4.830 58.100 5.680 58.950 ;
        RECT 23.780 61.050 24.630 61.900 ;
        RECT 24.830 61.050 25.680 61.900 ;
        RECT 20.430 60.100 21.280 60.950 ;
        RECT 21.380 60.100 22.230 60.950 ;
        RECT 22.830 60.100 23.680 60.950 ;
        RECT 23.780 60.100 24.630 60.950 ;
        RECT 24.830 60.100 25.680 60.950 ;
        RECT 25.780 60.100 26.630 60.950 ;
        RECT 27.230 60.100 28.080 60.950 ;
        RECT 28.180 60.100 29.030 60.950 ;
        RECT 20.430 59.050 21.280 59.900 ;
        RECT 21.380 59.050 22.230 59.900 ;
        RECT 22.830 59.050 23.680 59.900 ;
        RECT 23.780 59.050 24.630 59.900 ;
        RECT 24.830 59.050 25.680 59.900 ;
        RECT 25.780 59.050 26.630 59.900 ;
        RECT 27.230 59.050 28.080 59.900 ;
        RECT 28.180 59.050 29.030 59.900 ;
        RECT 23.780 58.100 24.630 58.950 ;
        RECT 24.830 58.100 25.680 58.950 ;
        RECT 43.780 61.050 44.630 61.900 ;
        RECT 44.830 61.050 45.680 61.900 ;
        RECT 40.430 60.100 41.280 60.950 ;
        RECT 41.380 60.100 42.230 60.950 ;
        RECT 42.830 60.100 43.680 60.950 ;
        RECT 43.780 60.100 44.630 60.950 ;
        RECT 44.830 60.100 45.680 60.950 ;
        RECT 45.780 60.100 46.630 60.950 ;
        RECT 47.230 60.100 48.080 60.950 ;
        RECT 48.180 60.100 49.030 60.950 ;
        RECT 40.430 59.050 41.280 59.900 ;
        RECT 41.380 59.050 42.230 59.900 ;
        RECT 42.830 59.050 43.680 59.900 ;
        RECT 43.780 59.050 44.630 59.900 ;
        RECT 44.830 59.050 45.680 59.900 ;
        RECT 45.780 59.050 46.630 59.900 ;
        RECT 47.230 59.050 48.080 59.900 ;
        RECT 48.180 59.050 49.030 59.900 ;
        RECT 43.780 58.100 44.630 58.950 ;
        RECT 44.830 58.100 45.680 58.950 ;
        RECT 63.780 61.050 64.630 61.900 ;
        RECT 64.830 61.050 65.680 61.900 ;
        RECT 60.430 60.100 61.280 60.950 ;
        RECT 61.380 60.100 62.230 60.950 ;
        RECT 62.830 60.100 63.680 60.950 ;
        RECT 63.780 60.100 64.630 60.950 ;
        RECT 64.830 60.100 65.680 60.950 ;
        RECT 65.780 60.100 66.630 60.950 ;
        RECT 67.230 60.100 68.080 60.950 ;
        RECT 68.180 60.100 69.030 60.950 ;
        RECT 60.430 59.050 61.280 59.900 ;
        RECT 61.380 59.050 62.230 59.900 ;
        RECT 62.830 59.050 63.680 59.900 ;
        RECT 63.780 59.050 64.630 59.900 ;
        RECT 64.830 59.050 65.680 59.900 ;
        RECT 65.780 59.050 66.630 59.900 ;
        RECT 67.230 59.050 68.080 59.900 ;
        RECT 68.180 59.050 69.030 59.900 ;
        RECT 63.780 58.100 64.630 58.950 ;
        RECT 64.830 58.100 65.680 58.950 ;
        RECT 83.780 61.050 84.630 61.900 ;
        RECT 84.830 61.050 85.680 61.900 ;
        RECT 80.430 60.100 81.280 60.950 ;
        RECT 81.380 60.100 82.230 60.950 ;
        RECT 82.830 60.100 83.680 60.950 ;
        RECT 83.780 60.100 84.630 60.950 ;
        RECT 84.830 60.100 85.680 60.950 ;
        RECT 85.780 60.100 86.630 60.950 ;
        RECT 87.230 60.100 88.080 60.950 ;
        RECT 88.180 60.100 89.030 60.950 ;
        RECT 80.430 59.050 81.280 59.900 ;
        RECT 81.380 59.050 82.230 59.900 ;
        RECT 82.830 59.050 83.680 59.900 ;
        RECT 83.780 59.050 84.630 59.900 ;
        RECT 84.830 59.050 85.680 59.900 ;
        RECT 85.780 59.050 86.630 59.900 ;
        RECT 87.230 59.050 88.080 59.900 ;
        RECT 88.180 59.050 89.030 59.900 ;
        RECT 83.780 58.100 84.630 58.950 ;
        RECT 84.830 58.100 85.680 58.950 ;
        RECT 103.780 61.050 104.630 61.900 ;
        RECT 104.830 61.050 105.680 61.900 ;
        RECT 100.430 60.100 101.280 60.950 ;
        RECT 101.380 60.100 102.230 60.950 ;
        RECT 102.830 60.100 103.680 60.950 ;
        RECT 103.780 60.100 104.630 60.950 ;
        RECT 104.830 60.100 105.680 60.950 ;
        RECT 105.780 60.100 106.630 60.950 ;
        RECT 107.230 60.100 108.080 60.950 ;
        RECT 108.180 60.100 109.030 60.950 ;
        RECT 100.430 59.050 101.280 59.900 ;
        RECT 101.380 59.050 102.230 59.900 ;
        RECT 102.830 59.050 103.680 59.900 ;
        RECT 103.780 59.050 104.630 59.900 ;
        RECT 104.830 59.050 105.680 59.900 ;
        RECT 105.780 59.050 106.630 59.900 ;
        RECT 107.230 59.050 108.080 59.900 ;
        RECT 108.180 59.050 109.030 59.900 ;
        RECT 103.780 58.100 104.630 58.950 ;
        RECT 104.830 58.100 105.680 58.950 ;
        RECT 123.780 61.050 124.630 61.900 ;
        RECT 120.430 60.100 121.280 60.950 ;
        RECT 121.380 60.100 122.230 60.950 ;
        RECT 122.830 60.100 123.680 60.950 ;
        RECT 123.780 60.100 124.630 60.950 ;
        RECT 120.430 59.050 121.280 59.900 ;
        RECT 121.380 59.050 122.230 59.900 ;
        RECT 122.830 59.050 123.680 59.900 ;
        RECT 123.780 59.050 124.630 59.900 ;
        RECT 123.780 58.100 124.630 58.950 ;
        RECT 2.515 57.050 2.875 57.430 ;
        RECT 3.145 57.050 3.505 57.430 ;
        RECT 3.745 57.050 4.105 57.430 ;
        RECT 2.515 56.460 2.875 56.840 ;
        RECT 3.145 56.460 3.505 56.840 ;
        RECT 3.745 56.460 4.105 56.840 ;
        RECT 4.830 56.650 5.680 57.500 ;
        RECT 23.780 56.650 24.630 57.500 ;
        RECT 24.830 56.650 25.680 57.500 ;
        RECT 43.780 56.650 44.630 57.500 ;
        RECT 44.830 56.650 45.680 57.500 ;
        RECT 63.780 56.650 64.630 57.500 ;
        RECT 64.830 56.650 65.680 57.500 ;
        RECT 83.780 56.650 84.630 57.500 ;
        RECT 84.830 56.650 85.680 57.500 ;
        RECT 103.780 56.650 104.630 57.500 ;
        RECT 104.830 56.650 105.680 57.500 ;
        RECT 123.780 56.650 124.630 57.500 ;
        RECT 4.830 55.700 5.680 56.550 ;
        RECT 23.780 55.700 24.630 56.550 ;
        RECT 24.830 55.700 25.680 56.550 ;
        RECT 43.780 55.700 44.630 56.550 ;
        RECT 44.830 55.700 45.680 56.550 ;
        RECT 63.780 55.700 64.630 56.550 ;
        RECT 64.830 55.700 65.680 56.550 ;
        RECT 83.780 55.700 84.630 56.550 ;
        RECT 84.830 55.700 85.680 56.550 ;
        RECT 103.780 55.700 104.630 56.550 ;
        RECT 104.830 55.700 105.680 56.550 ;
        RECT 123.780 55.700 124.630 56.550 ;
        RECT 125.340 56.805 125.700 57.185 ;
        RECT 125.970 56.805 126.330 57.185 ;
        RECT 126.570 56.805 126.930 57.185 ;
        RECT 125.340 56.215 125.700 56.595 ;
        RECT 125.970 56.215 126.330 56.595 ;
        RECT 126.570 56.215 126.930 56.595 ;
        RECT 2.520 54.920 2.880 55.300 ;
        RECT 3.130 54.920 3.490 55.300 ;
        RECT 3.760 54.920 4.120 55.300 ;
        RECT 2.520 54.185 2.880 54.565 ;
        RECT 3.130 54.185 3.490 54.565 ;
        RECT 3.760 54.185 4.120 54.565 ;
        RECT 2.520 53.500 2.880 53.880 ;
        RECT 3.130 53.500 3.490 53.880 ;
        RECT 3.760 53.500 4.120 53.880 ;
        RECT 2.520 46.120 2.880 46.500 ;
        RECT 3.130 46.120 3.490 46.500 ;
        RECT 3.760 46.120 4.120 46.500 ;
        RECT 2.520 45.385 2.880 45.765 ;
        RECT 3.130 45.385 3.490 45.765 ;
        RECT 3.760 45.385 4.120 45.765 ;
        RECT 2.520 44.700 2.880 45.080 ;
        RECT 3.130 44.700 3.490 45.080 ;
        RECT 3.760 44.700 4.120 45.080 ;
        RECT 4.830 43.450 5.680 44.300 ;
        RECT 23.780 43.450 24.630 44.300 ;
        RECT 24.830 43.450 25.680 44.300 ;
        RECT 43.780 43.450 44.630 44.300 ;
        RECT 44.830 43.450 45.680 44.300 ;
        RECT 63.780 43.450 64.630 44.300 ;
        RECT 64.830 43.450 65.680 44.300 ;
        RECT 83.780 43.450 84.630 44.300 ;
        RECT 84.830 43.450 85.680 44.300 ;
        RECT 103.780 43.450 104.630 44.300 ;
        RECT 104.830 43.450 105.680 44.300 ;
        RECT 123.780 43.450 124.630 44.300 ;
        RECT 2.515 42.725 2.875 43.105 ;
        RECT 3.145 42.725 3.505 43.105 ;
        RECT 3.745 42.725 4.105 43.105 ;
        RECT 2.515 42.135 2.875 42.515 ;
        RECT 3.145 42.135 3.505 42.515 ;
        RECT 3.745 42.135 4.105 42.515 ;
        RECT 4.830 42.500 5.680 43.350 ;
        RECT 23.780 42.500 24.630 43.350 ;
        RECT 24.830 42.500 25.680 43.350 ;
        RECT 43.780 42.500 44.630 43.350 ;
        RECT 44.830 42.500 45.680 43.350 ;
        RECT 63.780 42.500 64.630 43.350 ;
        RECT 64.830 42.500 65.680 43.350 ;
        RECT 83.780 42.500 84.630 43.350 ;
        RECT 84.830 42.500 85.680 43.350 ;
        RECT 103.780 42.500 104.630 43.350 ;
        RECT 104.830 42.500 105.680 43.350 ;
        RECT 123.780 42.500 124.630 43.350 ;
        RECT 4.830 41.050 5.680 41.900 ;
        RECT 4.830 40.100 5.680 40.950 ;
        RECT 5.780 40.100 6.630 40.950 ;
        RECT 7.230 40.100 8.080 40.950 ;
        RECT 8.180 40.100 9.030 40.950 ;
        RECT 4.830 39.050 5.680 39.900 ;
        RECT 5.780 39.050 6.630 39.900 ;
        RECT 7.230 39.050 8.080 39.900 ;
        RECT 8.180 39.050 9.030 39.900 ;
        RECT 4.830 38.100 5.680 38.950 ;
        RECT 23.780 41.050 24.630 41.900 ;
        RECT 24.830 41.050 25.680 41.900 ;
        RECT 20.430 40.100 21.280 40.950 ;
        RECT 21.380 40.100 22.230 40.950 ;
        RECT 22.830 40.100 23.680 40.950 ;
        RECT 23.780 40.100 24.630 40.950 ;
        RECT 24.830 40.100 25.680 40.950 ;
        RECT 25.780 40.100 26.630 40.950 ;
        RECT 27.230 40.100 28.080 40.950 ;
        RECT 28.180 40.100 29.030 40.950 ;
        RECT 20.430 39.050 21.280 39.900 ;
        RECT 21.380 39.050 22.230 39.900 ;
        RECT 22.830 39.050 23.680 39.900 ;
        RECT 23.780 39.050 24.630 39.900 ;
        RECT 24.830 39.050 25.680 39.900 ;
        RECT 25.780 39.050 26.630 39.900 ;
        RECT 27.230 39.050 28.080 39.900 ;
        RECT 28.180 39.050 29.030 39.900 ;
        RECT 23.780 38.100 24.630 38.950 ;
        RECT 24.830 38.100 25.680 38.950 ;
        RECT 43.780 41.050 44.630 41.900 ;
        RECT 44.830 41.050 45.680 41.900 ;
        RECT 40.430 40.100 41.280 40.950 ;
        RECT 41.380 40.100 42.230 40.950 ;
        RECT 42.830 40.100 43.680 40.950 ;
        RECT 43.780 40.100 44.630 40.950 ;
        RECT 44.830 40.100 45.680 40.950 ;
        RECT 45.780 40.100 46.630 40.950 ;
        RECT 47.230 40.100 48.080 40.950 ;
        RECT 48.180 40.100 49.030 40.950 ;
        RECT 40.430 39.050 41.280 39.900 ;
        RECT 41.380 39.050 42.230 39.900 ;
        RECT 42.830 39.050 43.680 39.900 ;
        RECT 43.780 39.050 44.630 39.900 ;
        RECT 44.830 39.050 45.680 39.900 ;
        RECT 45.780 39.050 46.630 39.900 ;
        RECT 47.230 39.050 48.080 39.900 ;
        RECT 48.180 39.050 49.030 39.900 ;
        RECT 43.780 38.100 44.630 38.950 ;
        RECT 44.830 38.100 45.680 38.950 ;
        RECT 63.780 41.050 64.630 41.900 ;
        RECT 64.830 41.050 65.680 41.900 ;
        RECT 60.430 40.100 61.280 40.950 ;
        RECT 61.380 40.100 62.230 40.950 ;
        RECT 62.830 40.100 63.680 40.950 ;
        RECT 63.780 40.100 64.630 40.950 ;
        RECT 64.830 40.100 65.680 40.950 ;
        RECT 65.780 40.100 66.630 40.950 ;
        RECT 67.230 40.100 68.080 40.950 ;
        RECT 68.180 40.100 69.030 40.950 ;
        RECT 60.430 39.050 61.280 39.900 ;
        RECT 61.380 39.050 62.230 39.900 ;
        RECT 62.830 39.050 63.680 39.900 ;
        RECT 63.780 39.050 64.630 39.900 ;
        RECT 64.830 39.050 65.680 39.900 ;
        RECT 65.780 39.050 66.630 39.900 ;
        RECT 67.230 39.050 68.080 39.900 ;
        RECT 68.180 39.050 69.030 39.900 ;
        RECT 63.780 38.100 64.630 38.950 ;
        RECT 64.830 38.100 65.680 38.950 ;
        RECT 83.780 41.050 84.630 41.900 ;
        RECT 84.830 41.050 85.680 41.900 ;
        RECT 80.430 40.100 81.280 40.950 ;
        RECT 81.380 40.100 82.230 40.950 ;
        RECT 82.830 40.100 83.680 40.950 ;
        RECT 83.780 40.100 84.630 40.950 ;
        RECT 84.830 40.100 85.680 40.950 ;
        RECT 85.780 40.100 86.630 40.950 ;
        RECT 87.230 40.100 88.080 40.950 ;
        RECT 88.180 40.100 89.030 40.950 ;
        RECT 80.430 39.050 81.280 39.900 ;
        RECT 81.380 39.050 82.230 39.900 ;
        RECT 82.830 39.050 83.680 39.900 ;
        RECT 83.780 39.050 84.630 39.900 ;
        RECT 84.830 39.050 85.680 39.900 ;
        RECT 85.780 39.050 86.630 39.900 ;
        RECT 87.230 39.050 88.080 39.900 ;
        RECT 88.180 39.050 89.030 39.900 ;
        RECT 83.780 38.100 84.630 38.950 ;
        RECT 84.830 38.100 85.680 38.950 ;
        RECT 103.780 41.050 104.630 41.900 ;
        RECT 104.830 41.050 105.680 41.900 ;
        RECT 100.430 40.100 101.280 40.950 ;
        RECT 101.380 40.100 102.230 40.950 ;
        RECT 102.830 40.100 103.680 40.950 ;
        RECT 103.780 40.100 104.630 40.950 ;
        RECT 104.830 40.100 105.680 40.950 ;
        RECT 105.780 40.100 106.630 40.950 ;
        RECT 107.230 40.100 108.080 40.950 ;
        RECT 108.180 40.100 109.030 40.950 ;
        RECT 100.430 39.050 101.280 39.900 ;
        RECT 101.380 39.050 102.230 39.900 ;
        RECT 102.830 39.050 103.680 39.900 ;
        RECT 103.780 39.050 104.630 39.900 ;
        RECT 104.830 39.050 105.680 39.900 ;
        RECT 105.780 39.050 106.630 39.900 ;
        RECT 107.230 39.050 108.080 39.900 ;
        RECT 108.180 39.050 109.030 39.900 ;
        RECT 103.780 38.100 104.630 38.950 ;
        RECT 104.830 38.100 105.680 38.950 ;
        RECT 123.780 41.050 124.630 41.900 ;
        RECT 125.340 42.590 125.700 42.970 ;
        RECT 125.970 42.590 126.330 42.970 ;
        RECT 126.570 42.590 126.930 42.970 ;
        RECT 125.340 42.000 125.700 42.380 ;
        RECT 125.970 42.000 126.330 42.380 ;
        RECT 126.570 42.000 126.930 42.380 ;
        RECT 120.430 40.100 121.280 40.950 ;
        RECT 121.380 40.100 122.230 40.950 ;
        RECT 122.830 40.100 123.680 40.950 ;
        RECT 123.780 40.100 124.630 40.950 ;
        RECT 120.430 39.050 121.280 39.900 ;
        RECT 121.380 39.050 122.230 39.900 ;
        RECT 122.830 39.050 123.680 39.900 ;
        RECT 123.780 39.050 124.630 39.900 ;
        RECT 123.780 38.100 124.630 38.950 ;
        RECT 2.515 37.115 2.875 37.495 ;
        RECT 3.145 37.115 3.505 37.495 ;
        RECT 3.745 37.115 4.105 37.495 ;
        RECT 2.515 36.525 2.875 36.905 ;
        RECT 3.145 36.525 3.505 36.905 ;
        RECT 3.745 36.525 4.105 36.905 ;
        RECT 4.830 36.650 5.680 37.500 ;
        RECT 23.780 36.650 24.630 37.500 ;
        RECT 24.830 36.650 25.680 37.500 ;
        RECT 43.780 36.650 44.630 37.500 ;
        RECT 44.830 36.650 45.680 37.500 ;
        RECT 63.780 36.650 64.630 37.500 ;
        RECT 64.830 36.650 65.680 37.500 ;
        RECT 83.780 36.650 84.630 37.500 ;
        RECT 84.830 36.650 85.680 37.500 ;
        RECT 103.780 36.650 104.630 37.500 ;
        RECT 104.830 36.650 105.680 37.500 ;
        RECT 123.780 36.650 124.630 37.500 ;
        RECT 4.830 35.700 5.680 36.550 ;
        RECT 23.780 35.700 24.630 36.550 ;
        RECT 24.830 35.700 25.680 36.550 ;
        RECT 43.780 35.700 44.630 36.550 ;
        RECT 44.830 35.700 45.680 36.550 ;
        RECT 63.780 35.700 64.630 36.550 ;
        RECT 64.830 35.700 65.680 36.550 ;
        RECT 83.780 35.700 84.630 36.550 ;
        RECT 84.830 35.700 85.680 36.550 ;
        RECT 103.780 35.700 104.630 36.550 ;
        RECT 104.830 35.700 105.680 36.550 ;
        RECT 123.780 35.700 124.630 36.550 ;
        RECT 125.340 36.805 125.700 37.185 ;
        RECT 125.970 36.805 126.330 37.185 ;
        RECT 126.570 36.805 126.930 37.185 ;
        RECT 125.340 36.215 125.700 36.595 ;
        RECT 125.970 36.215 126.330 36.595 ;
        RECT 126.570 36.215 126.930 36.595 ;
        RECT 2.520 34.925 2.880 35.305 ;
        RECT 3.130 34.925 3.490 35.305 ;
        RECT 3.760 34.925 4.120 35.305 ;
        RECT 2.520 34.190 2.880 34.570 ;
        RECT 3.130 34.190 3.490 34.570 ;
        RECT 3.760 34.190 4.120 34.570 ;
        RECT 2.520 33.505 2.880 33.885 ;
        RECT 3.130 33.505 3.490 33.885 ;
        RECT 3.760 33.505 4.120 33.885 ;
        RECT 2.520 26.115 2.880 26.495 ;
        RECT 3.130 26.115 3.490 26.495 ;
        RECT 3.760 26.115 4.120 26.495 ;
        RECT 2.520 25.380 2.880 25.760 ;
        RECT 3.130 25.380 3.490 25.760 ;
        RECT 3.760 25.380 4.120 25.760 ;
        RECT 2.520 24.695 2.880 25.075 ;
        RECT 3.130 24.695 3.490 25.075 ;
        RECT 3.760 24.695 4.120 25.075 ;
        RECT 4.830 23.450 5.680 24.300 ;
        RECT 23.780 23.450 24.630 24.300 ;
        RECT 24.830 23.450 25.680 24.300 ;
        RECT 43.780 23.450 44.630 24.300 ;
        RECT 44.830 23.450 45.680 24.300 ;
        RECT 63.780 23.450 64.630 24.300 ;
        RECT 64.830 23.450 65.680 24.300 ;
        RECT 83.780 23.450 84.630 24.300 ;
        RECT 84.830 23.450 85.680 24.300 ;
        RECT 103.780 23.450 104.630 24.300 ;
        RECT 104.830 23.450 105.680 24.300 ;
        RECT 123.780 23.450 124.630 24.300 ;
        RECT 2.515 22.815 2.875 23.195 ;
        RECT 3.145 22.815 3.505 23.195 ;
        RECT 3.745 22.815 4.105 23.195 ;
        RECT 2.515 22.225 2.875 22.605 ;
        RECT 3.145 22.225 3.505 22.605 ;
        RECT 3.745 22.225 4.105 22.605 ;
        RECT 4.830 22.500 5.680 23.350 ;
        RECT 23.780 22.500 24.630 23.350 ;
        RECT 24.830 22.500 25.680 23.350 ;
        RECT 43.780 22.500 44.630 23.350 ;
        RECT 44.830 22.500 45.680 23.350 ;
        RECT 63.780 22.500 64.630 23.350 ;
        RECT 64.830 22.500 65.680 23.350 ;
        RECT 83.780 22.500 84.630 23.350 ;
        RECT 84.830 22.500 85.680 23.350 ;
        RECT 103.780 22.500 104.630 23.350 ;
        RECT 104.830 22.500 105.680 23.350 ;
        RECT 123.780 22.500 124.630 23.350 ;
        RECT 4.830 21.050 5.680 21.900 ;
        RECT 4.830 20.100 5.680 20.950 ;
        RECT 5.780 20.100 6.630 20.950 ;
        RECT 7.230 20.100 8.080 20.950 ;
        RECT 8.180 20.100 9.030 20.950 ;
        RECT 4.830 19.050 5.680 19.900 ;
        RECT 5.780 19.050 6.630 19.900 ;
        RECT 7.230 19.050 8.080 19.900 ;
        RECT 8.180 19.050 9.030 19.900 ;
        RECT 4.830 18.100 5.680 18.950 ;
        RECT 23.780 21.050 24.630 21.900 ;
        RECT 24.830 21.050 25.680 21.900 ;
        RECT 20.430 20.100 21.280 20.950 ;
        RECT 21.380 20.100 22.230 20.950 ;
        RECT 22.830 20.100 23.680 20.950 ;
        RECT 23.780 20.100 24.630 20.950 ;
        RECT 24.830 20.100 25.680 20.950 ;
        RECT 25.780 20.100 26.630 20.950 ;
        RECT 27.230 20.100 28.080 20.950 ;
        RECT 28.180 20.100 29.030 20.950 ;
        RECT 20.430 19.050 21.280 19.900 ;
        RECT 21.380 19.050 22.230 19.900 ;
        RECT 22.830 19.050 23.680 19.900 ;
        RECT 23.780 19.050 24.630 19.900 ;
        RECT 24.830 19.050 25.680 19.900 ;
        RECT 25.780 19.050 26.630 19.900 ;
        RECT 27.230 19.050 28.080 19.900 ;
        RECT 28.180 19.050 29.030 19.900 ;
        RECT 23.780 18.100 24.630 18.950 ;
        RECT 24.830 18.100 25.680 18.950 ;
        RECT 43.780 21.050 44.630 21.900 ;
        RECT 44.830 21.050 45.680 21.900 ;
        RECT 40.430 20.100 41.280 20.950 ;
        RECT 41.380 20.100 42.230 20.950 ;
        RECT 42.830 20.100 43.680 20.950 ;
        RECT 43.780 20.100 44.630 20.950 ;
        RECT 44.830 20.100 45.680 20.950 ;
        RECT 45.780 20.100 46.630 20.950 ;
        RECT 47.230 20.100 48.080 20.950 ;
        RECT 48.180 20.100 49.030 20.950 ;
        RECT 40.430 19.050 41.280 19.900 ;
        RECT 41.380 19.050 42.230 19.900 ;
        RECT 42.830 19.050 43.680 19.900 ;
        RECT 43.780 19.050 44.630 19.900 ;
        RECT 44.830 19.050 45.680 19.900 ;
        RECT 45.780 19.050 46.630 19.900 ;
        RECT 47.230 19.050 48.080 19.900 ;
        RECT 48.180 19.050 49.030 19.900 ;
        RECT 43.780 18.100 44.630 18.950 ;
        RECT 44.830 18.100 45.680 18.950 ;
        RECT 63.780 21.050 64.630 21.900 ;
        RECT 64.830 21.050 65.680 21.900 ;
        RECT 60.430 20.100 61.280 20.950 ;
        RECT 61.380 20.100 62.230 20.950 ;
        RECT 62.830 20.100 63.680 20.950 ;
        RECT 63.780 20.100 64.630 20.950 ;
        RECT 64.830 20.100 65.680 20.950 ;
        RECT 65.780 20.100 66.630 20.950 ;
        RECT 67.230 20.100 68.080 20.950 ;
        RECT 68.180 20.100 69.030 20.950 ;
        RECT 60.430 19.050 61.280 19.900 ;
        RECT 61.380 19.050 62.230 19.900 ;
        RECT 62.830 19.050 63.680 19.900 ;
        RECT 63.780 19.050 64.630 19.900 ;
        RECT 64.830 19.050 65.680 19.900 ;
        RECT 65.780 19.050 66.630 19.900 ;
        RECT 67.230 19.050 68.080 19.900 ;
        RECT 68.180 19.050 69.030 19.900 ;
        RECT 63.780 18.100 64.630 18.950 ;
        RECT 64.830 18.100 65.680 18.950 ;
        RECT 83.780 21.050 84.630 21.900 ;
        RECT 84.830 21.050 85.680 21.900 ;
        RECT 80.430 20.100 81.280 20.950 ;
        RECT 81.380 20.100 82.230 20.950 ;
        RECT 82.830 20.100 83.680 20.950 ;
        RECT 83.780 20.100 84.630 20.950 ;
        RECT 84.830 20.100 85.680 20.950 ;
        RECT 85.780 20.100 86.630 20.950 ;
        RECT 87.230 20.100 88.080 20.950 ;
        RECT 88.180 20.100 89.030 20.950 ;
        RECT 80.430 19.050 81.280 19.900 ;
        RECT 81.380 19.050 82.230 19.900 ;
        RECT 82.830 19.050 83.680 19.900 ;
        RECT 83.780 19.050 84.630 19.900 ;
        RECT 84.830 19.050 85.680 19.900 ;
        RECT 85.780 19.050 86.630 19.900 ;
        RECT 87.230 19.050 88.080 19.900 ;
        RECT 88.180 19.050 89.030 19.900 ;
        RECT 83.780 18.100 84.630 18.950 ;
        RECT 84.830 18.100 85.680 18.950 ;
        RECT 103.780 21.050 104.630 21.900 ;
        RECT 104.830 21.050 105.680 21.900 ;
        RECT 100.430 20.100 101.280 20.950 ;
        RECT 101.380 20.100 102.230 20.950 ;
        RECT 102.830 20.100 103.680 20.950 ;
        RECT 103.780 20.100 104.630 20.950 ;
        RECT 104.830 20.100 105.680 20.950 ;
        RECT 105.780 20.100 106.630 20.950 ;
        RECT 107.230 20.100 108.080 20.950 ;
        RECT 108.180 20.100 109.030 20.950 ;
        RECT 100.430 19.050 101.280 19.900 ;
        RECT 101.380 19.050 102.230 19.900 ;
        RECT 102.830 19.050 103.680 19.900 ;
        RECT 103.780 19.050 104.630 19.900 ;
        RECT 104.830 19.050 105.680 19.900 ;
        RECT 105.780 19.050 106.630 19.900 ;
        RECT 107.230 19.050 108.080 19.900 ;
        RECT 108.180 19.050 109.030 19.900 ;
        RECT 103.780 18.100 104.630 18.950 ;
        RECT 104.830 18.100 105.680 18.950 ;
        RECT 123.780 21.050 124.630 21.900 ;
        RECT 125.340 22.590 125.700 22.970 ;
        RECT 125.970 22.590 126.330 22.970 ;
        RECT 126.570 22.590 126.930 22.970 ;
        RECT 125.340 22.000 125.700 22.380 ;
        RECT 125.970 22.000 126.330 22.380 ;
        RECT 126.570 22.000 126.930 22.380 ;
        RECT 120.430 20.100 121.280 20.950 ;
        RECT 121.380 20.100 122.230 20.950 ;
        RECT 122.830 20.100 123.680 20.950 ;
        RECT 123.780 20.100 124.630 20.950 ;
        RECT 120.430 19.050 121.280 19.900 ;
        RECT 121.380 19.050 122.230 19.900 ;
        RECT 122.830 19.050 123.680 19.900 ;
        RECT 123.780 19.050 124.630 19.900 ;
        RECT 123.780 18.100 124.630 18.950 ;
        RECT 2.515 17.260 2.875 17.640 ;
        RECT 3.145 17.260 3.505 17.640 ;
        RECT 3.745 17.260 4.105 17.640 ;
        RECT 2.515 16.670 2.875 17.050 ;
        RECT 3.145 16.670 3.505 17.050 ;
        RECT 3.745 16.670 4.105 17.050 ;
        RECT 4.830 16.650 5.680 17.500 ;
        RECT 23.780 16.650 24.630 17.500 ;
        RECT 24.830 16.650 25.680 17.500 ;
        RECT 43.780 16.650 44.630 17.500 ;
        RECT 44.830 16.650 45.680 17.500 ;
        RECT 63.780 16.650 64.630 17.500 ;
        RECT 64.830 16.650 65.680 17.500 ;
        RECT 83.780 16.650 84.630 17.500 ;
        RECT 84.830 16.650 85.680 17.500 ;
        RECT 103.780 16.650 104.630 17.500 ;
        RECT 104.830 16.650 105.680 17.500 ;
        RECT 123.780 16.650 124.630 17.500 ;
        RECT 4.830 15.700 5.680 16.550 ;
        RECT 23.780 15.700 24.630 16.550 ;
        RECT 24.830 15.700 25.680 16.550 ;
        RECT 43.780 15.700 44.630 16.550 ;
        RECT 44.830 15.700 45.680 16.550 ;
        RECT 63.780 15.700 64.630 16.550 ;
        RECT 64.830 15.700 65.680 16.550 ;
        RECT 83.780 15.700 84.630 16.550 ;
        RECT 84.830 15.700 85.680 16.550 ;
        RECT 103.780 15.700 104.630 16.550 ;
        RECT 104.830 15.700 105.680 16.550 ;
        RECT 123.780 15.700 124.630 16.550 ;
        RECT 125.340 16.805 125.700 17.185 ;
        RECT 125.970 16.805 126.330 17.185 ;
        RECT 126.570 16.805 126.930 17.185 ;
        RECT 125.340 16.215 125.700 16.595 ;
        RECT 125.970 16.215 126.330 16.595 ;
        RECT 126.570 16.215 126.930 16.595 ;
        RECT 2.520 14.925 2.880 15.305 ;
        RECT 3.130 14.925 3.490 15.305 ;
        RECT 3.760 14.925 4.120 15.305 ;
        RECT 2.520 14.190 2.880 14.570 ;
        RECT 3.130 14.190 3.490 14.570 ;
        RECT 3.760 14.190 4.120 14.570 ;
        RECT 2.520 13.505 2.880 13.885 ;
        RECT 3.130 13.505 3.490 13.885 ;
        RECT 3.760 13.505 4.120 13.885 ;
        RECT 2.520 6.120 2.880 6.500 ;
        RECT 3.130 6.120 3.490 6.500 ;
        RECT 3.760 6.120 4.120 6.500 ;
        RECT 2.520 5.385 2.880 5.765 ;
        RECT 3.130 5.385 3.490 5.765 ;
        RECT 3.760 5.385 4.120 5.765 ;
        RECT 2.520 4.700 2.880 5.080 ;
        RECT 3.130 4.700 3.490 5.080 ;
        RECT 3.760 4.700 4.120 5.080 ;
        RECT 2.515 3.145 2.875 3.525 ;
        RECT 3.145 3.145 3.505 3.525 ;
        RECT 3.745 3.145 4.105 3.525 ;
        RECT 2.515 2.555 2.875 2.935 ;
        RECT 3.145 2.555 3.505 2.935 ;
        RECT 3.745 2.555 4.105 2.935 ;
        RECT 4.830 3.450 5.680 4.300 ;
        RECT 23.780 3.450 24.630 4.300 ;
        RECT 24.830 3.450 25.680 4.300 ;
        RECT 43.780 3.450 44.630 4.300 ;
        RECT 44.830 3.450 45.680 4.300 ;
        RECT 63.780 3.450 64.630 4.300 ;
        RECT 64.830 3.450 65.680 4.300 ;
        RECT 83.780 3.450 84.630 4.300 ;
        RECT 84.830 3.450 85.680 4.300 ;
        RECT 103.780 3.450 104.630 4.300 ;
        RECT 104.830 3.450 105.680 4.300 ;
        RECT 123.780 3.450 124.630 4.300 ;
        RECT 4.830 2.500 5.680 3.350 ;
        RECT 23.780 2.500 24.630 3.350 ;
        RECT 24.830 2.500 25.680 3.350 ;
        RECT 43.780 2.500 44.630 3.350 ;
        RECT 44.830 2.500 45.680 3.350 ;
        RECT 63.780 2.500 64.630 3.350 ;
        RECT 64.830 2.500 65.680 3.350 ;
        RECT 83.780 2.500 84.630 3.350 ;
        RECT 84.830 2.500 85.680 3.350 ;
        RECT 103.780 2.500 104.630 3.350 ;
        RECT 104.830 2.500 105.680 3.350 ;
        RECT 123.780 2.500 124.630 3.350 ;
        RECT 4.830 1.050 5.680 1.900 ;
        RECT 4.830 0.100 5.680 0.950 ;
        RECT 5.780 0.100 6.630 0.950 ;
        RECT 7.230 0.100 8.080 0.950 ;
        RECT 8.180 0.100 9.030 0.950 ;
        RECT 23.780 1.050 24.630 1.900 ;
        RECT 24.830 1.050 25.680 1.900 ;
        RECT 20.430 0.100 21.280 0.950 ;
        RECT 21.380 0.100 22.230 0.950 ;
        RECT 22.830 0.100 23.680 0.950 ;
        RECT 23.780 0.100 24.630 0.950 ;
        RECT 24.830 0.100 25.680 0.950 ;
        RECT 25.780 0.100 26.630 0.950 ;
        RECT 27.230 0.100 28.080 0.950 ;
        RECT 28.180 0.100 29.030 0.950 ;
        RECT 43.780 1.050 44.630 1.900 ;
        RECT 44.830 1.050 45.680 1.900 ;
        RECT 40.430 0.100 41.280 0.950 ;
        RECT 41.380 0.100 42.230 0.950 ;
        RECT 42.830 0.100 43.680 0.950 ;
        RECT 43.780 0.100 44.630 0.950 ;
        RECT 44.830 0.100 45.680 0.950 ;
        RECT 45.780 0.100 46.630 0.950 ;
        RECT 47.230 0.100 48.080 0.950 ;
        RECT 48.180 0.100 49.030 0.950 ;
        RECT 63.780 1.050 64.630 1.900 ;
        RECT 64.830 1.050 65.680 1.900 ;
        RECT 60.430 0.100 61.280 0.950 ;
        RECT 61.380 0.100 62.230 0.950 ;
        RECT 62.830 0.100 63.680 0.950 ;
        RECT 63.780 0.100 64.630 0.950 ;
        RECT 64.830 0.100 65.680 0.950 ;
        RECT 65.780 0.100 66.630 0.950 ;
        RECT 67.230 0.100 68.080 0.950 ;
        RECT 68.180 0.100 69.030 0.950 ;
        RECT 83.780 1.050 84.630 1.900 ;
        RECT 84.830 1.050 85.680 1.900 ;
        RECT 80.430 0.100 81.280 0.950 ;
        RECT 81.380 0.100 82.230 0.950 ;
        RECT 82.830 0.100 83.680 0.950 ;
        RECT 83.780 0.100 84.630 0.950 ;
        RECT 84.830 0.100 85.680 0.950 ;
        RECT 85.780 0.100 86.630 0.950 ;
        RECT 87.230 0.100 88.080 0.950 ;
        RECT 88.180 0.100 89.030 0.950 ;
        RECT 103.780 1.050 104.630 1.900 ;
        RECT 104.830 1.050 105.680 1.900 ;
        RECT 100.430 0.100 101.280 0.950 ;
        RECT 101.380 0.100 102.230 0.950 ;
        RECT 102.830 0.100 103.680 0.950 ;
        RECT 103.780 0.100 104.630 0.950 ;
        RECT 104.830 0.100 105.680 0.950 ;
        RECT 105.780 0.100 106.630 0.950 ;
        RECT 107.230 0.100 108.080 0.950 ;
        RECT 108.180 0.100 109.030 0.950 ;
        RECT 123.780 1.050 124.630 1.900 ;
        RECT 125.340 2.590 125.700 2.970 ;
        RECT 125.970 2.590 126.330 2.970 ;
        RECT 126.570 2.590 126.930 2.970 ;
        RECT 125.340 2.000 125.700 2.380 ;
        RECT 125.970 2.000 126.330 2.380 ;
        RECT 126.570 2.000 126.930 2.380 ;
        RECT 120.430 0.100 121.280 0.950 ;
        RECT 121.380 0.100 122.230 0.950 ;
        RECT 122.830 0.100 123.680 0.950 ;
        RECT 123.780 0.100 124.630 0.950 ;
      LAYER met4 ;
        RECT 2.315 337.385 4.315 340.000 ;
        RECT 125.140 337.585 127.140 340.000 ;
        RECT 2.315 336.110 4.320 337.385 ;
        RECT 125.130 336.310 127.140 337.585 ;
        RECT 2.315 324.020 4.315 336.110 ;
        RECT 2.315 322.745 4.320 324.020 ;
        RECT 2.315 317.375 4.315 322.745 ;
        RECT 125.140 317.585 127.140 336.310 ;
        RECT 2.315 316.100 4.320 317.375 ;
        RECT 125.130 316.310 127.140 317.585 ;
        RECT 2.315 303.675 4.315 316.100 ;
        RECT 2.315 302.400 4.320 303.675 ;
        RECT 2.315 297.785 4.315 302.400 ;
        RECT 2.315 296.510 4.320 297.785 ;
        RECT 125.140 297.585 127.140 316.310 ;
        RECT 2.315 295.545 4.315 296.510 ;
        RECT 125.130 296.310 127.140 297.585 ;
        RECT 2.315 293.250 4.320 295.545 ;
        RECT 2.315 283.545 4.315 293.250 ;
        RECT 2.315 282.270 4.330 283.545 ;
        RECT 2.315 277.530 4.315 282.270 ;
        RECT 125.140 277.855 127.140 296.310 ;
        RECT 2.315 276.255 4.320 277.530 ;
        RECT 125.135 276.580 127.140 277.855 ;
        RECT 2.315 275.545 4.315 276.255 ;
        RECT 2.315 273.250 4.320 275.545 ;
        RECT 2.315 263.645 4.315 273.250 ;
        RECT 2.315 262.370 4.320 263.645 ;
        RECT 2.315 257.610 4.315 262.370 ;
        RECT 2.315 256.335 4.330 257.610 ;
        RECT 125.140 257.360 127.140 276.580 ;
        RECT 2.315 243.780 4.315 256.335 ;
        RECT 125.135 256.085 127.140 257.360 ;
        RECT 2.315 242.505 4.320 243.780 ;
        RECT 2.315 237.845 4.315 242.505 ;
        RECT 2.315 236.570 4.320 237.845 ;
        RECT 2.315 223.735 4.315 236.570 ;
        RECT 2.315 222.460 4.320 223.735 ;
        RECT 2.315 217.970 4.315 222.460 ;
        RECT 2.315 216.695 4.320 217.970 ;
        RECT 2.315 141.800 4.315 216.695 ;
        RECT 42.635 175.610 47.035 176.660 ;
        RECT 58.235 175.610 67.035 176.660 ;
        RECT 78.235 175.610 87.035 176.660 ;
        RECT 98.235 175.610 107.035 176.660 ;
        RECT 118.235 175.610 122.635 176.660 ;
        RECT 42.635 172.260 43.685 175.610 ;
        RECT 61.585 172.260 63.685 175.610 ;
        RECT 81.585 172.260 83.685 175.610 ;
        RECT 101.585 172.260 103.685 175.610 ;
        RECT 121.585 174.990 122.635 175.610 ;
        RECT 125.140 174.990 127.140 256.085 ;
        RECT 121.585 173.715 127.140 174.990 ;
        RECT 121.585 172.260 122.635 173.715 ;
        RECT 42.635 157.710 43.685 161.060 ;
        RECT 61.585 157.710 63.685 161.060 ;
        RECT 81.585 157.710 83.685 161.060 ;
        RECT 101.585 157.710 103.685 161.060 ;
        RECT 121.585 159.715 122.635 161.060 ;
        RECT 125.140 159.715 127.140 173.715 ;
        RECT 121.585 158.440 127.140 159.715 ;
        RECT 121.585 157.710 122.635 158.440 ;
        RECT 42.635 156.660 47.035 157.710 ;
        RECT 58.235 156.660 67.035 157.710 ;
        RECT 78.235 156.660 87.035 157.710 ;
        RECT 98.235 156.660 107.035 157.710 ;
        RECT 118.235 156.660 122.635 157.710 ;
        RECT 125.140 141.800 127.140 158.440 ;
        RECT 2.315 140.360 4.330 141.800 ;
        RECT 125.125 140.360 127.140 141.800 ;
        RECT 2.315 140.000 4.315 140.360 ;
        RECT 2.315 138.950 9.130 140.000 ;
        RECT 20.330 138.950 29.130 140.000 ;
        RECT 40.330 138.950 49.130 140.000 ;
        RECT 60.330 138.950 69.130 140.000 ;
        RECT 80.330 138.950 89.130 140.000 ;
        RECT 100.330 138.950 109.130 140.000 ;
        RECT 120.330 138.950 124.730 140.000 ;
        RECT 2.315 138.800 5.780 138.950 ;
        RECT 2.315 124.425 4.315 138.800 ;
        RECT 4.730 135.600 5.780 138.800 ;
        RECT 23.680 135.600 25.780 138.950 ;
        RECT 43.680 135.600 45.780 138.950 ;
        RECT 63.680 135.600 65.780 138.950 ;
        RECT 83.680 135.600 85.780 138.950 ;
        RECT 103.680 135.600 105.780 138.950 ;
        RECT 123.680 135.600 124.730 138.950 ;
        RECT 2.315 123.340 4.310 124.425 ;
        RECT 4.720 123.405 5.780 124.400 ;
        RECT 2.315 121.190 4.315 123.340 ;
        RECT 4.730 121.190 5.780 123.405 ;
        RECT 2.315 121.050 5.780 121.190 ;
        RECT 23.680 121.050 25.780 124.400 ;
        RECT 43.680 121.050 45.780 124.400 ;
        RECT 63.680 121.050 65.780 124.400 ;
        RECT 83.680 121.050 85.780 124.400 ;
        RECT 103.680 121.050 105.780 124.400 ;
        RECT 123.680 121.160 124.730 124.400 ;
        RECT 125.140 121.160 127.140 140.360 ;
        RECT 123.680 121.050 127.140 121.160 ;
        RECT 2.315 121.045 9.130 121.050 ;
        RECT 2.310 119.895 9.130 121.045 ;
        RECT 2.315 118.950 9.130 119.895 ;
        RECT 20.330 118.950 29.130 121.050 ;
        RECT 40.330 118.950 49.130 121.050 ;
        RECT 60.330 118.950 69.130 121.050 ;
        RECT 80.330 118.950 89.130 121.050 ;
        RECT 100.330 118.950 109.130 121.050 ;
        RECT 120.330 118.950 127.140 121.050 ;
        RECT 2.315 118.800 5.780 118.950 ;
        RECT 2.315 103.255 4.315 118.800 ;
        RECT 4.730 115.600 5.780 118.800 ;
        RECT 23.680 115.600 25.780 118.950 ;
        RECT 43.680 115.600 45.780 118.950 ;
        RECT 63.680 115.600 65.780 118.950 ;
        RECT 83.680 115.600 85.780 118.950 ;
        RECT 103.680 115.600 105.780 118.950 ;
        RECT 123.680 118.830 127.140 118.950 ;
        RECT 123.680 115.600 124.730 118.830 ;
        RECT 125.140 117.335 127.140 118.830 ;
        RECT 125.135 116.060 127.140 117.335 ;
        RECT 2.315 101.980 4.320 103.255 ;
        RECT 2.315 101.195 4.315 101.980 ;
        RECT 4.730 101.195 5.780 104.400 ;
        RECT 2.315 101.050 5.780 101.195 ;
        RECT 23.680 101.050 25.780 104.400 ;
        RECT 43.680 101.050 45.780 104.400 ;
        RECT 63.680 101.050 65.780 104.400 ;
        RECT 83.680 101.050 85.780 104.400 ;
        RECT 103.680 101.050 105.780 104.400 ;
        RECT 123.680 101.160 124.730 104.400 ;
        RECT 125.140 101.160 127.140 116.060 ;
        RECT 123.680 101.050 127.140 101.160 ;
        RECT 2.315 98.950 9.130 101.050 ;
        RECT 20.330 98.950 29.130 101.050 ;
        RECT 40.330 98.950 49.130 101.050 ;
        RECT 60.330 98.950 69.130 101.050 ;
        RECT 80.330 98.950 89.130 101.050 ;
        RECT 100.330 98.950 109.130 101.050 ;
        RECT 120.330 98.950 127.140 101.050 ;
        RECT 2.315 98.795 5.780 98.950 ;
        RECT 2.315 97.845 4.315 98.795 ;
        RECT 2.315 96.570 4.320 97.845 ;
        RECT 2.315 83.470 4.315 96.570 ;
        RECT 4.730 95.600 5.780 98.795 ;
        RECT 23.680 95.600 25.780 98.950 ;
        RECT 43.680 95.600 45.780 98.950 ;
        RECT 63.680 95.600 65.780 98.950 ;
        RECT 83.680 95.600 85.780 98.950 ;
        RECT 103.680 95.600 105.780 98.950 ;
        RECT 123.680 98.835 127.140 98.950 ;
        RECT 123.680 95.600 124.730 98.835 ;
        RECT 2.315 82.195 4.320 83.470 ;
        RECT 2.315 81.200 4.315 82.195 ;
        RECT 4.730 81.200 5.780 84.400 ;
        RECT 2.315 81.050 5.780 81.200 ;
        RECT 23.680 81.050 25.780 84.400 ;
        RECT 43.680 81.050 45.780 84.400 ;
        RECT 63.680 81.050 65.780 84.400 ;
        RECT 83.680 81.050 85.780 84.400 ;
        RECT 103.680 81.050 105.780 84.400 ;
        RECT 123.680 81.165 124.730 84.400 ;
        RECT 125.140 83.040 127.140 98.835 ;
        RECT 125.135 81.765 127.140 83.040 ;
        RECT 125.140 81.165 127.140 81.765 ;
        RECT 123.680 81.050 127.140 81.165 ;
        RECT 2.315 78.950 9.130 81.050 ;
        RECT 20.330 78.950 29.130 81.050 ;
        RECT 40.330 78.950 49.130 81.050 ;
        RECT 60.330 78.950 69.130 81.050 ;
        RECT 80.330 78.950 89.130 81.050 ;
        RECT 100.330 78.950 109.130 81.050 ;
        RECT 120.330 78.950 127.140 81.050 ;
        RECT 2.315 78.800 5.780 78.950 ;
        RECT 2.315 77.965 4.315 78.800 ;
        RECT 2.315 76.690 4.320 77.965 ;
        RECT 2.315 63.635 4.315 76.690 ;
        RECT 4.730 75.600 5.780 78.800 ;
        RECT 23.680 75.600 25.780 78.950 ;
        RECT 43.680 75.600 45.780 78.950 ;
        RECT 63.680 75.600 65.780 78.950 ;
        RECT 83.680 75.600 85.780 78.950 ;
        RECT 103.680 75.600 105.780 78.950 ;
        RECT 123.680 78.840 127.140 78.950 ;
        RECT 123.680 75.600 124.730 78.840 ;
        RECT 125.140 77.185 127.140 78.840 ;
        RECT 125.135 75.910 127.140 77.185 ;
        RECT 2.315 62.360 4.325 63.635 ;
        RECT 2.315 61.195 4.315 62.360 ;
        RECT 4.730 61.195 5.780 64.400 ;
        RECT 2.315 61.050 5.780 61.195 ;
        RECT 23.680 61.050 25.780 64.400 ;
        RECT 43.680 61.050 45.780 64.400 ;
        RECT 63.680 61.050 65.780 64.400 ;
        RECT 83.680 61.050 85.780 64.400 ;
        RECT 103.680 61.050 105.780 64.400 ;
        RECT 123.680 61.160 124.730 64.400 ;
        RECT 125.140 63.380 127.140 75.910 ;
        RECT 125.135 62.105 127.140 63.380 ;
        RECT 125.140 61.160 127.140 62.105 ;
        RECT 123.680 61.050 127.140 61.160 ;
        RECT 2.315 58.950 9.130 61.050 ;
        RECT 20.330 58.950 29.130 61.050 ;
        RECT 40.330 58.950 49.130 61.050 ;
        RECT 60.330 58.950 69.130 61.050 ;
        RECT 80.330 58.950 89.130 61.050 ;
        RECT 100.330 58.950 109.130 61.050 ;
        RECT 120.330 58.950 127.140 61.050 ;
        RECT 2.315 58.795 5.780 58.950 ;
        RECT 2.315 57.555 4.315 58.795 ;
        RECT 2.315 56.280 4.330 57.555 ;
        RECT 2.315 43.230 4.315 56.280 ;
        RECT 4.730 55.600 5.780 58.795 ;
        RECT 23.680 55.600 25.780 58.950 ;
        RECT 43.680 55.600 45.780 58.950 ;
        RECT 63.680 55.600 65.780 58.950 ;
        RECT 83.680 55.600 85.780 58.950 ;
        RECT 103.680 55.600 105.780 58.950 ;
        RECT 123.680 58.830 127.140 58.950 ;
        RECT 123.680 55.600 124.730 58.830 ;
        RECT 125.140 57.310 127.140 58.830 ;
        RECT 125.135 56.035 127.140 57.310 ;
        RECT 2.315 41.955 4.320 43.230 ;
        RECT 2.315 41.190 4.315 41.955 ;
        RECT 4.730 41.190 5.780 44.400 ;
        RECT 2.315 41.050 5.780 41.190 ;
        RECT 23.680 41.050 25.780 44.400 ;
        RECT 43.680 41.050 45.780 44.400 ;
        RECT 63.680 41.050 65.780 44.400 ;
        RECT 83.680 41.050 85.780 44.400 ;
        RECT 103.680 41.050 105.780 44.400 ;
        RECT 123.680 41.165 124.730 44.400 ;
        RECT 125.140 41.165 127.140 56.035 ;
        RECT 123.680 41.050 127.140 41.165 ;
        RECT 2.315 38.950 9.130 41.050 ;
        RECT 20.330 38.950 29.130 41.050 ;
        RECT 40.330 38.950 49.130 41.050 ;
        RECT 60.330 38.950 69.130 41.050 ;
        RECT 80.330 38.950 89.130 41.050 ;
        RECT 100.330 38.950 109.130 41.050 ;
        RECT 120.330 38.950 127.140 41.050 ;
        RECT 2.315 38.790 5.780 38.950 ;
        RECT 2.315 37.620 4.315 38.790 ;
        RECT 2.315 36.345 4.320 37.620 ;
        RECT 2.315 21.190 4.315 36.345 ;
        RECT 4.730 35.600 5.780 38.790 ;
        RECT 23.680 35.600 25.780 38.950 ;
        RECT 43.680 35.600 45.780 38.950 ;
        RECT 63.680 35.600 65.780 38.950 ;
        RECT 83.680 35.600 85.780 38.950 ;
        RECT 103.680 35.600 105.780 38.950 ;
        RECT 123.680 38.830 127.140 38.950 ;
        RECT 123.680 35.600 124.730 38.830 ;
        RECT 125.140 37.310 127.140 38.830 ;
        RECT 125.135 36.035 127.140 37.310 ;
        RECT 4.730 21.190 5.780 24.400 ;
        RECT 2.315 21.050 5.780 21.190 ;
        RECT 23.680 21.050 25.780 24.400 ;
        RECT 43.680 21.050 45.780 24.400 ;
        RECT 63.680 21.050 65.780 24.400 ;
        RECT 83.680 21.050 85.780 24.400 ;
        RECT 103.680 21.050 105.780 24.400 ;
        RECT 123.680 21.165 124.730 24.400 ;
        RECT 125.140 21.165 127.140 36.035 ;
        RECT 123.680 21.050 127.140 21.165 ;
        RECT 2.315 18.950 9.130 21.050 ;
        RECT 20.330 18.950 29.130 21.050 ;
        RECT 40.330 18.950 49.130 21.050 ;
        RECT 60.330 18.950 69.130 21.050 ;
        RECT 80.330 18.950 89.130 21.050 ;
        RECT 100.330 18.950 109.130 21.050 ;
        RECT 120.330 18.950 127.140 21.050 ;
        RECT 2.315 18.800 5.780 18.950 ;
        RECT 2.315 3.650 4.315 18.800 ;
        RECT 4.730 15.600 5.780 18.800 ;
        RECT 23.680 15.600 25.780 18.950 ;
        RECT 43.680 15.600 45.780 18.950 ;
        RECT 63.680 15.600 65.780 18.950 ;
        RECT 83.680 15.600 85.780 18.950 ;
        RECT 103.680 15.600 105.780 18.950 ;
        RECT 123.680 18.830 127.140 18.950 ;
        RECT 123.680 15.600 124.730 18.830 ;
        RECT 125.140 17.310 127.140 18.830 ;
        RECT 125.135 16.035 127.140 17.310 ;
        RECT 2.315 2.375 4.325 3.650 ;
        RECT 2.315 1.195 4.315 2.375 ;
        RECT 4.730 1.195 5.780 4.400 ;
        RECT 2.315 1.050 5.780 1.195 ;
        RECT 23.680 1.050 25.780 4.400 ;
        RECT 43.680 1.050 45.780 4.400 ;
        RECT 63.680 1.050 65.780 4.400 ;
        RECT 83.680 1.050 85.780 4.400 ;
        RECT 103.680 1.050 105.780 4.400 ;
        RECT 123.680 1.165 124.730 4.400 ;
        RECT 125.140 1.165 127.140 16.035 ;
        RECT 123.680 1.050 127.140 1.165 ;
        RECT 2.315 0.000 9.130 1.050 ;
        RECT 20.330 0.000 29.130 1.050 ;
        RECT 40.330 0.000 49.130 1.050 ;
        RECT 60.330 0.000 69.130 1.050 ;
        RECT 80.330 0.000 89.130 1.050 ;
        RECT 100.330 0.000 109.130 1.050 ;
        RECT 120.330 0.000 127.140 1.050 ;
    END
  END VSS
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 6.695 171.085 7.615 171.345 ;
        RECT 8.530 171.090 8.865 171.340 ;
        RECT 7.365 168.700 7.695 168.940 ;
      LAYER mcon ;
        RECT 7.395 171.125 7.575 171.300 ;
        RECT 8.575 171.120 8.745 171.290 ;
        RECT 7.405 168.740 7.575 168.910 ;
      LAYER met1 ;
        RECT 7.325 171.340 7.645 171.345 ;
        RECT 7.325 171.090 8.865 171.340 ;
        RECT 7.325 171.085 7.645 171.090 ;
        RECT 7.285 168.690 7.695 168.950 ;
      LAYER via ;
        RECT 7.355 171.085 7.615 171.345 ;
        RECT 7.315 168.690 7.575 168.950 ;
      LAYER met2 ;
        RECT 7.355 171.055 7.615 171.375 ;
        RECT 7.355 168.985 7.520 171.055 ;
        RECT 7.315 168.660 7.575 168.985 ;
    END
  END clk
  PIN vcm
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 22041.599609 ;
    ANTENNADIFFAREA 1.160000 ;
    PORT
      LAYER li1 ;
        RECT 5.930 337.600 9.930 337.800 ;
        RECT 5.930 337.000 6.330 337.600 ;
        RECT 5.930 336.800 9.930 337.000 ;
        RECT 5.930 336.200 6.330 336.800 ;
        RECT 5.930 336.000 9.930 336.200 ;
        RECT 5.930 335.400 6.330 336.000 ;
        RECT 5.930 335.200 9.930 335.400 ;
        RECT 5.930 334.600 6.330 335.200 ;
        RECT 5.930 334.400 9.930 334.600 ;
        RECT 5.930 333.800 6.330 334.400 ;
        RECT 5.930 333.600 9.930 333.800 ;
        RECT 5.930 333.000 6.330 333.600 ;
        RECT 5.930 332.800 9.930 333.000 ;
        RECT 5.930 332.200 6.330 332.800 ;
        RECT 5.930 332.000 9.930 332.200 ;
        RECT 5.930 331.400 6.330 332.000 ;
        RECT 5.930 331.200 9.930 331.400 ;
        RECT 5.930 330.600 6.330 331.200 ;
        RECT 5.930 330.400 9.930 330.600 ;
        RECT 5.930 330.200 6.330 330.400 ;
        RECT 10.680 330.200 10.880 337.800 ;
        RECT 11.480 330.200 11.680 337.800 ;
        RECT 12.280 330.200 12.480 337.800 ;
        RECT 13.080 330.200 13.280 337.800 ;
        RECT 13.880 330.200 14.080 337.800 ;
        RECT 5.930 329.800 14.080 330.200 ;
        RECT 5.930 329.600 6.330 329.800 ;
        RECT 5.930 329.400 9.930 329.600 ;
        RECT 5.930 328.800 6.330 329.400 ;
        RECT 5.930 328.600 9.930 328.800 ;
        RECT 5.930 328.000 6.330 328.600 ;
        RECT 5.930 327.800 9.930 328.000 ;
        RECT 5.930 327.200 6.330 327.800 ;
        RECT 5.930 327.000 9.930 327.200 ;
        RECT 5.930 326.400 6.330 327.000 ;
        RECT 5.930 326.200 9.930 326.400 ;
        RECT 5.930 325.600 6.330 326.200 ;
        RECT 5.930 325.400 9.930 325.600 ;
        RECT 5.930 324.800 6.330 325.400 ;
        RECT 5.930 324.600 9.930 324.800 ;
        RECT 5.930 324.000 6.330 324.600 ;
        RECT 5.930 323.800 9.930 324.000 ;
        RECT 5.930 323.200 6.330 323.800 ;
        RECT 5.930 323.000 9.930 323.200 ;
        RECT 5.930 322.400 6.330 323.000 ;
        RECT 5.930 322.200 9.930 322.400 ;
        RECT 10.680 322.200 10.880 329.800 ;
        RECT 11.480 322.200 11.680 329.800 ;
        RECT 12.280 322.200 12.480 329.800 ;
        RECT 13.080 322.200 13.280 329.800 ;
        RECT 13.880 322.200 14.080 329.800 ;
        RECT 15.380 330.200 15.580 337.800 ;
        RECT 16.180 330.200 16.380 337.800 ;
        RECT 16.980 330.200 17.180 337.800 ;
        RECT 17.780 330.200 17.980 337.800 ;
        RECT 18.580 330.200 18.780 337.800 ;
        RECT 19.530 337.600 23.530 337.800 ;
        RECT 23.130 337.000 23.530 337.600 ;
        RECT 19.530 336.800 23.530 337.000 ;
        RECT 23.130 336.200 23.530 336.800 ;
        RECT 19.530 336.000 23.530 336.200 ;
        RECT 23.130 335.400 23.530 336.000 ;
        RECT 19.530 335.200 23.530 335.400 ;
        RECT 23.130 334.600 23.530 335.200 ;
        RECT 19.530 334.400 23.530 334.600 ;
        RECT 23.130 333.800 23.530 334.400 ;
        RECT 19.530 333.600 23.530 333.800 ;
        RECT 23.130 333.000 23.530 333.600 ;
        RECT 19.530 332.800 23.530 333.000 ;
        RECT 23.130 332.200 23.530 332.800 ;
        RECT 19.530 332.000 23.530 332.200 ;
        RECT 23.130 331.400 23.530 332.000 ;
        RECT 19.530 331.200 23.530 331.400 ;
        RECT 23.130 330.600 23.530 331.200 ;
        RECT 19.530 330.400 23.530 330.600 ;
        RECT 23.130 330.200 23.530 330.400 ;
        RECT 15.380 329.800 23.530 330.200 ;
        RECT 15.380 322.200 15.580 329.800 ;
        RECT 16.180 322.200 16.380 329.800 ;
        RECT 16.980 322.200 17.180 329.800 ;
        RECT 17.780 322.200 17.980 329.800 ;
        RECT 18.580 322.200 18.780 329.800 ;
        RECT 23.130 329.600 23.530 329.800 ;
        RECT 19.530 329.400 23.530 329.600 ;
        RECT 23.130 328.800 23.530 329.400 ;
        RECT 19.530 328.600 23.530 328.800 ;
        RECT 23.130 328.000 23.530 328.600 ;
        RECT 19.530 327.800 23.530 328.000 ;
        RECT 23.130 327.200 23.530 327.800 ;
        RECT 19.530 327.000 23.530 327.200 ;
        RECT 23.130 326.400 23.530 327.000 ;
        RECT 19.530 326.200 23.530 326.400 ;
        RECT 23.130 325.600 23.530 326.200 ;
        RECT 19.530 325.400 23.530 325.600 ;
        RECT 23.130 324.800 23.530 325.400 ;
        RECT 19.530 324.600 23.530 324.800 ;
        RECT 23.130 324.000 23.530 324.600 ;
        RECT 19.530 323.800 23.530 324.000 ;
        RECT 23.130 323.200 23.530 323.800 ;
        RECT 19.530 323.000 23.530 323.200 ;
        RECT 23.130 322.400 23.530 323.000 ;
        RECT 19.530 322.200 23.530 322.400 ;
        RECT 25.930 337.600 29.930 337.800 ;
        RECT 25.930 337.000 26.330 337.600 ;
        RECT 25.930 336.800 29.930 337.000 ;
        RECT 25.930 336.200 26.330 336.800 ;
        RECT 25.930 336.000 29.930 336.200 ;
        RECT 25.930 335.400 26.330 336.000 ;
        RECT 25.930 335.200 29.930 335.400 ;
        RECT 25.930 334.600 26.330 335.200 ;
        RECT 25.930 334.400 29.930 334.600 ;
        RECT 25.930 333.800 26.330 334.400 ;
        RECT 25.930 333.600 29.930 333.800 ;
        RECT 25.930 333.000 26.330 333.600 ;
        RECT 25.930 332.800 29.930 333.000 ;
        RECT 25.930 332.200 26.330 332.800 ;
        RECT 25.930 332.000 29.930 332.200 ;
        RECT 25.930 331.400 26.330 332.000 ;
        RECT 25.930 331.200 29.930 331.400 ;
        RECT 25.930 330.600 26.330 331.200 ;
        RECT 25.930 330.400 29.930 330.600 ;
        RECT 25.930 330.200 26.330 330.400 ;
        RECT 30.680 330.200 30.880 337.800 ;
        RECT 31.480 330.200 31.680 337.800 ;
        RECT 32.280 330.200 32.480 337.800 ;
        RECT 33.080 330.200 33.280 337.800 ;
        RECT 33.880 330.200 34.080 337.800 ;
        RECT 25.930 329.800 34.080 330.200 ;
        RECT 25.930 329.600 26.330 329.800 ;
        RECT 25.930 329.400 29.930 329.600 ;
        RECT 25.930 328.800 26.330 329.400 ;
        RECT 25.930 328.600 29.930 328.800 ;
        RECT 25.930 328.000 26.330 328.600 ;
        RECT 25.930 327.800 29.930 328.000 ;
        RECT 25.930 327.200 26.330 327.800 ;
        RECT 25.930 327.000 29.930 327.200 ;
        RECT 25.930 326.400 26.330 327.000 ;
        RECT 25.930 326.200 29.930 326.400 ;
        RECT 25.930 325.600 26.330 326.200 ;
        RECT 25.930 325.400 29.930 325.600 ;
        RECT 25.930 324.800 26.330 325.400 ;
        RECT 25.930 324.600 29.930 324.800 ;
        RECT 25.930 324.000 26.330 324.600 ;
        RECT 25.930 323.800 29.930 324.000 ;
        RECT 25.930 323.200 26.330 323.800 ;
        RECT 25.930 323.000 29.930 323.200 ;
        RECT 25.930 322.400 26.330 323.000 ;
        RECT 25.930 322.200 29.930 322.400 ;
        RECT 30.680 322.200 30.880 329.800 ;
        RECT 31.480 322.200 31.680 329.800 ;
        RECT 32.280 322.200 32.480 329.800 ;
        RECT 33.080 322.200 33.280 329.800 ;
        RECT 33.880 322.200 34.080 329.800 ;
        RECT 35.380 330.200 35.580 337.800 ;
        RECT 36.180 330.200 36.380 337.800 ;
        RECT 36.980 330.200 37.180 337.800 ;
        RECT 37.780 330.200 37.980 337.800 ;
        RECT 38.580 330.200 38.780 337.800 ;
        RECT 39.530 337.600 43.530 337.800 ;
        RECT 43.130 337.000 43.530 337.600 ;
        RECT 39.530 336.800 43.530 337.000 ;
        RECT 43.130 336.200 43.530 336.800 ;
        RECT 39.530 336.000 43.530 336.200 ;
        RECT 43.130 335.400 43.530 336.000 ;
        RECT 39.530 335.200 43.530 335.400 ;
        RECT 43.130 334.600 43.530 335.200 ;
        RECT 39.530 334.400 43.530 334.600 ;
        RECT 43.130 333.800 43.530 334.400 ;
        RECT 39.530 333.600 43.530 333.800 ;
        RECT 43.130 333.000 43.530 333.600 ;
        RECT 39.530 332.800 43.530 333.000 ;
        RECT 43.130 332.200 43.530 332.800 ;
        RECT 39.530 332.000 43.530 332.200 ;
        RECT 43.130 331.400 43.530 332.000 ;
        RECT 39.530 331.200 43.530 331.400 ;
        RECT 43.130 330.600 43.530 331.200 ;
        RECT 39.530 330.400 43.530 330.600 ;
        RECT 43.130 330.200 43.530 330.400 ;
        RECT 35.380 329.800 43.530 330.200 ;
        RECT 35.380 322.200 35.580 329.800 ;
        RECT 36.180 322.200 36.380 329.800 ;
        RECT 36.980 322.200 37.180 329.800 ;
        RECT 37.780 322.200 37.980 329.800 ;
        RECT 38.580 322.200 38.780 329.800 ;
        RECT 43.130 329.600 43.530 329.800 ;
        RECT 39.530 329.400 43.530 329.600 ;
        RECT 43.130 328.800 43.530 329.400 ;
        RECT 39.530 328.600 43.530 328.800 ;
        RECT 43.130 328.000 43.530 328.600 ;
        RECT 39.530 327.800 43.530 328.000 ;
        RECT 43.130 327.200 43.530 327.800 ;
        RECT 39.530 327.000 43.530 327.200 ;
        RECT 43.130 326.400 43.530 327.000 ;
        RECT 39.530 326.200 43.530 326.400 ;
        RECT 43.130 325.600 43.530 326.200 ;
        RECT 39.530 325.400 43.530 325.600 ;
        RECT 43.130 324.800 43.530 325.400 ;
        RECT 39.530 324.600 43.530 324.800 ;
        RECT 43.130 324.000 43.530 324.600 ;
        RECT 39.530 323.800 43.530 324.000 ;
        RECT 43.130 323.200 43.530 323.800 ;
        RECT 39.530 323.000 43.530 323.200 ;
        RECT 43.130 322.400 43.530 323.000 ;
        RECT 39.530 322.200 43.530 322.400 ;
        RECT 45.930 337.600 49.930 337.800 ;
        RECT 45.930 337.000 46.330 337.600 ;
        RECT 45.930 336.800 49.930 337.000 ;
        RECT 45.930 336.200 46.330 336.800 ;
        RECT 45.930 336.000 49.930 336.200 ;
        RECT 45.930 335.400 46.330 336.000 ;
        RECT 45.930 335.200 49.930 335.400 ;
        RECT 45.930 334.600 46.330 335.200 ;
        RECT 45.930 334.400 49.930 334.600 ;
        RECT 45.930 333.800 46.330 334.400 ;
        RECT 45.930 333.600 49.930 333.800 ;
        RECT 45.930 333.000 46.330 333.600 ;
        RECT 45.930 332.800 49.930 333.000 ;
        RECT 45.930 332.200 46.330 332.800 ;
        RECT 45.930 332.000 49.930 332.200 ;
        RECT 45.930 331.400 46.330 332.000 ;
        RECT 45.930 331.200 49.930 331.400 ;
        RECT 45.930 330.600 46.330 331.200 ;
        RECT 45.930 330.400 49.930 330.600 ;
        RECT 45.930 330.200 46.330 330.400 ;
        RECT 50.680 330.200 50.880 337.800 ;
        RECT 51.480 330.200 51.680 337.800 ;
        RECT 52.280 330.200 52.480 337.800 ;
        RECT 53.080 330.200 53.280 337.800 ;
        RECT 53.880 330.200 54.080 337.800 ;
        RECT 45.930 329.800 54.080 330.200 ;
        RECT 45.930 329.600 46.330 329.800 ;
        RECT 45.930 329.400 49.930 329.600 ;
        RECT 45.930 328.800 46.330 329.400 ;
        RECT 45.930 328.600 49.930 328.800 ;
        RECT 45.930 328.000 46.330 328.600 ;
        RECT 45.930 327.800 49.930 328.000 ;
        RECT 45.930 327.200 46.330 327.800 ;
        RECT 45.930 327.000 49.930 327.200 ;
        RECT 45.930 326.400 46.330 327.000 ;
        RECT 45.930 326.200 49.930 326.400 ;
        RECT 45.930 325.600 46.330 326.200 ;
        RECT 45.930 325.400 49.930 325.600 ;
        RECT 45.930 324.800 46.330 325.400 ;
        RECT 45.930 324.600 49.930 324.800 ;
        RECT 45.930 324.000 46.330 324.600 ;
        RECT 45.930 323.800 49.930 324.000 ;
        RECT 45.930 323.200 46.330 323.800 ;
        RECT 45.930 323.000 49.930 323.200 ;
        RECT 45.930 322.400 46.330 323.000 ;
        RECT 45.930 322.200 49.930 322.400 ;
        RECT 50.680 322.200 50.880 329.800 ;
        RECT 51.480 322.200 51.680 329.800 ;
        RECT 52.280 322.200 52.480 329.800 ;
        RECT 53.080 322.200 53.280 329.800 ;
        RECT 53.880 322.200 54.080 329.800 ;
        RECT 55.380 330.200 55.580 337.800 ;
        RECT 56.180 330.200 56.380 337.800 ;
        RECT 56.980 330.200 57.180 337.800 ;
        RECT 57.780 330.200 57.980 337.800 ;
        RECT 58.580 330.200 58.780 337.800 ;
        RECT 59.530 337.600 63.530 337.800 ;
        RECT 63.130 337.000 63.530 337.600 ;
        RECT 59.530 336.800 63.530 337.000 ;
        RECT 63.130 336.200 63.530 336.800 ;
        RECT 59.530 336.000 63.530 336.200 ;
        RECT 63.130 335.400 63.530 336.000 ;
        RECT 59.530 335.200 63.530 335.400 ;
        RECT 63.130 334.600 63.530 335.200 ;
        RECT 59.530 334.400 63.530 334.600 ;
        RECT 63.130 333.800 63.530 334.400 ;
        RECT 59.530 333.600 63.530 333.800 ;
        RECT 63.130 333.000 63.530 333.600 ;
        RECT 59.530 332.800 63.530 333.000 ;
        RECT 63.130 332.200 63.530 332.800 ;
        RECT 59.530 332.000 63.530 332.200 ;
        RECT 63.130 331.400 63.530 332.000 ;
        RECT 59.530 331.200 63.530 331.400 ;
        RECT 63.130 330.600 63.530 331.200 ;
        RECT 59.530 330.400 63.530 330.600 ;
        RECT 63.130 330.200 63.530 330.400 ;
        RECT 55.380 329.800 63.530 330.200 ;
        RECT 55.380 322.200 55.580 329.800 ;
        RECT 56.180 322.200 56.380 329.800 ;
        RECT 56.980 322.200 57.180 329.800 ;
        RECT 57.780 322.200 57.980 329.800 ;
        RECT 58.580 322.200 58.780 329.800 ;
        RECT 63.130 329.600 63.530 329.800 ;
        RECT 59.530 329.400 63.530 329.600 ;
        RECT 63.130 328.800 63.530 329.400 ;
        RECT 59.530 328.600 63.530 328.800 ;
        RECT 63.130 328.000 63.530 328.600 ;
        RECT 59.530 327.800 63.530 328.000 ;
        RECT 63.130 327.200 63.530 327.800 ;
        RECT 59.530 327.000 63.530 327.200 ;
        RECT 63.130 326.400 63.530 327.000 ;
        RECT 59.530 326.200 63.530 326.400 ;
        RECT 63.130 325.600 63.530 326.200 ;
        RECT 59.530 325.400 63.530 325.600 ;
        RECT 63.130 324.800 63.530 325.400 ;
        RECT 59.530 324.600 63.530 324.800 ;
        RECT 63.130 324.000 63.530 324.600 ;
        RECT 59.530 323.800 63.530 324.000 ;
        RECT 63.130 323.200 63.530 323.800 ;
        RECT 59.530 323.000 63.530 323.200 ;
        RECT 63.130 322.400 63.530 323.000 ;
        RECT 59.530 322.200 63.530 322.400 ;
        RECT 65.930 337.600 69.930 337.800 ;
        RECT 65.930 337.000 66.330 337.600 ;
        RECT 65.930 336.800 69.930 337.000 ;
        RECT 65.930 336.200 66.330 336.800 ;
        RECT 65.930 336.000 69.930 336.200 ;
        RECT 65.930 335.400 66.330 336.000 ;
        RECT 65.930 335.200 69.930 335.400 ;
        RECT 65.930 334.600 66.330 335.200 ;
        RECT 65.930 334.400 69.930 334.600 ;
        RECT 65.930 333.800 66.330 334.400 ;
        RECT 65.930 333.600 69.930 333.800 ;
        RECT 65.930 333.000 66.330 333.600 ;
        RECT 65.930 332.800 69.930 333.000 ;
        RECT 65.930 332.200 66.330 332.800 ;
        RECT 65.930 332.000 69.930 332.200 ;
        RECT 65.930 331.400 66.330 332.000 ;
        RECT 65.930 331.200 69.930 331.400 ;
        RECT 65.930 330.600 66.330 331.200 ;
        RECT 65.930 330.400 69.930 330.600 ;
        RECT 65.930 330.200 66.330 330.400 ;
        RECT 70.680 330.200 70.880 337.800 ;
        RECT 71.480 330.200 71.680 337.800 ;
        RECT 72.280 330.200 72.480 337.800 ;
        RECT 73.080 330.200 73.280 337.800 ;
        RECT 73.880 330.200 74.080 337.800 ;
        RECT 65.930 329.800 74.080 330.200 ;
        RECT 65.930 329.600 66.330 329.800 ;
        RECT 65.930 329.400 69.930 329.600 ;
        RECT 65.930 328.800 66.330 329.400 ;
        RECT 65.930 328.600 69.930 328.800 ;
        RECT 65.930 328.000 66.330 328.600 ;
        RECT 65.930 327.800 69.930 328.000 ;
        RECT 65.930 327.200 66.330 327.800 ;
        RECT 65.930 327.000 69.930 327.200 ;
        RECT 65.930 326.400 66.330 327.000 ;
        RECT 65.930 326.200 69.930 326.400 ;
        RECT 65.930 325.600 66.330 326.200 ;
        RECT 65.930 325.400 69.930 325.600 ;
        RECT 65.930 324.800 66.330 325.400 ;
        RECT 65.930 324.600 69.930 324.800 ;
        RECT 65.930 324.000 66.330 324.600 ;
        RECT 65.930 323.800 69.930 324.000 ;
        RECT 65.930 323.200 66.330 323.800 ;
        RECT 65.930 323.000 69.930 323.200 ;
        RECT 65.930 322.400 66.330 323.000 ;
        RECT 65.930 322.200 69.930 322.400 ;
        RECT 70.680 322.200 70.880 329.800 ;
        RECT 71.480 322.200 71.680 329.800 ;
        RECT 72.280 322.200 72.480 329.800 ;
        RECT 73.080 322.200 73.280 329.800 ;
        RECT 73.880 322.200 74.080 329.800 ;
        RECT 75.380 330.200 75.580 337.800 ;
        RECT 76.180 330.200 76.380 337.800 ;
        RECT 76.980 330.200 77.180 337.800 ;
        RECT 77.780 330.200 77.980 337.800 ;
        RECT 78.580 330.200 78.780 337.800 ;
        RECT 79.530 337.600 83.530 337.800 ;
        RECT 83.130 337.000 83.530 337.600 ;
        RECT 79.530 336.800 83.530 337.000 ;
        RECT 83.130 336.200 83.530 336.800 ;
        RECT 79.530 336.000 83.530 336.200 ;
        RECT 83.130 335.400 83.530 336.000 ;
        RECT 79.530 335.200 83.530 335.400 ;
        RECT 83.130 334.600 83.530 335.200 ;
        RECT 79.530 334.400 83.530 334.600 ;
        RECT 83.130 333.800 83.530 334.400 ;
        RECT 79.530 333.600 83.530 333.800 ;
        RECT 83.130 333.000 83.530 333.600 ;
        RECT 79.530 332.800 83.530 333.000 ;
        RECT 83.130 332.200 83.530 332.800 ;
        RECT 79.530 332.000 83.530 332.200 ;
        RECT 83.130 331.400 83.530 332.000 ;
        RECT 79.530 331.200 83.530 331.400 ;
        RECT 83.130 330.600 83.530 331.200 ;
        RECT 79.530 330.400 83.530 330.600 ;
        RECT 83.130 330.200 83.530 330.400 ;
        RECT 75.380 329.800 83.530 330.200 ;
        RECT 75.380 322.200 75.580 329.800 ;
        RECT 76.180 322.200 76.380 329.800 ;
        RECT 76.980 322.200 77.180 329.800 ;
        RECT 77.780 322.200 77.980 329.800 ;
        RECT 78.580 322.200 78.780 329.800 ;
        RECT 83.130 329.600 83.530 329.800 ;
        RECT 79.530 329.400 83.530 329.600 ;
        RECT 83.130 328.800 83.530 329.400 ;
        RECT 79.530 328.600 83.530 328.800 ;
        RECT 83.130 328.000 83.530 328.600 ;
        RECT 79.530 327.800 83.530 328.000 ;
        RECT 83.130 327.200 83.530 327.800 ;
        RECT 79.530 327.000 83.530 327.200 ;
        RECT 83.130 326.400 83.530 327.000 ;
        RECT 79.530 326.200 83.530 326.400 ;
        RECT 83.130 325.600 83.530 326.200 ;
        RECT 79.530 325.400 83.530 325.600 ;
        RECT 83.130 324.800 83.530 325.400 ;
        RECT 79.530 324.600 83.530 324.800 ;
        RECT 83.130 324.000 83.530 324.600 ;
        RECT 79.530 323.800 83.530 324.000 ;
        RECT 83.130 323.200 83.530 323.800 ;
        RECT 79.530 323.000 83.530 323.200 ;
        RECT 83.130 322.400 83.530 323.000 ;
        RECT 79.530 322.200 83.530 322.400 ;
        RECT 85.930 337.600 89.930 337.800 ;
        RECT 85.930 337.000 86.330 337.600 ;
        RECT 85.930 336.800 89.930 337.000 ;
        RECT 85.930 336.200 86.330 336.800 ;
        RECT 85.930 336.000 89.930 336.200 ;
        RECT 85.930 335.400 86.330 336.000 ;
        RECT 85.930 335.200 89.930 335.400 ;
        RECT 85.930 334.600 86.330 335.200 ;
        RECT 85.930 334.400 89.930 334.600 ;
        RECT 85.930 333.800 86.330 334.400 ;
        RECT 85.930 333.600 89.930 333.800 ;
        RECT 85.930 333.000 86.330 333.600 ;
        RECT 85.930 332.800 89.930 333.000 ;
        RECT 85.930 332.200 86.330 332.800 ;
        RECT 85.930 332.000 89.930 332.200 ;
        RECT 85.930 331.400 86.330 332.000 ;
        RECT 85.930 331.200 89.930 331.400 ;
        RECT 85.930 330.600 86.330 331.200 ;
        RECT 85.930 330.400 89.930 330.600 ;
        RECT 85.930 330.200 86.330 330.400 ;
        RECT 90.680 330.200 90.880 337.800 ;
        RECT 91.480 330.200 91.680 337.800 ;
        RECT 92.280 330.200 92.480 337.800 ;
        RECT 93.080 330.200 93.280 337.800 ;
        RECT 93.880 330.200 94.080 337.800 ;
        RECT 85.930 329.800 94.080 330.200 ;
        RECT 85.930 329.600 86.330 329.800 ;
        RECT 85.930 329.400 89.930 329.600 ;
        RECT 85.930 328.800 86.330 329.400 ;
        RECT 85.930 328.600 89.930 328.800 ;
        RECT 85.930 328.000 86.330 328.600 ;
        RECT 85.930 327.800 89.930 328.000 ;
        RECT 85.930 327.200 86.330 327.800 ;
        RECT 85.930 327.000 89.930 327.200 ;
        RECT 85.930 326.400 86.330 327.000 ;
        RECT 85.930 326.200 89.930 326.400 ;
        RECT 85.930 325.600 86.330 326.200 ;
        RECT 85.930 325.400 89.930 325.600 ;
        RECT 85.930 324.800 86.330 325.400 ;
        RECT 85.930 324.600 89.930 324.800 ;
        RECT 85.930 324.000 86.330 324.600 ;
        RECT 85.930 323.800 89.930 324.000 ;
        RECT 85.930 323.200 86.330 323.800 ;
        RECT 85.930 323.000 89.930 323.200 ;
        RECT 85.930 322.400 86.330 323.000 ;
        RECT 85.930 322.200 89.930 322.400 ;
        RECT 90.680 322.200 90.880 329.800 ;
        RECT 91.480 322.200 91.680 329.800 ;
        RECT 92.280 322.200 92.480 329.800 ;
        RECT 93.080 322.200 93.280 329.800 ;
        RECT 93.880 322.200 94.080 329.800 ;
        RECT 95.380 330.200 95.580 337.800 ;
        RECT 96.180 330.200 96.380 337.800 ;
        RECT 96.980 330.200 97.180 337.800 ;
        RECT 97.780 330.200 97.980 337.800 ;
        RECT 98.580 330.200 98.780 337.800 ;
        RECT 99.530 337.600 103.530 337.800 ;
        RECT 103.130 337.000 103.530 337.600 ;
        RECT 99.530 336.800 103.530 337.000 ;
        RECT 103.130 336.200 103.530 336.800 ;
        RECT 99.530 336.000 103.530 336.200 ;
        RECT 103.130 335.400 103.530 336.000 ;
        RECT 99.530 335.200 103.530 335.400 ;
        RECT 103.130 334.600 103.530 335.200 ;
        RECT 99.530 334.400 103.530 334.600 ;
        RECT 103.130 333.800 103.530 334.400 ;
        RECT 99.530 333.600 103.530 333.800 ;
        RECT 103.130 333.000 103.530 333.600 ;
        RECT 99.530 332.800 103.530 333.000 ;
        RECT 103.130 332.200 103.530 332.800 ;
        RECT 99.530 332.000 103.530 332.200 ;
        RECT 103.130 331.400 103.530 332.000 ;
        RECT 99.530 331.200 103.530 331.400 ;
        RECT 103.130 330.600 103.530 331.200 ;
        RECT 99.530 330.400 103.530 330.600 ;
        RECT 103.130 330.200 103.530 330.400 ;
        RECT 95.380 329.800 103.530 330.200 ;
        RECT 95.380 322.200 95.580 329.800 ;
        RECT 96.180 322.200 96.380 329.800 ;
        RECT 96.980 322.200 97.180 329.800 ;
        RECT 97.780 322.200 97.980 329.800 ;
        RECT 98.580 322.200 98.780 329.800 ;
        RECT 103.130 329.600 103.530 329.800 ;
        RECT 99.530 329.400 103.530 329.600 ;
        RECT 103.130 328.800 103.530 329.400 ;
        RECT 99.530 328.600 103.530 328.800 ;
        RECT 103.130 328.000 103.530 328.600 ;
        RECT 99.530 327.800 103.530 328.000 ;
        RECT 103.130 327.200 103.530 327.800 ;
        RECT 99.530 327.000 103.530 327.200 ;
        RECT 103.130 326.400 103.530 327.000 ;
        RECT 99.530 326.200 103.530 326.400 ;
        RECT 103.130 325.600 103.530 326.200 ;
        RECT 99.530 325.400 103.530 325.600 ;
        RECT 103.130 324.800 103.530 325.400 ;
        RECT 99.530 324.600 103.530 324.800 ;
        RECT 103.130 324.000 103.530 324.600 ;
        RECT 99.530 323.800 103.530 324.000 ;
        RECT 103.130 323.200 103.530 323.800 ;
        RECT 99.530 323.000 103.530 323.200 ;
        RECT 103.130 322.400 103.530 323.000 ;
        RECT 99.530 322.200 103.530 322.400 ;
        RECT 105.930 337.600 109.930 337.800 ;
        RECT 105.930 337.000 106.330 337.600 ;
        RECT 105.930 336.800 109.930 337.000 ;
        RECT 105.930 336.200 106.330 336.800 ;
        RECT 105.930 336.000 109.930 336.200 ;
        RECT 105.930 335.400 106.330 336.000 ;
        RECT 105.930 335.200 109.930 335.400 ;
        RECT 105.930 334.600 106.330 335.200 ;
        RECT 105.930 334.400 109.930 334.600 ;
        RECT 105.930 333.800 106.330 334.400 ;
        RECT 105.930 333.600 109.930 333.800 ;
        RECT 105.930 333.000 106.330 333.600 ;
        RECT 105.930 332.800 109.930 333.000 ;
        RECT 105.930 332.200 106.330 332.800 ;
        RECT 105.930 332.000 109.930 332.200 ;
        RECT 105.930 331.400 106.330 332.000 ;
        RECT 105.930 331.200 109.930 331.400 ;
        RECT 105.930 330.600 106.330 331.200 ;
        RECT 105.930 330.400 109.930 330.600 ;
        RECT 105.930 330.200 106.330 330.400 ;
        RECT 110.680 330.200 110.880 337.800 ;
        RECT 111.480 330.200 111.680 337.800 ;
        RECT 112.280 330.200 112.480 337.800 ;
        RECT 113.080 330.200 113.280 337.800 ;
        RECT 113.880 330.200 114.080 337.800 ;
        RECT 105.930 329.800 114.080 330.200 ;
        RECT 105.930 329.600 106.330 329.800 ;
        RECT 105.930 329.400 109.930 329.600 ;
        RECT 105.930 328.800 106.330 329.400 ;
        RECT 105.930 328.600 109.930 328.800 ;
        RECT 105.930 328.000 106.330 328.600 ;
        RECT 105.930 327.800 109.930 328.000 ;
        RECT 105.930 327.200 106.330 327.800 ;
        RECT 105.930 327.000 109.930 327.200 ;
        RECT 105.930 326.400 106.330 327.000 ;
        RECT 105.930 326.200 109.930 326.400 ;
        RECT 105.930 325.600 106.330 326.200 ;
        RECT 105.930 325.400 109.930 325.600 ;
        RECT 105.930 324.800 106.330 325.400 ;
        RECT 105.930 324.600 109.930 324.800 ;
        RECT 105.930 324.000 106.330 324.600 ;
        RECT 105.930 323.800 109.930 324.000 ;
        RECT 105.930 323.200 106.330 323.800 ;
        RECT 105.930 323.000 109.930 323.200 ;
        RECT 105.930 322.400 106.330 323.000 ;
        RECT 105.930 322.200 109.930 322.400 ;
        RECT 110.680 322.200 110.880 329.800 ;
        RECT 111.480 322.200 111.680 329.800 ;
        RECT 112.280 322.200 112.480 329.800 ;
        RECT 113.080 322.200 113.280 329.800 ;
        RECT 113.880 322.200 114.080 329.800 ;
        RECT 115.380 330.200 115.580 337.800 ;
        RECT 116.180 330.200 116.380 337.800 ;
        RECT 116.980 330.200 117.180 337.800 ;
        RECT 117.780 330.200 117.980 337.800 ;
        RECT 118.580 330.200 118.780 337.800 ;
        RECT 119.530 337.600 123.530 337.800 ;
        RECT 123.130 337.000 123.530 337.600 ;
        RECT 119.530 336.800 123.530 337.000 ;
        RECT 123.130 336.200 123.530 336.800 ;
        RECT 119.530 336.000 123.530 336.200 ;
        RECT 123.130 335.400 123.530 336.000 ;
        RECT 119.530 335.200 123.530 335.400 ;
        RECT 123.130 334.600 123.530 335.200 ;
        RECT 119.530 334.400 123.530 334.600 ;
        RECT 123.130 333.800 123.530 334.400 ;
        RECT 119.530 333.600 123.530 333.800 ;
        RECT 123.130 333.000 123.530 333.600 ;
        RECT 119.530 332.800 123.530 333.000 ;
        RECT 123.130 332.200 123.530 332.800 ;
        RECT 119.530 332.000 123.530 332.200 ;
        RECT 123.130 331.400 123.530 332.000 ;
        RECT 119.530 331.200 123.530 331.400 ;
        RECT 123.130 330.600 123.530 331.200 ;
        RECT 119.530 330.400 123.530 330.600 ;
        RECT 123.130 330.200 123.530 330.400 ;
        RECT 115.380 329.800 123.530 330.200 ;
        RECT 130.050 329.975 130.410 330.355 ;
        RECT 130.680 329.975 131.040 330.355 ;
        RECT 131.280 329.975 131.640 330.355 ;
        RECT 115.380 322.200 115.580 329.800 ;
        RECT 116.180 322.200 116.380 329.800 ;
        RECT 116.980 322.200 117.180 329.800 ;
        RECT 117.780 322.200 117.980 329.800 ;
        RECT 118.580 322.200 118.780 329.800 ;
        RECT 123.130 329.600 123.530 329.800 ;
        RECT 119.530 329.400 123.530 329.600 ;
        RECT 123.130 328.800 123.530 329.400 ;
        RECT 130.050 329.385 130.410 329.765 ;
        RECT 130.680 329.385 131.040 329.765 ;
        RECT 131.280 329.385 131.640 329.765 ;
        RECT 119.530 328.600 123.530 328.800 ;
        RECT 123.130 328.000 123.530 328.600 ;
        RECT 119.530 327.800 123.530 328.000 ;
        RECT 123.130 327.200 123.530 327.800 ;
        RECT 119.530 327.000 123.530 327.200 ;
        RECT 123.130 326.400 123.530 327.000 ;
        RECT 119.530 326.200 123.530 326.400 ;
        RECT 123.130 325.600 123.530 326.200 ;
        RECT 119.530 325.400 123.530 325.600 ;
        RECT 123.130 324.800 123.530 325.400 ;
        RECT 119.530 324.600 123.530 324.800 ;
        RECT 123.130 324.000 123.530 324.600 ;
        RECT 119.530 323.800 123.530 324.000 ;
        RECT 123.130 323.200 123.530 323.800 ;
        RECT 119.530 323.000 123.530 323.200 ;
        RECT 123.130 322.400 123.530 323.000 ;
        RECT 119.530 322.200 123.530 322.400 ;
        RECT 5.930 317.600 9.930 317.800 ;
        RECT 5.930 317.000 6.330 317.600 ;
        RECT 5.930 316.800 9.930 317.000 ;
        RECT 5.930 316.200 6.330 316.800 ;
        RECT 5.930 316.000 9.930 316.200 ;
        RECT 5.930 315.400 6.330 316.000 ;
        RECT 5.930 315.200 9.930 315.400 ;
        RECT 5.930 314.600 6.330 315.200 ;
        RECT 5.930 314.400 9.930 314.600 ;
        RECT 5.930 313.800 6.330 314.400 ;
        RECT 5.930 313.600 9.930 313.800 ;
        RECT 5.930 313.000 6.330 313.600 ;
        RECT 5.930 312.800 9.930 313.000 ;
        RECT 5.930 312.200 6.330 312.800 ;
        RECT 5.930 312.000 9.930 312.200 ;
        RECT 5.930 311.400 6.330 312.000 ;
        RECT 5.930 311.200 9.930 311.400 ;
        RECT 5.930 310.600 6.330 311.200 ;
        RECT 5.930 310.400 9.930 310.600 ;
        RECT 5.930 310.200 6.330 310.400 ;
        RECT 10.680 310.200 10.880 317.800 ;
        RECT 11.480 310.200 11.680 317.800 ;
        RECT 12.280 310.200 12.480 317.800 ;
        RECT 13.080 310.200 13.280 317.800 ;
        RECT 13.880 310.200 14.080 317.800 ;
        RECT 5.930 309.800 14.080 310.200 ;
        RECT 5.930 309.600 6.330 309.800 ;
        RECT 5.930 309.400 9.930 309.600 ;
        RECT 5.930 308.800 6.330 309.400 ;
        RECT 5.930 308.600 9.930 308.800 ;
        RECT 5.930 308.000 6.330 308.600 ;
        RECT 5.930 307.800 9.930 308.000 ;
        RECT 5.930 307.200 6.330 307.800 ;
        RECT 5.930 307.000 9.930 307.200 ;
        RECT 5.930 306.400 6.330 307.000 ;
        RECT 5.930 306.200 9.930 306.400 ;
        RECT 5.930 305.600 6.330 306.200 ;
        RECT 5.930 305.400 9.930 305.600 ;
        RECT 5.930 304.800 6.330 305.400 ;
        RECT 5.930 304.600 9.930 304.800 ;
        RECT 5.930 304.000 6.330 304.600 ;
        RECT 5.930 303.800 9.930 304.000 ;
        RECT 5.930 303.200 6.330 303.800 ;
        RECT 5.930 303.000 9.930 303.200 ;
        RECT 5.930 302.400 6.330 303.000 ;
        RECT 5.930 302.200 9.930 302.400 ;
        RECT 10.680 302.200 10.880 309.800 ;
        RECT 11.480 302.200 11.680 309.800 ;
        RECT 12.280 302.200 12.480 309.800 ;
        RECT 13.080 302.200 13.280 309.800 ;
        RECT 13.880 302.200 14.080 309.800 ;
        RECT 15.380 310.200 15.580 317.800 ;
        RECT 16.180 310.200 16.380 317.800 ;
        RECT 16.980 310.200 17.180 317.800 ;
        RECT 17.780 310.200 17.980 317.800 ;
        RECT 18.580 310.200 18.780 317.800 ;
        RECT 19.530 317.600 23.530 317.800 ;
        RECT 23.130 317.000 23.530 317.600 ;
        RECT 19.530 316.800 23.530 317.000 ;
        RECT 23.130 316.200 23.530 316.800 ;
        RECT 19.530 316.000 23.530 316.200 ;
        RECT 23.130 315.400 23.530 316.000 ;
        RECT 19.530 315.200 23.530 315.400 ;
        RECT 23.130 314.600 23.530 315.200 ;
        RECT 19.530 314.400 23.530 314.600 ;
        RECT 23.130 313.800 23.530 314.400 ;
        RECT 19.530 313.600 23.530 313.800 ;
        RECT 23.130 313.000 23.530 313.600 ;
        RECT 19.530 312.800 23.530 313.000 ;
        RECT 23.130 312.200 23.530 312.800 ;
        RECT 19.530 312.000 23.530 312.200 ;
        RECT 23.130 311.400 23.530 312.000 ;
        RECT 19.530 311.200 23.530 311.400 ;
        RECT 23.130 310.600 23.530 311.200 ;
        RECT 19.530 310.400 23.530 310.600 ;
        RECT 23.130 310.200 23.530 310.400 ;
        RECT 15.380 309.800 23.530 310.200 ;
        RECT 15.380 302.200 15.580 309.800 ;
        RECT 16.180 302.200 16.380 309.800 ;
        RECT 16.980 302.200 17.180 309.800 ;
        RECT 17.780 302.200 17.980 309.800 ;
        RECT 18.580 302.200 18.780 309.800 ;
        RECT 23.130 309.600 23.530 309.800 ;
        RECT 19.530 309.400 23.530 309.600 ;
        RECT 23.130 308.800 23.530 309.400 ;
        RECT 19.530 308.600 23.530 308.800 ;
        RECT 23.130 308.000 23.530 308.600 ;
        RECT 19.530 307.800 23.530 308.000 ;
        RECT 23.130 307.200 23.530 307.800 ;
        RECT 19.530 307.000 23.530 307.200 ;
        RECT 23.130 306.400 23.530 307.000 ;
        RECT 19.530 306.200 23.530 306.400 ;
        RECT 23.130 305.600 23.530 306.200 ;
        RECT 19.530 305.400 23.530 305.600 ;
        RECT 23.130 304.800 23.530 305.400 ;
        RECT 19.530 304.600 23.530 304.800 ;
        RECT 23.130 304.000 23.530 304.600 ;
        RECT 19.530 303.800 23.530 304.000 ;
        RECT 23.130 303.200 23.530 303.800 ;
        RECT 19.530 303.000 23.530 303.200 ;
        RECT 23.130 302.400 23.530 303.000 ;
        RECT 19.530 302.200 23.530 302.400 ;
        RECT 25.930 317.600 29.930 317.800 ;
        RECT 25.930 317.000 26.330 317.600 ;
        RECT 25.930 316.800 29.930 317.000 ;
        RECT 25.930 316.200 26.330 316.800 ;
        RECT 25.930 316.000 29.930 316.200 ;
        RECT 25.930 315.400 26.330 316.000 ;
        RECT 25.930 315.200 29.930 315.400 ;
        RECT 25.930 314.600 26.330 315.200 ;
        RECT 25.930 314.400 29.930 314.600 ;
        RECT 25.930 313.800 26.330 314.400 ;
        RECT 25.930 313.600 29.930 313.800 ;
        RECT 25.930 313.000 26.330 313.600 ;
        RECT 25.930 312.800 29.930 313.000 ;
        RECT 25.930 312.200 26.330 312.800 ;
        RECT 25.930 312.000 29.930 312.200 ;
        RECT 25.930 311.400 26.330 312.000 ;
        RECT 25.930 311.200 29.930 311.400 ;
        RECT 25.930 310.600 26.330 311.200 ;
        RECT 25.930 310.400 29.930 310.600 ;
        RECT 25.930 310.200 26.330 310.400 ;
        RECT 30.680 310.200 30.880 317.800 ;
        RECT 31.480 310.200 31.680 317.800 ;
        RECT 32.280 310.200 32.480 317.800 ;
        RECT 33.080 310.200 33.280 317.800 ;
        RECT 33.880 310.200 34.080 317.800 ;
        RECT 25.930 309.800 34.080 310.200 ;
        RECT 25.930 309.600 26.330 309.800 ;
        RECT 25.930 309.400 29.930 309.600 ;
        RECT 25.930 308.800 26.330 309.400 ;
        RECT 25.930 308.600 29.930 308.800 ;
        RECT 25.930 308.000 26.330 308.600 ;
        RECT 25.930 307.800 29.930 308.000 ;
        RECT 25.930 307.200 26.330 307.800 ;
        RECT 25.930 307.000 29.930 307.200 ;
        RECT 25.930 306.400 26.330 307.000 ;
        RECT 25.930 306.200 29.930 306.400 ;
        RECT 25.930 305.600 26.330 306.200 ;
        RECT 25.930 305.400 29.930 305.600 ;
        RECT 25.930 304.800 26.330 305.400 ;
        RECT 25.930 304.600 29.930 304.800 ;
        RECT 25.930 304.000 26.330 304.600 ;
        RECT 25.930 303.800 29.930 304.000 ;
        RECT 25.930 303.200 26.330 303.800 ;
        RECT 25.930 303.000 29.930 303.200 ;
        RECT 25.930 302.400 26.330 303.000 ;
        RECT 25.930 302.200 29.930 302.400 ;
        RECT 30.680 302.200 30.880 309.800 ;
        RECT 31.480 302.200 31.680 309.800 ;
        RECT 32.280 302.200 32.480 309.800 ;
        RECT 33.080 302.200 33.280 309.800 ;
        RECT 33.880 302.200 34.080 309.800 ;
        RECT 35.380 310.200 35.580 317.800 ;
        RECT 36.180 310.200 36.380 317.800 ;
        RECT 36.980 310.200 37.180 317.800 ;
        RECT 37.780 310.200 37.980 317.800 ;
        RECT 38.580 310.200 38.780 317.800 ;
        RECT 39.530 317.600 43.530 317.800 ;
        RECT 43.130 317.000 43.530 317.600 ;
        RECT 39.530 316.800 43.530 317.000 ;
        RECT 43.130 316.200 43.530 316.800 ;
        RECT 39.530 316.000 43.530 316.200 ;
        RECT 43.130 315.400 43.530 316.000 ;
        RECT 39.530 315.200 43.530 315.400 ;
        RECT 43.130 314.600 43.530 315.200 ;
        RECT 39.530 314.400 43.530 314.600 ;
        RECT 43.130 313.800 43.530 314.400 ;
        RECT 39.530 313.600 43.530 313.800 ;
        RECT 43.130 313.000 43.530 313.600 ;
        RECT 39.530 312.800 43.530 313.000 ;
        RECT 43.130 312.200 43.530 312.800 ;
        RECT 39.530 312.000 43.530 312.200 ;
        RECT 43.130 311.400 43.530 312.000 ;
        RECT 39.530 311.200 43.530 311.400 ;
        RECT 43.130 310.600 43.530 311.200 ;
        RECT 39.530 310.400 43.530 310.600 ;
        RECT 43.130 310.200 43.530 310.400 ;
        RECT 35.380 309.800 43.530 310.200 ;
        RECT 35.380 302.200 35.580 309.800 ;
        RECT 36.180 302.200 36.380 309.800 ;
        RECT 36.980 302.200 37.180 309.800 ;
        RECT 37.780 302.200 37.980 309.800 ;
        RECT 38.580 302.200 38.780 309.800 ;
        RECT 43.130 309.600 43.530 309.800 ;
        RECT 39.530 309.400 43.530 309.600 ;
        RECT 43.130 308.800 43.530 309.400 ;
        RECT 39.530 308.600 43.530 308.800 ;
        RECT 43.130 308.000 43.530 308.600 ;
        RECT 39.530 307.800 43.530 308.000 ;
        RECT 43.130 307.200 43.530 307.800 ;
        RECT 39.530 307.000 43.530 307.200 ;
        RECT 43.130 306.400 43.530 307.000 ;
        RECT 39.530 306.200 43.530 306.400 ;
        RECT 43.130 305.600 43.530 306.200 ;
        RECT 39.530 305.400 43.530 305.600 ;
        RECT 43.130 304.800 43.530 305.400 ;
        RECT 39.530 304.600 43.530 304.800 ;
        RECT 43.130 304.000 43.530 304.600 ;
        RECT 39.530 303.800 43.530 304.000 ;
        RECT 43.130 303.200 43.530 303.800 ;
        RECT 39.530 303.000 43.530 303.200 ;
        RECT 43.130 302.400 43.530 303.000 ;
        RECT 39.530 302.200 43.530 302.400 ;
        RECT 45.930 317.600 49.930 317.800 ;
        RECT 45.930 317.000 46.330 317.600 ;
        RECT 45.930 316.800 49.930 317.000 ;
        RECT 45.930 316.200 46.330 316.800 ;
        RECT 45.930 316.000 49.930 316.200 ;
        RECT 45.930 315.400 46.330 316.000 ;
        RECT 45.930 315.200 49.930 315.400 ;
        RECT 45.930 314.600 46.330 315.200 ;
        RECT 45.930 314.400 49.930 314.600 ;
        RECT 45.930 313.800 46.330 314.400 ;
        RECT 45.930 313.600 49.930 313.800 ;
        RECT 45.930 313.000 46.330 313.600 ;
        RECT 45.930 312.800 49.930 313.000 ;
        RECT 45.930 312.200 46.330 312.800 ;
        RECT 45.930 312.000 49.930 312.200 ;
        RECT 45.930 311.400 46.330 312.000 ;
        RECT 45.930 311.200 49.930 311.400 ;
        RECT 45.930 310.600 46.330 311.200 ;
        RECT 45.930 310.400 49.930 310.600 ;
        RECT 45.930 310.200 46.330 310.400 ;
        RECT 50.680 310.200 50.880 317.800 ;
        RECT 51.480 310.200 51.680 317.800 ;
        RECT 52.280 310.200 52.480 317.800 ;
        RECT 53.080 310.200 53.280 317.800 ;
        RECT 53.880 310.200 54.080 317.800 ;
        RECT 45.930 309.800 54.080 310.200 ;
        RECT 45.930 309.600 46.330 309.800 ;
        RECT 45.930 309.400 49.930 309.600 ;
        RECT 45.930 308.800 46.330 309.400 ;
        RECT 45.930 308.600 49.930 308.800 ;
        RECT 45.930 308.000 46.330 308.600 ;
        RECT 45.930 307.800 49.930 308.000 ;
        RECT 45.930 307.200 46.330 307.800 ;
        RECT 45.930 307.000 49.930 307.200 ;
        RECT 45.930 306.400 46.330 307.000 ;
        RECT 45.930 306.200 49.930 306.400 ;
        RECT 45.930 305.600 46.330 306.200 ;
        RECT 45.930 305.400 49.930 305.600 ;
        RECT 45.930 304.800 46.330 305.400 ;
        RECT 45.930 304.600 49.930 304.800 ;
        RECT 45.930 304.000 46.330 304.600 ;
        RECT 45.930 303.800 49.930 304.000 ;
        RECT 45.930 303.200 46.330 303.800 ;
        RECT 45.930 303.000 49.930 303.200 ;
        RECT 45.930 302.400 46.330 303.000 ;
        RECT 45.930 302.200 49.930 302.400 ;
        RECT 50.680 302.200 50.880 309.800 ;
        RECT 51.480 302.200 51.680 309.800 ;
        RECT 52.280 302.200 52.480 309.800 ;
        RECT 53.080 302.200 53.280 309.800 ;
        RECT 53.880 302.200 54.080 309.800 ;
        RECT 55.380 310.200 55.580 317.800 ;
        RECT 56.180 310.200 56.380 317.800 ;
        RECT 56.980 310.200 57.180 317.800 ;
        RECT 57.780 310.200 57.980 317.800 ;
        RECT 58.580 310.200 58.780 317.800 ;
        RECT 59.530 317.600 63.530 317.800 ;
        RECT 63.130 317.000 63.530 317.600 ;
        RECT 59.530 316.800 63.530 317.000 ;
        RECT 63.130 316.200 63.530 316.800 ;
        RECT 59.530 316.000 63.530 316.200 ;
        RECT 63.130 315.400 63.530 316.000 ;
        RECT 59.530 315.200 63.530 315.400 ;
        RECT 63.130 314.600 63.530 315.200 ;
        RECT 59.530 314.400 63.530 314.600 ;
        RECT 63.130 313.800 63.530 314.400 ;
        RECT 59.530 313.600 63.530 313.800 ;
        RECT 63.130 313.000 63.530 313.600 ;
        RECT 59.530 312.800 63.530 313.000 ;
        RECT 63.130 312.200 63.530 312.800 ;
        RECT 59.530 312.000 63.530 312.200 ;
        RECT 63.130 311.400 63.530 312.000 ;
        RECT 59.530 311.200 63.530 311.400 ;
        RECT 63.130 310.600 63.530 311.200 ;
        RECT 59.530 310.400 63.530 310.600 ;
        RECT 63.130 310.200 63.530 310.400 ;
        RECT 55.380 309.800 63.530 310.200 ;
        RECT 55.380 302.200 55.580 309.800 ;
        RECT 56.180 302.200 56.380 309.800 ;
        RECT 56.980 302.200 57.180 309.800 ;
        RECT 57.780 302.200 57.980 309.800 ;
        RECT 58.580 302.200 58.780 309.800 ;
        RECT 63.130 309.600 63.530 309.800 ;
        RECT 59.530 309.400 63.530 309.600 ;
        RECT 63.130 308.800 63.530 309.400 ;
        RECT 59.530 308.600 63.530 308.800 ;
        RECT 63.130 308.000 63.530 308.600 ;
        RECT 59.530 307.800 63.530 308.000 ;
        RECT 63.130 307.200 63.530 307.800 ;
        RECT 59.530 307.000 63.530 307.200 ;
        RECT 63.130 306.400 63.530 307.000 ;
        RECT 59.530 306.200 63.530 306.400 ;
        RECT 63.130 305.600 63.530 306.200 ;
        RECT 59.530 305.400 63.530 305.600 ;
        RECT 63.130 304.800 63.530 305.400 ;
        RECT 59.530 304.600 63.530 304.800 ;
        RECT 63.130 304.000 63.530 304.600 ;
        RECT 59.530 303.800 63.530 304.000 ;
        RECT 63.130 303.200 63.530 303.800 ;
        RECT 59.530 303.000 63.530 303.200 ;
        RECT 63.130 302.400 63.530 303.000 ;
        RECT 59.530 302.200 63.530 302.400 ;
        RECT 65.930 317.600 69.930 317.800 ;
        RECT 65.930 317.000 66.330 317.600 ;
        RECT 65.930 316.800 69.930 317.000 ;
        RECT 65.930 316.200 66.330 316.800 ;
        RECT 65.930 316.000 69.930 316.200 ;
        RECT 65.930 315.400 66.330 316.000 ;
        RECT 65.930 315.200 69.930 315.400 ;
        RECT 65.930 314.600 66.330 315.200 ;
        RECT 65.930 314.400 69.930 314.600 ;
        RECT 65.930 313.800 66.330 314.400 ;
        RECT 65.930 313.600 69.930 313.800 ;
        RECT 65.930 313.000 66.330 313.600 ;
        RECT 65.930 312.800 69.930 313.000 ;
        RECT 65.930 312.200 66.330 312.800 ;
        RECT 65.930 312.000 69.930 312.200 ;
        RECT 65.930 311.400 66.330 312.000 ;
        RECT 65.930 311.200 69.930 311.400 ;
        RECT 65.930 310.600 66.330 311.200 ;
        RECT 65.930 310.400 69.930 310.600 ;
        RECT 65.930 310.200 66.330 310.400 ;
        RECT 70.680 310.200 70.880 317.800 ;
        RECT 71.480 310.200 71.680 317.800 ;
        RECT 72.280 310.200 72.480 317.800 ;
        RECT 73.080 310.200 73.280 317.800 ;
        RECT 73.880 310.200 74.080 317.800 ;
        RECT 65.930 309.800 74.080 310.200 ;
        RECT 65.930 309.600 66.330 309.800 ;
        RECT 65.930 309.400 69.930 309.600 ;
        RECT 65.930 308.800 66.330 309.400 ;
        RECT 65.930 308.600 69.930 308.800 ;
        RECT 65.930 308.000 66.330 308.600 ;
        RECT 65.930 307.800 69.930 308.000 ;
        RECT 65.930 307.200 66.330 307.800 ;
        RECT 65.930 307.000 69.930 307.200 ;
        RECT 65.930 306.400 66.330 307.000 ;
        RECT 65.930 306.200 69.930 306.400 ;
        RECT 65.930 305.600 66.330 306.200 ;
        RECT 65.930 305.400 69.930 305.600 ;
        RECT 65.930 304.800 66.330 305.400 ;
        RECT 65.930 304.600 69.930 304.800 ;
        RECT 65.930 304.000 66.330 304.600 ;
        RECT 65.930 303.800 69.930 304.000 ;
        RECT 65.930 303.200 66.330 303.800 ;
        RECT 65.930 303.000 69.930 303.200 ;
        RECT 65.930 302.400 66.330 303.000 ;
        RECT 65.930 302.200 69.930 302.400 ;
        RECT 70.680 302.200 70.880 309.800 ;
        RECT 71.480 302.200 71.680 309.800 ;
        RECT 72.280 302.200 72.480 309.800 ;
        RECT 73.080 302.200 73.280 309.800 ;
        RECT 73.880 302.200 74.080 309.800 ;
        RECT 75.380 310.200 75.580 317.800 ;
        RECT 76.180 310.200 76.380 317.800 ;
        RECT 76.980 310.200 77.180 317.800 ;
        RECT 77.780 310.200 77.980 317.800 ;
        RECT 78.580 310.200 78.780 317.800 ;
        RECT 79.530 317.600 83.530 317.800 ;
        RECT 83.130 317.000 83.530 317.600 ;
        RECT 79.530 316.800 83.530 317.000 ;
        RECT 83.130 316.200 83.530 316.800 ;
        RECT 79.530 316.000 83.530 316.200 ;
        RECT 83.130 315.400 83.530 316.000 ;
        RECT 79.530 315.200 83.530 315.400 ;
        RECT 83.130 314.600 83.530 315.200 ;
        RECT 79.530 314.400 83.530 314.600 ;
        RECT 83.130 313.800 83.530 314.400 ;
        RECT 79.530 313.600 83.530 313.800 ;
        RECT 83.130 313.000 83.530 313.600 ;
        RECT 79.530 312.800 83.530 313.000 ;
        RECT 83.130 312.200 83.530 312.800 ;
        RECT 79.530 312.000 83.530 312.200 ;
        RECT 83.130 311.400 83.530 312.000 ;
        RECT 79.530 311.200 83.530 311.400 ;
        RECT 83.130 310.600 83.530 311.200 ;
        RECT 79.530 310.400 83.530 310.600 ;
        RECT 83.130 310.200 83.530 310.400 ;
        RECT 75.380 309.800 83.530 310.200 ;
        RECT 75.380 302.200 75.580 309.800 ;
        RECT 76.180 302.200 76.380 309.800 ;
        RECT 76.980 302.200 77.180 309.800 ;
        RECT 77.780 302.200 77.980 309.800 ;
        RECT 78.580 302.200 78.780 309.800 ;
        RECT 83.130 309.600 83.530 309.800 ;
        RECT 79.530 309.400 83.530 309.600 ;
        RECT 83.130 308.800 83.530 309.400 ;
        RECT 79.530 308.600 83.530 308.800 ;
        RECT 83.130 308.000 83.530 308.600 ;
        RECT 79.530 307.800 83.530 308.000 ;
        RECT 83.130 307.200 83.530 307.800 ;
        RECT 79.530 307.000 83.530 307.200 ;
        RECT 83.130 306.400 83.530 307.000 ;
        RECT 79.530 306.200 83.530 306.400 ;
        RECT 83.130 305.600 83.530 306.200 ;
        RECT 79.530 305.400 83.530 305.600 ;
        RECT 83.130 304.800 83.530 305.400 ;
        RECT 79.530 304.600 83.530 304.800 ;
        RECT 83.130 304.000 83.530 304.600 ;
        RECT 79.530 303.800 83.530 304.000 ;
        RECT 83.130 303.200 83.530 303.800 ;
        RECT 79.530 303.000 83.530 303.200 ;
        RECT 83.130 302.400 83.530 303.000 ;
        RECT 79.530 302.200 83.530 302.400 ;
        RECT 85.930 317.600 89.930 317.800 ;
        RECT 85.930 317.000 86.330 317.600 ;
        RECT 85.930 316.800 89.930 317.000 ;
        RECT 85.930 316.200 86.330 316.800 ;
        RECT 85.930 316.000 89.930 316.200 ;
        RECT 85.930 315.400 86.330 316.000 ;
        RECT 85.930 315.200 89.930 315.400 ;
        RECT 85.930 314.600 86.330 315.200 ;
        RECT 85.930 314.400 89.930 314.600 ;
        RECT 85.930 313.800 86.330 314.400 ;
        RECT 85.930 313.600 89.930 313.800 ;
        RECT 85.930 313.000 86.330 313.600 ;
        RECT 85.930 312.800 89.930 313.000 ;
        RECT 85.930 312.200 86.330 312.800 ;
        RECT 85.930 312.000 89.930 312.200 ;
        RECT 85.930 311.400 86.330 312.000 ;
        RECT 85.930 311.200 89.930 311.400 ;
        RECT 85.930 310.600 86.330 311.200 ;
        RECT 85.930 310.400 89.930 310.600 ;
        RECT 85.930 310.200 86.330 310.400 ;
        RECT 90.680 310.200 90.880 317.800 ;
        RECT 91.480 310.200 91.680 317.800 ;
        RECT 92.280 310.200 92.480 317.800 ;
        RECT 93.080 310.200 93.280 317.800 ;
        RECT 93.880 310.200 94.080 317.800 ;
        RECT 85.930 309.800 94.080 310.200 ;
        RECT 85.930 309.600 86.330 309.800 ;
        RECT 85.930 309.400 89.930 309.600 ;
        RECT 85.930 308.800 86.330 309.400 ;
        RECT 85.930 308.600 89.930 308.800 ;
        RECT 85.930 308.000 86.330 308.600 ;
        RECT 85.930 307.800 89.930 308.000 ;
        RECT 85.930 307.200 86.330 307.800 ;
        RECT 85.930 307.000 89.930 307.200 ;
        RECT 85.930 306.400 86.330 307.000 ;
        RECT 85.930 306.200 89.930 306.400 ;
        RECT 85.930 305.600 86.330 306.200 ;
        RECT 85.930 305.400 89.930 305.600 ;
        RECT 85.930 304.800 86.330 305.400 ;
        RECT 85.930 304.600 89.930 304.800 ;
        RECT 85.930 304.000 86.330 304.600 ;
        RECT 85.930 303.800 89.930 304.000 ;
        RECT 85.930 303.200 86.330 303.800 ;
        RECT 85.930 303.000 89.930 303.200 ;
        RECT 85.930 302.400 86.330 303.000 ;
        RECT 85.930 302.200 89.930 302.400 ;
        RECT 90.680 302.200 90.880 309.800 ;
        RECT 91.480 302.200 91.680 309.800 ;
        RECT 92.280 302.200 92.480 309.800 ;
        RECT 93.080 302.200 93.280 309.800 ;
        RECT 93.880 302.200 94.080 309.800 ;
        RECT 95.380 310.200 95.580 317.800 ;
        RECT 96.180 310.200 96.380 317.800 ;
        RECT 96.980 310.200 97.180 317.800 ;
        RECT 97.780 310.200 97.980 317.800 ;
        RECT 98.580 310.200 98.780 317.800 ;
        RECT 99.530 317.600 103.530 317.800 ;
        RECT 103.130 317.000 103.530 317.600 ;
        RECT 99.530 316.800 103.530 317.000 ;
        RECT 103.130 316.200 103.530 316.800 ;
        RECT 99.530 316.000 103.530 316.200 ;
        RECT 103.130 315.400 103.530 316.000 ;
        RECT 99.530 315.200 103.530 315.400 ;
        RECT 103.130 314.600 103.530 315.200 ;
        RECT 99.530 314.400 103.530 314.600 ;
        RECT 103.130 313.800 103.530 314.400 ;
        RECT 99.530 313.600 103.530 313.800 ;
        RECT 103.130 313.000 103.530 313.600 ;
        RECT 99.530 312.800 103.530 313.000 ;
        RECT 103.130 312.200 103.530 312.800 ;
        RECT 99.530 312.000 103.530 312.200 ;
        RECT 103.130 311.400 103.530 312.000 ;
        RECT 99.530 311.200 103.530 311.400 ;
        RECT 103.130 310.600 103.530 311.200 ;
        RECT 99.530 310.400 103.530 310.600 ;
        RECT 103.130 310.200 103.530 310.400 ;
        RECT 95.380 309.800 103.530 310.200 ;
        RECT 95.380 302.200 95.580 309.800 ;
        RECT 96.180 302.200 96.380 309.800 ;
        RECT 96.980 302.200 97.180 309.800 ;
        RECT 97.780 302.200 97.980 309.800 ;
        RECT 98.580 302.200 98.780 309.800 ;
        RECT 103.130 309.600 103.530 309.800 ;
        RECT 99.530 309.400 103.530 309.600 ;
        RECT 103.130 308.800 103.530 309.400 ;
        RECT 99.530 308.600 103.530 308.800 ;
        RECT 103.130 308.000 103.530 308.600 ;
        RECT 99.530 307.800 103.530 308.000 ;
        RECT 103.130 307.200 103.530 307.800 ;
        RECT 99.530 307.000 103.530 307.200 ;
        RECT 103.130 306.400 103.530 307.000 ;
        RECT 99.530 306.200 103.530 306.400 ;
        RECT 103.130 305.600 103.530 306.200 ;
        RECT 99.530 305.400 103.530 305.600 ;
        RECT 103.130 304.800 103.530 305.400 ;
        RECT 99.530 304.600 103.530 304.800 ;
        RECT 103.130 304.000 103.530 304.600 ;
        RECT 99.530 303.800 103.530 304.000 ;
        RECT 103.130 303.200 103.530 303.800 ;
        RECT 99.530 303.000 103.530 303.200 ;
        RECT 103.130 302.400 103.530 303.000 ;
        RECT 99.530 302.200 103.530 302.400 ;
        RECT 105.930 317.600 109.930 317.800 ;
        RECT 105.930 317.000 106.330 317.600 ;
        RECT 105.930 316.800 109.930 317.000 ;
        RECT 105.930 316.200 106.330 316.800 ;
        RECT 105.930 316.000 109.930 316.200 ;
        RECT 105.930 315.400 106.330 316.000 ;
        RECT 105.930 315.200 109.930 315.400 ;
        RECT 105.930 314.600 106.330 315.200 ;
        RECT 105.930 314.400 109.930 314.600 ;
        RECT 105.930 313.800 106.330 314.400 ;
        RECT 105.930 313.600 109.930 313.800 ;
        RECT 105.930 313.000 106.330 313.600 ;
        RECT 105.930 312.800 109.930 313.000 ;
        RECT 105.930 312.200 106.330 312.800 ;
        RECT 105.930 312.000 109.930 312.200 ;
        RECT 105.930 311.400 106.330 312.000 ;
        RECT 105.930 311.200 109.930 311.400 ;
        RECT 105.930 310.600 106.330 311.200 ;
        RECT 105.930 310.400 109.930 310.600 ;
        RECT 105.930 310.200 106.330 310.400 ;
        RECT 110.680 310.200 110.880 317.800 ;
        RECT 111.480 310.200 111.680 317.800 ;
        RECT 112.280 310.200 112.480 317.800 ;
        RECT 113.080 310.200 113.280 317.800 ;
        RECT 113.880 310.200 114.080 317.800 ;
        RECT 105.930 309.800 114.080 310.200 ;
        RECT 105.930 309.600 106.330 309.800 ;
        RECT 105.930 309.400 109.930 309.600 ;
        RECT 105.930 308.800 106.330 309.400 ;
        RECT 105.930 308.600 109.930 308.800 ;
        RECT 105.930 308.000 106.330 308.600 ;
        RECT 105.930 307.800 109.930 308.000 ;
        RECT 105.930 307.200 106.330 307.800 ;
        RECT 105.930 307.000 109.930 307.200 ;
        RECT 105.930 306.400 106.330 307.000 ;
        RECT 105.930 306.200 109.930 306.400 ;
        RECT 105.930 305.600 106.330 306.200 ;
        RECT 105.930 305.400 109.930 305.600 ;
        RECT 105.930 304.800 106.330 305.400 ;
        RECT 105.930 304.600 109.930 304.800 ;
        RECT 105.930 304.000 106.330 304.600 ;
        RECT 105.930 303.800 109.930 304.000 ;
        RECT 105.930 303.200 106.330 303.800 ;
        RECT 105.930 303.000 109.930 303.200 ;
        RECT 105.930 302.400 106.330 303.000 ;
        RECT 105.930 302.200 109.930 302.400 ;
        RECT 110.680 302.200 110.880 309.800 ;
        RECT 111.480 302.200 111.680 309.800 ;
        RECT 112.280 302.200 112.480 309.800 ;
        RECT 113.080 302.200 113.280 309.800 ;
        RECT 113.880 302.200 114.080 309.800 ;
        RECT 115.380 310.200 115.580 317.800 ;
        RECT 116.180 310.200 116.380 317.800 ;
        RECT 116.980 310.200 117.180 317.800 ;
        RECT 117.780 310.200 117.980 317.800 ;
        RECT 118.580 310.200 118.780 317.800 ;
        RECT 119.530 317.600 123.530 317.800 ;
        RECT 123.130 317.000 123.530 317.600 ;
        RECT 119.530 316.800 123.530 317.000 ;
        RECT 123.130 316.200 123.530 316.800 ;
        RECT 119.530 316.000 123.530 316.200 ;
        RECT 123.130 315.400 123.530 316.000 ;
        RECT 119.530 315.200 123.530 315.400 ;
        RECT 123.130 314.600 123.530 315.200 ;
        RECT 119.530 314.400 123.530 314.600 ;
        RECT 123.130 313.800 123.530 314.400 ;
        RECT 119.530 313.600 123.530 313.800 ;
        RECT 123.130 313.000 123.530 313.600 ;
        RECT 119.530 312.800 123.530 313.000 ;
        RECT 123.130 312.200 123.530 312.800 ;
        RECT 119.530 312.000 123.530 312.200 ;
        RECT 123.130 311.400 123.530 312.000 ;
        RECT 119.530 311.200 123.530 311.400 ;
        RECT 123.130 310.600 123.530 311.200 ;
        RECT 119.530 310.400 123.530 310.600 ;
        RECT 123.130 310.200 123.530 310.400 ;
        RECT 115.380 309.800 123.530 310.200 ;
        RECT 130.050 309.910 130.410 310.290 ;
        RECT 130.680 309.910 131.040 310.290 ;
        RECT 131.280 309.910 131.640 310.290 ;
        RECT 115.380 302.200 115.580 309.800 ;
        RECT 116.180 302.200 116.380 309.800 ;
        RECT 116.980 302.200 117.180 309.800 ;
        RECT 117.780 302.200 117.980 309.800 ;
        RECT 118.580 302.200 118.780 309.800 ;
        RECT 123.130 309.600 123.530 309.800 ;
        RECT 119.530 309.400 123.530 309.600 ;
        RECT 123.130 308.800 123.530 309.400 ;
        RECT 130.050 309.320 130.410 309.700 ;
        RECT 130.680 309.320 131.040 309.700 ;
        RECT 131.280 309.320 131.640 309.700 ;
        RECT 119.530 308.600 123.530 308.800 ;
        RECT 123.130 308.000 123.530 308.600 ;
        RECT 119.530 307.800 123.530 308.000 ;
        RECT 123.130 307.200 123.530 307.800 ;
        RECT 119.530 307.000 123.530 307.200 ;
        RECT 123.130 306.400 123.530 307.000 ;
        RECT 119.530 306.200 123.530 306.400 ;
        RECT 123.130 305.600 123.530 306.200 ;
        RECT 119.530 305.400 123.530 305.600 ;
        RECT 123.130 304.800 123.530 305.400 ;
        RECT 119.530 304.600 123.530 304.800 ;
        RECT 123.130 304.000 123.530 304.600 ;
        RECT 119.530 303.800 123.530 304.000 ;
        RECT 123.130 303.200 123.530 303.800 ;
        RECT 119.530 303.000 123.530 303.200 ;
        RECT 123.130 302.400 123.530 303.000 ;
        RECT 119.530 302.200 123.530 302.400 ;
        RECT 5.930 297.600 9.930 297.800 ;
        RECT 5.930 297.000 6.330 297.600 ;
        RECT 5.930 296.800 9.930 297.000 ;
        RECT 5.930 296.200 6.330 296.800 ;
        RECT 5.930 296.000 9.930 296.200 ;
        RECT 5.930 295.400 6.330 296.000 ;
        RECT 5.930 295.200 9.930 295.400 ;
        RECT 5.930 294.600 6.330 295.200 ;
        RECT 5.930 294.400 9.930 294.600 ;
        RECT 5.930 293.800 6.330 294.400 ;
        RECT 5.930 293.600 9.930 293.800 ;
        RECT 5.930 293.000 6.330 293.600 ;
        RECT 5.930 292.800 9.930 293.000 ;
        RECT 5.930 292.200 6.330 292.800 ;
        RECT 5.930 292.000 9.930 292.200 ;
        RECT 5.930 291.400 6.330 292.000 ;
        RECT 5.930 291.200 9.930 291.400 ;
        RECT 5.930 290.600 6.330 291.200 ;
        RECT 5.930 290.400 9.930 290.600 ;
        RECT 5.930 290.200 6.330 290.400 ;
        RECT 10.680 290.200 10.880 297.800 ;
        RECT 11.480 290.200 11.680 297.800 ;
        RECT 12.280 290.200 12.480 297.800 ;
        RECT 13.080 290.200 13.280 297.800 ;
        RECT 13.880 290.200 14.080 297.800 ;
        RECT 5.930 289.800 14.080 290.200 ;
        RECT 5.930 289.600 6.330 289.800 ;
        RECT 5.930 289.400 9.930 289.600 ;
        RECT 5.930 288.800 6.330 289.400 ;
        RECT 5.930 288.600 9.930 288.800 ;
        RECT 5.930 288.000 6.330 288.600 ;
        RECT 5.930 287.800 9.930 288.000 ;
        RECT 5.930 287.200 6.330 287.800 ;
        RECT 5.930 287.000 9.930 287.200 ;
        RECT 5.930 286.400 6.330 287.000 ;
        RECT 5.930 286.200 9.930 286.400 ;
        RECT 5.930 285.600 6.330 286.200 ;
        RECT 5.930 285.400 9.930 285.600 ;
        RECT 5.930 284.800 6.330 285.400 ;
        RECT 5.930 284.600 9.930 284.800 ;
        RECT 5.930 284.000 6.330 284.600 ;
        RECT 5.930 283.800 9.930 284.000 ;
        RECT 5.930 283.200 6.330 283.800 ;
        RECT 5.930 283.000 9.930 283.200 ;
        RECT 5.930 282.400 6.330 283.000 ;
        RECT 5.930 282.200 9.930 282.400 ;
        RECT 10.680 282.200 10.880 289.800 ;
        RECT 11.480 282.200 11.680 289.800 ;
        RECT 12.280 282.200 12.480 289.800 ;
        RECT 13.080 282.200 13.280 289.800 ;
        RECT 13.880 282.200 14.080 289.800 ;
        RECT 15.380 290.200 15.580 297.800 ;
        RECT 16.180 290.200 16.380 297.800 ;
        RECT 16.980 290.200 17.180 297.800 ;
        RECT 17.780 290.200 17.980 297.800 ;
        RECT 18.580 290.200 18.780 297.800 ;
        RECT 19.530 297.600 23.530 297.800 ;
        RECT 23.130 297.000 23.530 297.600 ;
        RECT 19.530 296.800 23.530 297.000 ;
        RECT 23.130 296.200 23.530 296.800 ;
        RECT 19.530 296.000 23.530 296.200 ;
        RECT 23.130 295.400 23.530 296.000 ;
        RECT 19.530 295.200 23.530 295.400 ;
        RECT 23.130 294.600 23.530 295.200 ;
        RECT 19.530 294.400 23.530 294.600 ;
        RECT 23.130 293.800 23.530 294.400 ;
        RECT 19.530 293.600 23.530 293.800 ;
        RECT 23.130 293.000 23.530 293.600 ;
        RECT 19.530 292.800 23.530 293.000 ;
        RECT 23.130 292.200 23.530 292.800 ;
        RECT 19.530 292.000 23.530 292.200 ;
        RECT 23.130 291.400 23.530 292.000 ;
        RECT 19.530 291.200 23.530 291.400 ;
        RECT 23.130 290.600 23.530 291.200 ;
        RECT 19.530 290.400 23.530 290.600 ;
        RECT 23.130 290.200 23.530 290.400 ;
        RECT 15.380 289.800 23.530 290.200 ;
        RECT 15.380 282.200 15.580 289.800 ;
        RECT 16.180 282.200 16.380 289.800 ;
        RECT 16.980 282.200 17.180 289.800 ;
        RECT 17.780 282.200 17.980 289.800 ;
        RECT 18.580 282.200 18.780 289.800 ;
        RECT 23.130 289.600 23.530 289.800 ;
        RECT 19.530 289.400 23.530 289.600 ;
        RECT 23.130 288.800 23.530 289.400 ;
        RECT 19.530 288.600 23.530 288.800 ;
        RECT 23.130 288.000 23.530 288.600 ;
        RECT 19.530 287.800 23.530 288.000 ;
        RECT 23.130 287.200 23.530 287.800 ;
        RECT 19.530 287.000 23.530 287.200 ;
        RECT 23.130 286.400 23.530 287.000 ;
        RECT 19.530 286.200 23.530 286.400 ;
        RECT 23.130 285.600 23.530 286.200 ;
        RECT 19.530 285.400 23.530 285.600 ;
        RECT 23.130 284.800 23.530 285.400 ;
        RECT 19.530 284.600 23.530 284.800 ;
        RECT 23.130 284.000 23.530 284.600 ;
        RECT 19.530 283.800 23.530 284.000 ;
        RECT 23.130 283.200 23.530 283.800 ;
        RECT 19.530 283.000 23.530 283.200 ;
        RECT 23.130 282.400 23.530 283.000 ;
        RECT 19.530 282.200 23.530 282.400 ;
        RECT 25.930 297.600 29.930 297.800 ;
        RECT 25.930 297.000 26.330 297.600 ;
        RECT 25.930 296.800 29.930 297.000 ;
        RECT 25.930 296.200 26.330 296.800 ;
        RECT 25.930 296.000 29.930 296.200 ;
        RECT 25.930 295.400 26.330 296.000 ;
        RECT 25.930 295.200 29.930 295.400 ;
        RECT 25.930 294.600 26.330 295.200 ;
        RECT 25.930 294.400 29.930 294.600 ;
        RECT 25.930 293.800 26.330 294.400 ;
        RECT 25.930 293.600 29.930 293.800 ;
        RECT 25.930 293.000 26.330 293.600 ;
        RECT 25.930 292.800 29.930 293.000 ;
        RECT 25.930 292.200 26.330 292.800 ;
        RECT 25.930 292.000 29.930 292.200 ;
        RECT 25.930 291.400 26.330 292.000 ;
        RECT 25.930 291.200 29.930 291.400 ;
        RECT 25.930 290.600 26.330 291.200 ;
        RECT 25.930 290.400 29.930 290.600 ;
        RECT 25.930 290.200 26.330 290.400 ;
        RECT 30.680 290.200 30.880 297.800 ;
        RECT 31.480 290.200 31.680 297.800 ;
        RECT 32.280 290.200 32.480 297.800 ;
        RECT 33.080 290.200 33.280 297.800 ;
        RECT 33.880 290.200 34.080 297.800 ;
        RECT 25.930 289.800 34.080 290.200 ;
        RECT 25.930 289.600 26.330 289.800 ;
        RECT 25.930 289.400 29.930 289.600 ;
        RECT 25.930 288.800 26.330 289.400 ;
        RECT 25.930 288.600 29.930 288.800 ;
        RECT 25.930 288.000 26.330 288.600 ;
        RECT 25.930 287.800 29.930 288.000 ;
        RECT 25.930 287.200 26.330 287.800 ;
        RECT 25.930 287.000 29.930 287.200 ;
        RECT 25.930 286.400 26.330 287.000 ;
        RECT 25.930 286.200 29.930 286.400 ;
        RECT 25.930 285.600 26.330 286.200 ;
        RECT 25.930 285.400 29.930 285.600 ;
        RECT 25.930 284.800 26.330 285.400 ;
        RECT 25.930 284.600 29.930 284.800 ;
        RECT 25.930 284.000 26.330 284.600 ;
        RECT 25.930 283.800 29.930 284.000 ;
        RECT 25.930 283.200 26.330 283.800 ;
        RECT 25.930 283.000 29.930 283.200 ;
        RECT 25.930 282.400 26.330 283.000 ;
        RECT 25.930 282.200 29.930 282.400 ;
        RECT 30.680 282.200 30.880 289.800 ;
        RECT 31.480 282.200 31.680 289.800 ;
        RECT 32.280 282.200 32.480 289.800 ;
        RECT 33.080 282.200 33.280 289.800 ;
        RECT 33.880 282.200 34.080 289.800 ;
        RECT 35.380 290.200 35.580 297.800 ;
        RECT 36.180 290.200 36.380 297.800 ;
        RECT 36.980 290.200 37.180 297.800 ;
        RECT 37.780 290.200 37.980 297.800 ;
        RECT 38.580 290.200 38.780 297.800 ;
        RECT 39.530 297.600 43.530 297.800 ;
        RECT 43.130 297.000 43.530 297.600 ;
        RECT 39.530 296.800 43.530 297.000 ;
        RECT 43.130 296.200 43.530 296.800 ;
        RECT 39.530 296.000 43.530 296.200 ;
        RECT 43.130 295.400 43.530 296.000 ;
        RECT 39.530 295.200 43.530 295.400 ;
        RECT 43.130 294.600 43.530 295.200 ;
        RECT 39.530 294.400 43.530 294.600 ;
        RECT 43.130 293.800 43.530 294.400 ;
        RECT 39.530 293.600 43.530 293.800 ;
        RECT 43.130 293.000 43.530 293.600 ;
        RECT 39.530 292.800 43.530 293.000 ;
        RECT 43.130 292.200 43.530 292.800 ;
        RECT 39.530 292.000 43.530 292.200 ;
        RECT 43.130 291.400 43.530 292.000 ;
        RECT 39.530 291.200 43.530 291.400 ;
        RECT 43.130 290.600 43.530 291.200 ;
        RECT 39.530 290.400 43.530 290.600 ;
        RECT 43.130 290.200 43.530 290.400 ;
        RECT 35.380 289.800 43.530 290.200 ;
        RECT 35.380 282.200 35.580 289.800 ;
        RECT 36.180 282.200 36.380 289.800 ;
        RECT 36.980 282.200 37.180 289.800 ;
        RECT 37.780 282.200 37.980 289.800 ;
        RECT 38.580 282.200 38.780 289.800 ;
        RECT 43.130 289.600 43.530 289.800 ;
        RECT 39.530 289.400 43.530 289.600 ;
        RECT 43.130 288.800 43.530 289.400 ;
        RECT 39.530 288.600 43.530 288.800 ;
        RECT 43.130 288.000 43.530 288.600 ;
        RECT 39.530 287.800 43.530 288.000 ;
        RECT 43.130 287.200 43.530 287.800 ;
        RECT 39.530 287.000 43.530 287.200 ;
        RECT 43.130 286.400 43.530 287.000 ;
        RECT 39.530 286.200 43.530 286.400 ;
        RECT 43.130 285.600 43.530 286.200 ;
        RECT 39.530 285.400 43.530 285.600 ;
        RECT 43.130 284.800 43.530 285.400 ;
        RECT 39.530 284.600 43.530 284.800 ;
        RECT 43.130 284.000 43.530 284.600 ;
        RECT 39.530 283.800 43.530 284.000 ;
        RECT 43.130 283.200 43.530 283.800 ;
        RECT 39.530 283.000 43.530 283.200 ;
        RECT 43.130 282.400 43.530 283.000 ;
        RECT 39.530 282.200 43.530 282.400 ;
        RECT 45.930 297.600 49.930 297.800 ;
        RECT 45.930 297.000 46.330 297.600 ;
        RECT 45.930 296.800 49.930 297.000 ;
        RECT 45.930 296.200 46.330 296.800 ;
        RECT 45.930 296.000 49.930 296.200 ;
        RECT 45.930 295.400 46.330 296.000 ;
        RECT 45.930 295.200 49.930 295.400 ;
        RECT 45.930 294.600 46.330 295.200 ;
        RECT 45.930 294.400 49.930 294.600 ;
        RECT 45.930 293.800 46.330 294.400 ;
        RECT 45.930 293.600 49.930 293.800 ;
        RECT 45.930 293.000 46.330 293.600 ;
        RECT 45.930 292.800 49.930 293.000 ;
        RECT 45.930 292.200 46.330 292.800 ;
        RECT 45.930 292.000 49.930 292.200 ;
        RECT 45.930 291.400 46.330 292.000 ;
        RECT 45.930 291.200 49.930 291.400 ;
        RECT 45.930 290.600 46.330 291.200 ;
        RECT 45.930 290.400 49.930 290.600 ;
        RECT 45.930 290.200 46.330 290.400 ;
        RECT 50.680 290.200 50.880 297.800 ;
        RECT 51.480 290.200 51.680 297.800 ;
        RECT 52.280 290.200 52.480 297.800 ;
        RECT 53.080 290.200 53.280 297.800 ;
        RECT 53.880 290.200 54.080 297.800 ;
        RECT 45.930 289.800 54.080 290.200 ;
        RECT 45.930 289.600 46.330 289.800 ;
        RECT 45.930 289.400 49.930 289.600 ;
        RECT 45.930 288.800 46.330 289.400 ;
        RECT 45.930 288.600 49.930 288.800 ;
        RECT 45.930 288.000 46.330 288.600 ;
        RECT 45.930 287.800 49.930 288.000 ;
        RECT 45.930 287.200 46.330 287.800 ;
        RECT 45.930 287.000 49.930 287.200 ;
        RECT 45.930 286.400 46.330 287.000 ;
        RECT 45.930 286.200 49.930 286.400 ;
        RECT 45.930 285.600 46.330 286.200 ;
        RECT 45.930 285.400 49.930 285.600 ;
        RECT 45.930 284.800 46.330 285.400 ;
        RECT 45.930 284.600 49.930 284.800 ;
        RECT 45.930 284.000 46.330 284.600 ;
        RECT 45.930 283.800 49.930 284.000 ;
        RECT 45.930 283.200 46.330 283.800 ;
        RECT 45.930 283.000 49.930 283.200 ;
        RECT 45.930 282.400 46.330 283.000 ;
        RECT 45.930 282.200 49.930 282.400 ;
        RECT 50.680 282.200 50.880 289.800 ;
        RECT 51.480 282.200 51.680 289.800 ;
        RECT 52.280 282.200 52.480 289.800 ;
        RECT 53.080 282.200 53.280 289.800 ;
        RECT 53.880 282.200 54.080 289.800 ;
        RECT 55.380 290.200 55.580 297.800 ;
        RECT 56.180 290.200 56.380 297.800 ;
        RECT 56.980 290.200 57.180 297.800 ;
        RECT 57.780 290.200 57.980 297.800 ;
        RECT 58.580 290.200 58.780 297.800 ;
        RECT 59.530 297.600 63.530 297.800 ;
        RECT 63.130 297.000 63.530 297.600 ;
        RECT 59.530 296.800 63.530 297.000 ;
        RECT 63.130 296.200 63.530 296.800 ;
        RECT 59.530 296.000 63.530 296.200 ;
        RECT 63.130 295.400 63.530 296.000 ;
        RECT 59.530 295.200 63.530 295.400 ;
        RECT 63.130 294.600 63.530 295.200 ;
        RECT 59.530 294.400 63.530 294.600 ;
        RECT 63.130 293.800 63.530 294.400 ;
        RECT 59.530 293.600 63.530 293.800 ;
        RECT 63.130 293.000 63.530 293.600 ;
        RECT 59.530 292.800 63.530 293.000 ;
        RECT 63.130 292.200 63.530 292.800 ;
        RECT 59.530 292.000 63.530 292.200 ;
        RECT 63.130 291.400 63.530 292.000 ;
        RECT 59.530 291.200 63.530 291.400 ;
        RECT 63.130 290.600 63.530 291.200 ;
        RECT 59.530 290.400 63.530 290.600 ;
        RECT 63.130 290.200 63.530 290.400 ;
        RECT 55.380 289.800 63.530 290.200 ;
        RECT 55.380 282.200 55.580 289.800 ;
        RECT 56.180 282.200 56.380 289.800 ;
        RECT 56.980 282.200 57.180 289.800 ;
        RECT 57.780 282.200 57.980 289.800 ;
        RECT 58.580 282.200 58.780 289.800 ;
        RECT 63.130 289.600 63.530 289.800 ;
        RECT 59.530 289.400 63.530 289.600 ;
        RECT 63.130 288.800 63.530 289.400 ;
        RECT 59.530 288.600 63.530 288.800 ;
        RECT 63.130 288.000 63.530 288.600 ;
        RECT 59.530 287.800 63.530 288.000 ;
        RECT 63.130 287.200 63.530 287.800 ;
        RECT 59.530 287.000 63.530 287.200 ;
        RECT 63.130 286.400 63.530 287.000 ;
        RECT 59.530 286.200 63.530 286.400 ;
        RECT 63.130 285.600 63.530 286.200 ;
        RECT 59.530 285.400 63.530 285.600 ;
        RECT 63.130 284.800 63.530 285.400 ;
        RECT 59.530 284.600 63.530 284.800 ;
        RECT 63.130 284.000 63.530 284.600 ;
        RECT 59.530 283.800 63.530 284.000 ;
        RECT 63.130 283.200 63.530 283.800 ;
        RECT 59.530 283.000 63.530 283.200 ;
        RECT 63.130 282.400 63.530 283.000 ;
        RECT 59.530 282.200 63.530 282.400 ;
        RECT 65.930 297.600 69.930 297.800 ;
        RECT 65.930 297.000 66.330 297.600 ;
        RECT 65.930 296.800 69.930 297.000 ;
        RECT 65.930 296.200 66.330 296.800 ;
        RECT 65.930 296.000 69.930 296.200 ;
        RECT 65.930 295.400 66.330 296.000 ;
        RECT 65.930 295.200 69.930 295.400 ;
        RECT 65.930 294.600 66.330 295.200 ;
        RECT 65.930 294.400 69.930 294.600 ;
        RECT 65.930 293.800 66.330 294.400 ;
        RECT 65.930 293.600 69.930 293.800 ;
        RECT 65.930 293.000 66.330 293.600 ;
        RECT 65.930 292.800 69.930 293.000 ;
        RECT 65.930 292.200 66.330 292.800 ;
        RECT 65.930 292.000 69.930 292.200 ;
        RECT 65.930 291.400 66.330 292.000 ;
        RECT 65.930 291.200 69.930 291.400 ;
        RECT 65.930 290.600 66.330 291.200 ;
        RECT 65.930 290.400 69.930 290.600 ;
        RECT 65.930 290.200 66.330 290.400 ;
        RECT 70.680 290.200 70.880 297.800 ;
        RECT 71.480 290.200 71.680 297.800 ;
        RECT 72.280 290.200 72.480 297.800 ;
        RECT 73.080 290.200 73.280 297.800 ;
        RECT 73.880 290.200 74.080 297.800 ;
        RECT 65.930 289.800 74.080 290.200 ;
        RECT 65.930 289.600 66.330 289.800 ;
        RECT 65.930 289.400 69.930 289.600 ;
        RECT 65.930 288.800 66.330 289.400 ;
        RECT 65.930 288.600 69.930 288.800 ;
        RECT 65.930 288.000 66.330 288.600 ;
        RECT 65.930 287.800 69.930 288.000 ;
        RECT 65.930 287.200 66.330 287.800 ;
        RECT 65.930 287.000 69.930 287.200 ;
        RECT 65.930 286.400 66.330 287.000 ;
        RECT 65.930 286.200 69.930 286.400 ;
        RECT 65.930 285.600 66.330 286.200 ;
        RECT 65.930 285.400 69.930 285.600 ;
        RECT 65.930 284.800 66.330 285.400 ;
        RECT 65.930 284.600 69.930 284.800 ;
        RECT 65.930 284.000 66.330 284.600 ;
        RECT 65.930 283.800 69.930 284.000 ;
        RECT 65.930 283.200 66.330 283.800 ;
        RECT 65.930 283.000 69.930 283.200 ;
        RECT 65.930 282.400 66.330 283.000 ;
        RECT 65.930 282.200 69.930 282.400 ;
        RECT 70.680 282.200 70.880 289.800 ;
        RECT 71.480 282.200 71.680 289.800 ;
        RECT 72.280 282.200 72.480 289.800 ;
        RECT 73.080 282.200 73.280 289.800 ;
        RECT 73.880 282.200 74.080 289.800 ;
        RECT 75.380 290.200 75.580 297.800 ;
        RECT 76.180 290.200 76.380 297.800 ;
        RECT 76.980 290.200 77.180 297.800 ;
        RECT 77.780 290.200 77.980 297.800 ;
        RECT 78.580 290.200 78.780 297.800 ;
        RECT 79.530 297.600 83.530 297.800 ;
        RECT 83.130 297.000 83.530 297.600 ;
        RECT 79.530 296.800 83.530 297.000 ;
        RECT 83.130 296.200 83.530 296.800 ;
        RECT 79.530 296.000 83.530 296.200 ;
        RECT 83.130 295.400 83.530 296.000 ;
        RECT 79.530 295.200 83.530 295.400 ;
        RECT 83.130 294.600 83.530 295.200 ;
        RECT 79.530 294.400 83.530 294.600 ;
        RECT 83.130 293.800 83.530 294.400 ;
        RECT 79.530 293.600 83.530 293.800 ;
        RECT 83.130 293.000 83.530 293.600 ;
        RECT 79.530 292.800 83.530 293.000 ;
        RECT 83.130 292.200 83.530 292.800 ;
        RECT 79.530 292.000 83.530 292.200 ;
        RECT 83.130 291.400 83.530 292.000 ;
        RECT 79.530 291.200 83.530 291.400 ;
        RECT 83.130 290.600 83.530 291.200 ;
        RECT 79.530 290.400 83.530 290.600 ;
        RECT 83.130 290.200 83.530 290.400 ;
        RECT 75.380 289.800 83.530 290.200 ;
        RECT 75.380 282.200 75.580 289.800 ;
        RECT 76.180 282.200 76.380 289.800 ;
        RECT 76.980 282.200 77.180 289.800 ;
        RECT 77.780 282.200 77.980 289.800 ;
        RECT 78.580 282.200 78.780 289.800 ;
        RECT 83.130 289.600 83.530 289.800 ;
        RECT 79.530 289.400 83.530 289.600 ;
        RECT 83.130 288.800 83.530 289.400 ;
        RECT 79.530 288.600 83.530 288.800 ;
        RECT 83.130 288.000 83.530 288.600 ;
        RECT 79.530 287.800 83.530 288.000 ;
        RECT 83.130 287.200 83.530 287.800 ;
        RECT 79.530 287.000 83.530 287.200 ;
        RECT 83.130 286.400 83.530 287.000 ;
        RECT 79.530 286.200 83.530 286.400 ;
        RECT 83.130 285.600 83.530 286.200 ;
        RECT 79.530 285.400 83.530 285.600 ;
        RECT 83.130 284.800 83.530 285.400 ;
        RECT 79.530 284.600 83.530 284.800 ;
        RECT 83.130 284.000 83.530 284.600 ;
        RECT 79.530 283.800 83.530 284.000 ;
        RECT 83.130 283.200 83.530 283.800 ;
        RECT 79.530 283.000 83.530 283.200 ;
        RECT 83.130 282.400 83.530 283.000 ;
        RECT 79.530 282.200 83.530 282.400 ;
        RECT 85.930 297.600 89.930 297.800 ;
        RECT 85.930 297.000 86.330 297.600 ;
        RECT 85.930 296.800 89.930 297.000 ;
        RECT 85.930 296.200 86.330 296.800 ;
        RECT 85.930 296.000 89.930 296.200 ;
        RECT 85.930 295.400 86.330 296.000 ;
        RECT 85.930 295.200 89.930 295.400 ;
        RECT 85.930 294.600 86.330 295.200 ;
        RECT 85.930 294.400 89.930 294.600 ;
        RECT 85.930 293.800 86.330 294.400 ;
        RECT 85.930 293.600 89.930 293.800 ;
        RECT 85.930 293.000 86.330 293.600 ;
        RECT 85.930 292.800 89.930 293.000 ;
        RECT 85.930 292.200 86.330 292.800 ;
        RECT 85.930 292.000 89.930 292.200 ;
        RECT 85.930 291.400 86.330 292.000 ;
        RECT 85.930 291.200 89.930 291.400 ;
        RECT 85.930 290.600 86.330 291.200 ;
        RECT 85.930 290.400 89.930 290.600 ;
        RECT 85.930 290.200 86.330 290.400 ;
        RECT 90.680 290.200 90.880 297.800 ;
        RECT 91.480 290.200 91.680 297.800 ;
        RECT 92.280 290.200 92.480 297.800 ;
        RECT 93.080 290.200 93.280 297.800 ;
        RECT 93.880 290.200 94.080 297.800 ;
        RECT 85.930 289.800 94.080 290.200 ;
        RECT 85.930 289.600 86.330 289.800 ;
        RECT 85.930 289.400 89.930 289.600 ;
        RECT 85.930 288.800 86.330 289.400 ;
        RECT 85.930 288.600 89.930 288.800 ;
        RECT 85.930 288.000 86.330 288.600 ;
        RECT 85.930 287.800 89.930 288.000 ;
        RECT 85.930 287.200 86.330 287.800 ;
        RECT 85.930 287.000 89.930 287.200 ;
        RECT 85.930 286.400 86.330 287.000 ;
        RECT 85.930 286.200 89.930 286.400 ;
        RECT 85.930 285.600 86.330 286.200 ;
        RECT 85.930 285.400 89.930 285.600 ;
        RECT 85.930 284.800 86.330 285.400 ;
        RECT 85.930 284.600 89.930 284.800 ;
        RECT 85.930 284.000 86.330 284.600 ;
        RECT 85.930 283.800 89.930 284.000 ;
        RECT 85.930 283.200 86.330 283.800 ;
        RECT 85.930 283.000 89.930 283.200 ;
        RECT 85.930 282.400 86.330 283.000 ;
        RECT 85.930 282.200 89.930 282.400 ;
        RECT 90.680 282.200 90.880 289.800 ;
        RECT 91.480 282.200 91.680 289.800 ;
        RECT 92.280 282.200 92.480 289.800 ;
        RECT 93.080 282.200 93.280 289.800 ;
        RECT 93.880 282.200 94.080 289.800 ;
        RECT 95.380 290.200 95.580 297.800 ;
        RECT 96.180 290.200 96.380 297.800 ;
        RECT 96.980 290.200 97.180 297.800 ;
        RECT 97.780 290.200 97.980 297.800 ;
        RECT 98.580 290.200 98.780 297.800 ;
        RECT 99.530 297.600 103.530 297.800 ;
        RECT 103.130 297.000 103.530 297.600 ;
        RECT 99.530 296.800 103.530 297.000 ;
        RECT 103.130 296.200 103.530 296.800 ;
        RECT 99.530 296.000 103.530 296.200 ;
        RECT 103.130 295.400 103.530 296.000 ;
        RECT 99.530 295.200 103.530 295.400 ;
        RECT 103.130 294.600 103.530 295.200 ;
        RECT 99.530 294.400 103.530 294.600 ;
        RECT 103.130 293.800 103.530 294.400 ;
        RECT 99.530 293.600 103.530 293.800 ;
        RECT 103.130 293.000 103.530 293.600 ;
        RECT 99.530 292.800 103.530 293.000 ;
        RECT 103.130 292.200 103.530 292.800 ;
        RECT 99.530 292.000 103.530 292.200 ;
        RECT 103.130 291.400 103.530 292.000 ;
        RECT 99.530 291.200 103.530 291.400 ;
        RECT 103.130 290.600 103.530 291.200 ;
        RECT 99.530 290.400 103.530 290.600 ;
        RECT 103.130 290.200 103.530 290.400 ;
        RECT 95.380 289.800 103.530 290.200 ;
        RECT 95.380 282.200 95.580 289.800 ;
        RECT 96.180 282.200 96.380 289.800 ;
        RECT 96.980 282.200 97.180 289.800 ;
        RECT 97.780 282.200 97.980 289.800 ;
        RECT 98.580 282.200 98.780 289.800 ;
        RECT 103.130 289.600 103.530 289.800 ;
        RECT 99.530 289.400 103.530 289.600 ;
        RECT 103.130 288.800 103.530 289.400 ;
        RECT 99.530 288.600 103.530 288.800 ;
        RECT 103.130 288.000 103.530 288.600 ;
        RECT 99.530 287.800 103.530 288.000 ;
        RECT 103.130 287.200 103.530 287.800 ;
        RECT 99.530 287.000 103.530 287.200 ;
        RECT 103.130 286.400 103.530 287.000 ;
        RECT 99.530 286.200 103.530 286.400 ;
        RECT 103.130 285.600 103.530 286.200 ;
        RECT 99.530 285.400 103.530 285.600 ;
        RECT 103.130 284.800 103.530 285.400 ;
        RECT 99.530 284.600 103.530 284.800 ;
        RECT 103.130 284.000 103.530 284.600 ;
        RECT 99.530 283.800 103.530 284.000 ;
        RECT 103.130 283.200 103.530 283.800 ;
        RECT 99.530 283.000 103.530 283.200 ;
        RECT 103.130 282.400 103.530 283.000 ;
        RECT 99.530 282.200 103.530 282.400 ;
        RECT 105.930 297.600 109.930 297.800 ;
        RECT 105.930 297.000 106.330 297.600 ;
        RECT 105.930 296.800 109.930 297.000 ;
        RECT 105.930 296.200 106.330 296.800 ;
        RECT 105.930 296.000 109.930 296.200 ;
        RECT 105.930 295.400 106.330 296.000 ;
        RECT 105.930 295.200 109.930 295.400 ;
        RECT 105.930 294.600 106.330 295.200 ;
        RECT 105.930 294.400 109.930 294.600 ;
        RECT 105.930 293.800 106.330 294.400 ;
        RECT 105.930 293.600 109.930 293.800 ;
        RECT 105.930 293.000 106.330 293.600 ;
        RECT 105.930 292.800 109.930 293.000 ;
        RECT 105.930 292.200 106.330 292.800 ;
        RECT 105.930 292.000 109.930 292.200 ;
        RECT 105.930 291.400 106.330 292.000 ;
        RECT 105.930 291.200 109.930 291.400 ;
        RECT 105.930 290.600 106.330 291.200 ;
        RECT 105.930 290.400 109.930 290.600 ;
        RECT 105.930 290.200 106.330 290.400 ;
        RECT 110.680 290.200 110.880 297.800 ;
        RECT 111.480 290.200 111.680 297.800 ;
        RECT 112.280 290.200 112.480 297.800 ;
        RECT 113.080 290.200 113.280 297.800 ;
        RECT 113.880 290.200 114.080 297.800 ;
        RECT 105.930 289.800 114.080 290.200 ;
        RECT 105.930 289.600 106.330 289.800 ;
        RECT 105.930 289.400 109.930 289.600 ;
        RECT 105.930 288.800 106.330 289.400 ;
        RECT 105.930 288.600 109.930 288.800 ;
        RECT 105.930 288.000 106.330 288.600 ;
        RECT 105.930 287.800 109.930 288.000 ;
        RECT 105.930 287.200 106.330 287.800 ;
        RECT 105.930 287.000 109.930 287.200 ;
        RECT 105.930 286.400 106.330 287.000 ;
        RECT 105.930 286.200 109.930 286.400 ;
        RECT 105.930 285.600 106.330 286.200 ;
        RECT 105.930 285.400 109.930 285.600 ;
        RECT 105.930 284.800 106.330 285.400 ;
        RECT 105.930 284.600 109.930 284.800 ;
        RECT 105.930 284.000 106.330 284.600 ;
        RECT 105.930 283.800 109.930 284.000 ;
        RECT 105.930 283.200 106.330 283.800 ;
        RECT 105.930 283.000 109.930 283.200 ;
        RECT 105.930 282.400 106.330 283.000 ;
        RECT 105.930 282.200 109.930 282.400 ;
        RECT 110.680 282.200 110.880 289.800 ;
        RECT 111.480 282.200 111.680 289.800 ;
        RECT 112.280 282.200 112.480 289.800 ;
        RECT 113.080 282.200 113.280 289.800 ;
        RECT 113.880 282.200 114.080 289.800 ;
        RECT 115.380 290.200 115.580 297.800 ;
        RECT 116.180 290.200 116.380 297.800 ;
        RECT 116.980 290.200 117.180 297.800 ;
        RECT 117.780 290.200 117.980 297.800 ;
        RECT 118.580 290.200 118.780 297.800 ;
        RECT 119.530 297.600 123.530 297.800 ;
        RECT 123.130 297.000 123.530 297.600 ;
        RECT 119.530 296.800 123.530 297.000 ;
        RECT 123.130 296.200 123.530 296.800 ;
        RECT 119.530 296.000 123.530 296.200 ;
        RECT 123.130 295.400 123.530 296.000 ;
        RECT 119.530 295.200 123.530 295.400 ;
        RECT 123.130 294.600 123.530 295.200 ;
        RECT 119.530 294.400 123.530 294.600 ;
        RECT 123.130 293.800 123.530 294.400 ;
        RECT 119.530 293.600 123.530 293.800 ;
        RECT 123.130 293.000 123.530 293.600 ;
        RECT 119.530 292.800 123.530 293.000 ;
        RECT 123.130 292.200 123.530 292.800 ;
        RECT 119.530 292.000 123.530 292.200 ;
        RECT 123.130 291.400 123.530 292.000 ;
        RECT 119.530 291.200 123.530 291.400 ;
        RECT 123.130 290.600 123.530 291.200 ;
        RECT 119.530 290.400 123.530 290.600 ;
        RECT 123.130 290.200 123.530 290.400 ;
        RECT 115.380 289.800 123.530 290.200 ;
        RECT 130.050 289.905 130.410 290.285 ;
        RECT 130.680 289.905 131.040 290.285 ;
        RECT 131.280 289.905 131.640 290.285 ;
        RECT 115.380 282.200 115.580 289.800 ;
        RECT 116.180 282.200 116.380 289.800 ;
        RECT 116.980 282.200 117.180 289.800 ;
        RECT 117.780 282.200 117.980 289.800 ;
        RECT 118.580 282.200 118.780 289.800 ;
        RECT 123.130 289.600 123.530 289.800 ;
        RECT 119.530 289.400 123.530 289.600 ;
        RECT 123.130 288.800 123.530 289.400 ;
        RECT 130.050 289.315 130.410 289.695 ;
        RECT 130.680 289.315 131.040 289.695 ;
        RECT 131.280 289.315 131.640 289.695 ;
        RECT 119.530 288.600 123.530 288.800 ;
        RECT 123.130 288.000 123.530 288.600 ;
        RECT 119.530 287.800 123.530 288.000 ;
        RECT 123.130 287.200 123.530 287.800 ;
        RECT 119.530 287.000 123.530 287.200 ;
        RECT 123.130 286.400 123.530 287.000 ;
        RECT 119.530 286.200 123.530 286.400 ;
        RECT 123.130 285.600 123.530 286.200 ;
        RECT 119.530 285.400 123.530 285.600 ;
        RECT 123.130 284.800 123.530 285.400 ;
        RECT 119.530 284.600 123.530 284.800 ;
        RECT 123.130 284.000 123.530 284.600 ;
        RECT 119.530 283.800 123.530 284.000 ;
        RECT 123.130 283.200 123.530 283.800 ;
        RECT 119.530 283.000 123.530 283.200 ;
        RECT 123.130 282.400 123.530 283.000 ;
        RECT 119.530 282.200 123.530 282.400 ;
        RECT 5.930 277.600 9.930 277.800 ;
        RECT 5.930 277.000 6.330 277.600 ;
        RECT 5.930 276.800 9.930 277.000 ;
        RECT 5.930 276.200 6.330 276.800 ;
        RECT 5.930 276.000 9.930 276.200 ;
        RECT 5.930 275.400 6.330 276.000 ;
        RECT 5.930 275.200 9.930 275.400 ;
        RECT 5.930 274.600 6.330 275.200 ;
        RECT 5.930 274.400 9.930 274.600 ;
        RECT 5.930 273.800 6.330 274.400 ;
        RECT 5.930 273.600 9.930 273.800 ;
        RECT 5.930 273.000 6.330 273.600 ;
        RECT 5.930 272.800 9.930 273.000 ;
        RECT 5.930 272.200 6.330 272.800 ;
        RECT 5.930 272.000 9.930 272.200 ;
        RECT 5.930 271.400 6.330 272.000 ;
        RECT 5.930 271.200 9.930 271.400 ;
        RECT 5.930 270.600 6.330 271.200 ;
        RECT 5.930 270.400 9.930 270.600 ;
        RECT 5.930 270.200 6.330 270.400 ;
        RECT 10.680 270.200 10.880 277.800 ;
        RECT 11.480 270.200 11.680 277.800 ;
        RECT 12.280 270.200 12.480 277.800 ;
        RECT 13.080 270.200 13.280 277.800 ;
        RECT 13.880 270.200 14.080 277.800 ;
        RECT 5.930 269.800 14.080 270.200 ;
        RECT 5.930 269.600 6.330 269.800 ;
        RECT 5.930 269.400 9.930 269.600 ;
        RECT 5.930 268.800 6.330 269.400 ;
        RECT 5.930 268.600 9.930 268.800 ;
        RECT 5.930 268.000 6.330 268.600 ;
        RECT 5.930 267.800 9.930 268.000 ;
        RECT 5.930 267.200 6.330 267.800 ;
        RECT 5.930 267.000 9.930 267.200 ;
        RECT 5.930 266.400 6.330 267.000 ;
        RECT 5.930 266.200 9.930 266.400 ;
        RECT 5.930 265.600 6.330 266.200 ;
        RECT 5.930 265.400 9.930 265.600 ;
        RECT 5.930 264.800 6.330 265.400 ;
        RECT 5.930 264.600 9.930 264.800 ;
        RECT 5.930 264.000 6.330 264.600 ;
        RECT 5.930 263.800 9.930 264.000 ;
        RECT 5.930 263.200 6.330 263.800 ;
        RECT 5.930 263.000 9.930 263.200 ;
        RECT 5.930 262.400 6.330 263.000 ;
        RECT 5.930 262.200 9.930 262.400 ;
        RECT 10.680 262.200 10.880 269.800 ;
        RECT 11.480 262.200 11.680 269.800 ;
        RECT 12.280 262.200 12.480 269.800 ;
        RECT 13.080 262.200 13.280 269.800 ;
        RECT 13.880 262.200 14.080 269.800 ;
        RECT 15.380 270.200 15.580 277.800 ;
        RECT 16.180 270.200 16.380 277.800 ;
        RECT 16.980 270.200 17.180 277.800 ;
        RECT 17.780 270.200 17.980 277.800 ;
        RECT 18.580 270.200 18.780 277.800 ;
        RECT 19.530 277.600 23.530 277.800 ;
        RECT 23.130 277.000 23.530 277.600 ;
        RECT 19.530 276.800 23.530 277.000 ;
        RECT 23.130 276.200 23.530 276.800 ;
        RECT 19.530 276.000 23.530 276.200 ;
        RECT 23.130 275.400 23.530 276.000 ;
        RECT 19.530 275.200 23.530 275.400 ;
        RECT 23.130 274.600 23.530 275.200 ;
        RECT 19.530 274.400 23.530 274.600 ;
        RECT 23.130 273.800 23.530 274.400 ;
        RECT 19.530 273.600 23.530 273.800 ;
        RECT 23.130 273.000 23.530 273.600 ;
        RECT 19.530 272.800 23.530 273.000 ;
        RECT 23.130 272.200 23.530 272.800 ;
        RECT 19.530 272.000 23.530 272.200 ;
        RECT 23.130 271.400 23.530 272.000 ;
        RECT 19.530 271.200 23.530 271.400 ;
        RECT 23.130 270.600 23.530 271.200 ;
        RECT 19.530 270.400 23.530 270.600 ;
        RECT 23.130 270.200 23.530 270.400 ;
        RECT 15.380 269.800 23.530 270.200 ;
        RECT 15.380 262.200 15.580 269.800 ;
        RECT 16.180 262.200 16.380 269.800 ;
        RECT 16.980 262.200 17.180 269.800 ;
        RECT 17.780 262.200 17.980 269.800 ;
        RECT 18.580 262.200 18.780 269.800 ;
        RECT 23.130 269.600 23.530 269.800 ;
        RECT 19.530 269.400 23.530 269.600 ;
        RECT 23.130 268.800 23.530 269.400 ;
        RECT 19.530 268.600 23.530 268.800 ;
        RECT 23.130 268.000 23.530 268.600 ;
        RECT 19.530 267.800 23.530 268.000 ;
        RECT 23.130 267.200 23.530 267.800 ;
        RECT 19.530 267.000 23.530 267.200 ;
        RECT 23.130 266.400 23.530 267.000 ;
        RECT 19.530 266.200 23.530 266.400 ;
        RECT 23.130 265.600 23.530 266.200 ;
        RECT 19.530 265.400 23.530 265.600 ;
        RECT 23.130 264.800 23.530 265.400 ;
        RECT 19.530 264.600 23.530 264.800 ;
        RECT 23.130 264.000 23.530 264.600 ;
        RECT 19.530 263.800 23.530 264.000 ;
        RECT 23.130 263.200 23.530 263.800 ;
        RECT 19.530 263.000 23.530 263.200 ;
        RECT 23.130 262.400 23.530 263.000 ;
        RECT 19.530 262.200 23.530 262.400 ;
        RECT 25.930 277.600 29.930 277.800 ;
        RECT 25.930 277.000 26.330 277.600 ;
        RECT 25.930 276.800 29.930 277.000 ;
        RECT 25.930 276.200 26.330 276.800 ;
        RECT 25.930 276.000 29.930 276.200 ;
        RECT 25.930 275.400 26.330 276.000 ;
        RECT 25.930 275.200 29.930 275.400 ;
        RECT 25.930 274.600 26.330 275.200 ;
        RECT 25.930 274.400 29.930 274.600 ;
        RECT 25.930 273.800 26.330 274.400 ;
        RECT 25.930 273.600 29.930 273.800 ;
        RECT 25.930 273.000 26.330 273.600 ;
        RECT 25.930 272.800 29.930 273.000 ;
        RECT 25.930 272.200 26.330 272.800 ;
        RECT 25.930 272.000 29.930 272.200 ;
        RECT 25.930 271.400 26.330 272.000 ;
        RECT 25.930 271.200 29.930 271.400 ;
        RECT 25.930 270.600 26.330 271.200 ;
        RECT 25.930 270.400 29.930 270.600 ;
        RECT 25.930 270.200 26.330 270.400 ;
        RECT 30.680 270.200 30.880 277.800 ;
        RECT 31.480 270.200 31.680 277.800 ;
        RECT 32.280 270.200 32.480 277.800 ;
        RECT 33.080 270.200 33.280 277.800 ;
        RECT 33.880 270.200 34.080 277.800 ;
        RECT 25.930 269.800 34.080 270.200 ;
        RECT 25.930 269.600 26.330 269.800 ;
        RECT 25.930 269.400 29.930 269.600 ;
        RECT 25.930 268.800 26.330 269.400 ;
        RECT 25.930 268.600 29.930 268.800 ;
        RECT 25.930 268.000 26.330 268.600 ;
        RECT 25.930 267.800 29.930 268.000 ;
        RECT 25.930 267.200 26.330 267.800 ;
        RECT 25.930 267.000 29.930 267.200 ;
        RECT 25.930 266.400 26.330 267.000 ;
        RECT 25.930 266.200 29.930 266.400 ;
        RECT 25.930 265.600 26.330 266.200 ;
        RECT 25.930 265.400 29.930 265.600 ;
        RECT 25.930 264.800 26.330 265.400 ;
        RECT 25.930 264.600 29.930 264.800 ;
        RECT 25.930 264.000 26.330 264.600 ;
        RECT 25.930 263.800 29.930 264.000 ;
        RECT 25.930 263.200 26.330 263.800 ;
        RECT 25.930 263.000 29.930 263.200 ;
        RECT 25.930 262.400 26.330 263.000 ;
        RECT 25.930 262.200 29.930 262.400 ;
        RECT 30.680 262.200 30.880 269.800 ;
        RECT 31.480 262.200 31.680 269.800 ;
        RECT 32.280 262.200 32.480 269.800 ;
        RECT 33.080 262.200 33.280 269.800 ;
        RECT 33.880 262.200 34.080 269.800 ;
        RECT 35.380 270.200 35.580 277.800 ;
        RECT 36.180 270.200 36.380 277.800 ;
        RECT 36.980 270.200 37.180 277.800 ;
        RECT 37.780 270.200 37.980 277.800 ;
        RECT 38.580 270.200 38.780 277.800 ;
        RECT 39.530 277.600 43.530 277.800 ;
        RECT 43.130 277.000 43.530 277.600 ;
        RECT 39.530 276.800 43.530 277.000 ;
        RECT 43.130 276.200 43.530 276.800 ;
        RECT 39.530 276.000 43.530 276.200 ;
        RECT 43.130 275.400 43.530 276.000 ;
        RECT 39.530 275.200 43.530 275.400 ;
        RECT 43.130 274.600 43.530 275.200 ;
        RECT 39.530 274.400 43.530 274.600 ;
        RECT 43.130 273.800 43.530 274.400 ;
        RECT 39.530 273.600 43.530 273.800 ;
        RECT 43.130 273.000 43.530 273.600 ;
        RECT 39.530 272.800 43.530 273.000 ;
        RECT 43.130 272.200 43.530 272.800 ;
        RECT 39.530 272.000 43.530 272.200 ;
        RECT 43.130 271.400 43.530 272.000 ;
        RECT 39.530 271.200 43.530 271.400 ;
        RECT 43.130 270.600 43.530 271.200 ;
        RECT 39.530 270.400 43.530 270.600 ;
        RECT 43.130 270.200 43.530 270.400 ;
        RECT 35.380 269.800 43.530 270.200 ;
        RECT 35.380 262.200 35.580 269.800 ;
        RECT 36.180 262.200 36.380 269.800 ;
        RECT 36.980 262.200 37.180 269.800 ;
        RECT 37.780 262.200 37.980 269.800 ;
        RECT 38.580 262.200 38.780 269.800 ;
        RECT 43.130 269.600 43.530 269.800 ;
        RECT 39.530 269.400 43.530 269.600 ;
        RECT 43.130 268.800 43.530 269.400 ;
        RECT 39.530 268.600 43.530 268.800 ;
        RECT 43.130 268.000 43.530 268.600 ;
        RECT 39.530 267.800 43.530 268.000 ;
        RECT 43.130 267.200 43.530 267.800 ;
        RECT 39.530 267.000 43.530 267.200 ;
        RECT 43.130 266.400 43.530 267.000 ;
        RECT 39.530 266.200 43.530 266.400 ;
        RECT 43.130 265.600 43.530 266.200 ;
        RECT 39.530 265.400 43.530 265.600 ;
        RECT 43.130 264.800 43.530 265.400 ;
        RECT 39.530 264.600 43.530 264.800 ;
        RECT 43.130 264.000 43.530 264.600 ;
        RECT 39.530 263.800 43.530 264.000 ;
        RECT 43.130 263.200 43.530 263.800 ;
        RECT 39.530 263.000 43.530 263.200 ;
        RECT 43.130 262.400 43.530 263.000 ;
        RECT 39.530 262.200 43.530 262.400 ;
        RECT 45.930 277.600 49.930 277.800 ;
        RECT 45.930 277.000 46.330 277.600 ;
        RECT 45.930 276.800 49.930 277.000 ;
        RECT 45.930 276.200 46.330 276.800 ;
        RECT 45.930 276.000 49.930 276.200 ;
        RECT 45.930 275.400 46.330 276.000 ;
        RECT 45.930 275.200 49.930 275.400 ;
        RECT 45.930 274.600 46.330 275.200 ;
        RECT 45.930 274.400 49.930 274.600 ;
        RECT 45.930 273.800 46.330 274.400 ;
        RECT 45.930 273.600 49.930 273.800 ;
        RECT 45.930 273.000 46.330 273.600 ;
        RECT 45.930 272.800 49.930 273.000 ;
        RECT 45.930 272.200 46.330 272.800 ;
        RECT 45.930 272.000 49.930 272.200 ;
        RECT 45.930 271.400 46.330 272.000 ;
        RECT 45.930 271.200 49.930 271.400 ;
        RECT 45.930 270.600 46.330 271.200 ;
        RECT 45.930 270.400 49.930 270.600 ;
        RECT 45.930 270.200 46.330 270.400 ;
        RECT 50.680 270.200 50.880 277.800 ;
        RECT 51.480 270.200 51.680 277.800 ;
        RECT 52.280 270.200 52.480 277.800 ;
        RECT 53.080 270.200 53.280 277.800 ;
        RECT 53.880 270.200 54.080 277.800 ;
        RECT 45.930 269.800 54.080 270.200 ;
        RECT 45.930 269.600 46.330 269.800 ;
        RECT 45.930 269.400 49.930 269.600 ;
        RECT 45.930 268.800 46.330 269.400 ;
        RECT 45.930 268.600 49.930 268.800 ;
        RECT 45.930 268.000 46.330 268.600 ;
        RECT 45.930 267.800 49.930 268.000 ;
        RECT 45.930 267.200 46.330 267.800 ;
        RECT 45.930 267.000 49.930 267.200 ;
        RECT 45.930 266.400 46.330 267.000 ;
        RECT 45.930 266.200 49.930 266.400 ;
        RECT 45.930 265.600 46.330 266.200 ;
        RECT 45.930 265.400 49.930 265.600 ;
        RECT 45.930 264.800 46.330 265.400 ;
        RECT 45.930 264.600 49.930 264.800 ;
        RECT 45.930 264.000 46.330 264.600 ;
        RECT 45.930 263.800 49.930 264.000 ;
        RECT 45.930 263.200 46.330 263.800 ;
        RECT 45.930 263.000 49.930 263.200 ;
        RECT 45.930 262.400 46.330 263.000 ;
        RECT 45.930 262.200 49.930 262.400 ;
        RECT 50.680 262.200 50.880 269.800 ;
        RECT 51.480 262.200 51.680 269.800 ;
        RECT 52.280 262.200 52.480 269.800 ;
        RECT 53.080 262.200 53.280 269.800 ;
        RECT 53.880 262.200 54.080 269.800 ;
        RECT 55.380 270.200 55.580 277.800 ;
        RECT 56.180 270.200 56.380 277.800 ;
        RECT 56.980 270.200 57.180 277.800 ;
        RECT 57.780 270.200 57.980 277.800 ;
        RECT 58.580 270.200 58.780 277.800 ;
        RECT 59.530 277.600 63.530 277.800 ;
        RECT 63.130 277.000 63.530 277.600 ;
        RECT 59.530 276.800 63.530 277.000 ;
        RECT 63.130 276.200 63.530 276.800 ;
        RECT 59.530 276.000 63.530 276.200 ;
        RECT 63.130 275.400 63.530 276.000 ;
        RECT 59.530 275.200 63.530 275.400 ;
        RECT 63.130 274.600 63.530 275.200 ;
        RECT 59.530 274.400 63.530 274.600 ;
        RECT 63.130 273.800 63.530 274.400 ;
        RECT 59.530 273.600 63.530 273.800 ;
        RECT 63.130 273.000 63.530 273.600 ;
        RECT 59.530 272.800 63.530 273.000 ;
        RECT 63.130 272.200 63.530 272.800 ;
        RECT 59.530 272.000 63.530 272.200 ;
        RECT 63.130 271.400 63.530 272.000 ;
        RECT 59.530 271.200 63.530 271.400 ;
        RECT 63.130 270.600 63.530 271.200 ;
        RECT 59.530 270.400 63.530 270.600 ;
        RECT 63.130 270.200 63.530 270.400 ;
        RECT 55.380 269.800 63.530 270.200 ;
        RECT 55.380 262.200 55.580 269.800 ;
        RECT 56.180 262.200 56.380 269.800 ;
        RECT 56.980 262.200 57.180 269.800 ;
        RECT 57.780 262.200 57.980 269.800 ;
        RECT 58.580 262.200 58.780 269.800 ;
        RECT 63.130 269.600 63.530 269.800 ;
        RECT 59.530 269.400 63.530 269.600 ;
        RECT 63.130 268.800 63.530 269.400 ;
        RECT 59.530 268.600 63.530 268.800 ;
        RECT 63.130 268.000 63.530 268.600 ;
        RECT 59.530 267.800 63.530 268.000 ;
        RECT 63.130 267.200 63.530 267.800 ;
        RECT 59.530 267.000 63.530 267.200 ;
        RECT 63.130 266.400 63.530 267.000 ;
        RECT 59.530 266.200 63.530 266.400 ;
        RECT 63.130 265.600 63.530 266.200 ;
        RECT 59.530 265.400 63.530 265.600 ;
        RECT 63.130 264.800 63.530 265.400 ;
        RECT 59.530 264.600 63.530 264.800 ;
        RECT 63.130 264.000 63.530 264.600 ;
        RECT 59.530 263.800 63.530 264.000 ;
        RECT 63.130 263.200 63.530 263.800 ;
        RECT 59.530 263.000 63.530 263.200 ;
        RECT 63.130 262.400 63.530 263.000 ;
        RECT 59.530 262.200 63.530 262.400 ;
        RECT 65.930 277.600 69.930 277.800 ;
        RECT 65.930 277.000 66.330 277.600 ;
        RECT 65.930 276.800 69.930 277.000 ;
        RECT 65.930 276.200 66.330 276.800 ;
        RECT 65.930 276.000 69.930 276.200 ;
        RECT 65.930 275.400 66.330 276.000 ;
        RECT 65.930 275.200 69.930 275.400 ;
        RECT 65.930 274.600 66.330 275.200 ;
        RECT 65.930 274.400 69.930 274.600 ;
        RECT 65.930 273.800 66.330 274.400 ;
        RECT 65.930 273.600 69.930 273.800 ;
        RECT 65.930 273.000 66.330 273.600 ;
        RECT 65.930 272.800 69.930 273.000 ;
        RECT 65.930 272.200 66.330 272.800 ;
        RECT 65.930 272.000 69.930 272.200 ;
        RECT 65.930 271.400 66.330 272.000 ;
        RECT 65.930 271.200 69.930 271.400 ;
        RECT 65.930 270.600 66.330 271.200 ;
        RECT 65.930 270.400 69.930 270.600 ;
        RECT 65.930 270.200 66.330 270.400 ;
        RECT 70.680 270.200 70.880 277.800 ;
        RECT 71.480 270.200 71.680 277.800 ;
        RECT 72.280 270.200 72.480 277.800 ;
        RECT 73.080 270.200 73.280 277.800 ;
        RECT 73.880 270.200 74.080 277.800 ;
        RECT 65.930 269.800 74.080 270.200 ;
        RECT 65.930 269.600 66.330 269.800 ;
        RECT 65.930 269.400 69.930 269.600 ;
        RECT 65.930 268.800 66.330 269.400 ;
        RECT 65.930 268.600 69.930 268.800 ;
        RECT 65.930 268.000 66.330 268.600 ;
        RECT 65.930 267.800 69.930 268.000 ;
        RECT 65.930 267.200 66.330 267.800 ;
        RECT 65.930 267.000 69.930 267.200 ;
        RECT 65.930 266.400 66.330 267.000 ;
        RECT 65.930 266.200 69.930 266.400 ;
        RECT 65.930 265.600 66.330 266.200 ;
        RECT 65.930 265.400 69.930 265.600 ;
        RECT 65.930 264.800 66.330 265.400 ;
        RECT 65.930 264.600 69.930 264.800 ;
        RECT 65.930 264.000 66.330 264.600 ;
        RECT 65.930 263.800 69.930 264.000 ;
        RECT 65.930 263.200 66.330 263.800 ;
        RECT 65.930 263.000 69.930 263.200 ;
        RECT 65.930 262.400 66.330 263.000 ;
        RECT 65.930 262.200 69.930 262.400 ;
        RECT 70.680 262.200 70.880 269.800 ;
        RECT 71.480 262.200 71.680 269.800 ;
        RECT 72.280 262.200 72.480 269.800 ;
        RECT 73.080 262.200 73.280 269.800 ;
        RECT 73.880 262.200 74.080 269.800 ;
        RECT 75.380 270.200 75.580 277.800 ;
        RECT 76.180 270.200 76.380 277.800 ;
        RECT 76.980 270.200 77.180 277.800 ;
        RECT 77.780 270.200 77.980 277.800 ;
        RECT 78.580 270.200 78.780 277.800 ;
        RECT 79.530 277.600 83.530 277.800 ;
        RECT 83.130 277.000 83.530 277.600 ;
        RECT 79.530 276.800 83.530 277.000 ;
        RECT 83.130 276.200 83.530 276.800 ;
        RECT 79.530 276.000 83.530 276.200 ;
        RECT 83.130 275.400 83.530 276.000 ;
        RECT 79.530 275.200 83.530 275.400 ;
        RECT 83.130 274.600 83.530 275.200 ;
        RECT 79.530 274.400 83.530 274.600 ;
        RECT 83.130 273.800 83.530 274.400 ;
        RECT 79.530 273.600 83.530 273.800 ;
        RECT 83.130 273.000 83.530 273.600 ;
        RECT 79.530 272.800 83.530 273.000 ;
        RECT 83.130 272.200 83.530 272.800 ;
        RECT 79.530 272.000 83.530 272.200 ;
        RECT 83.130 271.400 83.530 272.000 ;
        RECT 79.530 271.200 83.530 271.400 ;
        RECT 83.130 270.600 83.530 271.200 ;
        RECT 79.530 270.400 83.530 270.600 ;
        RECT 83.130 270.200 83.530 270.400 ;
        RECT 75.380 269.800 83.530 270.200 ;
        RECT 75.380 262.200 75.580 269.800 ;
        RECT 76.180 262.200 76.380 269.800 ;
        RECT 76.980 262.200 77.180 269.800 ;
        RECT 77.780 262.200 77.980 269.800 ;
        RECT 78.580 262.200 78.780 269.800 ;
        RECT 83.130 269.600 83.530 269.800 ;
        RECT 79.530 269.400 83.530 269.600 ;
        RECT 83.130 268.800 83.530 269.400 ;
        RECT 79.530 268.600 83.530 268.800 ;
        RECT 83.130 268.000 83.530 268.600 ;
        RECT 79.530 267.800 83.530 268.000 ;
        RECT 83.130 267.200 83.530 267.800 ;
        RECT 79.530 267.000 83.530 267.200 ;
        RECT 83.130 266.400 83.530 267.000 ;
        RECT 79.530 266.200 83.530 266.400 ;
        RECT 83.130 265.600 83.530 266.200 ;
        RECT 79.530 265.400 83.530 265.600 ;
        RECT 83.130 264.800 83.530 265.400 ;
        RECT 79.530 264.600 83.530 264.800 ;
        RECT 83.130 264.000 83.530 264.600 ;
        RECT 79.530 263.800 83.530 264.000 ;
        RECT 83.130 263.200 83.530 263.800 ;
        RECT 79.530 263.000 83.530 263.200 ;
        RECT 83.130 262.400 83.530 263.000 ;
        RECT 79.530 262.200 83.530 262.400 ;
        RECT 85.930 277.600 89.930 277.800 ;
        RECT 85.930 277.000 86.330 277.600 ;
        RECT 85.930 276.800 89.930 277.000 ;
        RECT 85.930 276.200 86.330 276.800 ;
        RECT 85.930 276.000 89.930 276.200 ;
        RECT 85.930 275.400 86.330 276.000 ;
        RECT 85.930 275.200 89.930 275.400 ;
        RECT 85.930 274.600 86.330 275.200 ;
        RECT 85.930 274.400 89.930 274.600 ;
        RECT 85.930 273.800 86.330 274.400 ;
        RECT 85.930 273.600 89.930 273.800 ;
        RECT 85.930 273.000 86.330 273.600 ;
        RECT 85.930 272.800 89.930 273.000 ;
        RECT 85.930 272.200 86.330 272.800 ;
        RECT 85.930 272.000 89.930 272.200 ;
        RECT 85.930 271.400 86.330 272.000 ;
        RECT 85.930 271.200 89.930 271.400 ;
        RECT 85.930 270.600 86.330 271.200 ;
        RECT 85.930 270.400 89.930 270.600 ;
        RECT 85.930 270.200 86.330 270.400 ;
        RECT 90.680 270.200 90.880 277.800 ;
        RECT 91.480 270.200 91.680 277.800 ;
        RECT 92.280 270.200 92.480 277.800 ;
        RECT 93.080 270.200 93.280 277.800 ;
        RECT 93.880 270.200 94.080 277.800 ;
        RECT 85.930 269.800 94.080 270.200 ;
        RECT 85.930 269.600 86.330 269.800 ;
        RECT 85.930 269.400 89.930 269.600 ;
        RECT 85.930 268.800 86.330 269.400 ;
        RECT 85.930 268.600 89.930 268.800 ;
        RECT 85.930 268.000 86.330 268.600 ;
        RECT 85.930 267.800 89.930 268.000 ;
        RECT 85.930 267.200 86.330 267.800 ;
        RECT 85.930 267.000 89.930 267.200 ;
        RECT 85.930 266.400 86.330 267.000 ;
        RECT 85.930 266.200 89.930 266.400 ;
        RECT 85.930 265.600 86.330 266.200 ;
        RECT 85.930 265.400 89.930 265.600 ;
        RECT 85.930 264.800 86.330 265.400 ;
        RECT 85.930 264.600 89.930 264.800 ;
        RECT 85.930 264.000 86.330 264.600 ;
        RECT 85.930 263.800 89.930 264.000 ;
        RECT 85.930 263.200 86.330 263.800 ;
        RECT 85.930 263.000 89.930 263.200 ;
        RECT 85.930 262.400 86.330 263.000 ;
        RECT 85.930 262.200 89.930 262.400 ;
        RECT 90.680 262.200 90.880 269.800 ;
        RECT 91.480 262.200 91.680 269.800 ;
        RECT 92.280 262.200 92.480 269.800 ;
        RECT 93.080 262.200 93.280 269.800 ;
        RECT 93.880 262.200 94.080 269.800 ;
        RECT 95.380 270.200 95.580 277.800 ;
        RECT 96.180 270.200 96.380 277.800 ;
        RECT 96.980 270.200 97.180 277.800 ;
        RECT 97.780 270.200 97.980 277.800 ;
        RECT 98.580 270.200 98.780 277.800 ;
        RECT 99.530 277.600 103.530 277.800 ;
        RECT 103.130 277.000 103.530 277.600 ;
        RECT 99.530 276.800 103.530 277.000 ;
        RECT 103.130 276.200 103.530 276.800 ;
        RECT 99.530 276.000 103.530 276.200 ;
        RECT 103.130 275.400 103.530 276.000 ;
        RECT 99.530 275.200 103.530 275.400 ;
        RECT 103.130 274.600 103.530 275.200 ;
        RECT 99.530 274.400 103.530 274.600 ;
        RECT 103.130 273.800 103.530 274.400 ;
        RECT 99.530 273.600 103.530 273.800 ;
        RECT 103.130 273.000 103.530 273.600 ;
        RECT 99.530 272.800 103.530 273.000 ;
        RECT 103.130 272.200 103.530 272.800 ;
        RECT 99.530 272.000 103.530 272.200 ;
        RECT 103.130 271.400 103.530 272.000 ;
        RECT 99.530 271.200 103.530 271.400 ;
        RECT 103.130 270.600 103.530 271.200 ;
        RECT 99.530 270.400 103.530 270.600 ;
        RECT 103.130 270.200 103.530 270.400 ;
        RECT 95.380 269.800 103.530 270.200 ;
        RECT 95.380 262.200 95.580 269.800 ;
        RECT 96.180 262.200 96.380 269.800 ;
        RECT 96.980 262.200 97.180 269.800 ;
        RECT 97.780 262.200 97.980 269.800 ;
        RECT 98.580 262.200 98.780 269.800 ;
        RECT 103.130 269.600 103.530 269.800 ;
        RECT 99.530 269.400 103.530 269.600 ;
        RECT 103.130 268.800 103.530 269.400 ;
        RECT 99.530 268.600 103.530 268.800 ;
        RECT 103.130 268.000 103.530 268.600 ;
        RECT 99.530 267.800 103.530 268.000 ;
        RECT 103.130 267.200 103.530 267.800 ;
        RECT 99.530 267.000 103.530 267.200 ;
        RECT 103.130 266.400 103.530 267.000 ;
        RECT 99.530 266.200 103.530 266.400 ;
        RECT 103.130 265.600 103.530 266.200 ;
        RECT 99.530 265.400 103.530 265.600 ;
        RECT 103.130 264.800 103.530 265.400 ;
        RECT 99.530 264.600 103.530 264.800 ;
        RECT 103.130 264.000 103.530 264.600 ;
        RECT 99.530 263.800 103.530 264.000 ;
        RECT 103.130 263.200 103.530 263.800 ;
        RECT 99.530 263.000 103.530 263.200 ;
        RECT 103.130 262.400 103.530 263.000 ;
        RECT 99.530 262.200 103.530 262.400 ;
        RECT 105.930 277.600 109.930 277.800 ;
        RECT 105.930 277.000 106.330 277.600 ;
        RECT 105.930 276.800 109.930 277.000 ;
        RECT 105.930 276.200 106.330 276.800 ;
        RECT 105.930 276.000 109.930 276.200 ;
        RECT 105.930 275.400 106.330 276.000 ;
        RECT 105.930 275.200 109.930 275.400 ;
        RECT 105.930 274.600 106.330 275.200 ;
        RECT 105.930 274.400 109.930 274.600 ;
        RECT 105.930 273.800 106.330 274.400 ;
        RECT 105.930 273.600 109.930 273.800 ;
        RECT 105.930 273.000 106.330 273.600 ;
        RECT 105.930 272.800 109.930 273.000 ;
        RECT 105.930 272.200 106.330 272.800 ;
        RECT 105.930 272.000 109.930 272.200 ;
        RECT 105.930 271.400 106.330 272.000 ;
        RECT 105.930 271.200 109.930 271.400 ;
        RECT 105.930 270.600 106.330 271.200 ;
        RECT 105.930 270.400 109.930 270.600 ;
        RECT 105.930 270.200 106.330 270.400 ;
        RECT 110.680 270.200 110.880 277.800 ;
        RECT 111.480 270.200 111.680 277.800 ;
        RECT 112.280 270.200 112.480 277.800 ;
        RECT 113.080 270.200 113.280 277.800 ;
        RECT 113.880 270.200 114.080 277.800 ;
        RECT 105.930 269.800 114.080 270.200 ;
        RECT 105.930 269.600 106.330 269.800 ;
        RECT 105.930 269.400 109.930 269.600 ;
        RECT 105.930 268.800 106.330 269.400 ;
        RECT 105.930 268.600 109.930 268.800 ;
        RECT 105.930 268.000 106.330 268.600 ;
        RECT 105.930 267.800 109.930 268.000 ;
        RECT 105.930 267.200 106.330 267.800 ;
        RECT 105.930 267.000 109.930 267.200 ;
        RECT 105.930 266.400 106.330 267.000 ;
        RECT 105.930 266.200 109.930 266.400 ;
        RECT 105.930 265.600 106.330 266.200 ;
        RECT 105.930 265.400 109.930 265.600 ;
        RECT 105.930 264.800 106.330 265.400 ;
        RECT 105.930 264.600 109.930 264.800 ;
        RECT 105.930 264.000 106.330 264.600 ;
        RECT 105.930 263.800 109.930 264.000 ;
        RECT 105.930 263.200 106.330 263.800 ;
        RECT 105.930 263.000 109.930 263.200 ;
        RECT 105.930 262.400 106.330 263.000 ;
        RECT 105.930 262.200 109.930 262.400 ;
        RECT 110.680 262.200 110.880 269.800 ;
        RECT 111.480 262.200 111.680 269.800 ;
        RECT 112.280 262.200 112.480 269.800 ;
        RECT 113.080 262.200 113.280 269.800 ;
        RECT 113.880 262.200 114.080 269.800 ;
        RECT 115.380 270.200 115.580 277.800 ;
        RECT 116.180 270.200 116.380 277.800 ;
        RECT 116.980 270.200 117.180 277.800 ;
        RECT 117.780 270.200 117.980 277.800 ;
        RECT 118.580 270.200 118.780 277.800 ;
        RECT 119.530 277.600 123.530 277.800 ;
        RECT 123.130 277.000 123.530 277.600 ;
        RECT 119.530 276.800 123.530 277.000 ;
        RECT 123.130 276.200 123.530 276.800 ;
        RECT 119.530 276.000 123.530 276.200 ;
        RECT 123.130 275.400 123.530 276.000 ;
        RECT 119.530 275.200 123.530 275.400 ;
        RECT 123.130 274.600 123.530 275.200 ;
        RECT 119.530 274.400 123.530 274.600 ;
        RECT 123.130 273.800 123.530 274.400 ;
        RECT 119.530 273.600 123.530 273.800 ;
        RECT 123.130 273.000 123.530 273.600 ;
        RECT 119.530 272.800 123.530 273.000 ;
        RECT 123.130 272.200 123.530 272.800 ;
        RECT 119.530 272.000 123.530 272.200 ;
        RECT 123.130 271.400 123.530 272.000 ;
        RECT 119.530 271.200 123.530 271.400 ;
        RECT 123.130 270.600 123.530 271.200 ;
        RECT 119.530 270.400 123.530 270.600 ;
        RECT 123.130 270.200 123.530 270.400 ;
        RECT 115.380 269.800 123.530 270.200 ;
        RECT 130.050 270.100 130.410 270.480 ;
        RECT 130.680 270.100 131.040 270.480 ;
        RECT 131.280 270.100 131.640 270.480 ;
        RECT 115.380 262.200 115.580 269.800 ;
        RECT 116.180 262.200 116.380 269.800 ;
        RECT 116.980 262.200 117.180 269.800 ;
        RECT 117.780 262.200 117.980 269.800 ;
        RECT 118.580 262.200 118.780 269.800 ;
        RECT 123.130 269.600 123.530 269.800 ;
        RECT 119.530 269.400 123.530 269.600 ;
        RECT 130.050 269.510 130.410 269.890 ;
        RECT 130.680 269.510 131.040 269.890 ;
        RECT 131.280 269.510 131.640 269.890 ;
        RECT 123.130 268.800 123.530 269.400 ;
        RECT 119.530 268.600 123.530 268.800 ;
        RECT 123.130 268.000 123.530 268.600 ;
        RECT 119.530 267.800 123.530 268.000 ;
        RECT 123.130 267.200 123.530 267.800 ;
        RECT 119.530 267.000 123.530 267.200 ;
        RECT 123.130 266.400 123.530 267.000 ;
        RECT 119.530 266.200 123.530 266.400 ;
        RECT 123.130 265.600 123.530 266.200 ;
        RECT 119.530 265.400 123.530 265.600 ;
        RECT 123.130 264.800 123.530 265.400 ;
        RECT 119.530 264.600 123.530 264.800 ;
        RECT 123.130 264.000 123.530 264.600 ;
        RECT 119.530 263.800 123.530 264.000 ;
        RECT 123.130 263.200 123.530 263.800 ;
        RECT 119.530 263.000 123.530 263.200 ;
        RECT 123.130 262.400 123.530 263.000 ;
        RECT 119.530 262.200 123.530 262.400 ;
        RECT 5.930 257.600 9.930 257.800 ;
        RECT 5.930 257.000 6.330 257.600 ;
        RECT 5.930 256.800 9.930 257.000 ;
        RECT 5.930 256.200 6.330 256.800 ;
        RECT 5.930 256.000 9.930 256.200 ;
        RECT 5.930 255.400 6.330 256.000 ;
        RECT 5.930 255.200 9.930 255.400 ;
        RECT 5.930 254.600 6.330 255.200 ;
        RECT 5.930 254.400 9.930 254.600 ;
        RECT 5.930 253.800 6.330 254.400 ;
        RECT 5.930 253.600 9.930 253.800 ;
        RECT 5.930 253.000 6.330 253.600 ;
        RECT 5.930 252.800 9.930 253.000 ;
        RECT 5.930 252.200 6.330 252.800 ;
        RECT 5.930 252.000 9.930 252.200 ;
        RECT 5.930 251.400 6.330 252.000 ;
        RECT 5.930 251.200 9.930 251.400 ;
        RECT 5.930 250.600 6.330 251.200 ;
        RECT 5.930 250.400 9.930 250.600 ;
        RECT 5.930 250.200 6.330 250.400 ;
        RECT 10.680 250.200 10.880 257.800 ;
        RECT 11.480 250.200 11.680 257.800 ;
        RECT 12.280 250.200 12.480 257.800 ;
        RECT 13.080 250.200 13.280 257.800 ;
        RECT 13.880 250.200 14.080 257.800 ;
        RECT 5.930 249.800 14.080 250.200 ;
        RECT 5.930 249.600 6.330 249.800 ;
        RECT 5.930 249.400 9.930 249.600 ;
        RECT 5.930 248.800 6.330 249.400 ;
        RECT 5.930 248.600 9.930 248.800 ;
        RECT 5.930 248.000 6.330 248.600 ;
        RECT 5.930 247.800 9.930 248.000 ;
        RECT 5.930 247.200 6.330 247.800 ;
        RECT 5.930 247.000 9.930 247.200 ;
        RECT 5.930 246.400 6.330 247.000 ;
        RECT 5.930 246.200 9.930 246.400 ;
        RECT 5.930 245.600 6.330 246.200 ;
        RECT 5.930 245.400 9.930 245.600 ;
        RECT 5.930 244.800 6.330 245.400 ;
        RECT 5.930 244.600 9.930 244.800 ;
        RECT 5.930 244.000 6.330 244.600 ;
        RECT 5.930 243.800 9.930 244.000 ;
        RECT 5.930 243.200 6.330 243.800 ;
        RECT 5.930 243.000 9.930 243.200 ;
        RECT 5.930 242.400 6.330 243.000 ;
        RECT 5.930 242.200 9.930 242.400 ;
        RECT 10.680 242.200 10.880 249.800 ;
        RECT 11.480 242.200 11.680 249.800 ;
        RECT 12.280 242.200 12.480 249.800 ;
        RECT 13.080 242.200 13.280 249.800 ;
        RECT 13.880 242.200 14.080 249.800 ;
        RECT 15.380 250.200 15.580 257.800 ;
        RECT 16.180 250.200 16.380 257.800 ;
        RECT 16.980 250.200 17.180 257.800 ;
        RECT 17.780 250.200 17.980 257.800 ;
        RECT 18.580 250.200 18.780 257.800 ;
        RECT 19.530 257.600 23.530 257.800 ;
        RECT 23.130 257.000 23.530 257.600 ;
        RECT 19.530 256.800 23.530 257.000 ;
        RECT 23.130 256.200 23.530 256.800 ;
        RECT 19.530 256.000 23.530 256.200 ;
        RECT 23.130 255.400 23.530 256.000 ;
        RECT 19.530 255.200 23.530 255.400 ;
        RECT 23.130 254.600 23.530 255.200 ;
        RECT 19.530 254.400 23.530 254.600 ;
        RECT 23.130 253.800 23.530 254.400 ;
        RECT 19.530 253.600 23.530 253.800 ;
        RECT 23.130 253.000 23.530 253.600 ;
        RECT 19.530 252.800 23.530 253.000 ;
        RECT 23.130 252.200 23.530 252.800 ;
        RECT 19.530 252.000 23.530 252.200 ;
        RECT 23.130 251.400 23.530 252.000 ;
        RECT 19.530 251.200 23.530 251.400 ;
        RECT 23.130 250.600 23.530 251.200 ;
        RECT 19.530 250.400 23.530 250.600 ;
        RECT 23.130 250.200 23.530 250.400 ;
        RECT 15.380 249.800 23.530 250.200 ;
        RECT 15.380 242.200 15.580 249.800 ;
        RECT 16.180 242.200 16.380 249.800 ;
        RECT 16.980 242.200 17.180 249.800 ;
        RECT 17.780 242.200 17.980 249.800 ;
        RECT 18.580 242.200 18.780 249.800 ;
        RECT 23.130 249.600 23.530 249.800 ;
        RECT 19.530 249.400 23.530 249.600 ;
        RECT 23.130 248.800 23.530 249.400 ;
        RECT 19.530 248.600 23.530 248.800 ;
        RECT 23.130 248.000 23.530 248.600 ;
        RECT 19.530 247.800 23.530 248.000 ;
        RECT 23.130 247.200 23.530 247.800 ;
        RECT 19.530 247.000 23.530 247.200 ;
        RECT 23.130 246.400 23.530 247.000 ;
        RECT 19.530 246.200 23.530 246.400 ;
        RECT 23.130 245.600 23.530 246.200 ;
        RECT 19.530 245.400 23.530 245.600 ;
        RECT 23.130 244.800 23.530 245.400 ;
        RECT 19.530 244.600 23.530 244.800 ;
        RECT 23.130 244.000 23.530 244.600 ;
        RECT 19.530 243.800 23.530 244.000 ;
        RECT 23.130 243.200 23.530 243.800 ;
        RECT 19.530 243.000 23.530 243.200 ;
        RECT 23.130 242.400 23.530 243.000 ;
        RECT 19.530 242.200 23.530 242.400 ;
        RECT 25.930 257.600 29.930 257.800 ;
        RECT 25.930 257.000 26.330 257.600 ;
        RECT 25.930 256.800 29.930 257.000 ;
        RECT 25.930 256.200 26.330 256.800 ;
        RECT 25.930 256.000 29.930 256.200 ;
        RECT 25.930 255.400 26.330 256.000 ;
        RECT 25.930 255.200 29.930 255.400 ;
        RECT 25.930 254.600 26.330 255.200 ;
        RECT 25.930 254.400 29.930 254.600 ;
        RECT 25.930 253.800 26.330 254.400 ;
        RECT 25.930 253.600 29.930 253.800 ;
        RECT 25.930 253.000 26.330 253.600 ;
        RECT 25.930 252.800 29.930 253.000 ;
        RECT 25.930 252.200 26.330 252.800 ;
        RECT 25.930 252.000 29.930 252.200 ;
        RECT 25.930 251.400 26.330 252.000 ;
        RECT 25.930 251.200 29.930 251.400 ;
        RECT 25.930 250.600 26.330 251.200 ;
        RECT 25.930 250.400 29.930 250.600 ;
        RECT 25.930 250.200 26.330 250.400 ;
        RECT 30.680 250.200 30.880 257.800 ;
        RECT 31.480 250.200 31.680 257.800 ;
        RECT 32.280 250.200 32.480 257.800 ;
        RECT 33.080 250.200 33.280 257.800 ;
        RECT 33.880 250.200 34.080 257.800 ;
        RECT 25.930 249.800 34.080 250.200 ;
        RECT 25.930 249.600 26.330 249.800 ;
        RECT 25.930 249.400 29.930 249.600 ;
        RECT 25.930 248.800 26.330 249.400 ;
        RECT 25.930 248.600 29.930 248.800 ;
        RECT 25.930 248.000 26.330 248.600 ;
        RECT 25.930 247.800 29.930 248.000 ;
        RECT 25.930 247.200 26.330 247.800 ;
        RECT 25.930 247.000 29.930 247.200 ;
        RECT 25.930 246.400 26.330 247.000 ;
        RECT 25.930 246.200 29.930 246.400 ;
        RECT 25.930 245.600 26.330 246.200 ;
        RECT 25.930 245.400 29.930 245.600 ;
        RECT 25.930 244.800 26.330 245.400 ;
        RECT 25.930 244.600 29.930 244.800 ;
        RECT 25.930 244.000 26.330 244.600 ;
        RECT 25.930 243.800 29.930 244.000 ;
        RECT 25.930 243.200 26.330 243.800 ;
        RECT 25.930 243.000 29.930 243.200 ;
        RECT 25.930 242.400 26.330 243.000 ;
        RECT 25.930 242.200 29.930 242.400 ;
        RECT 30.680 242.200 30.880 249.800 ;
        RECT 31.480 242.200 31.680 249.800 ;
        RECT 32.280 242.200 32.480 249.800 ;
        RECT 33.080 242.200 33.280 249.800 ;
        RECT 33.880 242.200 34.080 249.800 ;
        RECT 35.380 250.200 35.580 257.800 ;
        RECT 36.180 250.200 36.380 257.800 ;
        RECT 36.980 250.200 37.180 257.800 ;
        RECT 37.780 250.200 37.980 257.800 ;
        RECT 38.580 250.200 38.780 257.800 ;
        RECT 39.530 257.600 43.530 257.800 ;
        RECT 43.130 257.000 43.530 257.600 ;
        RECT 39.530 256.800 43.530 257.000 ;
        RECT 43.130 256.200 43.530 256.800 ;
        RECT 39.530 256.000 43.530 256.200 ;
        RECT 43.130 255.400 43.530 256.000 ;
        RECT 39.530 255.200 43.530 255.400 ;
        RECT 43.130 254.600 43.530 255.200 ;
        RECT 39.530 254.400 43.530 254.600 ;
        RECT 43.130 253.800 43.530 254.400 ;
        RECT 39.530 253.600 43.530 253.800 ;
        RECT 43.130 253.000 43.530 253.600 ;
        RECT 39.530 252.800 43.530 253.000 ;
        RECT 43.130 252.200 43.530 252.800 ;
        RECT 39.530 252.000 43.530 252.200 ;
        RECT 43.130 251.400 43.530 252.000 ;
        RECT 39.530 251.200 43.530 251.400 ;
        RECT 43.130 250.600 43.530 251.200 ;
        RECT 39.530 250.400 43.530 250.600 ;
        RECT 43.130 250.200 43.530 250.400 ;
        RECT 35.380 249.800 43.530 250.200 ;
        RECT 35.380 242.200 35.580 249.800 ;
        RECT 36.180 242.200 36.380 249.800 ;
        RECT 36.980 242.200 37.180 249.800 ;
        RECT 37.780 242.200 37.980 249.800 ;
        RECT 38.580 242.200 38.780 249.800 ;
        RECT 43.130 249.600 43.530 249.800 ;
        RECT 39.530 249.400 43.530 249.600 ;
        RECT 43.130 248.800 43.530 249.400 ;
        RECT 39.530 248.600 43.530 248.800 ;
        RECT 43.130 248.000 43.530 248.600 ;
        RECT 39.530 247.800 43.530 248.000 ;
        RECT 43.130 247.200 43.530 247.800 ;
        RECT 39.530 247.000 43.530 247.200 ;
        RECT 43.130 246.400 43.530 247.000 ;
        RECT 39.530 246.200 43.530 246.400 ;
        RECT 43.130 245.600 43.530 246.200 ;
        RECT 39.530 245.400 43.530 245.600 ;
        RECT 43.130 244.800 43.530 245.400 ;
        RECT 39.530 244.600 43.530 244.800 ;
        RECT 43.130 244.000 43.530 244.600 ;
        RECT 39.530 243.800 43.530 244.000 ;
        RECT 43.130 243.200 43.530 243.800 ;
        RECT 39.530 243.000 43.530 243.200 ;
        RECT 43.130 242.400 43.530 243.000 ;
        RECT 39.530 242.200 43.530 242.400 ;
        RECT 45.930 257.600 49.930 257.800 ;
        RECT 45.930 257.000 46.330 257.600 ;
        RECT 45.930 256.800 49.930 257.000 ;
        RECT 45.930 256.200 46.330 256.800 ;
        RECT 45.930 256.000 49.930 256.200 ;
        RECT 45.930 255.400 46.330 256.000 ;
        RECT 45.930 255.200 49.930 255.400 ;
        RECT 45.930 254.600 46.330 255.200 ;
        RECT 45.930 254.400 49.930 254.600 ;
        RECT 45.930 253.800 46.330 254.400 ;
        RECT 45.930 253.600 49.930 253.800 ;
        RECT 45.930 253.000 46.330 253.600 ;
        RECT 45.930 252.800 49.930 253.000 ;
        RECT 45.930 252.200 46.330 252.800 ;
        RECT 45.930 252.000 49.930 252.200 ;
        RECT 45.930 251.400 46.330 252.000 ;
        RECT 45.930 251.200 49.930 251.400 ;
        RECT 45.930 250.600 46.330 251.200 ;
        RECT 45.930 250.400 49.930 250.600 ;
        RECT 45.930 250.200 46.330 250.400 ;
        RECT 50.680 250.200 50.880 257.800 ;
        RECT 51.480 250.200 51.680 257.800 ;
        RECT 52.280 250.200 52.480 257.800 ;
        RECT 53.080 250.200 53.280 257.800 ;
        RECT 53.880 250.200 54.080 257.800 ;
        RECT 45.930 249.800 54.080 250.200 ;
        RECT 45.930 249.600 46.330 249.800 ;
        RECT 45.930 249.400 49.930 249.600 ;
        RECT 45.930 248.800 46.330 249.400 ;
        RECT 45.930 248.600 49.930 248.800 ;
        RECT 45.930 248.000 46.330 248.600 ;
        RECT 45.930 247.800 49.930 248.000 ;
        RECT 45.930 247.200 46.330 247.800 ;
        RECT 45.930 247.000 49.930 247.200 ;
        RECT 45.930 246.400 46.330 247.000 ;
        RECT 45.930 246.200 49.930 246.400 ;
        RECT 45.930 245.600 46.330 246.200 ;
        RECT 45.930 245.400 49.930 245.600 ;
        RECT 45.930 244.800 46.330 245.400 ;
        RECT 45.930 244.600 49.930 244.800 ;
        RECT 45.930 244.000 46.330 244.600 ;
        RECT 45.930 243.800 49.930 244.000 ;
        RECT 45.930 243.200 46.330 243.800 ;
        RECT 45.930 243.000 49.930 243.200 ;
        RECT 45.930 242.400 46.330 243.000 ;
        RECT 45.930 242.200 49.930 242.400 ;
        RECT 50.680 242.200 50.880 249.800 ;
        RECT 51.480 242.200 51.680 249.800 ;
        RECT 52.280 242.200 52.480 249.800 ;
        RECT 53.080 242.200 53.280 249.800 ;
        RECT 53.880 242.200 54.080 249.800 ;
        RECT 55.380 250.200 55.580 257.800 ;
        RECT 56.180 250.200 56.380 257.800 ;
        RECT 56.980 250.200 57.180 257.800 ;
        RECT 57.780 250.200 57.980 257.800 ;
        RECT 58.580 250.200 58.780 257.800 ;
        RECT 59.530 257.600 63.530 257.800 ;
        RECT 63.130 257.000 63.530 257.600 ;
        RECT 59.530 256.800 63.530 257.000 ;
        RECT 63.130 256.200 63.530 256.800 ;
        RECT 59.530 256.000 63.530 256.200 ;
        RECT 63.130 255.400 63.530 256.000 ;
        RECT 59.530 255.200 63.530 255.400 ;
        RECT 63.130 254.600 63.530 255.200 ;
        RECT 59.530 254.400 63.530 254.600 ;
        RECT 63.130 253.800 63.530 254.400 ;
        RECT 59.530 253.600 63.530 253.800 ;
        RECT 63.130 253.000 63.530 253.600 ;
        RECT 59.530 252.800 63.530 253.000 ;
        RECT 63.130 252.200 63.530 252.800 ;
        RECT 59.530 252.000 63.530 252.200 ;
        RECT 63.130 251.400 63.530 252.000 ;
        RECT 59.530 251.200 63.530 251.400 ;
        RECT 63.130 250.600 63.530 251.200 ;
        RECT 59.530 250.400 63.530 250.600 ;
        RECT 63.130 250.200 63.530 250.400 ;
        RECT 55.380 249.800 63.530 250.200 ;
        RECT 55.380 242.200 55.580 249.800 ;
        RECT 56.180 242.200 56.380 249.800 ;
        RECT 56.980 242.200 57.180 249.800 ;
        RECT 57.780 242.200 57.980 249.800 ;
        RECT 58.580 242.200 58.780 249.800 ;
        RECT 63.130 249.600 63.530 249.800 ;
        RECT 59.530 249.400 63.530 249.600 ;
        RECT 63.130 248.800 63.530 249.400 ;
        RECT 59.530 248.600 63.530 248.800 ;
        RECT 63.130 248.000 63.530 248.600 ;
        RECT 59.530 247.800 63.530 248.000 ;
        RECT 63.130 247.200 63.530 247.800 ;
        RECT 59.530 247.000 63.530 247.200 ;
        RECT 63.130 246.400 63.530 247.000 ;
        RECT 59.530 246.200 63.530 246.400 ;
        RECT 63.130 245.600 63.530 246.200 ;
        RECT 59.530 245.400 63.530 245.600 ;
        RECT 63.130 244.800 63.530 245.400 ;
        RECT 59.530 244.600 63.530 244.800 ;
        RECT 63.130 244.000 63.530 244.600 ;
        RECT 59.530 243.800 63.530 244.000 ;
        RECT 63.130 243.200 63.530 243.800 ;
        RECT 59.530 243.000 63.530 243.200 ;
        RECT 63.130 242.400 63.530 243.000 ;
        RECT 59.530 242.200 63.530 242.400 ;
        RECT 65.930 257.600 69.930 257.800 ;
        RECT 65.930 257.000 66.330 257.600 ;
        RECT 65.930 256.800 69.930 257.000 ;
        RECT 65.930 256.200 66.330 256.800 ;
        RECT 65.930 256.000 69.930 256.200 ;
        RECT 65.930 255.400 66.330 256.000 ;
        RECT 65.930 255.200 69.930 255.400 ;
        RECT 65.930 254.600 66.330 255.200 ;
        RECT 65.930 254.400 69.930 254.600 ;
        RECT 65.930 253.800 66.330 254.400 ;
        RECT 65.930 253.600 69.930 253.800 ;
        RECT 65.930 253.000 66.330 253.600 ;
        RECT 65.930 252.800 69.930 253.000 ;
        RECT 65.930 252.200 66.330 252.800 ;
        RECT 65.930 252.000 69.930 252.200 ;
        RECT 65.930 251.400 66.330 252.000 ;
        RECT 65.930 251.200 69.930 251.400 ;
        RECT 65.930 250.600 66.330 251.200 ;
        RECT 65.930 250.400 69.930 250.600 ;
        RECT 65.930 250.200 66.330 250.400 ;
        RECT 70.680 250.200 70.880 257.800 ;
        RECT 71.480 250.200 71.680 257.800 ;
        RECT 72.280 250.200 72.480 257.800 ;
        RECT 73.080 250.200 73.280 257.800 ;
        RECT 73.880 250.200 74.080 257.800 ;
        RECT 65.930 249.800 74.080 250.200 ;
        RECT 65.930 249.600 66.330 249.800 ;
        RECT 65.930 249.400 69.930 249.600 ;
        RECT 65.930 248.800 66.330 249.400 ;
        RECT 65.930 248.600 69.930 248.800 ;
        RECT 65.930 248.000 66.330 248.600 ;
        RECT 65.930 247.800 69.930 248.000 ;
        RECT 65.930 247.200 66.330 247.800 ;
        RECT 65.930 247.000 69.930 247.200 ;
        RECT 65.930 246.400 66.330 247.000 ;
        RECT 65.930 246.200 69.930 246.400 ;
        RECT 65.930 245.600 66.330 246.200 ;
        RECT 65.930 245.400 69.930 245.600 ;
        RECT 65.930 244.800 66.330 245.400 ;
        RECT 65.930 244.600 69.930 244.800 ;
        RECT 65.930 244.000 66.330 244.600 ;
        RECT 65.930 243.800 69.930 244.000 ;
        RECT 65.930 243.200 66.330 243.800 ;
        RECT 65.930 243.000 69.930 243.200 ;
        RECT 65.930 242.400 66.330 243.000 ;
        RECT 65.930 242.200 69.930 242.400 ;
        RECT 70.680 242.200 70.880 249.800 ;
        RECT 71.480 242.200 71.680 249.800 ;
        RECT 72.280 242.200 72.480 249.800 ;
        RECT 73.080 242.200 73.280 249.800 ;
        RECT 73.880 242.200 74.080 249.800 ;
        RECT 75.380 250.200 75.580 257.800 ;
        RECT 76.180 250.200 76.380 257.800 ;
        RECT 76.980 250.200 77.180 257.800 ;
        RECT 77.780 250.200 77.980 257.800 ;
        RECT 78.580 250.200 78.780 257.800 ;
        RECT 79.530 257.600 83.530 257.800 ;
        RECT 83.130 257.000 83.530 257.600 ;
        RECT 79.530 256.800 83.530 257.000 ;
        RECT 83.130 256.200 83.530 256.800 ;
        RECT 79.530 256.000 83.530 256.200 ;
        RECT 83.130 255.400 83.530 256.000 ;
        RECT 79.530 255.200 83.530 255.400 ;
        RECT 83.130 254.600 83.530 255.200 ;
        RECT 79.530 254.400 83.530 254.600 ;
        RECT 83.130 253.800 83.530 254.400 ;
        RECT 79.530 253.600 83.530 253.800 ;
        RECT 83.130 253.000 83.530 253.600 ;
        RECT 79.530 252.800 83.530 253.000 ;
        RECT 83.130 252.200 83.530 252.800 ;
        RECT 79.530 252.000 83.530 252.200 ;
        RECT 83.130 251.400 83.530 252.000 ;
        RECT 79.530 251.200 83.530 251.400 ;
        RECT 83.130 250.600 83.530 251.200 ;
        RECT 79.530 250.400 83.530 250.600 ;
        RECT 83.130 250.200 83.530 250.400 ;
        RECT 75.380 249.800 83.530 250.200 ;
        RECT 75.380 242.200 75.580 249.800 ;
        RECT 76.180 242.200 76.380 249.800 ;
        RECT 76.980 242.200 77.180 249.800 ;
        RECT 77.780 242.200 77.980 249.800 ;
        RECT 78.580 242.200 78.780 249.800 ;
        RECT 83.130 249.600 83.530 249.800 ;
        RECT 79.530 249.400 83.530 249.600 ;
        RECT 83.130 248.800 83.530 249.400 ;
        RECT 79.530 248.600 83.530 248.800 ;
        RECT 83.130 248.000 83.530 248.600 ;
        RECT 79.530 247.800 83.530 248.000 ;
        RECT 83.130 247.200 83.530 247.800 ;
        RECT 79.530 247.000 83.530 247.200 ;
        RECT 83.130 246.400 83.530 247.000 ;
        RECT 79.530 246.200 83.530 246.400 ;
        RECT 83.130 245.600 83.530 246.200 ;
        RECT 79.530 245.400 83.530 245.600 ;
        RECT 83.130 244.800 83.530 245.400 ;
        RECT 79.530 244.600 83.530 244.800 ;
        RECT 83.130 244.000 83.530 244.600 ;
        RECT 79.530 243.800 83.530 244.000 ;
        RECT 83.130 243.200 83.530 243.800 ;
        RECT 79.530 243.000 83.530 243.200 ;
        RECT 83.130 242.400 83.530 243.000 ;
        RECT 79.530 242.200 83.530 242.400 ;
        RECT 85.930 257.600 89.930 257.800 ;
        RECT 85.930 257.000 86.330 257.600 ;
        RECT 85.930 256.800 89.930 257.000 ;
        RECT 85.930 256.200 86.330 256.800 ;
        RECT 85.930 256.000 89.930 256.200 ;
        RECT 85.930 255.400 86.330 256.000 ;
        RECT 85.930 255.200 89.930 255.400 ;
        RECT 85.930 254.600 86.330 255.200 ;
        RECT 85.930 254.400 89.930 254.600 ;
        RECT 85.930 253.800 86.330 254.400 ;
        RECT 85.930 253.600 89.930 253.800 ;
        RECT 85.930 253.000 86.330 253.600 ;
        RECT 85.930 252.800 89.930 253.000 ;
        RECT 85.930 252.200 86.330 252.800 ;
        RECT 85.930 252.000 89.930 252.200 ;
        RECT 85.930 251.400 86.330 252.000 ;
        RECT 85.930 251.200 89.930 251.400 ;
        RECT 85.930 250.600 86.330 251.200 ;
        RECT 85.930 250.400 89.930 250.600 ;
        RECT 85.930 250.200 86.330 250.400 ;
        RECT 90.680 250.200 90.880 257.800 ;
        RECT 91.480 250.200 91.680 257.800 ;
        RECT 92.280 250.200 92.480 257.800 ;
        RECT 93.080 250.200 93.280 257.800 ;
        RECT 93.880 250.200 94.080 257.800 ;
        RECT 85.930 249.800 94.080 250.200 ;
        RECT 85.930 249.600 86.330 249.800 ;
        RECT 85.930 249.400 89.930 249.600 ;
        RECT 85.930 248.800 86.330 249.400 ;
        RECT 85.930 248.600 89.930 248.800 ;
        RECT 85.930 248.000 86.330 248.600 ;
        RECT 85.930 247.800 89.930 248.000 ;
        RECT 85.930 247.200 86.330 247.800 ;
        RECT 85.930 247.000 89.930 247.200 ;
        RECT 85.930 246.400 86.330 247.000 ;
        RECT 85.930 246.200 89.930 246.400 ;
        RECT 85.930 245.600 86.330 246.200 ;
        RECT 85.930 245.400 89.930 245.600 ;
        RECT 85.930 244.800 86.330 245.400 ;
        RECT 85.930 244.600 89.930 244.800 ;
        RECT 85.930 244.000 86.330 244.600 ;
        RECT 85.930 243.800 89.930 244.000 ;
        RECT 85.930 243.200 86.330 243.800 ;
        RECT 85.930 243.000 89.930 243.200 ;
        RECT 85.930 242.400 86.330 243.000 ;
        RECT 85.930 242.200 89.930 242.400 ;
        RECT 90.680 242.200 90.880 249.800 ;
        RECT 91.480 242.200 91.680 249.800 ;
        RECT 92.280 242.200 92.480 249.800 ;
        RECT 93.080 242.200 93.280 249.800 ;
        RECT 93.880 242.200 94.080 249.800 ;
        RECT 95.380 250.200 95.580 257.800 ;
        RECT 96.180 250.200 96.380 257.800 ;
        RECT 96.980 250.200 97.180 257.800 ;
        RECT 97.780 250.200 97.980 257.800 ;
        RECT 98.580 250.200 98.780 257.800 ;
        RECT 99.530 257.600 103.530 257.800 ;
        RECT 103.130 257.000 103.530 257.600 ;
        RECT 99.530 256.800 103.530 257.000 ;
        RECT 103.130 256.200 103.530 256.800 ;
        RECT 99.530 256.000 103.530 256.200 ;
        RECT 103.130 255.400 103.530 256.000 ;
        RECT 99.530 255.200 103.530 255.400 ;
        RECT 103.130 254.600 103.530 255.200 ;
        RECT 99.530 254.400 103.530 254.600 ;
        RECT 103.130 253.800 103.530 254.400 ;
        RECT 99.530 253.600 103.530 253.800 ;
        RECT 103.130 253.000 103.530 253.600 ;
        RECT 99.530 252.800 103.530 253.000 ;
        RECT 103.130 252.200 103.530 252.800 ;
        RECT 99.530 252.000 103.530 252.200 ;
        RECT 103.130 251.400 103.530 252.000 ;
        RECT 99.530 251.200 103.530 251.400 ;
        RECT 103.130 250.600 103.530 251.200 ;
        RECT 99.530 250.400 103.530 250.600 ;
        RECT 103.130 250.200 103.530 250.400 ;
        RECT 95.380 249.800 103.530 250.200 ;
        RECT 95.380 242.200 95.580 249.800 ;
        RECT 96.180 242.200 96.380 249.800 ;
        RECT 96.980 242.200 97.180 249.800 ;
        RECT 97.780 242.200 97.980 249.800 ;
        RECT 98.580 242.200 98.780 249.800 ;
        RECT 103.130 249.600 103.530 249.800 ;
        RECT 99.530 249.400 103.530 249.600 ;
        RECT 103.130 248.800 103.530 249.400 ;
        RECT 99.530 248.600 103.530 248.800 ;
        RECT 103.130 248.000 103.530 248.600 ;
        RECT 99.530 247.800 103.530 248.000 ;
        RECT 103.130 247.200 103.530 247.800 ;
        RECT 99.530 247.000 103.530 247.200 ;
        RECT 103.130 246.400 103.530 247.000 ;
        RECT 99.530 246.200 103.530 246.400 ;
        RECT 103.130 245.600 103.530 246.200 ;
        RECT 99.530 245.400 103.530 245.600 ;
        RECT 103.130 244.800 103.530 245.400 ;
        RECT 99.530 244.600 103.530 244.800 ;
        RECT 103.130 244.000 103.530 244.600 ;
        RECT 99.530 243.800 103.530 244.000 ;
        RECT 103.130 243.200 103.530 243.800 ;
        RECT 99.530 243.000 103.530 243.200 ;
        RECT 103.130 242.400 103.530 243.000 ;
        RECT 99.530 242.200 103.530 242.400 ;
        RECT 105.930 257.600 109.930 257.800 ;
        RECT 105.930 257.000 106.330 257.600 ;
        RECT 105.930 256.800 109.930 257.000 ;
        RECT 105.930 256.200 106.330 256.800 ;
        RECT 105.930 256.000 109.930 256.200 ;
        RECT 105.930 255.400 106.330 256.000 ;
        RECT 105.930 255.200 109.930 255.400 ;
        RECT 105.930 254.600 106.330 255.200 ;
        RECT 105.930 254.400 109.930 254.600 ;
        RECT 105.930 253.800 106.330 254.400 ;
        RECT 105.930 253.600 109.930 253.800 ;
        RECT 105.930 253.000 106.330 253.600 ;
        RECT 105.930 252.800 109.930 253.000 ;
        RECT 105.930 252.200 106.330 252.800 ;
        RECT 105.930 252.000 109.930 252.200 ;
        RECT 105.930 251.400 106.330 252.000 ;
        RECT 105.930 251.200 109.930 251.400 ;
        RECT 105.930 250.600 106.330 251.200 ;
        RECT 105.930 250.400 109.930 250.600 ;
        RECT 105.930 250.200 106.330 250.400 ;
        RECT 110.680 250.200 110.880 257.800 ;
        RECT 111.480 250.200 111.680 257.800 ;
        RECT 112.280 250.200 112.480 257.800 ;
        RECT 113.080 250.200 113.280 257.800 ;
        RECT 113.880 250.200 114.080 257.800 ;
        RECT 105.930 249.800 114.080 250.200 ;
        RECT 105.930 249.600 106.330 249.800 ;
        RECT 105.930 249.400 109.930 249.600 ;
        RECT 105.930 248.800 106.330 249.400 ;
        RECT 105.930 248.600 109.930 248.800 ;
        RECT 105.930 248.000 106.330 248.600 ;
        RECT 105.930 247.800 109.930 248.000 ;
        RECT 105.930 247.200 106.330 247.800 ;
        RECT 105.930 247.000 109.930 247.200 ;
        RECT 105.930 246.400 106.330 247.000 ;
        RECT 105.930 246.200 109.930 246.400 ;
        RECT 105.930 245.600 106.330 246.200 ;
        RECT 105.930 245.400 109.930 245.600 ;
        RECT 105.930 244.800 106.330 245.400 ;
        RECT 105.930 244.600 109.930 244.800 ;
        RECT 105.930 244.000 106.330 244.600 ;
        RECT 105.930 243.800 109.930 244.000 ;
        RECT 105.930 243.200 106.330 243.800 ;
        RECT 105.930 243.000 109.930 243.200 ;
        RECT 105.930 242.400 106.330 243.000 ;
        RECT 105.930 242.200 109.930 242.400 ;
        RECT 110.680 242.200 110.880 249.800 ;
        RECT 111.480 242.200 111.680 249.800 ;
        RECT 112.280 242.200 112.480 249.800 ;
        RECT 113.080 242.200 113.280 249.800 ;
        RECT 113.880 242.200 114.080 249.800 ;
        RECT 115.380 250.200 115.580 257.800 ;
        RECT 116.180 250.200 116.380 257.800 ;
        RECT 116.980 250.200 117.180 257.800 ;
        RECT 117.780 250.200 117.980 257.800 ;
        RECT 118.580 250.200 118.780 257.800 ;
        RECT 119.530 257.600 123.530 257.800 ;
        RECT 123.130 257.000 123.530 257.600 ;
        RECT 119.530 256.800 123.530 257.000 ;
        RECT 123.130 256.200 123.530 256.800 ;
        RECT 119.530 256.000 123.530 256.200 ;
        RECT 123.130 255.400 123.530 256.000 ;
        RECT 119.530 255.200 123.530 255.400 ;
        RECT 123.130 254.600 123.530 255.200 ;
        RECT 119.530 254.400 123.530 254.600 ;
        RECT 123.130 253.800 123.530 254.400 ;
        RECT 119.530 253.600 123.530 253.800 ;
        RECT 123.130 253.000 123.530 253.600 ;
        RECT 119.530 252.800 123.530 253.000 ;
        RECT 123.130 252.200 123.530 252.800 ;
        RECT 119.530 252.000 123.530 252.200 ;
        RECT 123.130 251.400 123.530 252.000 ;
        RECT 119.530 251.200 123.530 251.400 ;
        RECT 123.130 250.600 123.530 251.200 ;
        RECT 119.530 250.400 123.530 250.600 ;
        RECT 123.130 250.200 123.530 250.400 ;
        RECT 115.380 249.800 123.530 250.200 ;
        RECT 130.050 250.015 130.410 250.395 ;
        RECT 130.680 250.015 131.040 250.395 ;
        RECT 131.280 250.015 131.640 250.395 ;
        RECT 115.380 242.200 115.580 249.800 ;
        RECT 116.180 242.200 116.380 249.800 ;
        RECT 116.980 242.200 117.180 249.800 ;
        RECT 117.780 242.200 117.980 249.800 ;
        RECT 118.580 242.200 118.780 249.800 ;
        RECT 123.130 249.600 123.530 249.800 ;
        RECT 119.530 249.400 123.530 249.600 ;
        RECT 130.050 249.425 130.410 249.805 ;
        RECT 130.680 249.425 131.040 249.805 ;
        RECT 131.280 249.425 131.640 249.805 ;
        RECT 123.130 248.800 123.530 249.400 ;
        RECT 119.530 248.600 123.530 248.800 ;
        RECT 123.130 248.000 123.530 248.600 ;
        RECT 119.530 247.800 123.530 248.000 ;
        RECT 123.130 247.200 123.530 247.800 ;
        RECT 119.530 247.000 123.530 247.200 ;
        RECT 123.130 246.400 123.530 247.000 ;
        RECT 119.530 246.200 123.530 246.400 ;
        RECT 123.130 245.600 123.530 246.200 ;
        RECT 119.530 245.400 123.530 245.600 ;
        RECT 123.130 244.800 123.530 245.400 ;
        RECT 119.530 244.600 123.530 244.800 ;
        RECT 123.130 244.000 123.530 244.600 ;
        RECT 119.530 243.800 123.530 244.000 ;
        RECT 123.130 243.200 123.530 243.800 ;
        RECT 119.530 243.000 123.530 243.200 ;
        RECT 123.130 242.400 123.530 243.000 ;
        RECT 119.530 242.200 123.530 242.400 ;
        RECT 5.930 237.600 9.930 237.800 ;
        RECT 5.930 237.000 6.330 237.600 ;
        RECT 5.930 236.800 9.930 237.000 ;
        RECT 5.930 236.200 6.330 236.800 ;
        RECT 5.930 236.000 9.930 236.200 ;
        RECT 5.930 235.400 6.330 236.000 ;
        RECT 5.930 235.200 9.930 235.400 ;
        RECT 5.930 234.600 6.330 235.200 ;
        RECT 5.930 234.400 9.930 234.600 ;
        RECT 5.930 233.800 6.330 234.400 ;
        RECT 5.930 233.600 9.930 233.800 ;
        RECT 5.930 233.000 6.330 233.600 ;
        RECT 5.930 232.800 9.930 233.000 ;
        RECT 5.930 232.200 6.330 232.800 ;
        RECT 5.930 232.000 9.930 232.200 ;
        RECT 5.930 231.400 6.330 232.000 ;
        RECT 5.930 231.200 9.930 231.400 ;
        RECT 5.930 230.600 6.330 231.200 ;
        RECT 5.930 230.400 9.930 230.600 ;
        RECT 5.930 230.200 6.330 230.400 ;
        RECT 10.680 230.200 10.880 237.800 ;
        RECT 11.480 230.200 11.680 237.800 ;
        RECT 12.280 230.200 12.480 237.800 ;
        RECT 13.080 230.200 13.280 237.800 ;
        RECT 13.880 230.200 14.080 237.800 ;
        RECT 5.930 229.800 14.080 230.200 ;
        RECT 5.930 229.600 6.330 229.800 ;
        RECT 5.930 229.400 9.930 229.600 ;
        RECT 5.930 228.800 6.330 229.400 ;
        RECT 5.930 228.600 9.930 228.800 ;
        RECT 5.930 228.000 6.330 228.600 ;
        RECT 5.930 227.800 9.930 228.000 ;
        RECT 5.930 227.200 6.330 227.800 ;
        RECT 5.930 227.000 9.930 227.200 ;
        RECT 5.930 226.400 6.330 227.000 ;
        RECT 5.930 226.200 9.930 226.400 ;
        RECT 5.930 225.600 6.330 226.200 ;
        RECT 5.930 225.400 9.930 225.600 ;
        RECT 5.930 224.800 6.330 225.400 ;
        RECT 5.930 224.600 9.930 224.800 ;
        RECT 5.930 224.000 6.330 224.600 ;
        RECT 5.930 223.800 9.930 224.000 ;
        RECT 5.930 223.200 6.330 223.800 ;
        RECT 5.930 223.000 9.930 223.200 ;
        RECT 5.930 222.400 6.330 223.000 ;
        RECT 5.930 222.200 9.930 222.400 ;
        RECT 10.680 222.200 10.880 229.800 ;
        RECT 11.480 222.200 11.680 229.800 ;
        RECT 12.280 222.200 12.480 229.800 ;
        RECT 13.080 222.200 13.280 229.800 ;
        RECT 13.880 222.200 14.080 229.800 ;
        RECT 15.380 230.200 15.580 237.800 ;
        RECT 16.180 230.200 16.380 237.800 ;
        RECT 16.980 230.200 17.180 237.800 ;
        RECT 17.780 230.200 17.980 237.800 ;
        RECT 18.580 230.200 18.780 237.800 ;
        RECT 19.530 237.600 23.530 237.800 ;
        RECT 23.130 237.000 23.530 237.600 ;
        RECT 19.530 236.800 23.530 237.000 ;
        RECT 23.130 236.200 23.530 236.800 ;
        RECT 19.530 236.000 23.530 236.200 ;
        RECT 23.130 235.400 23.530 236.000 ;
        RECT 19.530 235.200 23.530 235.400 ;
        RECT 23.130 234.600 23.530 235.200 ;
        RECT 19.530 234.400 23.530 234.600 ;
        RECT 23.130 233.800 23.530 234.400 ;
        RECT 19.530 233.600 23.530 233.800 ;
        RECT 23.130 233.000 23.530 233.600 ;
        RECT 19.530 232.800 23.530 233.000 ;
        RECT 23.130 232.200 23.530 232.800 ;
        RECT 19.530 232.000 23.530 232.200 ;
        RECT 23.130 231.400 23.530 232.000 ;
        RECT 19.530 231.200 23.530 231.400 ;
        RECT 23.130 230.600 23.530 231.200 ;
        RECT 19.530 230.400 23.530 230.600 ;
        RECT 23.130 230.200 23.530 230.400 ;
        RECT 15.380 229.800 23.530 230.200 ;
        RECT 15.380 222.200 15.580 229.800 ;
        RECT 16.180 222.200 16.380 229.800 ;
        RECT 16.980 222.200 17.180 229.800 ;
        RECT 17.780 222.200 17.980 229.800 ;
        RECT 18.580 222.200 18.780 229.800 ;
        RECT 23.130 229.600 23.530 229.800 ;
        RECT 19.530 229.400 23.530 229.600 ;
        RECT 23.130 228.800 23.530 229.400 ;
        RECT 19.530 228.600 23.530 228.800 ;
        RECT 23.130 228.000 23.530 228.600 ;
        RECT 19.530 227.800 23.530 228.000 ;
        RECT 23.130 227.200 23.530 227.800 ;
        RECT 19.530 227.000 23.530 227.200 ;
        RECT 23.130 226.400 23.530 227.000 ;
        RECT 19.530 226.200 23.530 226.400 ;
        RECT 23.130 225.600 23.530 226.200 ;
        RECT 19.530 225.400 23.530 225.600 ;
        RECT 23.130 224.800 23.530 225.400 ;
        RECT 19.530 224.600 23.530 224.800 ;
        RECT 23.130 224.000 23.530 224.600 ;
        RECT 19.530 223.800 23.530 224.000 ;
        RECT 23.130 223.200 23.530 223.800 ;
        RECT 19.530 223.000 23.530 223.200 ;
        RECT 23.130 222.400 23.530 223.000 ;
        RECT 19.530 222.200 23.530 222.400 ;
        RECT 25.930 237.600 29.930 237.800 ;
        RECT 25.930 237.000 26.330 237.600 ;
        RECT 25.930 236.800 29.930 237.000 ;
        RECT 25.930 236.200 26.330 236.800 ;
        RECT 25.930 236.000 29.930 236.200 ;
        RECT 25.930 235.400 26.330 236.000 ;
        RECT 25.930 235.200 29.930 235.400 ;
        RECT 25.930 234.600 26.330 235.200 ;
        RECT 25.930 234.400 29.930 234.600 ;
        RECT 25.930 233.800 26.330 234.400 ;
        RECT 25.930 233.600 29.930 233.800 ;
        RECT 25.930 233.000 26.330 233.600 ;
        RECT 25.930 232.800 29.930 233.000 ;
        RECT 25.930 232.200 26.330 232.800 ;
        RECT 25.930 232.000 29.930 232.200 ;
        RECT 25.930 231.400 26.330 232.000 ;
        RECT 25.930 231.200 29.930 231.400 ;
        RECT 25.930 230.600 26.330 231.200 ;
        RECT 25.930 230.400 29.930 230.600 ;
        RECT 25.930 230.200 26.330 230.400 ;
        RECT 30.680 230.200 30.880 237.800 ;
        RECT 31.480 230.200 31.680 237.800 ;
        RECT 32.280 230.200 32.480 237.800 ;
        RECT 33.080 230.200 33.280 237.800 ;
        RECT 33.880 230.200 34.080 237.800 ;
        RECT 25.930 229.800 34.080 230.200 ;
        RECT 25.930 229.600 26.330 229.800 ;
        RECT 25.930 229.400 29.930 229.600 ;
        RECT 25.930 228.800 26.330 229.400 ;
        RECT 25.930 228.600 29.930 228.800 ;
        RECT 25.930 228.000 26.330 228.600 ;
        RECT 25.930 227.800 29.930 228.000 ;
        RECT 25.930 227.200 26.330 227.800 ;
        RECT 25.930 227.000 29.930 227.200 ;
        RECT 25.930 226.400 26.330 227.000 ;
        RECT 25.930 226.200 29.930 226.400 ;
        RECT 25.930 225.600 26.330 226.200 ;
        RECT 25.930 225.400 29.930 225.600 ;
        RECT 25.930 224.800 26.330 225.400 ;
        RECT 25.930 224.600 29.930 224.800 ;
        RECT 25.930 224.000 26.330 224.600 ;
        RECT 25.930 223.800 29.930 224.000 ;
        RECT 25.930 223.200 26.330 223.800 ;
        RECT 25.930 223.000 29.930 223.200 ;
        RECT 25.930 222.400 26.330 223.000 ;
        RECT 25.930 222.200 29.930 222.400 ;
        RECT 30.680 222.200 30.880 229.800 ;
        RECT 31.480 222.200 31.680 229.800 ;
        RECT 32.280 222.200 32.480 229.800 ;
        RECT 33.080 222.200 33.280 229.800 ;
        RECT 33.880 222.200 34.080 229.800 ;
        RECT 35.380 230.200 35.580 237.800 ;
        RECT 36.180 230.200 36.380 237.800 ;
        RECT 36.980 230.200 37.180 237.800 ;
        RECT 37.780 230.200 37.980 237.800 ;
        RECT 38.580 230.200 38.780 237.800 ;
        RECT 39.530 237.600 43.530 237.800 ;
        RECT 43.130 237.000 43.530 237.600 ;
        RECT 39.530 236.800 43.530 237.000 ;
        RECT 43.130 236.200 43.530 236.800 ;
        RECT 39.530 236.000 43.530 236.200 ;
        RECT 43.130 235.400 43.530 236.000 ;
        RECT 39.530 235.200 43.530 235.400 ;
        RECT 43.130 234.600 43.530 235.200 ;
        RECT 39.530 234.400 43.530 234.600 ;
        RECT 43.130 233.800 43.530 234.400 ;
        RECT 39.530 233.600 43.530 233.800 ;
        RECT 43.130 233.000 43.530 233.600 ;
        RECT 39.530 232.800 43.530 233.000 ;
        RECT 43.130 232.200 43.530 232.800 ;
        RECT 39.530 232.000 43.530 232.200 ;
        RECT 43.130 231.400 43.530 232.000 ;
        RECT 39.530 231.200 43.530 231.400 ;
        RECT 43.130 230.600 43.530 231.200 ;
        RECT 39.530 230.400 43.530 230.600 ;
        RECT 43.130 230.200 43.530 230.400 ;
        RECT 35.380 229.800 43.530 230.200 ;
        RECT 35.380 222.200 35.580 229.800 ;
        RECT 36.180 222.200 36.380 229.800 ;
        RECT 36.980 222.200 37.180 229.800 ;
        RECT 37.780 222.200 37.980 229.800 ;
        RECT 38.580 222.200 38.780 229.800 ;
        RECT 43.130 229.600 43.530 229.800 ;
        RECT 39.530 229.400 43.530 229.600 ;
        RECT 43.130 228.800 43.530 229.400 ;
        RECT 39.530 228.600 43.530 228.800 ;
        RECT 43.130 228.000 43.530 228.600 ;
        RECT 39.530 227.800 43.530 228.000 ;
        RECT 43.130 227.200 43.530 227.800 ;
        RECT 39.530 227.000 43.530 227.200 ;
        RECT 43.130 226.400 43.530 227.000 ;
        RECT 39.530 226.200 43.530 226.400 ;
        RECT 43.130 225.600 43.530 226.200 ;
        RECT 39.530 225.400 43.530 225.600 ;
        RECT 43.130 224.800 43.530 225.400 ;
        RECT 39.530 224.600 43.530 224.800 ;
        RECT 43.130 224.000 43.530 224.600 ;
        RECT 39.530 223.800 43.530 224.000 ;
        RECT 43.130 223.200 43.530 223.800 ;
        RECT 39.530 223.000 43.530 223.200 ;
        RECT 43.130 222.400 43.530 223.000 ;
        RECT 39.530 222.200 43.530 222.400 ;
        RECT 45.930 237.600 49.930 237.800 ;
        RECT 45.930 237.000 46.330 237.600 ;
        RECT 45.930 236.800 49.930 237.000 ;
        RECT 45.930 236.200 46.330 236.800 ;
        RECT 45.930 236.000 49.930 236.200 ;
        RECT 45.930 235.400 46.330 236.000 ;
        RECT 45.930 235.200 49.930 235.400 ;
        RECT 45.930 234.600 46.330 235.200 ;
        RECT 45.930 234.400 49.930 234.600 ;
        RECT 45.930 233.800 46.330 234.400 ;
        RECT 45.930 233.600 49.930 233.800 ;
        RECT 45.930 233.000 46.330 233.600 ;
        RECT 45.930 232.800 49.930 233.000 ;
        RECT 45.930 232.200 46.330 232.800 ;
        RECT 45.930 232.000 49.930 232.200 ;
        RECT 45.930 231.400 46.330 232.000 ;
        RECT 45.930 231.200 49.930 231.400 ;
        RECT 45.930 230.600 46.330 231.200 ;
        RECT 45.930 230.400 49.930 230.600 ;
        RECT 45.930 230.200 46.330 230.400 ;
        RECT 50.680 230.200 50.880 237.800 ;
        RECT 51.480 230.200 51.680 237.800 ;
        RECT 52.280 230.200 52.480 237.800 ;
        RECT 53.080 230.200 53.280 237.800 ;
        RECT 53.880 230.200 54.080 237.800 ;
        RECT 45.930 229.800 54.080 230.200 ;
        RECT 45.930 229.600 46.330 229.800 ;
        RECT 45.930 229.400 49.930 229.600 ;
        RECT 45.930 228.800 46.330 229.400 ;
        RECT 45.930 228.600 49.930 228.800 ;
        RECT 45.930 228.000 46.330 228.600 ;
        RECT 45.930 227.800 49.930 228.000 ;
        RECT 45.930 227.200 46.330 227.800 ;
        RECT 45.930 227.000 49.930 227.200 ;
        RECT 45.930 226.400 46.330 227.000 ;
        RECT 45.930 226.200 49.930 226.400 ;
        RECT 45.930 225.600 46.330 226.200 ;
        RECT 45.930 225.400 49.930 225.600 ;
        RECT 45.930 224.800 46.330 225.400 ;
        RECT 45.930 224.600 49.930 224.800 ;
        RECT 45.930 224.000 46.330 224.600 ;
        RECT 45.930 223.800 49.930 224.000 ;
        RECT 45.930 223.200 46.330 223.800 ;
        RECT 45.930 223.000 49.930 223.200 ;
        RECT 45.930 222.400 46.330 223.000 ;
        RECT 45.930 222.200 49.930 222.400 ;
        RECT 50.680 222.200 50.880 229.800 ;
        RECT 51.480 222.200 51.680 229.800 ;
        RECT 52.280 222.200 52.480 229.800 ;
        RECT 53.080 222.200 53.280 229.800 ;
        RECT 53.880 222.200 54.080 229.800 ;
        RECT 55.380 230.200 55.580 237.800 ;
        RECT 56.180 230.200 56.380 237.800 ;
        RECT 56.980 230.200 57.180 237.800 ;
        RECT 57.780 230.200 57.980 237.800 ;
        RECT 58.580 230.200 58.780 237.800 ;
        RECT 59.530 237.600 63.530 237.800 ;
        RECT 63.130 237.000 63.530 237.600 ;
        RECT 59.530 236.800 63.530 237.000 ;
        RECT 63.130 236.200 63.530 236.800 ;
        RECT 59.530 236.000 63.530 236.200 ;
        RECT 63.130 235.400 63.530 236.000 ;
        RECT 59.530 235.200 63.530 235.400 ;
        RECT 63.130 234.600 63.530 235.200 ;
        RECT 59.530 234.400 63.530 234.600 ;
        RECT 63.130 233.800 63.530 234.400 ;
        RECT 59.530 233.600 63.530 233.800 ;
        RECT 63.130 233.000 63.530 233.600 ;
        RECT 59.530 232.800 63.530 233.000 ;
        RECT 63.130 232.200 63.530 232.800 ;
        RECT 59.530 232.000 63.530 232.200 ;
        RECT 63.130 231.400 63.530 232.000 ;
        RECT 59.530 231.200 63.530 231.400 ;
        RECT 63.130 230.600 63.530 231.200 ;
        RECT 59.530 230.400 63.530 230.600 ;
        RECT 63.130 230.200 63.530 230.400 ;
        RECT 55.380 229.800 63.530 230.200 ;
        RECT 55.380 222.200 55.580 229.800 ;
        RECT 56.180 222.200 56.380 229.800 ;
        RECT 56.980 222.200 57.180 229.800 ;
        RECT 57.780 222.200 57.980 229.800 ;
        RECT 58.580 222.200 58.780 229.800 ;
        RECT 63.130 229.600 63.530 229.800 ;
        RECT 59.530 229.400 63.530 229.600 ;
        RECT 63.130 228.800 63.530 229.400 ;
        RECT 59.530 228.600 63.530 228.800 ;
        RECT 63.130 228.000 63.530 228.600 ;
        RECT 59.530 227.800 63.530 228.000 ;
        RECT 63.130 227.200 63.530 227.800 ;
        RECT 59.530 227.000 63.530 227.200 ;
        RECT 63.130 226.400 63.530 227.000 ;
        RECT 59.530 226.200 63.530 226.400 ;
        RECT 63.130 225.600 63.530 226.200 ;
        RECT 59.530 225.400 63.530 225.600 ;
        RECT 63.130 224.800 63.530 225.400 ;
        RECT 59.530 224.600 63.530 224.800 ;
        RECT 63.130 224.000 63.530 224.600 ;
        RECT 59.530 223.800 63.530 224.000 ;
        RECT 63.130 223.200 63.530 223.800 ;
        RECT 59.530 223.000 63.530 223.200 ;
        RECT 63.130 222.400 63.530 223.000 ;
        RECT 59.530 222.200 63.530 222.400 ;
        RECT 65.930 237.600 69.930 237.800 ;
        RECT 65.930 237.000 66.330 237.600 ;
        RECT 65.930 236.800 69.930 237.000 ;
        RECT 65.930 236.200 66.330 236.800 ;
        RECT 65.930 236.000 69.930 236.200 ;
        RECT 65.930 235.400 66.330 236.000 ;
        RECT 65.930 235.200 69.930 235.400 ;
        RECT 65.930 234.600 66.330 235.200 ;
        RECT 65.930 234.400 69.930 234.600 ;
        RECT 65.930 233.800 66.330 234.400 ;
        RECT 65.930 233.600 69.930 233.800 ;
        RECT 65.930 233.000 66.330 233.600 ;
        RECT 65.930 232.800 69.930 233.000 ;
        RECT 65.930 232.200 66.330 232.800 ;
        RECT 65.930 232.000 69.930 232.200 ;
        RECT 65.930 231.400 66.330 232.000 ;
        RECT 65.930 231.200 69.930 231.400 ;
        RECT 65.930 230.600 66.330 231.200 ;
        RECT 65.930 230.400 69.930 230.600 ;
        RECT 65.930 230.200 66.330 230.400 ;
        RECT 70.680 230.200 70.880 237.800 ;
        RECT 71.480 230.200 71.680 237.800 ;
        RECT 72.280 230.200 72.480 237.800 ;
        RECT 73.080 230.200 73.280 237.800 ;
        RECT 73.880 230.200 74.080 237.800 ;
        RECT 65.930 229.800 74.080 230.200 ;
        RECT 65.930 229.600 66.330 229.800 ;
        RECT 65.930 229.400 69.930 229.600 ;
        RECT 65.930 228.800 66.330 229.400 ;
        RECT 65.930 228.600 69.930 228.800 ;
        RECT 65.930 228.000 66.330 228.600 ;
        RECT 65.930 227.800 69.930 228.000 ;
        RECT 65.930 227.200 66.330 227.800 ;
        RECT 65.930 227.000 69.930 227.200 ;
        RECT 65.930 226.400 66.330 227.000 ;
        RECT 65.930 226.200 69.930 226.400 ;
        RECT 65.930 225.600 66.330 226.200 ;
        RECT 65.930 225.400 69.930 225.600 ;
        RECT 65.930 224.800 66.330 225.400 ;
        RECT 65.930 224.600 69.930 224.800 ;
        RECT 65.930 224.000 66.330 224.600 ;
        RECT 65.930 223.800 69.930 224.000 ;
        RECT 65.930 223.200 66.330 223.800 ;
        RECT 65.930 223.000 69.930 223.200 ;
        RECT 65.930 222.400 66.330 223.000 ;
        RECT 65.930 222.200 69.930 222.400 ;
        RECT 70.680 222.200 70.880 229.800 ;
        RECT 71.480 222.200 71.680 229.800 ;
        RECT 72.280 222.200 72.480 229.800 ;
        RECT 73.080 222.200 73.280 229.800 ;
        RECT 73.880 222.200 74.080 229.800 ;
        RECT 75.380 230.200 75.580 237.800 ;
        RECT 76.180 230.200 76.380 237.800 ;
        RECT 76.980 230.200 77.180 237.800 ;
        RECT 77.780 230.200 77.980 237.800 ;
        RECT 78.580 230.200 78.780 237.800 ;
        RECT 79.530 237.600 83.530 237.800 ;
        RECT 83.130 237.000 83.530 237.600 ;
        RECT 79.530 236.800 83.530 237.000 ;
        RECT 83.130 236.200 83.530 236.800 ;
        RECT 79.530 236.000 83.530 236.200 ;
        RECT 83.130 235.400 83.530 236.000 ;
        RECT 79.530 235.200 83.530 235.400 ;
        RECT 83.130 234.600 83.530 235.200 ;
        RECT 79.530 234.400 83.530 234.600 ;
        RECT 83.130 233.800 83.530 234.400 ;
        RECT 79.530 233.600 83.530 233.800 ;
        RECT 83.130 233.000 83.530 233.600 ;
        RECT 79.530 232.800 83.530 233.000 ;
        RECT 83.130 232.200 83.530 232.800 ;
        RECT 79.530 232.000 83.530 232.200 ;
        RECT 83.130 231.400 83.530 232.000 ;
        RECT 79.530 231.200 83.530 231.400 ;
        RECT 83.130 230.600 83.530 231.200 ;
        RECT 79.530 230.400 83.530 230.600 ;
        RECT 83.130 230.200 83.530 230.400 ;
        RECT 75.380 229.800 83.530 230.200 ;
        RECT 75.380 222.200 75.580 229.800 ;
        RECT 76.180 222.200 76.380 229.800 ;
        RECT 76.980 222.200 77.180 229.800 ;
        RECT 77.780 222.200 77.980 229.800 ;
        RECT 78.580 222.200 78.780 229.800 ;
        RECT 83.130 229.600 83.530 229.800 ;
        RECT 79.530 229.400 83.530 229.600 ;
        RECT 83.130 228.800 83.530 229.400 ;
        RECT 79.530 228.600 83.530 228.800 ;
        RECT 83.130 228.000 83.530 228.600 ;
        RECT 79.530 227.800 83.530 228.000 ;
        RECT 83.130 227.200 83.530 227.800 ;
        RECT 79.530 227.000 83.530 227.200 ;
        RECT 83.130 226.400 83.530 227.000 ;
        RECT 79.530 226.200 83.530 226.400 ;
        RECT 83.130 225.600 83.530 226.200 ;
        RECT 79.530 225.400 83.530 225.600 ;
        RECT 83.130 224.800 83.530 225.400 ;
        RECT 79.530 224.600 83.530 224.800 ;
        RECT 83.130 224.000 83.530 224.600 ;
        RECT 79.530 223.800 83.530 224.000 ;
        RECT 83.130 223.200 83.530 223.800 ;
        RECT 79.530 223.000 83.530 223.200 ;
        RECT 83.130 222.400 83.530 223.000 ;
        RECT 79.530 222.200 83.530 222.400 ;
        RECT 85.930 237.600 89.930 237.800 ;
        RECT 85.930 237.000 86.330 237.600 ;
        RECT 85.930 236.800 89.930 237.000 ;
        RECT 85.930 236.200 86.330 236.800 ;
        RECT 85.930 236.000 89.930 236.200 ;
        RECT 85.930 235.400 86.330 236.000 ;
        RECT 85.930 235.200 89.930 235.400 ;
        RECT 85.930 234.600 86.330 235.200 ;
        RECT 85.930 234.400 89.930 234.600 ;
        RECT 85.930 233.800 86.330 234.400 ;
        RECT 85.930 233.600 89.930 233.800 ;
        RECT 85.930 233.000 86.330 233.600 ;
        RECT 85.930 232.800 89.930 233.000 ;
        RECT 85.930 232.200 86.330 232.800 ;
        RECT 85.930 232.000 89.930 232.200 ;
        RECT 85.930 231.400 86.330 232.000 ;
        RECT 85.930 231.200 89.930 231.400 ;
        RECT 85.930 230.600 86.330 231.200 ;
        RECT 85.930 230.400 89.930 230.600 ;
        RECT 85.930 230.200 86.330 230.400 ;
        RECT 90.680 230.200 90.880 237.800 ;
        RECT 91.480 230.200 91.680 237.800 ;
        RECT 92.280 230.200 92.480 237.800 ;
        RECT 93.080 230.200 93.280 237.800 ;
        RECT 93.880 230.200 94.080 237.800 ;
        RECT 85.930 229.800 94.080 230.200 ;
        RECT 85.930 229.600 86.330 229.800 ;
        RECT 85.930 229.400 89.930 229.600 ;
        RECT 85.930 228.800 86.330 229.400 ;
        RECT 85.930 228.600 89.930 228.800 ;
        RECT 85.930 228.000 86.330 228.600 ;
        RECT 85.930 227.800 89.930 228.000 ;
        RECT 85.930 227.200 86.330 227.800 ;
        RECT 85.930 227.000 89.930 227.200 ;
        RECT 85.930 226.400 86.330 227.000 ;
        RECT 85.930 226.200 89.930 226.400 ;
        RECT 85.930 225.600 86.330 226.200 ;
        RECT 85.930 225.400 89.930 225.600 ;
        RECT 85.930 224.800 86.330 225.400 ;
        RECT 85.930 224.600 89.930 224.800 ;
        RECT 85.930 224.000 86.330 224.600 ;
        RECT 85.930 223.800 89.930 224.000 ;
        RECT 85.930 223.200 86.330 223.800 ;
        RECT 85.930 223.000 89.930 223.200 ;
        RECT 85.930 222.400 86.330 223.000 ;
        RECT 85.930 222.200 89.930 222.400 ;
        RECT 90.680 222.200 90.880 229.800 ;
        RECT 91.480 222.200 91.680 229.800 ;
        RECT 92.280 222.200 92.480 229.800 ;
        RECT 93.080 222.200 93.280 229.800 ;
        RECT 93.880 222.200 94.080 229.800 ;
        RECT 95.380 230.200 95.580 237.800 ;
        RECT 96.180 230.200 96.380 237.800 ;
        RECT 96.980 230.200 97.180 237.800 ;
        RECT 97.780 230.200 97.980 237.800 ;
        RECT 98.580 230.200 98.780 237.800 ;
        RECT 99.530 237.600 103.530 237.800 ;
        RECT 103.130 237.000 103.530 237.600 ;
        RECT 99.530 236.800 103.530 237.000 ;
        RECT 103.130 236.200 103.530 236.800 ;
        RECT 99.530 236.000 103.530 236.200 ;
        RECT 103.130 235.400 103.530 236.000 ;
        RECT 99.530 235.200 103.530 235.400 ;
        RECT 103.130 234.600 103.530 235.200 ;
        RECT 99.530 234.400 103.530 234.600 ;
        RECT 103.130 233.800 103.530 234.400 ;
        RECT 99.530 233.600 103.530 233.800 ;
        RECT 103.130 233.000 103.530 233.600 ;
        RECT 99.530 232.800 103.530 233.000 ;
        RECT 103.130 232.200 103.530 232.800 ;
        RECT 99.530 232.000 103.530 232.200 ;
        RECT 103.130 231.400 103.530 232.000 ;
        RECT 99.530 231.200 103.530 231.400 ;
        RECT 103.130 230.600 103.530 231.200 ;
        RECT 99.530 230.400 103.530 230.600 ;
        RECT 103.130 230.200 103.530 230.400 ;
        RECT 95.380 229.800 103.530 230.200 ;
        RECT 95.380 222.200 95.580 229.800 ;
        RECT 96.180 222.200 96.380 229.800 ;
        RECT 96.980 222.200 97.180 229.800 ;
        RECT 97.780 222.200 97.980 229.800 ;
        RECT 98.580 222.200 98.780 229.800 ;
        RECT 103.130 229.600 103.530 229.800 ;
        RECT 99.530 229.400 103.530 229.600 ;
        RECT 103.130 228.800 103.530 229.400 ;
        RECT 99.530 228.600 103.530 228.800 ;
        RECT 103.130 228.000 103.530 228.600 ;
        RECT 99.530 227.800 103.530 228.000 ;
        RECT 103.130 227.200 103.530 227.800 ;
        RECT 99.530 227.000 103.530 227.200 ;
        RECT 103.130 226.400 103.530 227.000 ;
        RECT 99.530 226.200 103.530 226.400 ;
        RECT 103.130 225.600 103.530 226.200 ;
        RECT 99.530 225.400 103.530 225.600 ;
        RECT 103.130 224.800 103.530 225.400 ;
        RECT 99.530 224.600 103.530 224.800 ;
        RECT 103.130 224.000 103.530 224.600 ;
        RECT 99.530 223.800 103.530 224.000 ;
        RECT 103.130 223.200 103.530 223.800 ;
        RECT 99.530 223.000 103.530 223.200 ;
        RECT 103.130 222.400 103.530 223.000 ;
        RECT 99.530 222.200 103.530 222.400 ;
        RECT 105.930 237.600 109.930 237.800 ;
        RECT 105.930 237.000 106.330 237.600 ;
        RECT 105.930 236.800 109.930 237.000 ;
        RECT 105.930 236.200 106.330 236.800 ;
        RECT 105.930 236.000 109.930 236.200 ;
        RECT 105.930 235.400 106.330 236.000 ;
        RECT 105.930 235.200 109.930 235.400 ;
        RECT 105.930 234.600 106.330 235.200 ;
        RECT 105.930 234.400 109.930 234.600 ;
        RECT 105.930 233.800 106.330 234.400 ;
        RECT 105.930 233.600 109.930 233.800 ;
        RECT 105.930 233.000 106.330 233.600 ;
        RECT 105.930 232.800 109.930 233.000 ;
        RECT 105.930 232.200 106.330 232.800 ;
        RECT 105.930 232.000 109.930 232.200 ;
        RECT 105.930 231.400 106.330 232.000 ;
        RECT 105.930 231.200 109.930 231.400 ;
        RECT 105.930 230.600 106.330 231.200 ;
        RECT 105.930 230.400 109.930 230.600 ;
        RECT 105.930 230.200 106.330 230.400 ;
        RECT 110.680 230.200 110.880 237.800 ;
        RECT 111.480 230.200 111.680 237.800 ;
        RECT 112.280 230.200 112.480 237.800 ;
        RECT 113.080 230.200 113.280 237.800 ;
        RECT 113.880 230.200 114.080 237.800 ;
        RECT 105.930 229.800 114.080 230.200 ;
        RECT 105.930 229.600 106.330 229.800 ;
        RECT 105.930 229.400 109.930 229.600 ;
        RECT 105.930 228.800 106.330 229.400 ;
        RECT 105.930 228.600 109.930 228.800 ;
        RECT 105.930 228.000 106.330 228.600 ;
        RECT 105.930 227.800 109.930 228.000 ;
        RECT 105.930 227.200 106.330 227.800 ;
        RECT 105.930 227.000 109.930 227.200 ;
        RECT 105.930 226.400 106.330 227.000 ;
        RECT 105.930 226.200 109.930 226.400 ;
        RECT 105.930 225.600 106.330 226.200 ;
        RECT 105.930 225.400 109.930 225.600 ;
        RECT 105.930 224.800 106.330 225.400 ;
        RECT 105.930 224.600 109.930 224.800 ;
        RECT 105.930 224.000 106.330 224.600 ;
        RECT 105.930 223.800 109.930 224.000 ;
        RECT 105.930 223.200 106.330 223.800 ;
        RECT 105.930 223.000 109.930 223.200 ;
        RECT 105.930 222.400 106.330 223.000 ;
        RECT 105.930 222.200 109.930 222.400 ;
        RECT 110.680 222.200 110.880 229.800 ;
        RECT 111.480 222.200 111.680 229.800 ;
        RECT 112.280 222.200 112.480 229.800 ;
        RECT 113.080 222.200 113.280 229.800 ;
        RECT 113.880 222.200 114.080 229.800 ;
        RECT 115.380 230.200 115.580 237.800 ;
        RECT 116.180 230.200 116.380 237.800 ;
        RECT 116.980 230.200 117.180 237.800 ;
        RECT 117.780 230.200 117.980 237.800 ;
        RECT 118.580 230.200 118.780 237.800 ;
        RECT 119.530 237.600 123.530 237.800 ;
        RECT 123.130 237.000 123.530 237.600 ;
        RECT 119.530 236.800 123.530 237.000 ;
        RECT 123.130 236.200 123.530 236.800 ;
        RECT 119.530 236.000 123.530 236.200 ;
        RECT 123.130 235.400 123.530 236.000 ;
        RECT 119.530 235.200 123.530 235.400 ;
        RECT 123.130 234.600 123.530 235.200 ;
        RECT 119.530 234.400 123.530 234.600 ;
        RECT 123.130 233.800 123.530 234.400 ;
        RECT 119.530 233.600 123.530 233.800 ;
        RECT 123.130 233.000 123.530 233.600 ;
        RECT 119.530 232.800 123.530 233.000 ;
        RECT 123.130 232.200 123.530 232.800 ;
        RECT 119.530 232.000 123.530 232.200 ;
        RECT 123.130 231.400 123.530 232.000 ;
        RECT 119.530 231.200 123.530 231.400 ;
        RECT 123.130 230.600 123.530 231.200 ;
        RECT 119.530 230.400 123.530 230.600 ;
        RECT 130.050 230.410 130.410 230.790 ;
        RECT 130.680 230.410 131.040 230.790 ;
        RECT 131.280 230.410 131.640 230.790 ;
        RECT 123.130 230.200 123.530 230.400 ;
        RECT 115.380 229.800 123.530 230.200 ;
        RECT 130.050 229.820 130.410 230.200 ;
        RECT 130.680 229.820 131.040 230.200 ;
        RECT 131.280 229.820 131.640 230.200 ;
        RECT 115.380 222.200 115.580 229.800 ;
        RECT 116.180 222.200 116.380 229.800 ;
        RECT 116.980 222.200 117.180 229.800 ;
        RECT 117.780 222.200 117.980 229.800 ;
        RECT 118.580 222.200 118.780 229.800 ;
        RECT 123.130 229.600 123.530 229.800 ;
        RECT 119.530 229.400 123.530 229.600 ;
        RECT 123.130 228.800 123.530 229.400 ;
        RECT 119.530 228.600 123.530 228.800 ;
        RECT 123.130 228.000 123.530 228.600 ;
        RECT 119.530 227.800 123.530 228.000 ;
        RECT 123.130 227.200 123.530 227.800 ;
        RECT 119.530 227.000 123.530 227.200 ;
        RECT 123.130 226.400 123.530 227.000 ;
        RECT 119.530 226.200 123.530 226.400 ;
        RECT 123.130 225.600 123.530 226.200 ;
        RECT 119.530 225.400 123.530 225.600 ;
        RECT 123.130 224.800 123.530 225.400 ;
        RECT 119.530 224.600 123.530 224.800 ;
        RECT 123.130 224.000 123.530 224.600 ;
        RECT 119.530 223.800 123.530 224.000 ;
        RECT 123.130 223.200 123.530 223.800 ;
        RECT 119.530 223.000 123.530 223.200 ;
        RECT 123.130 222.400 123.530 223.000 ;
        RECT 119.530 222.200 123.530 222.400 ;
        RECT 5.930 217.600 9.930 217.800 ;
        RECT 5.930 217.000 6.330 217.600 ;
        RECT 5.930 216.800 9.930 217.000 ;
        RECT 5.930 216.200 6.330 216.800 ;
        RECT 5.930 216.000 9.930 216.200 ;
        RECT 5.930 215.400 6.330 216.000 ;
        RECT 5.930 215.200 9.930 215.400 ;
        RECT 5.930 214.600 6.330 215.200 ;
        RECT 5.930 214.400 9.930 214.600 ;
        RECT 5.930 213.800 6.330 214.400 ;
        RECT 5.930 213.600 9.930 213.800 ;
        RECT 5.930 213.000 6.330 213.600 ;
        RECT 5.930 212.800 9.930 213.000 ;
        RECT 5.930 212.200 6.330 212.800 ;
        RECT 5.930 212.000 9.930 212.200 ;
        RECT 5.930 211.400 6.330 212.000 ;
        RECT 5.930 211.200 9.930 211.400 ;
        RECT 5.930 210.600 6.330 211.200 ;
        RECT 5.930 210.400 9.930 210.600 ;
        RECT 5.930 210.200 6.330 210.400 ;
        RECT 10.680 210.200 10.880 217.800 ;
        RECT 11.480 210.200 11.680 217.800 ;
        RECT 12.280 210.200 12.480 217.800 ;
        RECT 13.080 210.200 13.280 217.800 ;
        RECT 13.880 210.200 14.080 217.800 ;
        RECT 5.930 209.800 14.080 210.200 ;
        RECT 5.930 209.600 6.330 209.800 ;
        RECT 5.930 209.400 9.930 209.600 ;
        RECT 5.930 208.800 6.330 209.400 ;
        RECT 5.930 208.600 9.930 208.800 ;
        RECT 5.930 208.000 6.330 208.600 ;
        RECT 5.930 207.800 9.930 208.000 ;
        RECT 5.930 207.200 6.330 207.800 ;
        RECT 5.930 207.000 9.930 207.200 ;
        RECT 5.930 206.400 6.330 207.000 ;
        RECT 5.930 206.200 9.930 206.400 ;
        RECT 5.930 205.600 6.330 206.200 ;
        RECT 5.930 205.400 9.930 205.600 ;
        RECT 5.930 204.800 6.330 205.400 ;
        RECT 5.930 204.600 9.930 204.800 ;
        RECT 5.930 204.000 6.330 204.600 ;
        RECT 5.930 203.800 9.930 204.000 ;
        RECT 5.930 203.200 6.330 203.800 ;
        RECT 5.930 203.000 9.930 203.200 ;
        RECT 5.930 202.400 6.330 203.000 ;
        RECT 5.930 202.200 9.930 202.400 ;
        RECT 10.680 202.200 10.880 209.800 ;
        RECT 11.480 202.200 11.680 209.800 ;
        RECT 12.280 202.200 12.480 209.800 ;
        RECT 13.080 202.200 13.280 209.800 ;
        RECT 13.880 202.200 14.080 209.800 ;
        RECT 15.380 210.200 15.580 217.800 ;
        RECT 16.180 210.200 16.380 217.800 ;
        RECT 16.980 210.200 17.180 217.800 ;
        RECT 17.780 210.200 17.980 217.800 ;
        RECT 18.580 210.200 18.780 217.800 ;
        RECT 19.530 217.600 23.530 217.800 ;
        RECT 23.130 217.000 23.530 217.600 ;
        RECT 19.530 216.800 23.530 217.000 ;
        RECT 23.130 216.200 23.530 216.800 ;
        RECT 19.530 216.000 23.530 216.200 ;
        RECT 23.130 215.400 23.530 216.000 ;
        RECT 19.530 215.200 23.530 215.400 ;
        RECT 23.130 214.600 23.530 215.200 ;
        RECT 19.530 214.400 23.530 214.600 ;
        RECT 23.130 213.800 23.530 214.400 ;
        RECT 19.530 213.600 23.530 213.800 ;
        RECT 23.130 213.000 23.530 213.600 ;
        RECT 19.530 212.800 23.530 213.000 ;
        RECT 23.130 212.200 23.530 212.800 ;
        RECT 19.530 212.000 23.530 212.200 ;
        RECT 23.130 211.400 23.530 212.000 ;
        RECT 19.530 211.200 23.530 211.400 ;
        RECT 23.130 210.600 23.530 211.200 ;
        RECT 19.530 210.400 23.530 210.600 ;
        RECT 23.130 210.200 23.530 210.400 ;
        RECT 15.380 209.800 23.530 210.200 ;
        RECT 15.380 202.200 15.580 209.800 ;
        RECT 16.180 202.200 16.380 209.800 ;
        RECT 16.980 202.200 17.180 209.800 ;
        RECT 17.780 202.200 17.980 209.800 ;
        RECT 18.580 202.200 18.780 209.800 ;
        RECT 23.130 209.600 23.530 209.800 ;
        RECT 19.530 209.400 23.530 209.600 ;
        RECT 23.130 208.800 23.530 209.400 ;
        RECT 19.530 208.600 23.530 208.800 ;
        RECT 23.130 208.000 23.530 208.600 ;
        RECT 19.530 207.800 23.530 208.000 ;
        RECT 23.130 207.200 23.530 207.800 ;
        RECT 19.530 207.000 23.530 207.200 ;
        RECT 23.130 206.400 23.530 207.000 ;
        RECT 19.530 206.200 23.530 206.400 ;
        RECT 23.130 205.600 23.530 206.200 ;
        RECT 19.530 205.400 23.530 205.600 ;
        RECT 23.130 204.800 23.530 205.400 ;
        RECT 19.530 204.600 23.530 204.800 ;
        RECT 23.130 204.000 23.530 204.600 ;
        RECT 19.530 203.800 23.530 204.000 ;
        RECT 23.130 203.200 23.530 203.800 ;
        RECT 19.530 203.000 23.530 203.200 ;
        RECT 23.130 202.400 23.530 203.000 ;
        RECT 19.530 202.200 23.530 202.400 ;
        RECT 25.930 217.600 29.930 217.800 ;
        RECT 25.930 217.000 26.330 217.600 ;
        RECT 25.930 216.800 29.930 217.000 ;
        RECT 25.930 216.200 26.330 216.800 ;
        RECT 25.930 216.000 29.930 216.200 ;
        RECT 25.930 215.400 26.330 216.000 ;
        RECT 25.930 215.200 29.930 215.400 ;
        RECT 25.930 214.600 26.330 215.200 ;
        RECT 25.930 214.400 29.930 214.600 ;
        RECT 25.930 213.800 26.330 214.400 ;
        RECT 25.930 213.600 29.930 213.800 ;
        RECT 25.930 213.000 26.330 213.600 ;
        RECT 25.930 212.800 29.930 213.000 ;
        RECT 25.930 212.200 26.330 212.800 ;
        RECT 25.930 212.000 29.930 212.200 ;
        RECT 25.930 211.400 26.330 212.000 ;
        RECT 25.930 211.200 29.930 211.400 ;
        RECT 25.930 210.600 26.330 211.200 ;
        RECT 25.930 210.400 29.930 210.600 ;
        RECT 25.930 210.200 26.330 210.400 ;
        RECT 30.680 210.200 30.880 217.800 ;
        RECT 31.480 210.200 31.680 217.800 ;
        RECT 32.280 210.200 32.480 217.800 ;
        RECT 33.080 210.200 33.280 217.800 ;
        RECT 33.880 210.200 34.080 217.800 ;
        RECT 25.930 209.800 34.080 210.200 ;
        RECT 25.930 209.600 26.330 209.800 ;
        RECT 25.930 209.400 29.930 209.600 ;
        RECT 25.930 208.800 26.330 209.400 ;
        RECT 25.930 208.600 29.930 208.800 ;
        RECT 25.930 208.000 26.330 208.600 ;
        RECT 25.930 207.800 29.930 208.000 ;
        RECT 25.930 207.200 26.330 207.800 ;
        RECT 25.930 207.000 29.930 207.200 ;
        RECT 25.930 206.400 26.330 207.000 ;
        RECT 25.930 206.200 29.930 206.400 ;
        RECT 25.930 205.600 26.330 206.200 ;
        RECT 25.930 205.400 29.930 205.600 ;
        RECT 25.930 204.800 26.330 205.400 ;
        RECT 25.930 204.600 29.930 204.800 ;
        RECT 25.930 204.000 26.330 204.600 ;
        RECT 25.930 203.800 29.930 204.000 ;
        RECT 25.930 203.200 26.330 203.800 ;
        RECT 25.930 203.000 29.930 203.200 ;
        RECT 25.930 202.400 26.330 203.000 ;
        RECT 25.930 202.200 29.930 202.400 ;
        RECT 30.680 202.200 30.880 209.800 ;
        RECT 31.480 202.200 31.680 209.800 ;
        RECT 32.280 202.200 32.480 209.800 ;
        RECT 33.080 202.200 33.280 209.800 ;
        RECT 33.880 202.200 34.080 209.800 ;
        RECT 35.380 210.200 35.580 217.800 ;
        RECT 36.180 210.200 36.380 217.800 ;
        RECT 36.980 210.200 37.180 217.800 ;
        RECT 37.780 210.200 37.980 217.800 ;
        RECT 38.580 210.200 38.780 217.800 ;
        RECT 39.530 217.600 43.530 217.800 ;
        RECT 43.130 217.000 43.530 217.600 ;
        RECT 39.530 216.800 43.530 217.000 ;
        RECT 43.130 216.200 43.530 216.800 ;
        RECT 39.530 216.000 43.530 216.200 ;
        RECT 43.130 215.400 43.530 216.000 ;
        RECT 39.530 215.200 43.530 215.400 ;
        RECT 43.130 214.600 43.530 215.200 ;
        RECT 39.530 214.400 43.530 214.600 ;
        RECT 43.130 213.800 43.530 214.400 ;
        RECT 39.530 213.600 43.530 213.800 ;
        RECT 43.130 213.000 43.530 213.600 ;
        RECT 39.530 212.800 43.530 213.000 ;
        RECT 43.130 212.200 43.530 212.800 ;
        RECT 39.530 212.000 43.530 212.200 ;
        RECT 43.130 211.400 43.530 212.000 ;
        RECT 39.530 211.200 43.530 211.400 ;
        RECT 43.130 210.600 43.530 211.200 ;
        RECT 39.530 210.400 43.530 210.600 ;
        RECT 43.130 210.200 43.530 210.400 ;
        RECT 35.380 209.800 43.530 210.200 ;
        RECT 35.380 202.200 35.580 209.800 ;
        RECT 36.180 202.200 36.380 209.800 ;
        RECT 36.980 202.200 37.180 209.800 ;
        RECT 37.780 202.200 37.980 209.800 ;
        RECT 38.580 202.200 38.780 209.800 ;
        RECT 43.130 209.600 43.530 209.800 ;
        RECT 39.530 209.400 43.530 209.600 ;
        RECT 43.130 208.800 43.530 209.400 ;
        RECT 39.530 208.600 43.530 208.800 ;
        RECT 43.130 208.000 43.530 208.600 ;
        RECT 39.530 207.800 43.530 208.000 ;
        RECT 43.130 207.200 43.530 207.800 ;
        RECT 39.530 207.000 43.530 207.200 ;
        RECT 43.130 206.400 43.530 207.000 ;
        RECT 39.530 206.200 43.530 206.400 ;
        RECT 43.130 205.600 43.530 206.200 ;
        RECT 39.530 205.400 43.530 205.600 ;
        RECT 43.130 204.800 43.530 205.400 ;
        RECT 39.530 204.600 43.530 204.800 ;
        RECT 43.130 204.000 43.530 204.600 ;
        RECT 39.530 203.800 43.530 204.000 ;
        RECT 43.130 203.200 43.530 203.800 ;
        RECT 39.530 203.000 43.530 203.200 ;
        RECT 43.130 202.400 43.530 203.000 ;
        RECT 39.530 202.200 43.530 202.400 ;
        RECT 45.930 217.600 49.930 217.800 ;
        RECT 45.930 217.000 46.330 217.600 ;
        RECT 45.930 216.800 49.930 217.000 ;
        RECT 45.930 216.200 46.330 216.800 ;
        RECT 45.930 216.000 49.930 216.200 ;
        RECT 45.930 215.400 46.330 216.000 ;
        RECT 45.930 215.200 49.930 215.400 ;
        RECT 45.930 214.600 46.330 215.200 ;
        RECT 45.930 214.400 49.930 214.600 ;
        RECT 45.930 213.800 46.330 214.400 ;
        RECT 45.930 213.600 49.930 213.800 ;
        RECT 45.930 213.000 46.330 213.600 ;
        RECT 45.930 212.800 49.930 213.000 ;
        RECT 45.930 212.200 46.330 212.800 ;
        RECT 45.930 212.000 49.930 212.200 ;
        RECT 45.930 211.400 46.330 212.000 ;
        RECT 45.930 211.200 49.930 211.400 ;
        RECT 45.930 210.600 46.330 211.200 ;
        RECT 45.930 210.400 49.930 210.600 ;
        RECT 45.930 210.200 46.330 210.400 ;
        RECT 50.680 210.200 50.880 217.800 ;
        RECT 51.480 210.200 51.680 217.800 ;
        RECT 52.280 210.200 52.480 217.800 ;
        RECT 53.080 210.200 53.280 217.800 ;
        RECT 53.880 210.200 54.080 217.800 ;
        RECT 45.930 209.800 54.080 210.200 ;
        RECT 45.930 209.600 46.330 209.800 ;
        RECT 45.930 209.400 49.930 209.600 ;
        RECT 45.930 208.800 46.330 209.400 ;
        RECT 45.930 208.600 49.930 208.800 ;
        RECT 45.930 208.000 46.330 208.600 ;
        RECT 45.930 207.800 49.930 208.000 ;
        RECT 45.930 207.200 46.330 207.800 ;
        RECT 45.930 207.000 49.930 207.200 ;
        RECT 45.930 206.400 46.330 207.000 ;
        RECT 45.930 206.200 49.930 206.400 ;
        RECT 45.930 205.600 46.330 206.200 ;
        RECT 45.930 205.400 49.930 205.600 ;
        RECT 45.930 204.800 46.330 205.400 ;
        RECT 45.930 204.600 49.930 204.800 ;
        RECT 45.930 204.000 46.330 204.600 ;
        RECT 45.930 203.800 49.930 204.000 ;
        RECT 45.930 203.200 46.330 203.800 ;
        RECT 45.930 203.000 49.930 203.200 ;
        RECT 45.930 202.400 46.330 203.000 ;
        RECT 45.930 202.200 49.930 202.400 ;
        RECT 50.680 202.200 50.880 209.800 ;
        RECT 51.480 202.200 51.680 209.800 ;
        RECT 52.280 202.200 52.480 209.800 ;
        RECT 53.080 202.200 53.280 209.800 ;
        RECT 53.880 202.200 54.080 209.800 ;
        RECT 55.380 210.200 55.580 217.800 ;
        RECT 56.180 210.200 56.380 217.800 ;
        RECT 56.980 210.200 57.180 217.800 ;
        RECT 57.780 210.200 57.980 217.800 ;
        RECT 58.580 210.200 58.780 217.800 ;
        RECT 59.530 217.600 63.530 217.800 ;
        RECT 63.130 217.000 63.530 217.600 ;
        RECT 59.530 216.800 63.530 217.000 ;
        RECT 63.130 216.200 63.530 216.800 ;
        RECT 59.530 216.000 63.530 216.200 ;
        RECT 63.130 215.400 63.530 216.000 ;
        RECT 59.530 215.200 63.530 215.400 ;
        RECT 63.130 214.600 63.530 215.200 ;
        RECT 59.530 214.400 63.530 214.600 ;
        RECT 63.130 213.800 63.530 214.400 ;
        RECT 59.530 213.600 63.530 213.800 ;
        RECT 63.130 213.000 63.530 213.600 ;
        RECT 59.530 212.800 63.530 213.000 ;
        RECT 63.130 212.200 63.530 212.800 ;
        RECT 59.530 212.000 63.530 212.200 ;
        RECT 63.130 211.400 63.530 212.000 ;
        RECT 59.530 211.200 63.530 211.400 ;
        RECT 63.130 210.600 63.530 211.200 ;
        RECT 59.530 210.400 63.530 210.600 ;
        RECT 63.130 210.200 63.530 210.400 ;
        RECT 55.380 209.800 63.530 210.200 ;
        RECT 55.380 202.200 55.580 209.800 ;
        RECT 56.180 202.200 56.380 209.800 ;
        RECT 56.980 202.200 57.180 209.800 ;
        RECT 57.780 202.200 57.980 209.800 ;
        RECT 58.580 202.200 58.780 209.800 ;
        RECT 63.130 209.600 63.530 209.800 ;
        RECT 59.530 209.400 63.530 209.600 ;
        RECT 63.130 208.800 63.530 209.400 ;
        RECT 59.530 208.600 63.530 208.800 ;
        RECT 63.130 208.000 63.530 208.600 ;
        RECT 59.530 207.800 63.530 208.000 ;
        RECT 63.130 207.200 63.530 207.800 ;
        RECT 59.530 207.000 63.530 207.200 ;
        RECT 63.130 206.400 63.530 207.000 ;
        RECT 59.530 206.200 63.530 206.400 ;
        RECT 63.130 205.600 63.530 206.200 ;
        RECT 59.530 205.400 63.530 205.600 ;
        RECT 63.130 204.800 63.530 205.400 ;
        RECT 59.530 204.600 63.530 204.800 ;
        RECT 63.130 204.000 63.530 204.600 ;
        RECT 59.530 203.800 63.530 204.000 ;
        RECT 63.130 203.200 63.530 203.800 ;
        RECT 59.530 203.000 63.530 203.200 ;
        RECT 63.130 202.400 63.530 203.000 ;
        RECT 59.530 202.200 63.530 202.400 ;
        RECT 65.930 217.600 69.930 217.800 ;
        RECT 65.930 217.000 66.330 217.600 ;
        RECT 65.930 216.800 69.930 217.000 ;
        RECT 65.930 216.200 66.330 216.800 ;
        RECT 65.930 216.000 69.930 216.200 ;
        RECT 65.930 215.400 66.330 216.000 ;
        RECT 65.930 215.200 69.930 215.400 ;
        RECT 65.930 214.600 66.330 215.200 ;
        RECT 65.930 214.400 69.930 214.600 ;
        RECT 65.930 213.800 66.330 214.400 ;
        RECT 65.930 213.600 69.930 213.800 ;
        RECT 65.930 213.000 66.330 213.600 ;
        RECT 65.930 212.800 69.930 213.000 ;
        RECT 65.930 212.200 66.330 212.800 ;
        RECT 65.930 212.000 69.930 212.200 ;
        RECT 65.930 211.400 66.330 212.000 ;
        RECT 65.930 211.200 69.930 211.400 ;
        RECT 65.930 210.600 66.330 211.200 ;
        RECT 65.930 210.400 69.930 210.600 ;
        RECT 65.930 210.200 66.330 210.400 ;
        RECT 70.680 210.200 70.880 217.800 ;
        RECT 71.480 210.200 71.680 217.800 ;
        RECT 72.280 210.200 72.480 217.800 ;
        RECT 73.080 210.200 73.280 217.800 ;
        RECT 73.880 210.200 74.080 217.800 ;
        RECT 65.930 209.800 74.080 210.200 ;
        RECT 65.930 209.600 66.330 209.800 ;
        RECT 65.930 209.400 69.930 209.600 ;
        RECT 65.930 208.800 66.330 209.400 ;
        RECT 65.930 208.600 69.930 208.800 ;
        RECT 65.930 208.000 66.330 208.600 ;
        RECT 65.930 207.800 69.930 208.000 ;
        RECT 65.930 207.200 66.330 207.800 ;
        RECT 65.930 207.000 69.930 207.200 ;
        RECT 65.930 206.400 66.330 207.000 ;
        RECT 65.930 206.200 69.930 206.400 ;
        RECT 65.930 205.600 66.330 206.200 ;
        RECT 65.930 205.400 69.930 205.600 ;
        RECT 65.930 204.800 66.330 205.400 ;
        RECT 65.930 204.600 69.930 204.800 ;
        RECT 65.930 204.000 66.330 204.600 ;
        RECT 65.930 203.800 69.930 204.000 ;
        RECT 65.930 203.200 66.330 203.800 ;
        RECT 65.930 203.000 69.930 203.200 ;
        RECT 65.930 202.400 66.330 203.000 ;
        RECT 65.930 202.200 69.930 202.400 ;
        RECT 70.680 202.200 70.880 209.800 ;
        RECT 71.480 202.200 71.680 209.800 ;
        RECT 72.280 202.200 72.480 209.800 ;
        RECT 73.080 202.200 73.280 209.800 ;
        RECT 73.880 202.200 74.080 209.800 ;
        RECT 75.380 210.200 75.580 217.800 ;
        RECT 76.180 210.200 76.380 217.800 ;
        RECT 76.980 210.200 77.180 217.800 ;
        RECT 77.780 210.200 77.980 217.800 ;
        RECT 78.580 210.200 78.780 217.800 ;
        RECT 79.530 217.600 83.530 217.800 ;
        RECT 83.130 217.000 83.530 217.600 ;
        RECT 79.530 216.800 83.530 217.000 ;
        RECT 83.130 216.200 83.530 216.800 ;
        RECT 79.530 216.000 83.530 216.200 ;
        RECT 83.130 215.400 83.530 216.000 ;
        RECT 79.530 215.200 83.530 215.400 ;
        RECT 83.130 214.600 83.530 215.200 ;
        RECT 79.530 214.400 83.530 214.600 ;
        RECT 83.130 213.800 83.530 214.400 ;
        RECT 79.530 213.600 83.530 213.800 ;
        RECT 83.130 213.000 83.530 213.600 ;
        RECT 79.530 212.800 83.530 213.000 ;
        RECT 83.130 212.200 83.530 212.800 ;
        RECT 79.530 212.000 83.530 212.200 ;
        RECT 83.130 211.400 83.530 212.000 ;
        RECT 79.530 211.200 83.530 211.400 ;
        RECT 83.130 210.600 83.530 211.200 ;
        RECT 79.530 210.400 83.530 210.600 ;
        RECT 83.130 210.200 83.530 210.400 ;
        RECT 75.380 209.800 83.530 210.200 ;
        RECT 75.380 202.200 75.580 209.800 ;
        RECT 76.180 202.200 76.380 209.800 ;
        RECT 76.980 202.200 77.180 209.800 ;
        RECT 77.780 202.200 77.980 209.800 ;
        RECT 78.580 202.200 78.780 209.800 ;
        RECT 83.130 209.600 83.530 209.800 ;
        RECT 79.530 209.400 83.530 209.600 ;
        RECT 83.130 208.800 83.530 209.400 ;
        RECT 79.530 208.600 83.530 208.800 ;
        RECT 83.130 208.000 83.530 208.600 ;
        RECT 79.530 207.800 83.530 208.000 ;
        RECT 83.130 207.200 83.530 207.800 ;
        RECT 79.530 207.000 83.530 207.200 ;
        RECT 83.130 206.400 83.530 207.000 ;
        RECT 79.530 206.200 83.530 206.400 ;
        RECT 83.130 205.600 83.530 206.200 ;
        RECT 79.530 205.400 83.530 205.600 ;
        RECT 83.130 204.800 83.530 205.400 ;
        RECT 79.530 204.600 83.530 204.800 ;
        RECT 83.130 204.000 83.530 204.600 ;
        RECT 79.530 203.800 83.530 204.000 ;
        RECT 83.130 203.200 83.530 203.800 ;
        RECT 79.530 203.000 83.530 203.200 ;
        RECT 83.130 202.400 83.530 203.000 ;
        RECT 79.530 202.200 83.530 202.400 ;
        RECT 85.930 217.600 89.930 217.800 ;
        RECT 85.930 217.000 86.330 217.600 ;
        RECT 85.930 216.800 89.930 217.000 ;
        RECT 85.930 216.200 86.330 216.800 ;
        RECT 85.930 216.000 89.930 216.200 ;
        RECT 85.930 215.400 86.330 216.000 ;
        RECT 85.930 215.200 89.930 215.400 ;
        RECT 85.930 214.600 86.330 215.200 ;
        RECT 85.930 214.400 89.930 214.600 ;
        RECT 85.930 213.800 86.330 214.400 ;
        RECT 85.930 213.600 89.930 213.800 ;
        RECT 85.930 213.000 86.330 213.600 ;
        RECT 85.930 212.800 89.930 213.000 ;
        RECT 85.930 212.200 86.330 212.800 ;
        RECT 85.930 212.000 89.930 212.200 ;
        RECT 85.930 211.400 86.330 212.000 ;
        RECT 85.930 211.200 89.930 211.400 ;
        RECT 85.930 210.600 86.330 211.200 ;
        RECT 85.930 210.400 89.930 210.600 ;
        RECT 85.930 210.200 86.330 210.400 ;
        RECT 90.680 210.200 90.880 217.800 ;
        RECT 91.480 210.200 91.680 217.800 ;
        RECT 92.280 210.200 92.480 217.800 ;
        RECT 93.080 210.200 93.280 217.800 ;
        RECT 93.880 210.200 94.080 217.800 ;
        RECT 85.930 209.800 94.080 210.200 ;
        RECT 85.930 209.600 86.330 209.800 ;
        RECT 85.930 209.400 89.930 209.600 ;
        RECT 85.930 208.800 86.330 209.400 ;
        RECT 85.930 208.600 89.930 208.800 ;
        RECT 85.930 208.000 86.330 208.600 ;
        RECT 85.930 207.800 89.930 208.000 ;
        RECT 85.930 207.200 86.330 207.800 ;
        RECT 85.930 207.000 89.930 207.200 ;
        RECT 85.930 206.400 86.330 207.000 ;
        RECT 85.930 206.200 89.930 206.400 ;
        RECT 85.930 205.600 86.330 206.200 ;
        RECT 85.930 205.400 89.930 205.600 ;
        RECT 85.930 204.800 86.330 205.400 ;
        RECT 85.930 204.600 89.930 204.800 ;
        RECT 85.930 204.000 86.330 204.600 ;
        RECT 85.930 203.800 89.930 204.000 ;
        RECT 85.930 203.200 86.330 203.800 ;
        RECT 85.930 203.000 89.930 203.200 ;
        RECT 85.930 202.400 86.330 203.000 ;
        RECT 85.930 202.200 89.930 202.400 ;
        RECT 90.680 202.200 90.880 209.800 ;
        RECT 91.480 202.200 91.680 209.800 ;
        RECT 92.280 202.200 92.480 209.800 ;
        RECT 93.080 202.200 93.280 209.800 ;
        RECT 93.880 202.200 94.080 209.800 ;
        RECT 95.380 210.200 95.580 217.800 ;
        RECT 96.180 210.200 96.380 217.800 ;
        RECT 96.980 210.200 97.180 217.800 ;
        RECT 97.780 210.200 97.980 217.800 ;
        RECT 98.580 210.200 98.780 217.800 ;
        RECT 99.530 217.600 103.530 217.800 ;
        RECT 103.130 217.000 103.530 217.600 ;
        RECT 99.530 216.800 103.530 217.000 ;
        RECT 103.130 216.200 103.530 216.800 ;
        RECT 99.530 216.000 103.530 216.200 ;
        RECT 103.130 215.400 103.530 216.000 ;
        RECT 99.530 215.200 103.530 215.400 ;
        RECT 103.130 214.600 103.530 215.200 ;
        RECT 99.530 214.400 103.530 214.600 ;
        RECT 103.130 213.800 103.530 214.400 ;
        RECT 99.530 213.600 103.530 213.800 ;
        RECT 103.130 213.000 103.530 213.600 ;
        RECT 99.530 212.800 103.530 213.000 ;
        RECT 103.130 212.200 103.530 212.800 ;
        RECT 99.530 212.000 103.530 212.200 ;
        RECT 103.130 211.400 103.530 212.000 ;
        RECT 99.530 211.200 103.530 211.400 ;
        RECT 103.130 210.600 103.530 211.200 ;
        RECT 99.530 210.400 103.530 210.600 ;
        RECT 103.130 210.200 103.530 210.400 ;
        RECT 95.380 209.800 103.530 210.200 ;
        RECT 95.380 202.200 95.580 209.800 ;
        RECT 96.180 202.200 96.380 209.800 ;
        RECT 96.980 202.200 97.180 209.800 ;
        RECT 97.780 202.200 97.980 209.800 ;
        RECT 98.580 202.200 98.780 209.800 ;
        RECT 103.130 209.600 103.530 209.800 ;
        RECT 99.530 209.400 103.530 209.600 ;
        RECT 103.130 208.800 103.530 209.400 ;
        RECT 99.530 208.600 103.530 208.800 ;
        RECT 103.130 208.000 103.530 208.600 ;
        RECT 99.530 207.800 103.530 208.000 ;
        RECT 103.130 207.200 103.530 207.800 ;
        RECT 99.530 207.000 103.530 207.200 ;
        RECT 103.130 206.400 103.530 207.000 ;
        RECT 99.530 206.200 103.530 206.400 ;
        RECT 103.130 205.600 103.530 206.200 ;
        RECT 99.530 205.400 103.530 205.600 ;
        RECT 103.130 204.800 103.530 205.400 ;
        RECT 99.530 204.600 103.530 204.800 ;
        RECT 103.130 204.000 103.530 204.600 ;
        RECT 99.530 203.800 103.530 204.000 ;
        RECT 103.130 203.200 103.530 203.800 ;
        RECT 99.530 203.000 103.530 203.200 ;
        RECT 103.130 202.400 103.530 203.000 ;
        RECT 99.530 202.200 103.530 202.400 ;
        RECT 105.930 217.600 109.930 217.800 ;
        RECT 105.930 217.000 106.330 217.600 ;
        RECT 105.930 216.800 109.930 217.000 ;
        RECT 105.930 216.200 106.330 216.800 ;
        RECT 105.930 216.000 109.930 216.200 ;
        RECT 105.930 215.400 106.330 216.000 ;
        RECT 105.930 215.200 109.930 215.400 ;
        RECT 105.930 214.600 106.330 215.200 ;
        RECT 105.930 214.400 109.930 214.600 ;
        RECT 105.930 213.800 106.330 214.400 ;
        RECT 105.930 213.600 109.930 213.800 ;
        RECT 105.930 213.000 106.330 213.600 ;
        RECT 105.930 212.800 109.930 213.000 ;
        RECT 105.930 212.200 106.330 212.800 ;
        RECT 105.930 212.000 109.930 212.200 ;
        RECT 105.930 211.400 106.330 212.000 ;
        RECT 105.930 211.200 109.930 211.400 ;
        RECT 105.930 210.600 106.330 211.200 ;
        RECT 105.930 210.400 109.930 210.600 ;
        RECT 105.930 210.200 106.330 210.400 ;
        RECT 110.680 210.200 110.880 217.800 ;
        RECT 111.480 210.200 111.680 217.800 ;
        RECT 112.280 210.200 112.480 217.800 ;
        RECT 113.080 210.200 113.280 217.800 ;
        RECT 113.880 210.200 114.080 217.800 ;
        RECT 105.930 209.800 114.080 210.200 ;
        RECT 105.930 209.600 106.330 209.800 ;
        RECT 105.930 209.400 109.930 209.600 ;
        RECT 105.930 208.800 106.330 209.400 ;
        RECT 105.930 208.600 109.930 208.800 ;
        RECT 105.930 208.000 106.330 208.600 ;
        RECT 105.930 207.800 109.930 208.000 ;
        RECT 105.930 207.200 106.330 207.800 ;
        RECT 105.930 207.000 109.930 207.200 ;
        RECT 105.930 206.400 106.330 207.000 ;
        RECT 105.930 206.200 109.930 206.400 ;
        RECT 105.930 205.600 106.330 206.200 ;
        RECT 105.930 205.400 109.930 205.600 ;
        RECT 105.930 204.800 106.330 205.400 ;
        RECT 105.930 204.600 109.930 204.800 ;
        RECT 105.930 204.000 106.330 204.600 ;
        RECT 105.930 203.800 109.930 204.000 ;
        RECT 105.930 203.200 106.330 203.800 ;
        RECT 105.930 203.000 109.930 203.200 ;
        RECT 105.930 202.400 106.330 203.000 ;
        RECT 105.930 202.200 109.930 202.400 ;
        RECT 110.680 202.200 110.880 209.800 ;
        RECT 111.480 202.200 111.680 209.800 ;
        RECT 112.280 202.200 112.480 209.800 ;
        RECT 113.080 202.200 113.280 209.800 ;
        RECT 113.880 202.200 114.080 209.800 ;
        RECT 115.380 210.200 115.580 217.800 ;
        RECT 116.180 210.200 116.380 217.800 ;
        RECT 116.980 210.200 117.180 217.800 ;
        RECT 117.780 210.200 117.980 217.800 ;
        RECT 118.580 210.200 118.780 217.800 ;
        RECT 119.530 217.600 123.530 217.800 ;
        RECT 123.130 217.000 123.530 217.600 ;
        RECT 119.530 216.800 123.530 217.000 ;
        RECT 123.130 216.200 123.530 216.800 ;
        RECT 119.530 216.000 123.530 216.200 ;
        RECT 123.130 215.400 123.530 216.000 ;
        RECT 119.530 215.200 123.530 215.400 ;
        RECT 123.130 214.600 123.530 215.200 ;
        RECT 119.530 214.400 123.530 214.600 ;
        RECT 123.130 213.800 123.530 214.400 ;
        RECT 119.530 213.600 123.530 213.800 ;
        RECT 123.130 213.000 123.530 213.600 ;
        RECT 119.530 212.800 123.530 213.000 ;
        RECT 123.130 212.200 123.530 212.800 ;
        RECT 119.530 212.000 123.530 212.200 ;
        RECT 123.130 211.400 123.530 212.000 ;
        RECT 119.530 211.200 123.530 211.400 ;
        RECT 123.130 210.600 123.530 211.200 ;
        RECT 119.530 210.400 123.530 210.600 ;
        RECT 123.130 210.200 123.530 210.400 ;
        RECT 115.380 209.800 123.530 210.200 ;
        RECT 115.380 202.200 115.580 209.800 ;
        RECT 116.180 202.200 116.380 209.800 ;
        RECT 116.980 202.200 117.180 209.800 ;
        RECT 117.780 202.200 117.980 209.800 ;
        RECT 118.580 202.200 118.780 209.800 ;
        RECT 123.130 209.600 123.530 209.800 ;
        RECT 119.530 209.400 123.530 209.600 ;
        RECT 123.130 208.800 123.530 209.400 ;
        RECT 130.050 209.120 130.410 209.500 ;
        RECT 130.680 209.120 131.040 209.500 ;
        RECT 131.280 209.120 131.640 209.500 ;
        RECT 119.530 208.600 123.530 208.800 ;
        RECT 123.130 208.000 123.530 208.600 ;
        RECT 130.050 208.530 130.410 208.910 ;
        RECT 130.680 208.530 131.040 208.910 ;
        RECT 131.280 208.530 131.640 208.910 ;
        RECT 119.530 207.800 123.530 208.000 ;
        RECT 123.130 207.200 123.530 207.800 ;
        RECT 119.530 207.000 123.530 207.200 ;
        RECT 123.130 206.400 123.530 207.000 ;
        RECT 119.530 206.200 123.530 206.400 ;
        RECT 123.130 205.600 123.530 206.200 ;
        RECT 119.530 205.400 123.530 205.600 ;
        RECT 123.130 204.800 123.530 205.400 ;
        RECT 119.530 204.600 123.530 204.800 ;
        RECT 123.130 204.000 123.530 204.600 ;
        RECT 119.530 203.800 123.530 204.000 ;
        RECT 123.130 203.200 123.530 203.800 ;
        RECT 119.530 203.000 123.530 203.200 ;
        RECT 123.130 202.400 123.530 203.000 ;
        RECT 119.530 202.200 123.530 202.400 ;
        RECT 9.340 176.355 12.515 177.050 ;
        RECT 9.340 176.350 10.045 176.355 ;
        RECT 11.755 175.425 12.515 176.355 ;
        RECT 10.175 173.440 10.345 175.425 ;
        RECT 11.755 174.885 12.570 175.425 ;
        RECT 13.965 174.885 14.155 175.425 ;
        RECT 11.755 173.440 11.925 174.885 ;
        RECT 12.395 174.255 12.570 174.885 ;
        RECT 12.400 173.445 12.570 174.255 ;
        RECT 13.980 174.255 14.155 174.885 ;
        RECT 13.980 173.445 14.150 174.255 ;
        RECT 5.930 137.600 9.930 137.800 ;
        RECT 5.930 137.000 6.330 137.600 ;
        RECT 5.930 136.800 9.930 137.000 ;
        RECT 5.930 136.200 6.330 136.800 ;
        RECT 5.930 136.000 9.930 136.200 ;
        RECT 5.930 135.400 6.330 136.000 ;
        RECT 5.930 135.200 9.930 135.400 ;
        RECT 5.930 134.600 6.330 135.200 ;
        RECT 5.930 134.400 9.930 134.600 ;
        RECT 5.930 133.800 6.330 134.400 ;
        RECT 5.930 133.600 9.930 133.800 ;
        RECT 5.930 133.000 6.330 133.600 ;
        RECT 5.930 132.800 9.930 133.000 ;
        RECT 5.930 132.200 6.330 132.800 ;
        RECT 5.930 132.000 9.930 132.200 ;
        RECT 5.930 131.400 6.330 132.000 ;
        RECT 5.930 131.200 9.930 131.400 ;
        RECT 5.930 130.600 6.330 131.200 ;
        RECT 5.930 130.400 9.930 130.600 ;
        RECT 5.930 130.200 6.330 130.400 ;
        RECT 10.680 130.200 10.880 137.800 ;
        RECT 11.480 130.200 11.680 137.800 ;
        RECT 12.280 130.200 12.480 137.800 ;
        RECT 13.080 130.200 13.280 137.800 ;
        RECT 13.880 130.200 14.080 137.800 ;
        RECT 5.930 129.800 14.080 130.200 ;
        RECT 5.930 129.600 6.330 129.800 ;
        RECT 5.930 129.400 9.930 129.600 ;
        RECT 5.930 128.800 6.330 129.400 ;
        RECT 5.930 128.600 9.930 128.800 ;
        RECT 5.930 128.000 6.330 128.600 ;
        RECT 5.930 127.800 9.930 128.000 ;
        RECT 5.930 127.200 6.330 127.800 ;
        RECT 5.930 127.000 9.930 127.200 ;
        RECT 5.930 126.400 6.330 127.000 ;
        RECT 5.930 126.200 9.930 126.400 ;
        RECT 5.930 125.600 6.330 126.200 ;
        RECT 5.930 125.400 9.930 125.600 ;
        RECT 5.930 124.800 6.330 125.400 ;
        RECT 5.930 124.600 9.930 124.800 ;
        RECT 5.930 124.000 6.330 124.600 ;
        RECT 5.930 123.800 9.930 124.000 ;
        RECT 5.930 123.200 6.330 123.800 ;
        RECT 5.930 123.000 9.930 123.200 ;
        RECT 5.930 122.400 6.330 123.000 ;
        RECT 5.930 122.200 9.930 122.400 ;
        RECT 10.680 122.200 10.880 129.800 ;
        RECT 11.480 122.200 11.680 129.800 ;
        RECT 12.280 122.200 12.480 129.800 ;
        RECT 13.080 122.200 13.280 129.800 ;
        RECT 13.880 122.200 14.080 129.800 ;
        RECT 15.380 130.200 15.580 137.800 ;
        RECT 16.180 130.200 16.380 137.800 ;
        RECT 16.980 130.200 17.180 137.800 ;
        RECT 17.780 130.200 17.980 137.800 ;
        RECT 18.580 130.200 18.780 137.800 ;
        RECT 19.530 137.600 23.530 137.800 ;
        RECT 23.130 137.000 23.530 137.600 ;
        RECT 19.530 136.800 23.530 137.000 ;
        RECT 23.130 136.200 23.530 136.800 ;
        RECT 19.530 136.000 23.530 136.200 ;
        RECT 23.130 135.400 23.530 136.000 ;
        RECT 19.530 135.200 23.530 135.400 ;
        RECT 23.130 134.600 23.530 135.200 ;
        RECT 19.530 134.400 23.530 134.600 ;
        RECT 23.130 133.800 23.530 134.400 ;
        RECT 19.530 133.600 23.530 133.800 ;
        RECT 23.130 133.000 23.530 133.600 ;
        RECT 19.530 132.800 23.530 133.000 ;
        RECT 23.130 132.200 23.530 132.800 ;
        RECT 19.530 132.000 23.530 132.200 ;
        RECT 23.130 131.400 23.530 132.000 ;
        RECT 19.530 131.200 23.530 131.400 ;
        RECT 23.130 130.600 23.530 131.200 ;
        RECT 19.530 130.400 23.530 130.600 ;
        RECT 23.130 130.200 23.530 130.400 ;
        RECT 15.380 129.800 23.530 130.200 ;
        RECT 15.380 122.200 15.580 129.800 ;
        RECT 16.180 122.200 16.380 129.800 ;
        RECT 16.980 122.200 17.180 129.800 ;
        RECT 17.780 122.200 17.980 129.800 ;
        RECT 18.580 122.200 18.780 129.800 ;
        RECT 23.130 129.600 23.530 129.800 ;
        RECT 19.530 129.400 23.530 129.600 ;
        RECT 23.130 128.800 23.530 129.400 ;
        RECT 19.530 128.600 23.530 128.800 ;
        RECT 23.130 128.000 23.530 128.600 ;
        RECT 19.530 127.800 23.530 128.000 ;
        RECT 23.130 127.200 23.530 127.800 ;
        RECT 19.530 127.000 23.530 127.200 ;
        RECT 23.130 126.400 23.530 127.000 ;
        RECT 19.530 126.200 23.530 126.400 ;
        RECT 23.130 125.600 23.530 126.200 ;
        RECT 19.530 125.400 23.530 125.600 ;
        RECT 23.130 124.800 23.530 125.400 ;
        RECT 19.530 124.600 23.530 124.800 ;
        RECT 23.130 124.000 23.530 124.600 ;
        RECT 19.530 123.800 23.530 124.000 ;
        RECT 23.130 123.200 23.530 123.800 ;
        RECT 19.530 123.000 23.530 123.200 ;
        RECT 23.130 122.400 23.530 123.000 ;
        RECT 19.530 122.200 23.530 122.400 ;
        RECT 25.930 137.600 29.930 137.800 ;
        RECT 25.930 137.000 26.330 137.600 ;
        RECT 25.930 136.800 29.930 137.000 ;
        RECT 25.930 136.200 26.330 136.800 ;
        RECT 25.930 136.000 29.930 136.200 ;
        RECT 25.930 135.400 26.330 136.000 ;
        RECT 25.930 135.200 29.930 135.400 ;
        RECT 25.930 134.600 26.330 135.200 ;
        RECT 25.930 134.400 29.930 134.600 ;
        RECT 25.930 133.800 26.330 134.400 ;
        RECT 25.930 133.600 29.930 133.800 ;
        RECT 25.930 133.000 26.330 133.600 ;
        RECT 25.930 132.800 29.930 133.000 ;
        RECT 25.930 132.200 26.330 132.800 ;
        RECT 25.930 132.000 29.930 132.200 ;
        RECT 25.930 131.400 26.330 132.000 ;
        RECT 25.930 131.200 29.930 131.400 ;
        RECT 25.930 130.600 26.330 131.200 ;
        RECT 25.930 130.400 29.930 130.600 ;
        RECT 25.930 130.200 26.330 130.400 ;
        RECT 30.680 130.200 30.880 137.800 ;
        RECT 31.480 130.200 31.680 137.800 ;
        RECT 32.280 130.200 32.480 137.800 ;
        RECT 33.080 130.200 33.280 137.800 ;
        RECT 33.880 130.200 34.080 137.800 ;
        RECT 25.930 129.800 34.080 130.200 ;
        RECT 25.930 129.600 26.330 129.800 ;
        RECT 25.930 129.400 29.930 129.600 ;
        RECT 25.930 128.800 26.330 129.400 ;
        RECT 25.930 128.600 29.930 128.800 ;
        RECT 25.930 128.000 26.330 128.600 ;
        RECT 25.930 127.800 29.930 128.000 ;
        RECT 25.930 127.200 26.330 127.800 ;
        RECT 25.930 127.000 29.930 127.200 ;
        RECT 25.930 126.400 26.330 127.000 ;
        RECT 25.930 126.200 29.930 126.400 ;
        RECT 25.930 125.600 26.330 126.200 ;
        RECT 25.930 125.400 29.930 125.600 ;
        RECT 25.930 124.800 26.330 125.400 ;
        RECT 25.930 124.600 29.930 124.800 ;
        RECT 25.930 124.000 26.330 124.600 ;
        RECT 25.930 123.800 29.930 124.000 ;
        RECT 25.930 123.200 26.330 123.800 ;
        RECT 25.930 123.000 29.930 123.200 ;
        RECT 25.930 122.400 26.330 123.000 ;
        RECT 25.930 122.200 29.930 122.400 ;
        RECT 30.680 122.200 30.880 129.800 ;
        RECT 31.480 122.200 31.680 129.800 ;
        RECT 32.280 122.200 32.480 129.800 ;
        RECT 33.080 122.200 33.280 129.800 ;
        RECT 33.880 122.200 34.080 129.800 ;
        RECT 35.380 130.200 35.580 137.800 ;
        RECT 36.180 130.200 36.380 137.800 ;
        RECT 36.980 130.200 37.180 137.800 ;
        RECT 37.780 130.200 37.980 137.800 ;
        RECT 38.580 130.200 38.780 137.800 ;
        RECT 39.530 137.600 43.530 137.800 ;
        RECT 43.130 137.000 43.530 137.600 ;
        RECT 39.530 136.800 43.530 137.000 ;
        RECT 43.130 136.200 43.530 136.800 ;
        RECT 39.530 136.000 43.530 136.200 ;
        RECT 43.130 135.400 43.530 136.000 ;
        RECT 39.530 135.200 43.530 135.400 ;
        RECT 43.130 134.600 43.530 135.200 ;
        RECT 39.530 134.400 43.530 134.600 ;
        RECT 43.130 133.800 43.530 134.400 ;
        RECT 39.530 133.600 43.530 133.800 ;
        RECT 43.130 133.000 43.530 133.600 ;
        RECT 39.530 132.800 43.530 133.000 ;
        RECT 43.130 132.200 43.530 132.800 ;
        RECT 39.530 132.000 43.530 132.200 ;
        RECT 43.130 131.400 43.530 132.000 ;
        RECT 39.530 131.200 43.530 131.400 ;
        RECT 43.130 130.600 43.530 131.200 ;
        RECT 39.530 130.400 43.530 130.600 ;
        RECT 43.130 130.200 43.530 130.400 ;
        RECT 35.380 129.800 43.530 130.200 ;
        RECT 35.380 122.200 35.580 129.800 ;
        RECT 36.180 122.200 36.380 129.800 ;
        RECT 36.980 122.200 37.180 129.800 ;
        RECT 37.780 122.200 37.980 129.800 ;
        RECT 38.580 122.200 38.780 129.800 ;
        RECT 43.130 129.600 43.530 129.800 ;
        RECT 39.530 129.400 43.530 129.600 ;
        RECT 43.130 128.800 43.530 129.400 ;
        RECT 39.530 128.600 43.530 128.800 ;
        RECT 43.130 128.000 43.530 128.600 ;
        RECT 39.530 127.800 43.530 128.000 ;
        RECT 43.130 127.200 43.530 127.800 ;
        RECT 39.530 127.000 43.530 127.200 ;
        RECT 43.130 126.400 43.530 127.000 ;
        RECT 39.530 126.200 43.530 126.400 ;
        RECT 43.130 125.600 43.530 126.200 ;
        RECT 39.530 125.400 43.530 125.600 ;
        RECT 43.130 124.800 43.530 125.400 ;
        RECT 39.530 124.600 43.530 124.800 ;
        RECT 43.130 124.000 43.530 124.600 ;
        RECT 39.530 123.800 43.530 124.000 ;
        RECT 43.130 123.200 43.530 123.800 ;
        RECT 39.530 123.000 43.530 123.200 ;
        RECT 43.130 122.400 43.530 123.000 ;
        RECT 39.530 122.200 43.530 122.400 ;
        RECT 45.930 137.600 49.930 137.800 ;
        RECT 45.930 137.000 46.330 137.600 ;
        RECT 45.930 136.800 49.930 137.000 ;
        RECT 45.930 136.200 46.330 136.800 ;
        RECT 45.930 136.000 49.930 136.200 ;
        RECT 45.930 135.400 46.330 136.000 ;
        RECT 45.930 135.200 49.930 135.400 ;
        RECT 45.930 134.600 46.330 135.200 ;
        RECT 45.930 134.400 49.930 134.600 ;
        RECT 45.930 133.800 46.330 134.400 ;
        RECT 45.930 133.600 49.930 133.800 ;
        RECT 45.930 133.000 46.330 133.600 ;
        RECT 45.930 132.800 49.930 133.000 ;
        RECT 45.930 132.200 46.330 132.800 ;
        RECT 45.930 132.000 49.930 132.200 ;
        RECT 45.930 131.400 46.330 132.000 ;
        RECT 45.930 131.200 49.930 131.400 ;
        RECT 45.930 130.600 46.330 131.200 ;
        RECT 45.930 130.400 49.930 130.600 ;
        RECT 45.930 130.200 46.330 130.400 ;
        RECT 50.680 130.200 50.880 137.800 ;
        RECT 51.480 130.200 51.680 137.800 ;
        RECT 52.280 130.200 52.480 137.800 ;
        RECT 53.080 130.200 53.280 137.800 ;
        RECT 53.880 130.200 54.080 137.800 ;
        RECT 45.930 129.800 54.080 130.200 ;
        RECT 45.930 129.600 46.330 129.800 ;
        RECT 45.930 129.400 49.930 129.600 ;
        RECT 45.930 128.800 46.330 129.400 ;
        RECT 45.930 128.600 49.930 128.800 ;
        RECT 45.930 128.000 46.330 128.600 ;
        RECT 45.930 127.800 49.930 128.000 ;
        RECT 45.930 127.200 46.330 127.800 ;
        RECT 45.930 127.000 49.930 127.200 ;
        RECT 45.930 126.400 46.330 127.000 ;
        RECT 45.930 126.200 49.930 126.400 ;
        RECT 45.930 125.600 46.330 126.200 ;
        RECT 45.930 125.400 49.930 125.600 ;
        RECT 45.930 124.800 46.330 125.400 ;
        RECT 45.930 124.600 49.930 124.800 ;
        RECT 45.930 124.000 46.330 124.600 ;
        RECT 45.930 123.800 49.930 124.000 ;
        RECT 45.930 123.200 46.330 123.800 ;
        RECT 45.930 123.000 49.930 123.200 ;
        RECT 45.930 122.400 46.330 123.000 ;
        RECT 45.930 122.200 49.930 122.400 ;
        RECT 50.680 122.200 50.880 129.800 ;
        RECT 51.480 122.200 51.680 129.800 ;
        RECT 52.280 122.200 52.480 129.800 ;
        RECT 53.080 122.200 53.280 129.800 ;
        RECT 53.880 122.200 54.080 129.800 ;
        RECT 55.380 130.200 55.580 137.800 ;
        RECT 56.180 130.200 56.380 137.800 ;
        RECT 56.980 130.200 57.180 137.800 ;
        RECT 57.780 130.200 57.980 137.800 ;
        RECT 58.580 130.200 58.780 137.800 ;
        RECT 59.530 137.600 63.530 137.800 ;
        RECT 63.130 137.000 63.530 137.600 ;
        RECT 59.530 136.800 63.530 137.000 ;
        RECT 63.130 136.200 63.530 136.800 ;
        RECT 59.530 136.000 63.530 136.200 ;
        RECT 63.130 135.400 63.530 136.000 ;
        RECT 59.530 135.200 63.530 135.400 ;
        RECT 63.130 134.600 63.530 135.200 ;
        RECT 59.530 134.400 63.530 134.600 ;
        RECT 63.130 133.800 63.530 134.400 ;
        RECT 59.530 133.600 63.530 133.800 ;
        RECT 63.130 133.000 63.530 133.600 ;
        RECT 59.530 132.800 63.530 133.000 ;
        RECT 63.130 132.200 63.530 132.800 ;
        RECT 59.530 132.000 63.530 132.200 ;
        RECT 63.130 131.400 63.530 132.000 ;
        RECT 59.530 131.200 63.530 131.400 ;
        RECT 63.130 130.600 63.530 131.200 ;
        RECT 59.530 130.400 63.530 130.600 ;
        RECT 63.130 130.200 63.530 130.400 ;
        RECT 55.380 129.800 63.530 130.200 ;
        RECT 55.380 122.200 55.580 129.800 ;
        RECT 56.180 122.200 56.380 129.800 ;
        RECT 56.980 122.200 57.180 129.800 ;
        RECT 57.780 122.200 57.980 129.800 ;
        RECT 58.580 122.200 58.780 129.800 ;
        RECT 63.130 129.600 63.530 129.800 ;
        RECT 59.530 129.400 63.530 129.600 ;
        RECT 63.130 128.800 63.530 129.400 ;
        RECT 59.530 128.600 63.530 128.800 ;
        RECT 63.130 128.000 63.530 128.600 ;
        RECT 59.530 127.800 63.530 128.000 ;
        RECT 63.130 127.200 63.530 127.800 ;
        RECT 59.530 127.000 63.530 127.200 ;
        RECT 63.130 126.400 63.530 127.000 ;
        RECT 59.530 126.200 63.530 126.400 ;
        RECT 63.130 125.600 63.530 126.200 ;
        RECT 59.530 125.400 63.530 125.600 ;
        RECT 63.130 124.800 63.530 125.400 ;
        RECT 59.530 124.600 63.530 124.800 ;
        RECT 63.130 124.000 63.530 124.600 ;
        RECT 59.530 123.800 63.530 124.000 ;
        RECT 63.130 123.200 63.530 123.800 ;
        RECT 59.530 123.000 63.530 123.200 ;
        RECT 63.130 122.400 63.530 123.000 ;
        RECT 59.530 122.200 63.530 122.400 ;
        RECT 65.930 137.600 69.930 137.800 ;
        RECT 65.930 137.000 66.330 137.600 ;
        RECT 65.930 136.800 69.930 137.000 ;
        RECT 65.930 136.200 66.330 136.800 ;
        RECT 65.930 136.000 69.930 136.200 ;
        RECT 65.930 135.400 66.330 136.000 ;
        RECT 65.930 135.200 69.930 135.400 ;
        RECT 65.930 134.600 66.330 135.200 ;
        RECT 65.930 134.400 69.930 134.600 ;
        RECT 65.930 133.800 66.330 134.400 ;
        RECT 65.930 133.600 69.930 133.800 ;
        RECT 65.930 133.000 66.330 133.600 ;
        RECT 65.930 132.800 69.930 133.000 ;
        RECT 65.930 132.200 66.330 132.800 ;
        RECT 65.930 132.000 69.930 132.200 ;
        RECT 65.930 131.400 66.330 132.000 ;
        RECT 65.930 131.200 69.930 131.400 ;
        RECT 65.930 130.600 66.330 131.200 ;
        RECT 65.930 130.400 69.930 130.600 ;
        RECT 65.930 130.200 66.330 130.400 ;
        RECT 70.680 130.200 70.880 137.800 ;
        RECT 71.480 130.200 71.680 137.800 ;
        RECT 72.280 130.200 72.480 137.800 ;
        RECT 73.080 130.200 73.280 137.800 ;
        RECT 73.880 130.200 74.080 137.800 ;
        RECT 65.930 129.800 74.080 130.200 ;
        RECT 65.930 129.600 66.330 129.800 ;
        RECT 65.930 129.400 69.930 129.600 ;
        RECT 65.930 128.800 66.330 129.400 ;
        RECT 65.930 128.600 69.930 128.800 ;
        RECT 65.930 128.000 66.330 128.600 ;
        RECT 65.930 127.800 69.930 128.000 ;
        RECT 65.930 127.200 66.330 127.800 ;
        RECT 65.930 127.000 69.930 127.200 ;
        RECT 65.930 126.400 66.330 127.000 ;
        RECT 65.930 126.200 69.930 126.400 ;
        RECT 65.930 125.600 66.330 126.200 ;
        RECT 65.930 125.400 69.930 125.600 ;
        RECT 65.930 124.800 66.330 125.400 ;
        RECT 65.930 124.600 69.930 124.800 ;
        RECT 65.930 124.000 66.330 124.600 ;
        RECT 65.930 123.800 69.930 124.000 ;
        RECT 65.930 123.200 66.330 123.800 ;
        RECT 65.930 123.000 69.930 123.200 ;
        RECT 65.930 122.400 66.330 123.000 ;
        RECT 65.930 122.200 69.930 122.400 ;
        RECT 70.680 122.200 70.880 129.800 ;
        RECT 71.480 122.200 71.680 129.800 ;
        RECT 72.280 122.200 72.480 129.800 ;
        RECT 73.080 122.200 73.280 129.800 ;
        RECT 73.880 122.200 74.080 129.800 ;
        RECT 75.380 130.200 75.580 137.800 ;
        RECT 76.180 130.200 76.380 137.800 ;
        RECT 76.980 130.200 77.180 137.800 ;
        RECT 77.780 130.200 77.980 137.800 ;
        RECT 78.580 130.200 78.780 137.800 ;
        RECT 79.530 137.600 83.530 137.800 ;
        RECT 83.130 137.000 83.530 137.600 ;
        RECT 79.530 136.800 83.530 137.000 ;
        RECT 83.130 136.200 83.530 136.800 ;
        RECT 79.530 136.000 83.530 136.200 ;
        RECT 83.130 135.400 83.530 136.000 ;
        RECT 79.530 135.200 83.530 135.400 ;
        RECT 83.130 134.600 83.530 135.200 ;
        RECT 79.530 134.400 83.530 134.600 ;
        RECT 83.130 133.800 83.530 134.400 ;
        RECT 79.530 133.600 83.530 133.800 ;
        RECT 83.130 133.000 83.530 133.600 ;
        RECT 79.530 132.800 83.530 133.000 ;
        RECT 83.130 132.200 83.530 132.800 ;
        RECT 79.530 132.000 83.530 132.200 ;
        RECT 83.130 131.400 83.530 132.000 ;
        RECT 79.530 131.200 83.530 131.400 ;
        RECT 83.130 130.600 83.530 131.200 ;
        RECT 79.530 130.400 83.530 130.600 ;
        RECT 83.130 130.200 83.530 130.400 ;
        RECT 75.380 129.800 83.530 130.200 ;
        RECT 75.380 122.200 75.580 129.800 ;
        RECT 76.180 122.200 76.380 129.800 ;
        RECT 76.980 122.200 77.180 129.800 ;
        RECT 77.780 122.200 77.980 129.800 ;
        RECT 78.580 122.200 78.780 129.800 ;
        RECT 83.130 129.600 83.530 129.800 ;
        RECT 79.530 129.400 83.530 129.600 ;
        RECT 83.130 128.800 83.530 129.400 ;
        RECT 79.530 128.600 83.530 128.800 ;
        RECT 83.130 128.000 83.530 128.600 ;
        RECT 79.530 127.800 83.530 128.000 ;
        RECT 83.130 127.200 83.530 127.800 ;
        RECT 79.530 127.000 83.530 127.200 ;
        RECT 83.130 126.400 83.530 127.000 ;
        RECT 79.530 126.200 83.530 126.400 ;
        RECT 83.130 125.600 83.530 126.200 ;
        RECT 79.530 125.400 83.530 125.600 ;
        RECT 83.130 124.800 83.530 125.400 ;
        RECT 79.530 124.600 83.530 124.800 ;
        RECT 83.130 124.000 83.530 124.600 ;
        RECT 79.530 123.800 83.530 124.000 ;
        RECT 83.130 123.200 83.530 123.800 ;
        RECT 79.530 123.000 83.530 123.200 ;
        RECT 83.130 122.400 83.530 123.000 ;
        RECT 79.530 122.200 83.530 122.400 ;
        RECT 85.930 137.600 89.930 137.800 ;
        RECT 85.930 137.000 86.330 137.600 ;
        RECT 85.930 136.800 89.930 137.000 ;
        RECT 85.930 136.200 86.330 136.800 ;
        RECT 85.930 136.000 89.930 136.200 ;
        RECT 85.930 135.400 86.330 136.000 ;
        RECT 85.930 135.200 89.930 135.400 ;
        RECT 85.930 134.600 86.330 135.200 ;
        RECT 85.930 134.400 89.930 134.600 ;
        RECT 85.930 133.800 86.330 134.400 ;
        RECT 85.930 133.600 89.930 133.800 ;
        RECT 85.930 133.000 86.330 133.600 ;
        RECT 85.930 132.800 89.930 133.000 ;
        RECT 85.930 132.200 86.330 132.800 ;
        RECT 85.930 132.000 89.930 132.200 ;
        RECT 85.930 131.400 86.330 132.000 ;
        RECT 85.930 131.200 89.930 131.400 ;
        RECT 85.930 130.600 86.330 131.200 ;
        RECT 85.930 130.400 89.930 130.600 ;
        RECT 85.930 130.200 86.330 130.400 ;
        RECT 90.680 130.200 90.880 137.800 ;
        RECT 91.480 130.200 91.680 137.800 ;
        RECT 92.280 130.200 92.480 137.800 ;
        RECT 93.080 130.200 93.280 137.800 ;
        RECT 93.880 130.200 94.080 137.800 ;
        RECT 85.930 129.800 94.080 130.200 ;
        RECT 85.930 129.600 86.330 129.800 ;
        RECT 85.930 129.400 89.930 129.600 ;
        RECT 85.930 128.800 86.330 129.400 ;
        RECT 85.930 128.600 89.930 128.800 ;
        RECT 85.930 128.000 86.330 128.600 ;
        RECT 85.930 127.800 89.930 128.000 ;
        RECT 85.930 127.200 86.330 127.800 ;
        RECT 85.930 127.000 89.930 127.200 ;
        RECT 85.930 126.400 86.330 127.000 ;
        RECT 85.930 126.200 89.930 126.400 ;
        RECT 85.930 125.600 86.330 126.200 ;
        RECT 85.930 125.400 89.930 125.600 ;
        RECT 85.930 124.800 86.330 125.400 ;
        RECT 85.930 124.600 89.930 124.800 ;
        RECT 85.930 124.000 86.330 124.600 ;
        RECT 85.930 123.800 89.930 124.000 ;
        RECT 85.930 123.200 86.330 123.800 ;
        RECT 85.930 123.000 89.930 123.200 ;
        RECT 85.930 122.400 86.330 123.000 ;
        RECT 85.930 122.200 89.930 122.400 ;
        RECT 90.680 122.200 90.880 129.800 ;
        RECT 91.480 122.200 91.680 129.800 ;
        RECT 92.280 122.200 92.480 129.800 ;
        RECT 93.080 122.200 93.280 129.800 ;
        RECT 93.880 122.200 94.080 129.800 ;
        RECT 95.380 130.200 95.580 137.800 ;
        RECT 96.180 130.200 96.380 137.800 ;
        RECT 96.980 130.200 97.180 137.800 ;
        RECT 97.780 130.200 97.980 137.800 ;
        RECT 98.580 130.200 98.780 137.800 ;
        RECT 99.530 137.600 103.530 137.800 ;
        RECT 103.130 137.000 103.530 137.600 ;
        RECT 99.530 136.800 103.530 137.000 ;
        RECT 103.130 136.200 103.530 136.800 ;
        RECT 99.530 136.000 103.530 136.200 ;
        RECT 103.130 135.400 103.530 136.000 ;
        RECT 99.530 135.200 103.530 135.400 ;
        RECT 103.130 134.600 103.530 135.200 ;
        RECT 99.530 134.400 103.530 134.600 ;
        RECT 103.130 133.800 103.530 134.400 ;
        RECT 99.530 133.600 103.530 133.800 ;
        RECT 103.130 133.000 103.530 133.600 ;
        RECT 99.530 132.800 103.530 133.000 ;
        RECT 103.130 132.200 103.530 132.800 ;
        RECT 99.530 132.000 103.530 132.200 ;
        RECT 103.130 131.400 103.530 132.000 ;
        RECT 99.530 131.200 103.530 131.400 ;
        RECT 103.130 130.600 103.530 131.200 ;
        RECT 99.530 130.400 103.530 130.600 ;
        RECT 103.130 130.200 103.530 130.400 ;
        RECT 95.380 129.800 103.530 130.200 ;
        RECT 95.380 122.200 95.580 129.800 ;
        RECT 96.180 122.200 96.380 129.800 ;
        RECT 96.980 122.200 97.180 129.800 ;
        RECT 97.780 122.200 97.980 129.800 ;
        RECT 98.580 122.200 98.780 129.800 ;
        RECT 103.130 129.600 103.530 129.800 ;
        RECT 99.530 129.400 103.530 129.600 ;
        RECT 103.130 128.800 103.530 129.400 ;
        RECT 99.530 128.600 103.530 128.800 ;
        RECT 103.130 128.000 103.530 128.600 ;
        RECT 99.530 127.800 103.530 128.000 ;
        RECT 103.130 127.200 103.530 127.800 ;
        RECT 99.530 127.000 103.530 127.200 ;
        RECT 103.130 126.400 103.530 127.000 ;
        RECT 99.530 126.200 103.530 126.400 ;
        RECT 103.130 125.600 103.530 126.200 ;
        RECT 99.530 125.400 103.530 125.600 ;
        RECT 103.130 124.800 103.530 125.400 ;
        RECT 99.530 124.600 103.530 124.800 ;
        RECT 103.130 124.000 103.530 124.600 ;
        RECT 99.530 123.800 103.530 124.000 ;
        RECT 103.130 123.200 103.530 123.800 ;
        RECT 99.530 123.000 103.530 123.200 ;
        RECT 103.130 122.400 103.530 123.000 ;
        RECT 99.530 122.200 103.530 122.400 ;
        RECT 105.930 137.600 109.930 137.800 ;
        RECT 105.930 137.000 106.330 137.600 ;
        RECT 105.930 136.800 109.930 137.000 ;
        RECT 105.930 136.200 106.330 136.800 ;
        RECT 105.930 136.000 109.930 136.200 ;
        RECT 105.930 135.400 106.330 136.000 ;
        RECT 105.930 135.200 109.930 135.400 ;
        RECT 105.930 134.600 106.330 135.200 ;
        RECT 105.930 134.400 109.930 134.600 ;
        RECT 105.930 133.800 106.330 134.400 ;
        RECT 105.930 133.600 109.930 133.800 ;
        RECT 105.930 133.000 106.330 133.600 ;
        RECT 105.930 132.800 109.930 133.000 ;
        RECT 105.930 132.200 106.330 132.800 ;
        RECT 105.930 132.000 109.930 132.200 ;
        RECT 105.930 131.400 106.330 132.000 ;
        RECT 105.930 131.200 109.930 131.400 ;
        RECT 105.930 130.600 106.330 131.200 ;
        RECT 105.930 130.400 109.930 130.600 ;
        RECT 105.930 130.200 106.330 130.400 ;
        RECT 110.680 130.200 110.880 137.800 ;
        RECT 111.480 130.200 111.680 137.800 ;
        RECT 112.280 130.200 112.480 137.800 ;
        RECT 113.080 130.200 113.280 137.800 ;
        RECT 113.880 130.200 114.080 137.800 ;
        RECT 105.930 129.800 114.080 130.200 ;
        RECT 105.930 129.600 106.330 129.800 ;
        RECT 105.930 129.400 109.930 129.600 ;
        RECT 105.930 128.800 106.330 129.400 ;
        RECT 105.930 128.600 109.930 128.800 ;
        RECT 105.930 128.000 106.330 128.600 ;
        RECT 105.930 127.800 109.930 128.000 ;
        RECT 105.930 127.200 106.330 127.800 ;
        RECT 105.930 127.000 109.930 127.200 ;
        RECT 105.930 126.400 106.330 127.000 ;
        RECT 105.930 126.200 109.930 126.400 ;
        RECT 105.930 125.600 106.330 126.200 ;
        RECT 105.930 125.400 109.930 125.600 ;
        RECT 105.930 124.800 106.330 125.400 ;
        RECT 105.930 124.600 109.930 124.800 ;
        RECT 105.930 124.000 106.330 124.600 ;
        RECT 105.930 123.800 109.930 124.000 ;
        RECT 105.930 123.200 106.330 123.800 ;
        RECT 105.930 123.000 109.930 123.200 ;
        RECT 105.930 122.400 106.330 123.000 ;
        RECT 105.930 122.200 109.930 122.400 ;
        RECT 110.680 122.200 110.880 129.800 ;
        RECT 111.480 122.200 111.680 129.800 ;
        RECT 112.280 122.200 112.480 129.800 ;
        RECT 113.080 122.200 113.280 129.800 ;
        RECT 113.880 122.200 114.080 129.800 ;
        RECT 115.380 130.200 115.580 137.800 ;
        RECT 116.180 130.200 116.380 137.800 ;
        RECT 116.980 130.200 117.180 137.800 ;
        RECT 117.780 130.200 117.980 137.800 ;
        RECT 118.580 130.200 118.780 137.800 ;
        RECT 119.530 137.600 123.530 137.800 ;
        RECT 123.130 137.000 123.530 137.600 ;
        RECT 119.530 136.800 123.530 137.000 ;
        RECT 123.130 136.200 123.530 136.800 ;
        RECT 119.530 136.000 123.530 136.200 ;
        RECT 123.130 135.400 123.530 136.000 ;
        RECT 119.530 135.200 123.530 135.400 ;
        RECT 123.130 134.600 123.530 135.200 ;
        RECT 119.530 134.400 123.530 134.600 ;
        RECT 123.130 133.800 123.530 134.400 ;
        RECT 119.530 133.600 123.530 133.800 ;
        RECT 123.130 133.000 123.530 133.600 ;
        RECT 119.530 132.800 123.530 133.000 ;
        RECT 123.130 132.200 123.530 132.800 ;
        RECT 119.530 132.000 123.530 132.200 ;
        RECT 123.130 131.400 123.530 132.000 ;
        RECT 119.530 131.200 123.530 131.400 ;
        RECT 123.130 130.600 123.530 131.200 ;
        RECT 119.530 130.400 123.530 130.600 ;
        RECT 123.130 130.200 123.530 130.400 ;
        RECT 130.050 130.270 130.410 130.650 ;
        RECT 130.680 130.270 131.040 130.650 ;
        RECT 131.280 130.270 131.640 130.650 ;
        RECT 115.380 129.800 123.530 130.200 ;
        RECT 115.380 122.200 115.580 129.800 ;
        RECT 116.180 122.200 116.380 129.800 ;
        RECT 116.980 122.200 117.180 129.800 ;
        RECT 117.780 122.200 117.980 129.800 ;
        RECT 118.580 122.200 118.780 129.800 ;
        RECT 123.130 129.600 123.530 129.800 ;
        RECT 130.050 129.680 130.410 130.060 ;
        RECT 130.680 129.680 131.040 130.060 ;
        RECT 131.280 129.680 131.640 130.060 ;
        RECT 119.530 129.400 123.530 129.600 ;
        RECT 123.130 128.800 123.530 129.400 ;
        RECT 119.530 128.600 123.530 128.800 ;
        RECT 123.130 128.000 123.530 128.600 ;
        RECT 119.530 127.800 123.530 128.000 ;
        RECT 123.130 127.200 123.530 127.800 ;
        RECT 119.530 127.000 123.530 127.200 ;
        RECT 123.130 126.400 123.530 127.000 ;
        RECT 119.530 126.200 123.530 126.400 ;
        RECT 123.130 125.600 123.530 126.200 ;
        RECT 119.530 125.400 123.530 125.600 ;
        RECT 123.130 124.800 123.530 125.400 ;
        RECT 119.530 124.600 123.530 124.800 ;
        RECT 123.130 124.000 123.530 124.600 ;
        RECT 119.530 123.800 123.530 124.000 ;
        RECT 123.130 123.200 123.530 123.800 ;
        RECT 119.530 123.000 123.530 123.200 ;
        RECT 123.130 122.400 123.530 123.000 ;
        RECT 119.530 122.200 123.530 122.400 ;
        RECT 5.930 117.600 9.930 117.800 ;
        RECT 5.930 117.000 6.330 117.600 ;
        RECT 5.930 116.800 9.930 117.000 ;
        RECT 5.930 116.200 6.330 116.800 ;
        RECT 5.930 116.000 9.930 116.200 ;
        RECT 5.930 115.400 6.330 116.000 ;
        RECT 5.930 115.200 9.930 115.400 ;
        RECT 5.930 114.600 6.330 115.200 ;
        RECT 5.930 114.400 9.930 114.600 ;
        RECT 5.930 113.800 6.330 114.400 ;
        RECT 5.930 113.600 9.930 113.800 ;
        RECT 5.930 113.000 6.330 113.600 ;
        RECT 5.930 112.800 9.930 113.000 ;
        RECT 5.930 112.200 6.330 112.800 ;
        RECT 5.930 112.000 9.930 112.200 ;
        RECT 5.930 111.400 6.330 112.000 ;
        RECT 5.930 111.200 9.930 111.400 ;
        RECT 5.930 110.600 6.330 111.200 ;
        RECT 5.930 110.400 9.930 110.600 ;
        RECT 5.930 110.200 6.330 110.400 ;
        RECT 10.680 110.200 10.880 117.800 ;
        RECT 11.480 110.200 11.680 117.800 ;
        RECT 12.280 110.200 12.480 117.800 ;
        RECT 13.080 110.200 13.280 117.800 ;
        RECT 13.880 110.200 14.080 117.800 ;
        RECT 5.930 109.800 14.080 110.200 ;
        RECT 5.930 109.600 6.330 109.800 ;
        RECT 5.930 109.400 9.930 109.600 ;
        RECT 5.930 108.800 6.330 109.400 ;
        RECT 5.930 108.600 9.930 108.800 ;
        RECT 5.930 108.000 6.330 108.600 ;
        RECT 5.930 107.800 9.930 108.000 ;
        RECT 5.930 107.200 6.330 107.800 ;
        RECT 5.930 107.000 9.930 107.200 ;
        RECT 5.930 106.400 6.330 107.000 ;
        RECT 5.930 106.200 9.930 106.400 ;
        RECT 5.930 105.600 6.330 106.200 ;
        RECT 5.930 105.400 9.930 105.600 ;
        RECT 5.930 104.800 6.330 105.400 ;
        RECT 5.930 104.600 9.930 104.800 ;
        RECT 5.930 104.000 6.330 104.600 ;
        RECT 5.930 103.800 9.930 104.000 ;
        RECT 5.930 103.200 6.330 103.800 ;
        RECT 5.930 103.000 9.930 103.200 ;
        RECT 5.930 102.400 6.330 103.000 ;
        RECT 5.930 102.200 9.930 102.400 ;
        RECT 10.680 102.200 10.880 109.800 ;
        RECT 11.480 102.200 11.680 109.800 ;
        RECT 12.280 102.200 12.480 109.800 ;
        RECT 13.080 102.200 13.280 109.800 ;
        RECT 13.880 102.200 14.080 109.800 ;
        RECT 15.380 110.200 15.580 117.800 ;
        RECT 16.180 110.200 16.380 117.800 ;
        RECT 16.980 110.200 17.180 117.800 ;
        RECT 17.780 110.200 17.980 117.800 ;
        RECT 18.580 110.200 18.780 117.800 ;
        RECT 19.530 117.600 23.530 117.800 ;
        RECT 23.130 117.000 23.530 117.600 ;
        RECT 19.530 116.800 23.530 117.000 ;
        RECT 23.130 116.200 23.530 116.800 ;
        RECT 19.530 116.000 23.530 116.200 ;
        RECT 23.130 115.400 23.530 116.000 ;
        RECT 19.530 115.200 23.530 115.400 ;
        RECT 23.130 114.600 23.530 115.200 ;
        RECT 19.530 114.400 23.530 114.600 ;
        RECT 23.130 113.800 23.530 114.400 ;
        RECT 19.530 113.600 23.530 113.800 ;
        RECT 23.130 113.000 23.530 113.600 ;
        RECT 19.530 112.800 23.530 113.000 ;
        RECT 23.130 112.200 23.530 112.800 ;
        RECT 19.530 112.000 23.530 112.200 ;
        RECT 23.130 111.400 23.530 112.000 ;
        RECT 19.530 111.200 23.530 111.400 ;
        RECT 23.130 110.600 23.530 111.200 ;
        RECT 19.530 110.400 23.530 110.600 ;
        RECT 23.130 110.200 23.530 110.400 ;
        RECT 15.380 109.800 23.530 110.200 ;
        RECT 15.380 102.200 15.580 109.800 ;
        RECT 16.180 102.200 16.380 109.800 ;
        RECT 16.980 102.200 17.180 109.800 ;
        RECT 17.780 102.200 17.980 109.800 ;
        RECT 18.580 102.200 18.780 109.800 ;
        RECT 23.130 109.600 23.530 109.800 ;
        RECT 19.530 109.400 23.530 109.600 ;
        RECT 23.130 108.800 23.530 109.400 ;
        RECT 19.530 108.600 23.530 108.800 ;
        RECT 23.130 108.000 23.530 108.600 ;
        RECT 19.530 107.800 23.530 108.000 ;
        RECT 23.130 107.200 23.530 107.800 ;
        RECT 19.530 107.000 23.530 107.200 ;
        RECT 23.130 106.400 23.530 107.000 ;
        RECT 19.530 106.200 23.530 106.400 ;
        RECT 23.130 105.600 23.530 106.200 ;
        RECT 19.530 105.400 23.530 105.600 ;
        RECT 23.130 104.800 23.530 105.400 ;
        RECT 19.530 104.600 23.530 104.800 ;
        RECT 23.130 104.000 23.530 104.600 ;
        RECT 19.530 103.800 23.530 104.000 ;
        RECT 23.130 103.200 23.530 103.800 ;
        RECT 19.530 103.000 23.530 103.200 ;
        RECT 23.130 102.400 23.530 103.000 ;
        RECT 19.530 102.200 23.530 102.400 ;
        RECT 25.930 117.600 29.930 117.800 ;
        RECT 25.930 117.000 26.330 117.600 ;
        RECT 25.930 116.800 29.930 117.000 ;
        RECT 25.930 116.200 26.330 116.800 ;
        RECT 25.930 116.000 29.930 116.200 ;
        RECT 25.930 115.400 26.330 116.000 ;
        RECT 25.930 115.200 29.930 115.400 ;
        RECT 25.930 114.600 26.330 115.200 ;
        RECT 25.930 114.400 29.930 114.600 ;
        RECT 25.930 113.800 26.330 114.400 ;
        RECT 25.930 113.600 29.930 113.800 ;
        RECT 25.930 113.000 26.330 113.600 ;
        RECT 25.930 112.800 29.930 113.000 ;
        RECT 25.930 112.200 26.330 112.800 ;
        RECT 25.930 112.000 29.930 112.200 ;
        RECT 25.930 111.400 26.330 112.000 ;
        RECT 25.930 111.200 29.930 111.400 ;
        RECT 25.930 110.600 26.330 111.200 ;
        RECT 25.930 110.400 29.930 110.600 ;
        RECT 25.930 110.200 26.330 110.400 ;
        RECT 30.680 110.200 30.880 117.800 ;
        RECT 31.480 110.200 31.680 117.800 ;
        RECT 32.280 110.200 32.480 117.800 ;
        RECT 33.080 110.200 33.280 117.800 ;
        RECT 33.880 110.200 34.080 117.800 ;
        RECT 25.930 109.800 34.080 110.200 ;
        RECT 25.930 109.600 26.330 109.800 ;
        RECT 25.930 109.400 29.930 109.600 ;
        RECT 25.930 108.800 26.330 109.400 ;
        RECT 25.930 108.600 29.930 108.800 ;
        RECT 25.930 108.000 26.330 108.600 ;
        RECT 25.930 107.800 29.930 108.000 ;
        RECT 25.930 107.200 26.330 107.800 ;
        RECT 25.930 107.000 29.930 107.200 ;
        RECT 25.930 106.400 26.330 107.000 ;
        RECT 25.930 106.200 29.930 106.400 ;
        RECT 25.930 105.600 26.330 106.200 ;
        RECT 25.930 105.400 29.930 105.600 ;
        RECT 25.930 104.800 26.330 105.400 ;
        RECT 25.930 104.600 29.930 104.800 ;
        RECT 25.930 104.000 26.330 104.600 ;
        RECT 25.930 103.800 29.930 104.000 ;
        RECT 25.930 103.200 26.330 103.800 ;
        RECT 25.930 103.000 29.930 103.200 ;
        RECT 25.930 102.400 26.330 103.000 ;
        RECT 25.930 102.200 29.930 102.400 ;
        RECT 30.680 102.200 30.880 109.800 ;
        RECT 31.480 102.200 31.680 109.800 ;
        RECT 32.280 102.200 32.480 109.800 ;
        RECT 33.080 102.200 33.280 109.800 ;
        RECT 33.880 102.200 34.080 109.800 ;
        RECT 35.380 110.200 35.580 117.800 ;
        RECT 36.180 110.200 36.380 117.800 ;
        RECT 36.980 110.200 37.180 117.800 ;
        RECT 37.780 110.200 37.980 117.800 ;
        RECT 38.580 110.200 38.780 117.800 ;
        RECT 39.530 117.600 43.530 117.800 ;
        RECT 43.130 117.000 43.530 117.600 ;
        RECT 39.530 116.800 43.530 117.000 ;
        RECT 43.130 116.200 43.530 116.800 ;
        RECT 39.530 116.000 43.530 116.200 ;
        RECT 43.130 115.400 43.530 116.000 ;
        RECT 39.530 115.200 43.530 115.400 ;
        RECT 43.130 114.600 43.530 115.200 ;
        RECT 39.530 114.400 43.530 114.600 ;
        RECT 43.130 113.800 43.530 114.400 ;
        RECT 39.530 113.600 43.530 113.800 ;
        RECT 43.130 113.000 43.530 113.600 ;
        RECT 39.530 112.800 43.530 113.000 ;
        RECT 43.130 112.200 43.530 112.800 ;
        RECT 39.530 112.000 43.530 112.200 ;
        RECT 43.130 111.400 43.530 112.000 ;
        RECT 39.530 111.200 43.530 111.400 ;
        RECT 43.130 110.600 43.530 111.200 ;
        RECT 39.530 110.400 43.530 110.600 ;
        RECT 43.130 110.200 43.530 110.400 ;
        RECT 35.380 109.800 43.530 110.200 ;
        RECT 35.380 102.200 35.580 109.800 ;
        RECT 36.180 102.200 36.380 109.800 ;
        RECT 36.980 102.200 37.180 109.800 ;
        RECT 37.780 102.200 37.980 109.800 ;
        RECT 38.580 102.200 38.780 109.800 ;
        RECT 43.130 109.600 43.530 109.800 ;
        RECT 39.530 109.400 43.530 109.600 ;
        RECT 43.130 108.800 43.530 109.400 ;
        RECT 39.530 108.600 43.530 108.800 ;
        RECT 43.130 108.000 43.530 108.600 ;
        RECT 39.530 107.800 43.530 108.000 ;
        RECT 43.130 107.200 43.530 107.800 ;
        RECT 39.530 107.000 43.530 107.200 ;
        RECT 43.130 106.400 43.530 107.000 ;
        RECT 39.530 106.200 43.530 106.400 ;
        RECT 43.130 105.600 43.530 106.200 ;
        RECT 39.530 105.400 43.530 105.600 ;
        RECT 43.130 104.800 43.530 105.400 ;
        RECT 39.530 104.600 43.530 104.800 ;
        RECT 43.130 104.000 43.530 104.600 ;
        RECT 39.530 103.800 43.530 104.000 ;
        RECT 43.130 103.200 43.530 103.800 ;
        RECT 39.530 103.000 43.530 103.200 ;
        RECT 43.130 102.400 43.530 103.000 ;
        RECT 39.530 102.200 43.530 102.400 ;
        RECT 45.930 117.600 49.930 117.800 ;
        RECT 45.930 117.000 46.330 117.600 ;
        RECT 45.930 116.800 49.930 117.000 ;
        RECT 45.930 116.200 46.330 116.800 ;
        RECT 45.930 116.000 49.930 116.200 ;
        RECT 45.930 115.400 46.330 116.000 ;
        RECT 45.930 115.200 49.930 115.400 ;
        RECT 45.930 114.600 46.330 115.200 ;
        RECT 45.930 114.400 49.930 114.600 ;
        RECT 45.930 113.800 46.330 114.400 ;
        RECT 45.930 113.600 49.930 113.800 ;
        RECT 45.930 113.000 46.330 113.600 ;
        RECT 45.930 112.800 49.930 113.000 ;
        RECT 45.930 112.200 46.330 112.800 ;
        RECT 45.930 112.000 49.930 112.200 ;
        RECT 45.930 111.400 46.330 112.000 ;
        RECT 45.930 111.200 49.930 111.400 ;
        RECT 45.930 110.600 46.330 111.200 ;
        RECT 45.930 110.400 49.930 110.600 ;
        RECT 45.930 110.200 46.330 110.400 ;
        RECT 50.680 110.200 50.880 117.800 ;
        RECT 51.480 110.200 51.680 117.800 ;
        RECT 52.280 110.200 52.480 117.800 ;
        RECT 53.080 110.200 53.280 117.800 ;
        RECT 53.880 110.200 54.080 117.800 ;
        RECT 45.930 109.800 54.080 110.200 ;
        RECT 45.930 109.600 46.330 109.800 ;
        RECT 45.930 109.400 49.930 109.600 ;
        RECT 45.930 108.800 46.330 109.400 ;
        RECT 45.930 108.600 49.930 108.800 ;
        RECT 45.930 108.000 46.330 108.600 ;
        RECT 45.930 107.800 49.930 108.000 ;
        RECT 45.930 107.200 46.330 107.800 ;
        RECT 45.930 107.000 49.930 107.200 ;
        RECT 45.930 106.400 46.330 107.000 ;
        RECT 45.930 106.200 49.930 106.400 ;
        RECT 45.930 105.600 46.330 106.200 ;
        RECT 45.930 105.400 49.930 105.600 ;
        RECT 45.930 104.800 46.330 105.400 ;
        RECT 45.930 104.600 49.930 104.800 ;
        RECT 45.930 104.000 46.330 104.600 ;
        RECT 45.930 103.800 49.930 104.000 ;
        RECT 45.930 103.200 46.330 103.800 ;
        RECT 45.930 103.000 49.930 103.200 ;
        RECT 45.930 102.400 46.330 103.000 ;
        RECT 45.930 102.200 49.930 102.400 ;
        RECT 50.680 102.200 50.880 109.800 ;
        RECT 51.480 102.200 51.680 109.800 ;
        RECT 52.280 102.200 52.480 109.800 ;
        RECT 53.080 102.200 53.280 109.800 ;
        RECT 53.880 102.200 54.080 109.800 ;
        RECT 55.380 110.200 55.580 117.800 ;
        RECT 56.180 110.200 56.380 117.800 ;
        RECT 56.980 110.200 57.180 117.800 ;
        RECT 57.780 110.200 57.980 117.800 ;
        RECT 58.580 110.200 58.780 117.800 ;
        RECT 59.530 117.600 63.530 117.800 ;
        RECT 63.130 117.000 63.530 117.600 ;
        RECT 59.530 116.800 63.530 117.000 ;
        RECT 63.130 116.200 63.530 116.800 ;
        RECT 59.530 116.000 63.530 116.200 ;
        RECT 63.130 115.400 63.530 116.000 ;
        RECT 59.530 115.200 63.530 115.400 ;
        RECT 63.130 114.600 63.530 115.200 ;
        RECT 59.530 114.400 63.530 114.600 ;
        RECT 63.130 113.800 63.530 114.400 ;
        RECT 59.530 113.600 63.530 113.800 ;
        RECT 63.130 113.000 63.530 113.600 ;
        RECT 59.530 112.800 63.530 113.000 ;
        RECT 63.130 112.200 63.530 112.800 ;
        RECT 59.530 112.000 63.530 112.200 ;
        RECT 63.130 111.400 63.530 112.000 ;
        RECT 59.530 111.200 63.530 111.400 ;
        RECT 63.130 110.600 63.530 111.200 ;
        RECT 59.530 110.400 63.530 110.600 ;
        RECT 63.130 110.200 63.530 110.400 ;
        RECT 55.380 109.800 63.530 110.200 ;
        RECT 55.380 102.200 55.580 109.800 ;
        RECT 56.180 102.200 56.380 109.800 ;
        RECT 56.980 102.200 57.180 109.800 ;
        RECT 57.780 102.200 57.980 109.800 ;
        RECT 58.580 102.200 58.780 109.800 ;
        RECT 63.130 109.600 63.530 109.800 ;
        RECT 59.530 109.400 63.530 109.600 ;
        RECT 63.130 108.800 63.530 109.400 ;
        RECT 59.530 108.600 63.530 108.800 ;
        RECT 63.130 108.000 63.530 108.600 ;
        RECT 59.530 107.800 63.530 108.000 ;
        RECT 63.130 107.200 63.530 107.800 ;
        RECT 59.530 107.000 63.530 107.200 ;
        RECT 63.130 106.400 63.530 107.000 ;
        RECT 59.530 106.200 63.530 106.400 ;
        RECT 63.130 105.600 63.530 106.200 ;
        RECT 59.530 105.400 63.530 105.600 ;
        RECT 63.130 104.800 63.530 105.400 ;
        RECT 59.530 104.600 63.530 104.800 ;
        RECT 63.130 104.000 63.530 104.600 ;
        RECT 59.530 103.800 63.530 104.000 ;
        RECT 63.130 103.200 63.530 103.800 ;
        RECT 59.530 103.000 63.530 103.200 ;
        RECT 63.130 102.400 63.530 103.000 ;
        RECT 59.530 102.200 63.530 102.400 ;
        RECT 65.930 117.600 69.930 117.800 ;
        RECT 65.930 117.000 66.330 117.600 ;
        RECT 65.930 116.800 69.930 117.000 ;
        RECT 65.930 116.200 66.330 116.800 ;
        RECT 65.930 116.000 69.930 116.200 ;
        RECT 65.930 115.400 66.330 116.000 ;
        RECT 65.930 115.200 69.930 115.400 ;
        RECT 65.930 114.600 66.330 115.200 ;
        RECT 65.930 114.400 69.930 114.600 ;
        RECT 65.930 113.800 66.330 114.400 ;
        RECT 65.930 113.600 69.930 113.800 ;
        RECT 65.930 113.000 66.330 113.600 ;
        RECT 65.930 112.800 69.930 113.000 ;
        RECT 65.930 112.200 66.330 112.800 ;
        RECT 65.930 112.000 69.930 112.200 ;
        RECT 65.930 111.400 66.330 112.000 ;
        RECT 65.930 111.200 69.930 111.400 ;
        RECT 65.930 110.600 66.330 111.200 ;
        RECT 65.930 110.400 69.930 110.600 ;
        RECT 65.930 110.200 66.330 110.400 ;
        RECT 70.680 110.200 70.880 117.800 ;
        RECT 71.480 110.200 71.680 117.800 ;
        RECT 72.280 110.200 72.480 117.800 ;
        RECT 73.080 110.200 73.280 117.800 ;
        RECT 73.880 110.200 74.080 117.800 ;
        RECT 65.930 109.800 74.080 110.200 ;
        RECT 65.930 109.600 66.330 109.800 ;
        RECT 65.930 109.400 69.930 109.600 ;
        RECT 65.930 108.800 66.330 109.400 ;
        RECT 65.930 108.600 69.930 108.800 ;
        RECT 65.930 108.000 66.330 108.600 ;
        RECT 65.930 107.800 69.930 108.000 ;
        RECT 65.930 107.200 66.330 107.800 ;
        RECT 65.930 107.000 69.930 107.200 ;
        RECT 65.930 106.400 66.330 107.000 ;
        RECT 65.930 106.200 69.930 106.400 ;
        RECT 65.930 105.600 66.330 106.200 ;
        RECT 65.930 105.400 69.930 105.600 ;
        RECT 65.930 104.800 66.330 105.400 ;
        RECT 65.930 104.600 69.930 104.800 ;
        RECT 65.930 104.000 66.330 104.600 ;
        RECT 65.930 103.800 69.930 104.000 ;
        RECT 65.930 103.200 66.330 103.800 ;
        RECT 65.930 103.000 69.930 103.200 ;
        RECT 65.930 102.400 66.330 103.000 ;
        RECT 65.930 102.200 69.930 102.400 ;
        RECT 70.680 102.200 70.880 109.800 ;
        RECT 71.480 102.200 71.680 109.800 ;
        RECT 72.280 102.200 72.480 109.800 ;
        RECT 73.080 102.200 73.280 109.800 ;
        RECT 73.880 102.200 74.080 109.800 ;
        RECT 75.380 110.200 75.580 117.800 ;
        RECT 76.180 110.200 76.380 117.800 ;
        RECT 76.980 110.200 77.180 117.800 ;
        RECT 77.780 110.200 77.980 117.800 ;
        RECT 78.580 110.200 78.780 117.800 ;
        RECT 79.530 117.600 83.530 117.800 ;
        RECT 83.130 117.000 83.530 117.600 ;
        RECT 79.530 116.800 83.530 117.000 ;
        RECT 83.130 116.200 83.530 116.800 ;
        RECT 79.530 116.000 83.530 116.200 ;
        RECT 83.130 115.400 83.530 116.000 ;
        RECT 79.530 115.200 83.530 115.400 ;
        RECT 83.130 114.600 83.530 115.200 ;
        RECT 79.530 114.400 83.530 114.600 ;
        RECT 83.130 113.800 83.530 114.400 ;
        RECT 79.530 113.600 83.530 113.800 ;
        RECT 83.130 113.000 83.530 113.600 ;
        RECT 79.530 112.800 83.530 113.000 ;
        RECT 83.130 112.200 83.530 112.800 ;
        RECT 79.530 112.000 83.530 112.200 ;
        RECT 83.130 111.400 83.530 112.000 ;
        RECT 79.530 111.200 83.530 111.400 ;
        RECT 83.130 110.600 83.530 111.200 ;
        RECT 79.530 110.400 83.530 110.600 ;
        RECT 83.130 110.200 83.530 110.400 ;
        RECT 75.380 109.800 83.530 110.200 ;
        RECT 75.380 102.200 75.580 109.800 ;
        RECT 76.180 102.200 76.380 109.800 ;
        RECT 76.980 102.200 77.180 109.800 ;
        RECT 77.780 102.200 77.980 109.800 ;
        RECT 78.580 102.200 78.780 109.800 ;
        RECT 83.130 109.600 83.530 109.800 ;
        RECT 79.530 109.400 83.530 109.600 ;
        RECT 83.130 108.800 83.530 109.400 ;
        RECT 79.530 108.600 83.530 108.800 ;
        RECT 83.130 108.000 83.530 108.600 ;
        RECT 79.530 107.800 83.530 108.000 ;
        RECT 83.130 107.200 83.530 107.800 ;
        RECT 79.530 107.000 83.530 107.200 ;
        RECT 83.130 106.400 83.530 107.000 ;
        RECT 79.530 106.200 83.530 106.400 ;
        RECT 83.130 105.600 83.530 106.200 ;
        RECT 79.530 105.400 83.530 105.600 ;
        RECT 83.130 104.800 83.530 105.400 ;
        RECT 79.530 104.600 83.530 104.800 ;
        RECT 83.130 104.000 83.530 104.600 ;
        RECT 79.530 103.800 83.530 104.000 ;
        RECT 83.130 103.200 83.530 103.800 ;
        RECT 79.530 103.000 83.530 103.200 ;
        RECT 83.130 102.400 83.530 103.000 ;
        RECT 79.530 102.200 83.530 102.400 ;
        RECT 85.930 117.600 89.930 117.800 ;
        RECT 85.930 117.000 86.330 117.600 ;
        RECT 85.930 116.800 89.930 117.000 ;
        RECT 85.930 116.200 86.330 116.800 ;
        RECT 85.930 116.000 89.930 116.200 ;
        RECT 85.930 115.400 86.330 116.000 ;
        RECT 85.930 115.200 89.930 115.400 ;
        RECT 85.930 114.600 86.330 115.200 ;
        RECT 85.930 114.400 89.930 114.600 ;
        RECT 85.930 113.800 86.330 114.400 ;
        RECT 85.930 113.600 89.930 113.800 ;
        RECT 85.930 113.000 86.330 113.600 ;
        RECT 85.930 112.800 89.930 113.000 ;
        RECT 85.930 112.200 86.330 112.800 ;
        RECT 85.930 112.000 89.930 112.200 ;
        RECT 85.930 111.400 86.330 112.000 ;
        RECT 85.930 111.200 89.930 111.400 ;
        RECT 85.930 110.600 86.330 111.200 ;
        RECT 85.930 110.400 89.930 110.600 ;
        RECT 85.930 110.200 86.330 110.400 ;
        RECT 90.680 110.200 90.880 117.800 ;
        RECT 91.480 110.200 91.680 117.800 ;
        RECT 92.280 110.200 92.480 117.800 ;
        RECT 93.080 110.200 93.280 117.800 ;
        RECT 93.880 110.200 94.080 117.800 ;
        RECT 85.930 109.800 94.080 110.200 ;
        RECT 85.930 109.600 86.330 109.800 ;
        RECT 85.930 109.400 89.930 109.600 ;
        RECT 85.930 108.800 86.330 109.400 ;
        RECT 85.930 108.600 89.930 108.800 ;
        RECT 85.930 108.000 86.330 108.600 ;
        RECT 85.930 107.800 89.930 108.000 ;
        RECT 85.930 107.200 86.330 107.800 ;
        RECT 85.930 107.000 89.930 107.200 ;
        RECT 85.930 106.400 86.330 107.000 ;
        RECT 85.930 106.200 89.930 106.400 ;
        RECT 85.930 105.600 86.330 106.200 ;
        RECT 85.930 105.400 89.930 105.600 ;
        RECT 85.930 104.800 86.330 105.400 ;
        RECT 85.930 104.600 89.930 104.800 ;
        RECT 85.930 104.000 86.330 104.600 ;
        RECT 85.930 103.800 89.930 104.000 ;
        RECT 85.930 103.200 86.330 103.800 ;
        RECT 85.930 103.000 89.930 103.200 ;
        RECT 85.930 102.400 86.330 103.000 ;
        RECT 85.930 102.200 89.930 102.400 ;
        RECT 90.680 102.200 90.880 109.800 ;
        RECT 91.480 102.200 91.680 109.800 ;
        RECT 92.280 102.200 92.480 109.800 ;
        RECT 93.080 102.200 93.280 109.800 ;
        RECT 93.880 102.200 94.080 109.800 ;
        RECT 95.380 110.200 95.580 117.800 ;
        RECT 96.180 110.200 96.380 117.800 ;
        RECT 96.980 110.200 97.180 117.800 ;
        RECT 97.780 110.200 97.980 117.800 ;
        RECT 98.580 110.200 98.780 117.800 ;
        RECT 99.530 117.600 103.530 117.800 ;
        RECT 103.130 117.000 103.530 117.600 ;
        RECT 99.530 116.800 103.530 117.000 ;
        RECT 103.130 116.200 103.530 116.800 ;
        RECT 99.530 116.000 103.530 116.200 ;
        RECT 103.130 115.400 103.530 116.000 ;
        RECT 99.530 115.200 103.530 115.400 ;
        RECT 103.130 114.600 103.530 115.200 ;
        RECT 99.530 114.400 103.530 114.600 ;
        RECT 103.130 113.800 103.530 114.400 ;
        RECT 99.530 113.600 103.530 113.800 ;
        RECT 103.130 113.000 103.530 113.600 ;
        RECT 99.530 112.800 103.530 113.000 ;
        RECT 103.130 112.200 103.530 112.800 ;
        RECT 99.530 112.000 103.530 112.200 ;
        RECT 103.130 111.400 103.530 112.000 ;
        RECT 99.530 111.200 103.530 111.400 ;
        RECT 103.130 110.600 103.530 111.200 ;
        RECT 99.530 110.400 103.530 110.600 ;
        RECT 103.130 110.200 103.530 110.400 ;
        RECT 95.380 109.800 103.530 110.200 ;
        RECT 95.380 102.200 95.580 109.800 ;
        RECT 96.180 102.200 96.380 109.800 ;
        RECT 96.980 102.200 97.180 109.800 ;
        RECT 97.780 102.200 97.980 109.800 ;
        RECT 98.580 102.200 98.780 109.800 ;
        RECT 103.130 109.600 103.530 109.800 ;
        RECT 99.530 109.400 103.530 109.600 ;
        RECT 103.130 108.800 103.530 109.400 ;
        RECT 99.530 108.600 103.530 108.800 ;
        RECT 103.130 108.000 103.530 108.600 ;
        RECT 99.530 107.800 103.530 108.000 ;
        RECT 103.130 107.200 103.530 107.800 ;
        RECT 99.530 107.000 103.530 107.200 ;
        RECT 103.130 106.400 103.530 107.000 ;
        RECT 99.530 106.200 103.530 106.400 ;
        RECT 103.130 105.600 103.530 106.200 ;
        RECT 99.530 105.400 103.530 105.600 ;
        RECT 103.130 104.800 103.530 105.400 ;
        RECT 99.530 104.600 103.530 104.800 ;
        RECT 103.130 104.000 103.530 104.600 ;
        RECT 99.530 103.800 103.530 104.000 ;
        RECT 103.130 103.200 103.530 103.800 ;
        RECT 99.530 103.000 103.530 103.200 ;
        RECT 103.130 102.400 103.530 103.000 ;
        RECT 99.530 102.200 103.530 102.400 ;
        RECT 105.930 117.600 109.930 117.800 ;
        RECT 105.930 117.000 106.330 117.600 ;
        RECT 105.930 116.800 109.930 117.000 ;
        RECT 105.930 116.200 106.330 116.800 ;
        RECT 105.930 116.000 109.930 116.200 ;
        RECT 105.930 115.400 106.330 116.000 ;
        RECT 105.930 115.200 109.930 115.400 ;
        RECT 105.930 114.600 106.330 115.200 ;
        RECT 105.930 114.400 109.930 114.600 ;
        RECT 105.930 113.800 106.330 114.400 ;
        RECT 105.930 113.600 109.930 113.800 ;
        RECT 105.930 113.000 106.330 113.600 ;
        RECT 105.930 112.800 109.930 113.000 ;
        RECT 105.930 112.200 106.330 112.800 ;
        RECT 105.930 112.000 109.930 112.200 ;
        RECT 105.930 111.400 106.330 112.000 ;
        RECT 105.930 111.200 109.930 111.400 ;
        RECT 105.930 110.600 106.330 111.200 ;
        RECT 105.930 110.400 109.930 110.600 ;
        RECT 105.930 110.200 106.330 110.400 ;
        RECT 110.680 110.200 110.880 117.800 ;
        RECT 111.480 110.200 111.680 117.800 ;
        RECT 112.280 110.200 112.480 117.800 ;
        RECT 113.080 110.200 113.280 117.800 ;
        RECT 113.880 110.200 114.080 117.800 ;
        RECT 105.930 109.800 114.080 110.200 ;
        RECT 105.930 109.600 106.330 109.800 ;
        RECT 105.930 109.400 109.930 109.600 ;
        RECT 105.930 108.800 106.330 109.400 ;
        RECT 105.930 108.600 109.930 108.800 ;
        RECT 105.930 108.000 106.330 108.600 ;
        RECT 105.930 107.800 109.930 108.000 ;
        RECT 105.930 107.200 106.330 107.800 ;
        RECT 105.930 107.000 109.930 107.200 ;
        RECT 105.930 106.400 106.330 107.000 ;
        RECT 105.930 106.200 109.930 106.400 ;
        RECT 105.930 105.600 106.330 106.200 ;
        RECT 105.930 105.400 109.930 105.600 ;
        RECT 105.930 104.800 106.330 105.400 ;
        RECT 105.930 104.600 109.930 104.800 ;
        RECT 105.930 104.000 106.330 104.600 ;
        RECT 105.930 103.800 109.930 104.000 ;
        RECT 105.930 103.200 106.330 103.800 ;
        RECT 105.930 103.000 109.930 103.200 ;
        RECT 105.930 102.400 106.330 103.000 ;
        RECT 105.930 102.200 109.930 102.400 ;
        RECT 110.680 102.200 110.880 109.800 ;
        RECT 111.480 102.200 111.680 109.800 ;
        RECT 112.280 102.200 112.480 109.800 ;
        RECT 113.080 102.200 113.280 109.800 ;
        RECT 113.880 102.200 114.080 109.800 ;
        RECT 115.380 110.200 115.580 117.800 ;
        RECT 116.180 110.200 116.380 117.800 ;
        RECT 116.980 110.200 117.180 117.800 ;
        RECT 117.780 110.200 117.980 117.800 ;
        RECT 118.580 110.200 118.780 117.800 ;
        RECT 119.530 117.600 123.530 117.800 ;
        RECT 123.130 117.000 123.530 117.600 ;
        RECT 119.530 116.800 123.530 117.000 ;
        RECT 123.130 116.200 123.530 116.800 ;
        RECT 119.530 116.000 123.530 116.200 ;
        RECT 123.130 115.400 123.530 116.000 ;
        RECT 119.530 115.200 123.530 115.400 ;
        RECT 123.130 114.600 123.530 115.200 ;
        RECT 119.530 114.400 123.530 114.600 ;
        RECT 123.130 113.800 123.530 114.400 ;
        RECT 119.530 113.600 123.530 113.800 ;
        RECT 123.130 113.000 123.530 113.600 ;
        RECT 119.530 112.800 123.530 113.000 ;
        RECT 123.130 112.200 123.530 112.800 ;
        RECT 119.530 112.000 123.530 112.200 ;
        RECT 123.130 111.400 123.530 112.000 ;
        RECT 119.530 111.200 123.530 111.400 ;
        RECT 123.130 110.600 123.530 111.200 ;
        RECT 119.530 110.400 123.530 110.600 ;
        RECT 123.130 110.200 123.530 110.400 ;
        RECT 115.380 109.800 123.530 110.200 ;
        RECT 115.380 102.200 115.580 109.800 ;
        RECT 116.180 102.200 116.380 109.800 ;
        RECT 116.980 102.200 117.180 109.800 ;
        RECT 117.780 102.200 117.980 109.800 ;
        RECT 118.580 102.200 118.780 109.800 ;
        RECT 123.130 109.600 123.530 109.800 ;
        RECT 119.530 109.400 123.530 109.600 ;
        RECT 130.050 109.475 130.410 109.855 ;
        RECT 130.680 109.475 131.040 109.855 ;
        RECT 131.280 109.475 131.640 109.855 ;
        RECT 123.130 108.800 123.530 109.400 ;
        RECT 130.050 108.885 130.410 109.265 ;
        RECT 130.680 108.885 131.040 109.265 ;
        RECT 131.280 108.885 131.640 109.265 ;
        RECT 119.530 108.600 123.530 108.800 ;
        RECT 123.130 108.000 123.530 108.600 ;
        RECT 119.530 107.800 123.530 108.000 ;
        RECT 123.130 107.200 123.530 107.800 ;
        RECT 119.530 107.000 123.530 107.200 ;
        RECT 123.130 106.400 123.530 107.000 ;
        RECT 119.530 106.200 123.530 106.400 ;
        RECT 123.130 105.600 123.530 106.200 ;
        RECT 119.530 105.400 123.530 105.600 ;
        RECT 123.130 104.800 123.530 105.400 ;
        RECT 119.530 104.600 123.530 104.800 ;
        RECT 123.130 104.000 123.530 104.600 ;
        RECT 119.530 103.800 123.530 104.000 ;
        RECT 123.130 103.200 123.530 103.800 ;
        RECT 119.530 103.000 123.530 103.200 ;
        RECT 123.130 102.400 123.530 103.000 ;
        RECT 119.530 102.200 123.530 102.400 ;
        RECT 5.930 97.600 9.930 97.800 ;
        RECT 5.930 97.000 6.330 97.600 ;
        RECT 5.930 96.800 9.930 97.000 ;
        RECT 5.930 96.200 6.330 96.800 ;
        RECT 5.930 96.000 9.930 96.200 ;
        RECT 5.930 95.400 6.330 96.000 ;
        RECT 5.930 95.200 9.930 95.400 ;
        RECT 5.930 94.600 6.330 95.200 ;
        RECT 5.930 94.400 9.930 94.600 ;
        RECT 5.930 93.800 6.330 94.400 ;
        RECT 5.930 93.600 9.930 93.800 ;
        RECT 5.930 93.000 6.330 93.600 ;
        RECT 5.930 92.800 9.930 93.000 ;
        RECT 5.930 92.200 6.330 92.800 ;
        RECT 5.930 92.000 9.930 92.200 ;
        RECT 5.930 91.400 6.330 92.000 ;
        RECT 5.930 91.200 9.930 91.400 ;
        RECT 5.930 90.600 6.330 91.200 ;
        RECT 5.930 90.400 9.930 90.600 ;
        RECT 5.930 90.200 6.330 90.400 ;
        RECT 10.680 90.200 10.880 97.800 ;
        RECT 11.480 90.200 11.680 97.800 ;
        RECT 12.280 90.200 12.480 97.800 ;
        RECT 13.080 90.200 13.280 97.800 ;
        RECT 13.880 90.200 14.080 97.800 ;
        RECT 5.930 89.800 14.080 90.200 ;
        RECT 5.930 89.600 6.330 89.800 ;
        RECT 5.930 89.400 9.930 89.600 ;
        RECT 5.930 88.800 6.330 89.400 ;
        RECT 5.930 88.600 9.930 88.800 ;
        RECT 5.930 88.000 6.330 88.600 ;
        RECT 5.930 87.800 9.930 88.000 ;
        RECT 5.930 87.200 6.330 87.800 ;
        RECT 5.930 87.000 9.930 87.200 ;
        RECT 5.930 86.400 6.330 87.000 ;
        RECT 5.930 86.200 9.930 86.400 ;
        RECT 5.930 85.600 6.330 86.200 ;
        RECT 5.930 85.400 9.930 85.600 ;
        RECT 5.930 84.800 6.330 85.400 ;
        RECT 5.930 84.600 9.930 84.800 ;
        RECT 5.930 84.000 6.330 84.600 ;
        RECT 5.930 83.800 9.930 84.000 ;
        RECT 5.930 83.200 6.330 83.800 ;
        RECT 5.930 83.000 9.930 83.200 ;
        RECT 5.930 82.400 6.330 83.000 ;
        RECT 5.930 82.200 9.930 82.400 ;
        RECT 10.680 82.200 10.880 89.800 ;
        RECT 11.480 82.200 11.680 89.800 ;
        RECT 12.280 82.200 12.480 89.800 ;
        RECT 13.080 82.200 13.280 89.800 ;
        RECT 13.880 82.200 14.080 89.800 ;
        RECT 15.380 90.200 15.580 97.800 ;
        RECT 16.180 90.200 16.380 97.800 ;
        RECT 16.980 90.200 17.180 97.800 ;
        RECT 17.780 90.200 17.980 97.800 ;
        RECT 18.580 90.200 18.780 97.800 ;
        RECT 19.530 97.600 23.530 97.800 ;
        RECT 23.130 97.000 23.530 97.600 ;
        RECT 19.530 96.800 23.530 97.000 ;
        RECT 23.130 96.200 23.530 96.800 ;
        RECT 19.530 96.000 23.530 96.200 ;
        RECT 23.130 95.400 23.530 96.000 ;
        RECT 19.530 95.200 23.530 95.400 ;
        RECT 23.130 94.600 23.530 95.200 ;
        RECT 19.530 94.400 23.530 94.600 ;
        RECT 23.130 93.800 23.530 94.400 ;
        RECT 19.530 93.600 23.530 93.800 ;
        RECT 23.130 93.000 23.530 93.600 ;
        RECT 19.530 92.800 23.530 93.000 ;
        RECT 23.130 92.200 23.530 92.800 ;
        RECT 19.530 92.000 23.530 92.200 ;
        RECT 23.130 91.400 23.530 92.000 ;
        RECT 19.530 91.200 23.530 91.400 ;
        RECT 23.130 90.600 23.530 91.200 ;
        RECT 19.530 90.400 23.530 90.600 ;
        RECT 23.130 90.200 23.530 90.400 ;
        RECT 15.380 89.800 23.530 90.200 ;
        RECT 15.380 82.200 15.580 89.800 ;
        RECT 16.180 82.200 16.380 89.800 ;
        RECT 16.980 82.200 17.180 89.800 ;
        RECT 17.780 82.200 17.980 89.800 ;
        RECT 18.580 82.200 18.780 89.800 ;
        RECT 23.130 89.600 23.530 89.800 ;
        RECT 19.530 89.400 23.530 89.600 ;
        RECT 23.130 88.800 23.530 89.400 ;
        RECT 19.530 88.600 23.530 88.800 ;
        RECT 23.130 88.000 23.530 88.600 ;
        RECT 19.530 87.800 23.530 88.000 ;
        RECT 23.130 87.200 23.530 87.800 ;
        RECT 19.530 87.000 23.530 87.200 ;
        RECT 23.130 86.400 23.530 87.000 ;
        RECT 19.530 86.200 23.530 86.400 ;
        RECT 23.130 85.600 23.530 86.200 ;
        RECT 19.530 85.400 23.530 85.600 ;
        RECT 23.130 84.800 23.530 85.400 ;
        RECT 19.530 84.600 23.530 84.800 ;
        RECT 23.130 84.000 23.530 84.600 ;
        RECT 19.530 83.800 23.530 84.000 ;
        RECT 23.130 83.200 23.530 83.800 ;
        RECT 19.530 83.000 23.530 83.200 ;
        RECT 23.130 82.400 23.530 83.000 ;
        RECT 19.530 82.200 23.530 82.400 ;
        RECT 25.930 97.600 29.930 97.800 ;
        RECT 25.930 97.000 26.330 97.600 ;
        RECT 25.930 96.800 29.930 97.000 ;
        RECT 25.930 96.200 26.330 96.800 ;
        RECT 25.930 96.000 29.930 96.200 ;
        RECT 25.930 95.400 26.330 96.000 ;
        RECT 25.930 95.200 29.930 95.400 ;
        RECT 25.930 94.600 26.330 95.200 ;
        RECT 25.930 94.400 29.930 94.600 ;
        RECT 25.930 93.800 26.330 94.400 ;
        RECT 25.930 93.600 29.930 93.800 ;
        RECT 25.930 93.000 26.330 93.600 ;
        RECT 25.930 92.800 29.930 93.000 ;
        RECT 25.930 92.200 26.330 92.800 ;
        RECT 25.930 92.000 29.930 92.200 ;
        RECT 25.930 91.400 26.330 92.000 ;
        RECT 25.930 91.200 29.930 91.400 ;
        RECT 25.930 90.600 26.330 91.200 ;
        RECT 25.930 90.400 29.930 90.600 ;
        RECT 25.930 90.200 26.330 90.400 ;
        RECT 30.680 90.200 30.880 97.800 ;
        RECT 31.480 90.200 31.680 97.800 ;
        RECT 32.280 90.200 32.480 97.800 ;
        RECT 33.080 90.200 33.280 97.800 ;
        RECT 33.880 90.200 34.080 97.800 ;
        RECT 25.930 89.800 34.080 90.200 ;
        RECT 25.930 89.600 26.330 89.800 ;
        RECT 25.930 89.400 29.930 89.600 ;
        RECT 25.930 88.800 26.330 89.400 ;
        RECT 25.930 88.600 29.930 88.800 ;
        RECT 25.930 88.000 26.330 88.600 ;
        RECT 25.930 87.800 29.930 88.000 ;
        RECT 25.930 87.200 26.330 87.800 ;
        RECT 25.930 87.000 29.930 87.200 ;
        RECT 25.930 86.400 26.330 87.000 ;
        RECT 25.930 86.200 29.930 86.400 ;
        RECT 25.930 85.600 26.330 86.200 ;
        RECT 25.930 85.400 29.930 85.600 ;
        RECT 25.930 84.800 26.330 85.400 ;
        RECT 25.930 84.600 29.930 84.800 ;
        RECT 25.930 84.000 26.330 84.600 ;
        RECT 25.930 83.800 29.930 84.000 ;
        RECT 25.930 83.200 26.330 83.800 ;
        RECT 25.930 83.000 29.930 83.200 ;
        RECT 25.930 82.400 26.330 83.000 ;
        RECT 25.930 82.200 29.930 82.400 ;
        RECT 30.680 82.200 30.880 89.800 ;
        RECT 31.480 82.200 31.680 89.800 ;
        RECT 32.280 82.200 32.480 89.800 ;
        RECT 33.080 82.200 33.280 89.800 ;
        RECT 33.880 82.200 34.080 89.800 ;
        RECT 35.380 90.200 35.580 97.800 ;
        RECT 36.180 90.200 36.380 97.800 ;
        RECT 36.980 90.200 37.180 97.800 ;
        RECT 37.780 90.200 37.980 97.800 ;
        RECT 38.580 90.200 38.780 97.800 ;
        RECT 39.530 97.600 43.530 97.800 ;
        RECT 43.130 97.000 43.530 97.600 ;
        RECT 39.530 96.800 43.530 97.000 ;
        RECT 43.130 96.200 43.530 96.800 ;
        RECT 39.530 96.000 43.530 96.200 ;
        RECT 43.130 95.400 43.530 96.000 ;
        RECT 39.530 95.200 43.530 95.400 ;
        RECT 43.130 94.600 43.530 95.200 ;
        RECT 39.530 94.400 43.530 94.600 ;
        RECT 43.130 93.800 43.530 94.400 ;
        RECT 39.530 93.600 43.530 93.800 ;
        RECT 43.130 93.000 43.530 93.600 ;
        RECT 39.530 92.800 43.530 93.000 ;
        RECT 43.130 92.200 43.530 92.800 ;
        RECT 39.530 92.000 43.530 92.200 ;
        RECT 43.130 91.400 43.530 92.000 ;
        RECT 39.530 91.200 43.530 91.400 ;
        RECT 43.130 90.600 43.530 91.200 ;
        RECT 39.530 90.400 43.530 90.600 ;
        RECT 43.130 90.200 43.530 90.400 ;
        RECT 35.380 89.800 43.530 90.200 ;
        RECT 35.380 82.200 35.580 89.800 ;
        RECT 36.180 82.200 36.380 89.800 ;
        RECT 36.980 82.200 37.180 89.800 ;
        RECT 37.780 82.200 37.980 89.800 ;
        RECT 38.580 82.200 38.780 89.800 ;
        RECT 43.130 89.600 43.530 89.800 ;
        RECT 39.530 89.400 43.530 89.600 ;
        RECT 43.130 88.800 43.530 89.400 ;
        RECT 39.530 88.600 43.530 88.800 ;
        RECT 43.130 88.000 43.530 88.600 ;
        RECT 39.530 87.800 43.530 88.000 ;
        RECT 43.130 87.200 43.530 87.800 ;
        RECT 39.530 87.000 43.530 87.200 ;
        RECT 43.130 86.400 43.530 87.000 ;
        RECT 39.530 86.200 43.530 86.400 ;
        RECT 43.130 85.600 43.530 86.200 ;
        RECT 39.530 85.400 43.530 85.600 ;
        RECT 43.130 84.800 43.530 85.400 ;
        RECT 39.530 84.600 43.530 84.800 ;
        RECT 43.130 84.000 43.530 84.600 ;
        RECT 39.530 83.800 43.530 84.000 ;
        RECT 43.130 83.200 43.530 83.800 ;
        RECT 39.530 83.000 43.530 83.200 ;
        RECT 43.130 82.400 43.530 83.000 ;
        RECT 39.530 82.200 43.530 82.400 ;
        RECT 45.930 97.600 49.930 97.800 ;
        RECT 45.930 97.000 46.330 97.600 ;
        RECT 45.930 96.800 49.930 97.000 ;
        RECT 45.930 96.200 46.330 96.800 ;
        RECT 45.930 96.000 49.930 96.200 ;
        RECT 45.930 95.400 46.330 96.000 ;
        RECT 45.930 95.200 49.930 95.400 ;
        RECT 45.930 94.600 46.330 95.200 ;
        RECT 45.930 94.400 49.930 94.600 ;
        RECT 45.930 93.800 46.330 94.400 ;
        RECT 45.930 93.600 49.930 93.800 ;
        RECT 45.930 93.000 46.330 93.600 ;
        RECT 45.930 92.800 49.930 93.000 ;
        RECT 45.930 92.200 46.330 92.800 ;
        RECT 45.930 92.000 49.930 92.200 ;
        RECT 45.930 91.400 46.330 92.000 ;
        RECT 45.930 91.200 49.930 91.400 ;
        RECT 45.930 90.600 46.330 91.200 ;
        RECT 45.930 90.400 49.930 90.600 ;
        RECT 45.930 90.200 46.330 90.400 ;
        RECT 50.680 90.200 50.880 97.800 ;
        RECT 51.480 90.200 51.680 97.800 ;
        RECT 52.280 90.200 52.480 97.800 ;
        RECT 53.080 90.200 53.280 97.800 ;
        RECT 53.880 90.200 54.080 97.800 ;
        RECT 45.930 89.800 54.080 90.200 ;
        RECT 45.930 89.600 46.330 89.800 ;
        RECT 45.930 89.400 49.930 89.600 ;
        RECT 45.930 88.800 46.330 89.400 ;
        RECT 45.930 88.600 49.930 88.800 ;
        RECT 45.930 88.000 46.330 88.600 ;
        RECT 45.930 87.800 49.930 88.000 ;
        RECT 45.930 87.200 46.330 87.800 ;
        RECT 45.930 87.000 49.930 87.200 ;
        RECT 45.930 86.400 46.330 87.000 ;
        RECT 45.930 86.200 49.930 86.400 ;
        RECT 45.930 85.600 46.330 86.200 ;
        RECT 45.930 85.400 49.930 85.600 ;
        RECT 45.930 84.800 46.330 85.400 ;
        RECT 45.930 84.600 49.930 84.800 ;
        RECT 45.930 84.000 46.330 84.600 ;
        RECT 45.930 83.800 49.930 84.000 ;
        RECT 45.930 83.200 46.330 83.800 ;
        RECT 45.930 83.000 49.930 83.200 ;
        RECT 45.930 82.400 46.330 83.000 ;
        RECT 45.930 82.200 49.930 82.400 ;
        RECT 50.680 82.200 50.880 89.800 ;
        RECT 51.480 82.200 51.680 89.800 ;
        RECT 52.280 82.200 52.480 89.800 ;
        RECT 53.080 82.200 53.280 89.800 ;
        RECT 53.880 82.200 54.080 89.800 ;
        RECT 55.380 90.200 55.580 97.800 ;
        RECT 56.180 90.200 56.380 97.800 ;
        RECT 56.980 90.200 57.180 97.800 ;
        RECT 57.780 90.200 57.980 97.800 ;
        RECT 58.580 90.200 58.780 97.800 ;
        RECT 59.530 97.600 63.530 97.800 ;
        RECT 63.130 97.000 63.530 97.600 ;
        RECT 59.530 96.800 63.530 97.000 ;
        RECT 63.130 96.200 63.530 96.800 ;
        RECT 59.530 96.000 63.530 96.200 ;
        RECT 63.130 95.400 63.530 96.000 ;
        RECT 59.530 95.200 63.530 95.400 ;
        RECT 63.130 94.600 63.530 95.200 ;
        RECT 59.530 94.400 63.530 94.600 ;
        RECT 63.130 93.800 63.530 94.400 ;
        RECT 59.530 93.600 63.530 93.800 ;
        RECT 63.130 93.000 63.530 93.600 ;
        RECT 59.530 92.800 63.530 93.000 ;
        RECT 63.130 92.200 63.530 92.800 ;
        RECT 59.530 92.000 63.530 92.200 ;
        RECT 63.130 91.400 63.530 92.000 ;
        RECT 59.530 91.200 63.530 91.400 ;
        RECT 63.130 90.600 63.530 91.200 ;
        RECT 59.530 90.400 63.530 90.600 ;
        RECT 63.130 90.200 63.530 90.400 ;
        RECT 55.380 89.800 63.530 90.200 ;
        RECT 55.380 82.200 55.580 89.800 ;
        RECT 56.180 82.200 56.380 89.800 ;
        RECT 56.980 82.200 57.180 89.800 ;
        RECT 57.780 82.200 57.980 89.800 ;
        RECT 58.580 82.200 58.780 89.800 ;
        RECT 63.130 89.600 63.530 89.800 ;
        RECT 59.530 89.400 63.530 89.600 ;
        RECT 63.130 88.800 63.530 89.400 ;
        RECT 59.530 88.600 63.530 88.800 ;
        RECT 63.130 88.000 63.530 88.600 ;
        RECT 59.530 87.800 63.530 88.000 ;
        RECT 63.130 87.200 63.530 87.800 ;
        RECT 59.530 87.000 63.530 87.200 ;
        RECT 63.130 86.400 63.530 87.000 ;
        RECT 59.530 86.200 63.530 86.400 ;
        RECT 63.130 85.600 63.530 86.200 ;
        RECT 59.530 85.400 63.530 85.600 ;
        RECT 63.130 84.800 63.530 85.400 ;
        RECT 59.530 84.600 63.530 84.800 ;
        RECT 63.130 84.000 63.530 84.600 ;
        RECT 59.530 83.800 63.530 84.000 ;
        RECT 63.130 83.200 63.530 83.800 ;
        RECT 59.530 83.000 63.530 83.200 ;
        RECT 63.130 82.400 63.530 83.000 ;
        RECT 59.530 82.200 63.530 82.400 ;
        RECT 65.930 97.600 69.930 97.800 ;
        RECT 65.930 97.000 66.330 97.600 ;
        RECT 65.930 96.800 69.930 97.000 ;
        RECT 65.930 96.200 66.330 96.800 ;
        RECT 65.930 96.000 69.930 96.200 ;
        RECT 65.930 95.400 66.330 96.000 ;
        RECT 65.930 95.200 69.930 95.400 ;
        RECT 65.930 94.600 66.330 95.200 ;
        RECT 65.930 94.400 69.930 94.600 ;
        RECT 65.930 93.800 66.330 94.400 ;
        RECT 65.930 93.600 69.930 93.800 ;
        RECT 65.930 93.000 66.330 93.600 ;
        RECT 65.930 92.800 69.930 93.000 ;
        RECT 65.930 92.200 66.330 92.800 ;
        RECT 65.930 92.000 69.930 92.200 ;
        RECT 65.930 91.400 66.330 92.000 ;
        RECT 65.930 91.200 69.930 91.400 ;
        RECT 65.930 90.600 66.330 91.200 ;
        RECT 65.930 90.400 69.930 90.600 ;
        RECT 65.930 90.200 66.330 90.400 ;
        RECT 70.680 90.200 70.880 97.800 ;
        RECT 71.480 90.200 71.680 97.800 ;
        RECT 72.280 90.200 72.480 97.800 ;
        RECT 73.080 90.200 73.280 97.800 ;
        RECT 73.880 90.200 74.080 97.800 ;
        RECT 65.930 89.800 74.080 90.200 ;
        RECT 65.930 89.600 66.330 89.800 ;
        RECT 65.930 89.400 69.930 89.600 ;
        RECT 65.930 88.800 66.330 89.400 ;
        RECT 65.930 88.600 69.930 88.800 ;
        RECT 65.930 88.000 66.330 88.600 ;
        RECT 65.930 87.800 69.930 88.000 ;
        RECT 65.930 87.200 66.330 87.800 ;
        RECT 65.930 87.000 69.930 87.200 ;
        RECT 65.930 86.400 66.330 87.000 ;
        RECT 65.930 86.200 69.930 86.400 ;
        RECT 65.930 85.600 66.330 86.200 ;
        RECT 65.930 85.400 69.930 85.600 ;
        RECT 65.930 84.800 66.330 85.400 ;
        RECT 65.930 84.600 69.930 84.800 ;
        RECT 65.930 84.000 66.330 84.600 ;
        RECT 65.930 83.800 69.930 84.000 ;
        RECT 65.930 83.200 66.330 83.800 ;
        RECT 65.930 83.000 69.930 83.200 ;
        RECT 65.930 82.400 66.330 83.000 ;
        RECT 65.930 82.200 69.930 82.400 ;
        RECT 70.680 82.200 70.880 89.800 ;
        RECT 71.480 82.200 71.680 89.800 ;
        RECT 72.280 82.200 72.480 89.800 ;
        RECT 73.080 82.200 73.280 89.800 ;
        RECT 73.880 82.200 74.080 89.800 ;
        RECT 75.380 90.200 75.580 97.800 ;
        RECT 76.180 90.200 76.380 97.800 ;
        RECT 76.980 90.200 77.180 97.800 ;
        RECT 77.780 90.200 77.980 97.800 ;
        RECT 78.580 90.200 78.780 97.800 ;
        RECT 79.530 97.600 83.530 97.800 ;
        RECT 83.130 97.000 83.530 97.600 ;
        RECT 79.530 96.800 83.530 97.000 ;
        RECT 83.130 96.200 83.530 96.800 ;
        RECT 79.530 96.000 83.530 96.200 ;
        RECT 83.130 95.400 83.530 96.000 ;
        RECT 79.530 95.200 83.530 95.400 ;
        RECT 83.130 94.600 83.530 95.200 ;
        RECT 79.530 94.400 83.530 94.600 ;
        RECT 83.130 93.800 83.530 94.400 ;
        RECT 79.530 93.600 83.530 93.800 ;
        RECT 83.130 93.000 83.530 93.600 ;
        RECT 79.530 92.800 83.530 93.000 ;
        RECT 83.130 92.200 83.530 92.800 ;
        RECT 79.530 92.000 83.530 92.200 ;
        RECT 83.130 91.400 83.530 92.000 ;
        RECT 79.530 91.200 83.530 91.400 ;
        RECT 83.130 90.600 83.530 91.200 ;
        RECT 79.530 90.400 83.530 90.600 ;
        RECT 83.130 90.200 83.530 90.400 ;
        RECT 75.380 89.800 83.530 90.200 ;
        RECT 75.380 82.200 75.580 89.800 ;
        RECT 76.180 82.200 76.380 89.800 ;
        RECT 76.980 82.200 77.180 89.800 ;
        RECT 77.780 82.200 77.980 89.800 ;
        RECT 78.580 82.200 78.780 89.800 ;
        RECT 83.130 89.600 83.530 89.800 ;
        RECT 79.530 89.400 83.530 89.600 ;
        RECT 83.130 88.800 83.530 89.400 ;
        RECT 79.530 88.600 83.530 88.800 ;
        RECT 83.130 88.000 83.530 88.600 ;
        RECT 79.530 87.800 83.530 88.000 ;
        RECT 83.130 87.200 83.530 87.800 ;
        RECT 79.530 87.000 83.530 87.200 ;
        RECT 83.130 86.400 83.530 87.000 ;
        RECT 79.530 86.200 83.530 86.400 ;
        RECT 83.130 85.600 83.530 86.200 ;
        RECT 79.530 85.400 83.530 85.600 ;
        RECT 83.130 84.800 83.530 85.400 ;
        RECT 79.530 84.600 83.530 84.800 ;
        RECT 83.130 84.000 83.530 84.600 ;
        RECT 79.530 83.800 83.530 84.000 ;
        RECT 83.130 83.200 83.530 83.800 ;
        RECT 79.530 83.000 83.530 83.200 ;
        RECT 83.130 82.400 83.530 83.000 ;
        RECT 79.530 82.200 83.530 82.400 ;
        RECT 85.930 97.600 89.930 97.800 ;
        RECT 85.930 97.000 86.330 97.600 ;
        RECT 85.930 96.800 89.930 97.000 ;
        RECT 85.930 96.200 86.330 96.800 ;
        RECT 85.930 96.000 89.930 96.200 ;
        RECT 85.930 95.400 86.330 96.000 ;
        RECT 85.930 95.200 89.930 95.400 ;
        RECT 85.930 94.600 86.330 95.200 ;
        RECT 85.930 94.400 89.930 94.600 ;
        RECT 85.930 93.800 86.330 94.400 ;
        RECT 85.930 93.600 89.930 93.800 ;
        RECT 85.930 93.000 86.330 93.600 ;
        RECT 85.930 92.800 89.930 93.000 ;
        RECT 85.930 92.200 86.330 92.800 ;
        RECT 85.930 92.000 89.930 92.200 ;
        RECT 85.930 91.400 86.330 92.000 ;
        RECT 85.930 91.200 89.930 91.400 ;
        RECT 85.930 90.600 86.330 91.200 ;
        RECT 85.930 90.400 89.930 90.600 ;
        RECT 85.930 90.200 86.330 90.400 ;
        RECT 90.680 90.200 90.880 97.800 ;
        RECT 91.480 90.200 91.680 97.800 ;
        RECT 92.280 90.200 92.480 97.800 ;
        RECT 93.080 90.200 93.280 97.800 ;
        RECT 93.880 90.200 94.080 97.800 ;
        RECT 85.930 89.800 94.080 90.200 ;
        RECT 85.930 89.600 86.330 89.800 ;
        RECT 85.930 89.400 89.930 89.600 ;
        RECT 85.930 88.800 86.330 89.400 ;
        RECT 85.930 88.600 89.930 88.800 ;
        RECT 85.930 88.000 86.330 88.600 ;
        RECT 85.930 87.800 89.930 88.000 ;
        RECT 85.930 87.200 86.330 87.800 ;
        RECT 85.930 87.000 89.930 87.200 ;
        RECT 85.930 86.400 86.330 87.000 ;
        RECT 85.930 86.200 89.930 86.400 ;
        RECT 85.930 85.600 86.330 86.200 ;
        RECT 85.930 85.400 89.930 85.600 ;
        RECT 85.930 84.800 86.330 85.400 ;
        RECT 85.930 84.600 89.930 84.800 ;
        RECT 85.930 84.000 86.330 84.600 ;
        RECT 85.930 83.800 89.930 84.000 ;
        RECT 85.930 83.200 86.330 83.800 ;
        RECT 85.930 83.000 89.930 83.200 ;
        RECT 85.930 82.400 86.330 83.000 ;
        RECT 85.930 82.200 89.930 82.400 ;
        RECT 90.680 82.200 90.880 89.800 ;
        RECT 91.480 82.200 91.680 89.800 ;
        RECT 92.280 82.200 92.480 89.800 ;
        RECT 93.080 82.200 93.280 89.800 ;
        RECT 93.880 82.200 94.080 89.800 ;
        RECT 95.380 90.200 95.580 97.800 ;
        RECT 96.180 90.200 96.380 97.800 ;
        RECT 96.980 90.200 97.180 97.800 ;
        RECT 97.780 90.200 97.980 97.800 ;
        RECT 98.580 90.200 98.780 97.800 ;
        RECT 99.530 97.600 103.530 97.800 ;
        RECT 103.130 97.000 103.530 97.600 ;
        RECT 99.530 96.800 103.530 97.000 ;
        RECT 103.130 96.200 103.530 96.800 ;
        RECT 99.530 96.000 103.530 96.200 ;
        RECT 103.130 95.400 103.530 96.000 ;
        RECT 99.530 95.200 103.530 95.400 ;
        RECT 103.130 94.600 103.530 95.200 ;
        RECT 99.530 94.400 103.530 94.600 ;
        RECT 103.130 93.800 103.530 94.400 ;
        RECT 99.530 93.600 103.530 93.800 ;
        RECT 103.130 93.000 103.530 93.600 ;
        RECT 99.530 92.800 103.530 93.000 ;
        RECT 103.130 92.200 103.530 92.800 ;
        RECT 99.530 92.000 103.530 92.200 ;
        RECT 103.130 91.400 103.530 92.000 ;
        RECT 99.530 91.200 103.530 91.400 ;
        RECT 103.130 90.600 103.530 91.200 ;
        RECT 99.530 90.400 103.530 90.600 ;
        RECT 103.130 90.200 103.530 90.400 ;
        RECT 95.380 89.800 103.530 90.200 ;
        RECT 95.380 82.200 95.580 89.800 ;
        RECT 96.180 82.200 96.380 89.800 ;
        RECT 96.980 82.200 97.180 89.800 ;
        RECT 97.780 82.200 97.980 89.800 ;
        RECT 98.580 82.200 98.780 89.800 ;
        RECT 103.130 89.600 103.530 89.800 ;
        RECT 99.530 89.400 103.530 89.600 ;
        RECT 103.130 88.800 103.530 89.400 ;
        RECT 99.530 88.600 103.530 88.800 ;
        RECT 103.130 88.000 103.530 88.600 ;
        RECT 99.530 87.800 103.530 88.000 ;
        RECT 103.130 87.200 103.530 87.800 ;
        RECT 99.530 87.000 103.530 87.200 ;
        RECT 103.130 86.400 103.530 87.000 ;
        RECT 99.530 86.200 103.530 86.400 ;
        RECT 103.130 85.600 103.530 86.200 ;
        RECT 99.530 85.400 103.530 85.600 ;
        RECT 103.130 84.800 103.530 85.400 ;
        RECT 99.530 84.600 103.530 84.800 ;
        RECT 103.130 84.000 103.530 84.600 ;
        RECT 99.530 83.800 103.530 84.000 ;
        RECT 103.130 83.200 103.530 83.800 ;
        RECT 99.530 83.000 103.530 83.200 ;
        RECT 103.130 82.400 103.530 83.000 ;
        RECT 99.530 82.200 103.530 82.400 ;
        RECT 105.930 97.600 109.930 97.800 ;
        RECT 105.930 97.000 106.330 97.600 ;
        RECT 105.930 96.800 109.930 97.000 ;
        RECT 105.930 96.200 106.330 96.800 ;
        RECT 105.930 96.000 109.930 96.200 ;
        RECT 105.930 95.400 106.330 96.000 ;
        RECT 105.930 95.200 109.930 95.400 ;
        RECT 105.930 94.600 106.330 95.200 ;
        RECT 105.930 94.400 109.930 94.600 ;
        RECT 105.930 93.800 106.330 94.400 ;
        RECT 105.930 93.600 109.930 93.800 ;
        RECT 105.930 93.000 106.330 93.600 ;
        RECT 105.930 92.800 109.930 93.000 ;
        RECT 105.930 92.200 106.330 92.800 ;
        RECT 105.930 92.000 109.930 92.200 ;
        RECT 105.930 91.400 106.330 92.000 ;
        RECT 105.930 91.200 109.930 91.400 ;
        RECT 105.930 90.600 106.330 91.200 ;
        RECT 105.930 90.400 109.930 90.600 ;
        RECT 105.930 90.200 106.330 90.400 ;
        RECT 110.680 90.200 110.880 97.800 ;
        RECT 111.480 90.200 111.680 97.800 ;
        RECT 112.280 90.200 112.480 97.800 ;
        RECT 113.080 90.200 113.280 97.800 ;
        RECT 113.880 90.200 114.080 97.800 ;
        RECT 105.930 89.800 114.080 90.200 ;
        RECT 105.930 89.600 106.330 89.800 ;
        RECT 105.930 89.400 109.930 89.600 ;
        RECT 105.930 88.800 106.330 89.400 ;
        RECT 105.930 88.600 109.930 88.800 ;
        RECT 105.930 88.000 106.330 88.600 ;
        RECT 105.930 87.800 109.930 88.000 ;
        RECT 105.930 87.200 106.330 87.800 ;
        RECT 105.930 87.000 109.930 87.200 ;
        RECT 105.930 86.400 106.330 87.000 ;
        RECT 105.930 86.200 109.930 86.400 ;
        RECT 105.930 85.600 106.330 86.200 ;
        RECT 105.930 85.400 109.930 85.600 ;
        RECT 105.930 84.800 106.330 85.400 ;
        RECT 105.930 84.600 109.930 84.800 ;
        RECT 105.930 84.000 106.330 84.600 ;
        RECT 105.930 83.800 109.930 84.000 ;
        RECT 105.930 83.200 106.330 83.800 ;
        RECT 105.930 83.000 109.930 83.200 ;
        RECT 105.930 82.400 106.330 83.000 ;
        RECT 105.930 82.200 109.930 82.400 ;
        RECT 110.680 82.200 110.880 89.800 ;
        RECT 111.480 82.200 111.680 89.800 ;
        RECT 112.280 82.200 112.480 89.800 ;
        RECT 113.080 82.200 113.280 89.800 ;
        RECT 113.880 82.200 114.080 89.800 ;
        RECT 115.380 90.200 115.580 97.800 ;
        RECT 116.180 90.200 116.380 97.800 ;
        RECT 116.980 90.200 117.180 97.800 ;
        RECT 117.780 90.200 117.980 97.800 ;
        RECT 118.580 90.200 118.780 97.800 ;
        RECT 119.530 97.600 123.530 97.800 ;
        RECT 123.130 97.000 123.530 97.600 ;
        RECT 119.530 96.800 123.530 97.000 ;
        RECT 123.130 96.200 123.530 96.800 ;
        RECT 119.530 96.000 123.530 96.200 ;
        RECT 123.130 95.400 123.530 96.000 ;
        RECT 119.530 95.200 123.530 95.400 ;
        RECT 123.130 94.600 123.530 95.200 ;
        RECT 119.530 94.400 123.530 94.600 ;
        RECT 123.130 93.800 123.530 94.400 ;
        RECT 119.530 93.600 123.530 93.800 ;
        RECT 123.130 93.000 123.530 93.600 ;
        RECT 119.530 92.800 123.530 93.000 ;
        RECT 123.130 92.200 123.530 92.800 ;
        RECT 119.530 92.000 123.530 92.200 ;
        RECT 123.130 91.400 123.530 92.000 ;
        RECT 119.530 91.200 123.530 91.400 ;
        RECT 123.130 90.600 123.530 91.200 ;
        RECT 119.530 90.400 123.530 90.600 ;
        RECT 130.050 90.525 130.410 90.905 ;
        RECT 130.680 90.525 131.040 90.905 ;
        RECT 131.280 90.525 131.640 90.905 ;
        RECT 123.130 90.200 123.530 90.400 ;
        RECT 115.380 89.800 123.530 90.200 ;
        RECT 130.050 89.935 130.410 90.315 ;
        RECT 130.680 89.935 131.040 90.315 ;
        RECT 131.280 89.935 131.640 90.315 ;
        RECT 115.380 82.200 115.580 89.800 ;
        RECT 116.180 82.200 116.380 89.800 ;
        RECT 116.980 82.200 117.180 89.800 ;
        RECT 117.780 82.200 117.980 89.800 ;
        RECT 118.580 82.200 118.780 89.800 ;
        RECT 123.130 89.600 123.530 89.800 ;
        RECT 119.530 89.400 123.530 89.600 ;
        RECT 123.130 88.800 123.530 89.400 ;
        RECT 119.530 88.600 123.530 88.800 ;
        RECT 123.130 88.000 123.530 88.600 ;
        RECT 119.530 87.800 123.530 88.000 ;
        RECT 123.130 87.200 123.530 87.800 ;
        RECT 119.530 87.000 123.530 87.200 ;
        RECT 123.130 86.400 123.530 87.000 ;
        RECT 119.530 86.200 123.530 86.400 ;
        RECT 123.130 85.600 123.530 86.200 ;
        RECT 119.530 85.400 123.530 85.600 ;
        RECT 123.130 84.800 123.530 85.400 ;
        RECT 119.530 84.600 123.530 84.800 ;
        RECT 123.130 84.000 123.530 84.600 ;
        RECT 119.530 83.800 123.530 84.000 ;
        RECT 123.130 83.200 123.530 83.800 ;
        RECT 119.530 83.000 123.530 83.200 ;
        RECT 123.130 82.400 123.530 83.000 ;
        RECT 119.530 82.200 123.530 82.400 ;
        RECT 5.930 77.600 9.930 77.800 ;
        RECT 5.930 77.000 6.330 77.600 ;
        RECT 5.930 76.800 9.930 77.000 ;
        RECT 5.930 76.200 6.330 76.800 ;
        RECT 5.930 76.000 9.930 76.200 ;
        RECT 5.930 75.400 6.330 76.000 ;
        RECT 5.930 75.200 9.930 75.400 ;
        RECT 5.930 74.600 6.330 75.200 ;
        RECT 5.930 74.400 9.930 74.600 ;
        RECT 5.930 73.800 6.330 74.400 ;
        RECT 5.930 73.600 9.930 73.800 ;
        RECT 5.930 73.000 6.330 73.600 ;
        RECT 5.930 72.800 9.930 73.000 ;
        RECT 5.930 72.200 6.330 72.800 ;
        RECT 5.930 72.000 9.930 72.200 ;
        RECT 5.930 71.400 6.330 72.000 ;
        RECT 5.930 71.200 9.930 71.400 ;
        RECT 5.930 70.600 6.330 71.200 ;
        RECT 5.930 70.400 9.930 70.600 ;
        RECT 5.930 70.200 6.330 70.400 ;
        RECT 10.680 70.200 10.880 77.800 ;
        RECT 11.480 70.200 11.680 77.800 ;
        RECT 12.280 70.200 12.480 77.800 ;
        RECT 13.080 70.200 13.280 77.800 ;
        RECT 13.880 70.200 14.080 77.800 ;
        RECT 5.930 69.800 14.080 70.200 ;
        RECT 5.930 69.600 6.330 69.800 ;
        RECT 5.930 69.400 9.930 69.600 ;
        RECT 5.930 68.800 6.330 69.400 ;
        RECT 5.930 68.600 9.930 68.800 ;
        RECT 5.930 68.000 6.330 68.600 ;
        RECT 5.930 67.800 9.930 68.000 ;
        RECT 5.930 67.200 6.330 67.800 ;
        RECT 5.930 67.000 9.930 67.200 ;
        RECT 5.930 66.400 6.330 67.000 ;
        RECT 5.930 66.200 9.930 66.400 ;
        RECT 5.930 65.600 6.330 66.200 ;
        RECT 5.930 65.400 9.930 65.600 ;
        RECT 5.930 64.800 6.330 65.400 ;
        RECT 5.930 64.600 9.930 64.800 ;
        RECT 5.930 64.000 6.330 64.600 ;
        RECT 5.930 63.800 9.930 64.000 ;
        RECT 5.930 63.200 6.330 63.800 ;
        RECT 5.930 63.000 9.930 63.200 ;
        RECT 5.930 62.400 6.330 63.000 ;
        RECT 5.930 62.200 9.930 62.400 ;
        RECT 10.680 62.200 10.880 69.800 ;
        RECT 11.480 62.200 11.680 69.800 ;
        RECT 12.280 62.200 12.480 69.800 ;
        RECT 13.080 62.200 13.280 69.800 ;
        RECT 13.880 62.200 14.080 69.800 ;
        RECT 15.380 70.200 15.580 77.800 ;
        RECT 16.180 70.200 16.380 77.800 ;
        RECT 16.980 70.200 17.180 77.800 ;
        RECT 17.780 70.200 17.980 77.800 ;
        RECT 18.580 70.200 18.780 77.800 ;
        RECT 19.530 77.600 23.530 77.800 ;
        RECT 23.130 77.000 23.530 77.600 ;
        RECT 19.530 76.800 23.530 77.000 ;
        RECT 23.130 76.200 23.530 76.800 ;
        RECT 19.530 76.000 23.530 76.200 ;
        RECT 23.130 75.400 23.530 76.000 ;
        RECT 19.530 75.200 23.530 75.400 ;
        RECT 23.130 74.600 23.530 75.200 ;
        RECT 19.530 74.400 23.530 74.600 ;
        RECT 23.130 73.800 23.530 74.400 ;
        RECT 19.530 73.600 23.530 73.800 ;
        RECT 23.130 73.000 23.530 73.600 ;
        RECT 19.530 72.800 23.530 73.000 ;
        RECT 23.130 72.200 23.530 72.800 ;
        RECT 19.530 72.000 23.530 72.200 ;
        RECT 23.130 71.400 23.530 72.000 ;
        RECT 19.530 71.200 23.530 71.400 ;
        RECT 23.130 70.600 23.530 71.200 ;
        RECT 19.530 70.400 23.530 70.600 ;
        RECT 23.130 70.200 23.530 70.400 ;
        RECT 15.380 69.800 23.530 70.200 ;
        RECT 15.380 62.200 15.580 69.800 ;
        RECT 16.180 62.200 16.380 69.800 ;
        RECT 16.980 62.200 17.180 69.800 ;
        RECT 17.780 62.200 17.980 69.800 ;
        RECT 18.580 62.200 18.780 69.800 ;
        RECT 23.130 69.600 23.530 69.800 ;
        RECT 19.530 69.400 23.530 69.600 ;
        RECT 23.130 68.800 23.530 69.400 ;
        RECT 19.530 68.600 23.530 68.800 ;
        RECT 23.130 68.000 23.530 68.600 ;
        RECT 19.530 67.800 23.530 68.000 ;
        RECT 23.130 67.200 23.530 67.800 ;
        RECT 19.530 67.000 23.530 67.200 ;
        RECT 23.130 66.400 23.530 67.000 ;
        RECT 19.530 66.200 23.530 66.400 ;
        RECT 23.130 65.600 23.530 66.200 ;
        RECT 19.530 65.400 23.530 65.600 ;
        RECT 23.130 64.800 23.530 65.400 ;
        RECT 19.530 64.600 23.530 64.800 ;
        RECT 23.130 64.000 23.530 64.600 ;
        RECT 19.530 63.800 23.530 64.000 ;
        RECT 23.130 63.200 23.530 63.800 ;
        RECT 19.530 63.000 23.530 63.200 ;
        RECT 23.130 62.400 23.530 63.000 ;
        RECT 19.530 62.200 23.530 62.400 ;
        RECT 25.930 77.600 29.930 77.800 ;
        RECT 25.930 77.000 26.330 77.600 ;
        RECT 25.930 76.800 29.930 77.000 ;
        RECT 25.930 76.200 26.330 76.800 ;
        RECT 25.930 76.000 29.930 76.200 ;
        RECT 25.930 75.400 26.330 76.000 ;
        RECT 25.930 75.200 29.930 75.400 ;
        RECT 25.930 74.600 26.330 75.200 ;
        RECT 25.930 74.400 29.930 74.600 ;
        RECT 25.930 73.800 26.330 74.400 ;
        RECT 25.930 73.600 29.930 73.800 ;
        RECT 25.930 73.000 26.330 73.600 ;
        RECT 25.930 72.800 29.930 73.000 ;
        RECT 25.930 72.200 26.330 72.800 ;
        RECT 25.930 72.000 29.930 72.200 ;
        RECT 25.930 71.400 26.330 72.000 ;
        RECT 25.930 71.200 29.930 71.400 ;
        RECT 25.930 70.600 26.330 71.200 ;
        RECT 25.930 70.400 29.930 70.600 ;
        RECT 25.930 70.200 26.330 70.400 ;
        RECT 30.680 70.200 30.880 77.800 ;
        RECT 31.480 70.200 31.680 77.800 ;
        RECT 32.280 70.200 32.480 77.800 ;
        RECT 33.080 70.200 33.280 77.800 ;
        RECT 33.880 70.200 34.080 77.800 ;
        RECT 25.930 69.800 34.080 70.200 ;
        RECT 25.930 69.600 26.330 69.800 ;
        RECT 25.930 69.400 29.930 69.600 ;
        RECT 25.930 68.800 26.330 69.400 ;
        RECT 25.930 68.600 29.930 68.800 ;
        RECT 25.930 68.000 26.330 68.600 ;
        RECT 25.930 67.800 29.930 68.000 ;
        RECT 25.930 67.200 26.330 67.800 ;
        RECT 25.930 67.000 29.930 67.200 ;
        RECT 25.930 66.400 26.330 67.000 ;
        RECT 25.930 66.200 29.930 66.400 ;
        RECT 25.930 65.600 26.330 66.200 ;
        RECT 25.930 65.400 29.930 65.600 ;
        RECT 25.930 64.800 26.330 65.400 ;
        RECT 25.930 64.600 29.930 64.800 ;
        RECT 25.930 64.000 26.330 64.600 ;
        RECT 25.930 63.800 29.930 64.000 ;
        RECT 25.930 63.200 26.330 63.800 ;
        RECT 25.930 63.000 29.930 63.200 ;
        RECT 25.930 62.400 26.330 63.000 ;
        RECT 25.930 62.200 29.930 62.400 ;
        RECT 30.680 62.200 30.880 69.800 ;
        RECT 31.480 62.200 31.680 69.800 ;
        RECT 32.280 62.200 32.480 69.800 ;
        RECT 33.080 62.200 33.280 69.800 ;
        RECT 33.880 62.200 34.080 69.800 ;
        RECT 35.380 70.200 35.580 77.800 ;
        RECT 36.180 70.200 36.380 77.800 ;
        RECT 36.980 70.200 37.180 77.800 ;
        RECT 37.780 70.200 37.980 77.800 ;
        RECT 38.580 70.200 38.780 77.800 ;
        RECT 39.530 77.600 43.530 77.800 ;
        RECT 43.130 77.000 43.530 77.600 ;
        RECT 39.530 76.800 43.530 77.000 ;
        RECT 43.130 76.200 43.530 76.800 ;
        RECT 39.530 76.000 43.530 76.200 ;
        RECT 43.130 75.400 43.530 76.000 ;
        RECT 39.530 75.200 43.530 75.400 ;
        RECT 43.130 74.600 43.530 75.200 ;
        RECT 39.530 74.400 43.530 74.600 ;
        RECT 43.130 73.800 43.530 74.400 ;
        RECT 39.530 73.600 43.530 73.800 ;
        RECT 43.130 73.000 43.530 73.600 ;
        RECT 39.530 72.800 43.530 73.000 ;
        RECT 43.130 72.200 43.530 72.800 ;
        RECT 39.530 72.000 43.530 72.200 ;
        RECT 43.130 71.400 43.530 72.000 ;
        RECT 39.530 71.200 43.530 71.400 ;
        RECT 43.130 70.600 43.530 71.200 ;
        RECT 39.530 70.400 43.530 70.600 ;
        RECT 43.130 70.200 43.530 70.400 ;
        RECT 35.380 69.800 43.530 70.200 ;
        RECT 35.380 62.200 35.580 69.800 ;
        RECT 36.180 62.200 36.380 69.800 ;
        RECT 36.980 62.200 37.180 69.800 ;
        RECT 37.780 62.200 37.980 69.800 ;
        RECT 38.580 62.200 38.780 69.800 ;
        RECT 43.130 69.600 43.530 69.800 ;
        RECT 39.530 69.400 43.530 69.600 ;
        RECT 43.130 68.800 43.530 69.400 ;
        RECT 39.530 68.600 43.530 68.800 ;
        RECT 43.130 68.000 43.530 68.600 ;
        RECT 39.530 67.800 43.530 68.000 ;
        RECT 43.130 67.200 43.530 67.800 ;
        RECT 39.530 67.000 43.530 67.200 ;
        RECT 43.130 66.400 43.530 67.000 ;
        RECT 39.530 66.200 43.530 66.400 ;
        RECT 43.130 65.600 43.530 66.200 ;
        RECT 39.530 65.400 43.530 65.600 ;
        RECT 43.130 64.800 43.530 65.400 ;
        RECT 39.530 64.600 43.530 64.800 ;
        RECT 43.130 64.000 43.530 64.600 ;
        RECT 39.530 63.800 43.530 64.000 ;
        RECT 43.130 63.200 43.530 63.800 ;
        RECT 39.530 63.000 43.530 63.200 ;
        RECT 43.130 62.400 43.530 63.000 ;
        RECT 39.530 62.200 43.530 62.400 ;
        RECT 45.930 77.600 49.930 77.800 ;
        RECT 45.930 77.000 46.330 77.600 ;
        RECT 45.930 76.800 49.930 77.000 ;
        RECT 45.930 76.200 46.330 76.800 ;
        RECT 45.930 76.000 49.930 76.200 ;
        RECT 45.930 75.400 46.330 76.000 ;
        RECT 45.930 75.200 49.930 75.400 ;
        RECT 45.930 74.600 46.330 75.200 ;
        RECT 45.930 74.400 49.930 74.600 ;
        RECT 45.930 73.800 46.330 74.400 ;
        RECT 45.930 73.600 49.930 73.800 ;
        RECT 45.930 73.000 46.330 73.600 ;
        RECT 45.930 72.800 49.930 73.000 ;
        RECT 45.930 72.200 46.330 72.800 ;
        RECT 45.930 72.000 49.930 72.200 ;
        RECT 45.930 71.400 46.330 72.000 ;
        RECT 45.930 71.200 49.930 71.400 ;
        RECT 45.930 70.600 46.330 71.200 ;
        RECT 45.930 70.400 49.930 70.600 ;
        RECT 45.930 70.200 46.330 70.400 ;
        RECT 50.680 70.200 50.880 77.800 ;
        RECT 51.480 70.200 51.680 77.800 ;
        RECT 52.280 70.200 52.480 77.800 ;
        RECT 53.080 70.200 53.280 77.800 ;
        RECT 53.880 70.200 54.080 77.800 ;
        RECT 45.930 69.800 54.080 70.200 ;
        RECT 45.930 69.600 46.330 69.800 ;
        RECT 45.930 69.400 49.930 69.600 ;
        RECT 45.930 68.800 46.330 69.400 ;
        RECT 45.930 68.600 49.930 68.800 ;
        RECT 45.930 68.000 46.330 68.600 ;
        RECT 45.930 67.800 49.930 68.000 ;
        RECT 45.930 67.200 46.330 67.800 ;
        RECT 45.930 67.000 49.930 67.200 ;
        RECT 45.930 66.400 46.330 67.000 ;
        RECT 45.930 66.200 49.930 66.400 ;
        RECT 45.930 65.600 46.330 66.200 ;
        RECT 45.930 65.400 49.930 65.600 ;
        RECT 45.930 64.800 46.330 65.400 ;
        RECT 45.930 64.600 49.930 64.800 ;
        RECT 45.930 64.000 46.330 64.600 ;
        RECT 45.930 63.800 49.930 64.000 ;
        RECT 45.930 63.200 46.330 63.800 ;
        RECT 45.930 63.000 49.930 63.200 ;
        RECT 45.930 62.400 46.330 63.000 ;
        RECT 45.930 62.200 49.930 62.400 ;
        RECT 50.680 62.200 50.880 69.800 ;
        RECT 51.480 62.200 51.680 69.800 ;
        RECT 52.280 62.200 52.480 69.800 ;
        RECT 53.080 62.200 53.280 69.800 ;
        RECT 53.880 62.200 54.080 69.800 ;
        RECT 55.380 70.200 55.580 77.800 ;
        RECT 56.180 70.200 56.380 77.800 ;
        RECT 56.980 70.200 57.180 77.800 ;
        RECT 57.780 70.200 57.980 77.800 ;
        RECT 58.580 70.200 58.780 77.800 ;
        RECT 59.530 77.600 63.530 77.800 ;
        RECT 63.130 77.000 63.530 77.600 ;
        RECT 59.530 76.800 63.530 77.000 ;
        RECT 63.130 76.200 63.530 76.800 ;
        RECT 59.530 76.000 63.530 76.200 ;
        RECT 63.130 75.400 63.530 76.000 ;
        RECT 59.530 75.200 63.530 75.400 ;
        RECT 63.130 74.600 63.530 75.200 ;
        RECT 59.530 74.400 63.530 74.600 ;
        RECT 63.130 73.800 63.530 74.400 ;
        RECT 59.530 73.600 63.530 73.800 ;
        RECT 63.130 73.000 63.530 73.600 ;
        RECT 59.530 72.800 63.530 73.000 ;
        RECT 63.130 72.200 63.530 72.800 ;
        RECT 59.530 72.000 63.530 72.200 ;
        RECT 63.130 71.400 63.530 72.000 ;
        RECT 59.530 71.200 63.530 71.400 ;
        RECT 63.130 70.600 63.530 71.200 ;
        RECT 59.530 70.400 63.530 70.600 ;
        RECT 63.130 70.200 63.530 70.400 ;
        RECT 55.380 69.800 63.530 70.200 ;
        RECT 55.380 62.200 55.580 69.800 ;
        RECT 56.180 62.200 56.380 69.800 ;
        RECT 56.980 62.200 57.180 69.800 ;
        RECT 57.780 62.200 57.980 69.800 ;
        RECT 58.580 62.200 58.780 69.800 ;
        RECT 63.130 69.600 63.530 69.800 ;
        RECT 59.530 69.400 63.530 69.600 ;
        RECT 63.130 68.800 63.530 69.400 ;
        RECT 59.530 68.600 63.530 68.800 ;
        RECT 63.130 68.000 63.530 68.600 ;
        RECT 59.530 67.800 63.530 68.000 ;
        RECT 63.130 67.200 63.530 67.800 ;
        RECT 59.530 67.000 63.530 67.200 ;
        RECT 63.130 66.400 63.530 67.000 ;
        RECT 59.530 66.200 63.530 66.400 ;
        RECT 63.130 65.600 63.530 66.200 ;
        RECT 59.530 65.400 63.530 65.600 ;
        RECT 63.130 64.800 63.530 65.400 ;
        RECT 59.530 64.600 63.530 64.800 ;
        RECT 63.130 64.000 63.530 64.600 ;
        RECT 59.530 63.800 63.530 64.000 ;
        RECT 63.130 63.200 63.530 63.800 ;
        RECT 59.530 63.000 63.530 63.200 ;
        RECT 63.130 62.400 63.530 63.000 ;
        RECT 59.530 62.200 63.530 62.400 ;
        RECT 65.930 77.600 69.930 77.800 ;
        RECT 65.930 77.000 66.330 77.600 ;
        RECT 65.930 76.800 69.930 77.000 ;
        RECT 65.930 76.200 66.330 76.800 ;
        RECT 65.930 76.000 69.930 76.200 ;
        RECT 65.930 75.400 66.330 76.000 ;
        RECT 65.930 75.200 69.930 75.400 ;
        RECT 65.930 74.600 66.330 75.200 ;
        RECT 65.930 74.400 69.930 74.600 ;
        RECT 65.930 73.800 66.330 74.400 ;
        RECT 65.930 73.600 69.930 73.800 ;
        RECT 65.930 73.000 66.330 73.600 ;
        RECT 65.930 72.800 69.930 73.000 ;
        RECT 65.930 72.200 66.330 72.800 ;
        RECT 65.930 72.000 69.930 72.200 ;
        RECT 65.930 71.400 66.330 72.000 ;
        RECT 65.930 71.200 69.930 71.400 ;
        RECT 65.930 70.600 66.330 71.200 ;
        RECT 65.930 70.400 69.930 70.600 ;
        RECT 65.930 70.200 66.330 70.400 ;
        RECT 70.680 70.200 70.880 77.800 ;
        RECT 71.480 70.200 71.680 77.800 ;
        RECT 72.280 70.200 72.480 77.800 ;
        RECT 73.080 70.200 73.280 77.800 ;
        RECT 73.880 70.200 74.080 77.800 ;
        RECT 65.930 69.800 74.080 70.200 ;
        RECT 65.930 69.600 66.330 69.800 ;
        RECT 65.930 69.400 69.930 69.600 ;
        RECT 65.930 68.800 66.330 69.400 ;
        RECT 65.930 68.600 69.930 68.800 ;
        RECT 65.930 68.000 66.330 68.600 ;
        RECT 65.930 67.800 69.930 68.000 ;
        RECT 65.930 67.200 66.330 67.800 ;
        RECT 65.930 67.000 69.930 67.200 ;
        RECT 65.930 66.400 66.330 67.000 ;
        RECT 65.930 66.200 69.930 66.400 ;
        RECT 65.930 65.600 66.330 66.200 ;
        RECT 65.930 65.400 69.930 65.600 ;
        RECT 65.930 64.800 66.330 65.400 ;
        RECT 65.930 64.600 69.930 64.800 ;
        RECT 65.930 64.000 66.330 64.600 ;
        RECT 65.930 63.800 69.930 64.000 ;
        RECT 65.930 63.200 66.330 63.800 ;
        RECT 65.930 63.000 69.930 63.200 ;
        RECT 65.930 62.400 66.330 63.000 ;
        RECT 65.930 62.200 69.930 62.400 ;
        RECT 70.680 62.200 70.880 69.800 ;
        RECT 71.480 62.200 71.680 69.800 ;
        RECT 72.280 62.200 72.480 69.800 ;
        RECT 73.080 62.200 73.280 69.800 ;
        RECT 73.880 62.200 74.080 69.800 ;
        RECT 75.380 70.200 75.580 77.800 ;
        RECT 76.180 70.200 76.380 77.800 ;
        RECT 76.980 70.200 77.180 77.800 ;
        RECT 77.780 70.200 77.980 77.800 ;
        RECT 78.580 70.200 78.780 77.800 ;
        RECT 79.530 77.600 83.530 77.800 ;
        RECT 83.130 77.000 83.530 77.600 ;
        RECT 79.530 76.800 83.530 77.000 ;
        RECT 83.130 76.200 83.530 76.800 ;
        RECT 79.530 76.000 83.530 76.200 ;
        RECT 83.130 75.400 83.530 76.000 ;
        RECT 79.530 75.200 83.530 75.400 ;
        RECT 83.130 74.600 83.530 75.200 ;
        RECT 79.530 74.400 83.530 74.600 ;
        RECT 83.130 73.800 83.530 74.400 ;
        RECT 79.530 73.600 83.530 73.800 ;
        RECT 83.130 73.000 83.530 73.600 ;
        RECT 79.530 72.800 83.530 73.000 ;
        RECT 83.130 72.200 83.530 72.800 ;
        RECT 79.530 72.000 83.530 72.200 ;
        RECT 83.130 71.400 83.530 72.000 ;
        RECT 79.530 71.200 83.530 71.400 ;
        RECT 83.130 70.600 83.530 71.200 ;
        RECT 79.530 70.400 83.530 70.600 ;
        RECT 83.130 70.200 83.530 70.400 ;
        RECT 75.380 69.800 83.530 70.200 ;
        RECT 75.380 62.200 75.580 69.800 ;
        RECT 76.180 62.200 76.380 69.800 ;
        RECT 76.980 62.200 77.180 69.800 ;
        RECT 77.780 62.200 77.980 69.800 ;
        RECT 78.580 62.200 78.780 69.800 ;
        RECT 83.130 69.600 83.530 69.800 ;
        RECT 79.530 69.400 83.530 69.600 ;
        RECT 83.130 68.800 83.530 69.400 ;
        RECT 79.530 68.600 83.530 68.800 ;
        RECT 83.130 68.000 83.530 68.600 ;
        RECT 79.530 67.800 83.530 68.000 ;
        RECT 83.130 67.200 83.530 67.800 ;
        RECT 79.530 67.000 83.530 67.200 ;
        RECT 83.130 66.400 83.530 67.000 ;
        RECT 79.530 66.200 83.530 66.400 ;
        RECT 83.130 65.600 83.530 66.200 ;
        RECT 79.530 65.400 83.530 65.600 ;
        RECT 83.130 64.800 83.530 65.400 ;
        RECT 79.530 64.600 83.530 64.800 ;
        RECT 83.130 64.000 83.530 64.600 ;
        RECT 79.530 63.800 83.530 64.000 ;
        RECT 83.130 63.200 83.530 63.800 ;
        RECT 79.530 63.000 83.530 63.200 ;
        RECT 83.130 62.400 83.530 63.000 ;
        RECT 79.530 62.200 83.530 62.400 ;
        RECT 85.930 77.600 89.930 77.800 ;
        RECT 85.930 77.000 86.330 77.600 ;
        RECT 85.930 76.800 89.930 77.000 ;
        RECT 85.930 76.200 86.330 76.800 ;
        RECT 85.930 76.000 89.930 76.200 ;
        RECT 85.930 75.400 86.330 76.000 ;
        RECT 85.930 75.200 89.930 75.400 ;
        RECT 85.930 74.600 86.330 75.200 ;
        RECT 85.930 74.400 89.930 74.600 ;
        RECT 85.930 73.800 86.330 74.400 ;
        RECT 85.930 73.600 89.930 73.800 ;
        RECT 85.930 73.000 86.330 73.600 ;
        RECT 85.930 72.800 89.930 73.000 ;
        RECT 85.930 72.200 86.330 72.800 ;
        RECT 85.930 72.000 89.930 72.200 ;
        RECT 85.930 71.400 86.330 72.000 ;
        RECT 85.930 71.200 89.930 71.400 ;
        RECT 85.930 70.600 86.330 71.200 ;
        RECT 85.930 70.400 89.930 70.600 ;
        RECT 85.930 70.200 86.330 70.400 ;
        RECT 90.680 70.200 90.880 77.800 ;
        RECT 91.480 70.200 91.680 77.800 ;
        RECT 92.280 70.200 92.480 77.800 ;
        RECT 93.080 70.200 93.280 77.800 ;
        RECT 93.880 70.200 94.080 77.800 ;
        RECT 85.930 69.800 94.080 70.200 ;
        RECT 85.930 69.600 86.330 69.800 ;
        RECT 85.930 69.400 89.930 69.600 ;
        RECT 85.930 68.800 86.330 69.400 ;
        RECT 85.930 68.600 89.930 68.800 ;
        RECT 85.930 68.000 86.330 68.600 ;
        RECT 85.930 67.800 89.930 68.000 ;
        RECT 85.930 67.200 86.330 67.800 ;
        RECT 85.930 67.000 89.930 67.200 ;
        RECT 85.930 66.400 86.330 67.000 ;
        RECT 85.930 66.200 89.930 66.400 ;
        RECT 85.930 65.600 86.330 66.200 ;
        RECT 85.930 65.400 89.930 65.600 ;
        RECT 85.930 64.800 86.330 65.400 ;
        RECT 85.930 64.600 89.930 64.800 ;
        RECT 85.930 64.000 86.330 64.600 ;
        RECT 85.930 63.800 89.930 64.000 ;
        RECT 85.930 63.200 86.330 63.800 ;
        RECT 85.930 63.000 89.930 63.200 ;
        RECT 85.930 62.400 86.330 63.000 ;
        RECT 85.930 62.200 89.930 62.400 ;
        RECT 90.680 62.200 90.880 69.800 ;
        RECT 91.480 62.200 91.680 69.800 ;
        RECT 92.280 62.200 92.480 69.800 ;
        RECT 93.080 62.200 93.280 69.800 ;
        RECT 93.880 62.200 94.080 69.800 ;
        RECT 95.380 70.200 95.580 77.800 ;
        RECT 96.180 70.200 96.380 77.800 ;
        RECT 96.980 70.200 97.180 77.800 ;
        RECT 97.780 70.200 97.980 77.800 ;
        RECT 98.580 70.200 98.780 77.800 ;
        RECT 99.530 77.600 103.530 77.800 ;
        RECT 103.130 77.000 103.530 77.600 ;
        RECT 99.530 76.800 103.530 77.000 ;
        RECT 103.130 76.200 103.530 76.800 ;
        RECT 99.530 76.000 103.530 76.200 ;
        RECT 103.130 75.400 103.530 76.000 ;
        RECT 99.530 75.200 103.530 75.400 ;
        RECT 103.130 74.600 103.530 75.200 ;
        RECT 99.530 74.400 103.530 74.600 ;
        RECT 103.130 73.800 103.530 74.400 ;
        RECT 99.530 73.600 103.530 73.800 ;
        RECT 103.130 73.000 103.530 73.600 ;
        RECT 99.530 72.800 103.530 73.000 ;
        RECT 103.130 72.200 103.530 72.800 ;
        RECT 99.530 72.000 103.530 72.200 ;
        RECT 103.130 71.400 103.530 72.000 ;
        RECT 99.530 71.200 103.530 71.400 ;
        RECT 103.130 70.600 103.530 71.200 ;
        RECT 99.530 70.400 103.530 70.600 ;
        RECT 103.130 70.200 103.530 70.400 ;
        RECT 95.380 69.800 103.530 70.200 ;
        RECT 95.380 62.200 95.580 69.800 ;
        RECT 96.180 62.200 96.380 69.800 ;
        RECT 96.980 62.200 97.180 69.800 ;
        RECT 97.780 62.200 97.980 69.800 ;
        RECT 98.580 62.200 98.780 69.800 ;
        RECT 103.130 69.600 103.530 69.800 ;
        RECT 99.530 69.400 103.530 69.600 ;
        RECT 103.130 68.800 103.530 69.400 ;
        RECT 99.530 68.600 103.530 68.800 ;
        RECT 103.130 68.000 103.530 68.600 ;
        RECT 99.530 67.800 103.530 68.000 ;
        RECT 103.130 67.200 103.530 67.800 ;
        RECT 99.530 67.000 103.530 67.200 ;
        RECT 103.130 66.400 103.530 67.000 ;
        RECT 99.530 66.200 103.530 66.400 ;
        RECT 103.130 65.600 103.530 66.200 ;
        RECT 99.530 65.400 103.530 65.600 ;
        RECT 103.130 64.800 103.530 65.400 ;
        RECT 99.530 64.600 103.530 64.800 ;
        RECT 103.130 64.000 103.530 64.600 ;
        RECT 99.530 63.800 103.530 64.000 ;
        RECT 103.130 63.200 103.530 63.800 ;
        RECT 99.530 63.000 103.530 63.200 ;
        RECT 103.130 62.400 103.530 63.000 ;
        RECT 99.530 62.200 103.530 62.400 ;
        RECT 105.930 77.600 109.930 77.800 ;
        RECT 105.930 77.000 106.330 77.600 ;
        RECT 105.930 76.800 109.930 77.000 ;
        RECT 105.930 76.200 106.330 76.800 ;
        RECT 105.930 76.000 109.930 76.200 ;
        RECT 105.930 75.400 106.330 76.000 ;
        RECT 105.930 75.200 109.930 75.400 ;
        RECT 105.930 74.600 106.330 75.200 ;
        RECT 105.930 74.400 109.930 74.600 ;
        RECT 105.930 73.800 106.330 74.400 ;
        RECT 105.930 73.600 109.930 73.800 ;
        RECT 105.930 73.000 106.330 73.600 ;
        RECT 105.930 72.800 109.930 73.000 ;
        RECT 105.930 72.200 106.330 72.800 ;
        RECT 105.930 72.000 109.930 72.200 ;
        RECT 105.930 71.400 106.330 72.000 ;
        RECT 105.930 71.200 109.930 71.400 ;
        RECT 105.930 70.600 106.330 71.200 ;
        RECT 105.930 70.400 109.930 70.600 ;
        RECT 105.930 70.200 106.330 70.400 ;
        RECT 110.680 70.200 110.880 77.800 ;
        RECT 111.480 70.200 111.680 77.800 ;
        RECT 112.280 70.200 112.480 77.800 ;
        RECT 113.080 70.200 113.280 77.800 ;
        RECT 113.880 70.200 114.080 77.800 ;
        RECT 105.930 69.800 114.080 70.200 ;
        RECT 105.930 69.600 106.330 69.800 ;
        RECT 105.930 69.400 109.930 69.600 ;
        RECT 105.930 68.800 106.330 69.400 ;
        RECT 105.930 68.600 109.930 68.800 ;
        RECT 105.930 68.000 106.330 68.600 ;
        RECT 105.930 67.800 109.930 68.000 ;
        RECT 105.930 67.200 106.330 67.800 ;
        RECT 105.930 67.000 109.930 67.200 ;
        RECT 105.930 66.400 106.330 67.000 ;
        RECT 105.930 66.200 109.930 66.400 ;
        RECT 105.930 65.600 106.330 66.200 ;
        RECT 105.930 65.400 109.930 65.600 ;
        RECT 105.930 64.800 106.330 65.400 ;
        RECT 105.930 64.600 109.930 64.800 ;
        RECT 105.930 64.000 106.330 64.600 ;
        RECT 105.930 63.800 109.930 64.000 ;
        RECT 105.930 63.200 106.330 63.800 ;
        RECT 105.930 63.000 109.930 63.200 ;
        RECT 105.930 62.400 106.330 63.000 ;
        RECT 105.930 62.200 109.930 62.400 ;
        RECT 110.680 62.200 110.880 69.800 ;
        RECT 111.480 62.200 111.680 69.800 ;
        RECT 112.280 62.200 112.480 69.800 ;
        RECT 113.080 62.200 113.280 69.800 ;
        RECT 113.880 62.200 114.080 69.800 ;
        RECT 115.380 70.200 115.580 77.800 ;
        RECT 116.180 70.200 116.380 77.800 ;
        RECT 116.980 70.200 117.180 77.800 ;
        RECT 117.780 70.200 117.980 77.800 ;
        RECT 118.580 70.200 118.780 77.800 ;
        RECT 119.530 77.600 123.530 77.800 ;
        RECT 123.130 77.000 123.530 77.600 ;
        RECT 119.530 76.800 123.530 77.000 ;
        RECT 123.130 76.200 123.530 76.800 ;
        RECT 119.530 76.000 123.530 76.200 ;
        RECT 123.130 75.400 123.530 76.000 ;
        RECT 119.530 75.200 123.530 75.400 ;
        RECT 123.130 74.600 123.530 75.200 ;
        RECT 119.530 74.400 123.530 74.600 ;
        RECT 123.130 73.800 123.530 74.400 ;
        RECT 119.530 73.600 123.530 73.800 ;
        RECT 123.130 73.000 123.530 73.600 ;
        RECT 119.530 72.800 123.530 73.000 ;
        RECT 123.130 72.200 123.530 72.800 ;
        RECT 119.530 72.000 123.530 72.200 ;
        RECT 123.130 71.400 123.530 72.000 ;
        RECT 119.530 71.200 123.530 71.400 ;
        RECT 123.130 70.600 123.530 71.200 ;
        RECT 119.530 70.400 123.530 70.600 ;
        RECT 123.130 70.200 123.530 70.400 ;
        RECT 115.380 69.800 123.530 70.200 ;
        RECT 130.050 69.990 130.410 70.370 ;
        RECT 130.680 69.990 131.040 70.370 ;
        RECT 131.280 69.990 131.640 70.370 ;
        RECT 115.380 62.200 115.580 69.800 ;
        RECT 116.180 62.200 116.380 69.800 ;
        RECT 116.980 62.200 117.180 69.800 ;
        RECT 117.780 62.200 117.980 69.800 ;
        RECT 118.580 62.200 118.780 69.800 ;
        RECT 123.130 69.600 123.530 69.800 ;
        RECT 119.530 69.400 123.530 69.600 ;
        RECT 130.050 69.400 130.410 69.780 ;
        RECT 130.680 69.400 131.040 69.780 ;
        RECT 131.280 69.400 131.640 69.780 ;
        RECT 123.130 68.800 123.530 69.400 ;
        RECT 119.530 68.600 123.530 68.800 ;
        RECT 123.130 68.000 123.530 68.600 ;
        RECT 119.530 67.800 123.530 68.000 ;
        RECT 123.130 67.200 123.530 67.800 ;
        RECT 119.530 67.000 123.530 67.200 ;
        RECT 123.130 66.400 123.530 67.000 ;
        RECT 119.530 66.200 123.530 66.400 ;
        RECT 123.130 65.600 123.530 66.200 ;
        RECT 119.530 65.400 123.530 65.600 ;
        RECT 123.130 64.800 123.530 65.400 ;
        RECT 119.530 64.600 123.530 64.800 ;
        RECT 123.130 64.000 123.530 64.600 ;
        RECT 119.530 63.800 123.530 64.000 ;
        RECT 123.130 63.200 123.530 63.800 ;
        RECT 119.530 63.000 123.530 63.200 ;
        RECT 123.130 62.400 123.530 63.000 ;
        RECT 119.530 62.200 123.530 62.400 ;
        RECT 5.930 57.600 9.930 57.800 ;
        RECT 5.930 57.000 6.330 57.600 ;
        RECT 5.930 56.800 9.930 57.000 ;
        RECT 5.930 56.200 6.330 56.800 ;
        RECT 5.930 56.000 9.930 56.200 ;
        RECT 5.930 55.400 6.330 56.000 ;
        RECT 5.930 55.200 9.930 55.400 ;
        RECT 5.930 54.600 6.330 55.200 ;
        RECT 5.930 54.400 9.930 54.600 ;
        RECT 5.930 53.800 6.330 54.400 ;
        RECT 5.930 53.600 9.930 53.800 ;
        RECT 5.930 53.000 6.330 53.600 ;
        RECT 5.930 52.800 9.930 53.000 ;
        RECT 5.930 52.200 6.330 52.800 ;
        RECT 5.930 52.000 9.930 52.200 ;
        RECT 5.930 51.400 6.330 52.000 ;
        RECT 5.930 51.200 9.930 51.400 ;
        RECT 5.930 50.600 6.330 51.200 ;
        RECT 5.930 50.400 9.930 50.600 ;
        RECT 5.930 50.200 6.330 50.400 ;
        RECT 10.680 50.200 10.880 57.800 ;
        RECT 11.480 50.200 11.680 57.800 ;
        RECT 12.280 50.200 12.480 57.800 ;
        RECT 13.080 50.200 13.280 57.800 ;
        RECT 13.880 50.200 14.080 57.800 ;
        RECT 5.930 49.800 14.080 50.200 ;
        RECT 5.930 49.600 6.330 49.800 ;
        RECT 5.930 49.400 9.930 49.600 ;
        RECT 5.930 48.800 6.330 49.400 ;
        RECT 5.930 48.600 9.930 48.800 ;
        RECT 5.930 48.000 6.330 48.600 ;
        RECT 5.930 47.800 9.930 48.000 ;
        RECT 5.930 47.200 6.330 47.800 ;
        RECT 5.930 47.000 9.930 47.200 ;
        RECT 5.930 46.400 6.330 47.000 ;
        RECT 5.930 46.200 9.930 46.400 ;
        RECT 5.930 45.600 6.330 46.200 ;
        RECT 5.930 45.400 9.930 45.600 ;
        RECT 5.930 44.800 6.330 45.400 ;
        RECT 5.930 44.600 9.930 44.800 ;
        RECT 5.930 44.000 6.330 44.600 ;
        RECT 5.930 43.800 9.930 44.000 ;
        RECT 5.930 43.200 6.330 43.800 ;
        RECT 5.930 43.000 9.930 43.200 ;
        RECT 5.930 42.400 6.330 43.000 ;
        RECT 5.930 42.200 9.930 42.400 ;
        RECT 10.680 42.200 10.880 49.800 ;
        RECT 11.480 42.200 11.680 49.800 ;
        RECT 12.280 42.200 12.480 49.800 ;
        RECT 13.080 42.200 13.280 49.800 ;
        RECT 13.880 42.200 14.080 49.800 ;
        RECT 15.380 50.200 15.580 57.800 ;
        RECT 16.180 50.200 16.380 57.800 ;
        RECT 16.980 50.200 17.180 57.800 ;
        RECT 17.780 50.200 17.980 57.800 ;
        RECT 18.580 50.200 18.780 57.800 ;
        RECT 19.530 57.600 23.530 57.800 ;
        RECT 23.130 57.000 23.530 57.600 ;
        RECT 19.530 56.800 23.530 57.000 ;
        RECT 23.130 56.200 23.530 56.800 ;
        RECT 19.530 56.000 23.530 56.200 ;
        RECT 23.130 55.400 23.530 56.000 ;
        RECT 19.530 55.200 23.530 55.400 ;
        RECT 23.130 54.600 23.530 55.200 ;
        RECT 19.530 54.400 23.530 54.600 ;
        RECT 23.130 53.800 23.530 54.400 ;
        RECT 19.530 53.600 23.530 53.800 ;
        RECT 23.130 53.000 23.530 53.600 ;
        RECT 19.530 52.800 23.530 53.000 ;
        RECT 23.130 52.200 23.530 52.800 ;
        RECT 19.530 52.000 23.530 52.200 ;
        RECT 23.130 51.400 23.530 52.000 ;
        RECT 19.530 51.200 23.530 51.400 ;
        RECT 23.130 50.600 23.530 51.200 ;
        RECT 19.530 50.400 23.530 50.600 ;
        RECT 23.130 50.200 23.530 50.400 ;
        RECT 15.380 49.800 23.530 50.200 ;
        RECT 15.380 42.200 15.580 49.800 ;
        RECT 16.180 42.200 16.380 49.800 ;
        RECT 16.980 42.200 17.180 49.800 ;
        RECT 17.780 42.200 17.980 49.800 ;
        RECT 18.580 42.200 18.780 49.800 ;
        RECT 23.130 49.600 23.530 49.800 ;
        RECT 19.530 49.400 23.530 49.600 ;
        RECT 23.130 48.800 23.530 49.400 ;
        RECT 19.530 48.600 23.530 48.800 ;
        RECT 23.130 48.000 23.530 48.600 ;
        RECT 19.530 47.800 23.530 48.000 ;
        RECT 23.130 47.200 23.530 47.800 ;
        RECT 19.530 47.000 23.530 47.200 ;
        RECT 23.130 46.400 23.530 47.000 ;
        RECT 19.530 46.200 23.530 46.400 ;
        RECT 23.130 45.600 23.530 46.200 ;
        RECT 19.530 45.400 23.530 45.600 ;
        RECT 23.130 44.800 23.530 45.400 ;
        RECT 19.530 44.600 23.530 44.800 ;
        RECT 23.130 44.000 23.530 44.600 ;
        RECT 19.530 43.800 23.530 44.000 ;
        RECT 23.130 43.200 23.530 43.800 ;
        RECT 19.530 43.000 23.530 43.200 ;
        RECT 23.130 42.400 23.530 43.000 ;
        RECT 19.530 42.200 23.530 42.400 ;
        RECT 25.930 57.600 29.930 57.800 ;
        RECT 25.930 57.000 26.330 57.600 ;
        RECT 25.930 56.800 29.930 57.000 ;
        RECT 25.930 56.200 26.330 56.800 ;
        RECT 25.930 56.000 29.930 56.200 ;
        RECT 25.930 55.400 26.330 56.000 ;
        RECT 25.930 55.200 29.930 55.400 ;
        RECT 25.930 54.600 26.330 55.200 ;
        RECT 25.930 54.400 29.930 54.600 ;
        RECT 25.930 53.800 26.330 54.400 ;
        RECT 25.930 53.600 29.930 53.800 ;
        RECT 25.930 53.000 26.330 53.600 ;
        RECT 25.930 52.800 29.930 53.000 ;
        RECT 25.930 52.200 26.330 52.800 ;
        RECT 25.930 52.000 29.930 52.200 ;
        RECT 25.930 51.400 26.330 52.000 ;
        RECT 25.930 51.200 29.930 51.400 ;
        RECT 25.930 50.600 26.330 51.200 ;
        RECT 25.930 50.400 29.930 50.600 ;
        RECT 25.930 50.200 26.330 50.400 ;
        RECT 30.680 50.200 30.880 57.800 ;
        RECT 31.480 50.200 31.680 57.800 ;
        RECT 32.280 50.200 32.480 57.800 ;
        RECT 33.080 50.200 33.280 57.800 ;
        RECT 33.880 50.200 34.080 57.800 ;
        RECT 25.930 49.800 34.080 50.200 ;
        RECT 25.930 49.600 26.330 49.800 ;
        RECT 25.930 49.400 29.930 49.600 ;
        RECT 25.930 48.800 26.330 49.400 ;
        RECT 25.930 48.600 29.930 48.800 ;
        RECT 25.930 48.000 26.330 48.600 ;
        RECT 25.930 47.800 29.930 48.000 ;
        RECT 25.930 47.200 26.330 47.800 ;
        RECT 25.930 47.000 29.930 47.200 ;
        RECT 25.930 46.400 26.330 47.000 ;
        RECT 25.930 46.200 29.930 46.400 ;
        RECT 25.930 45.600 26.330 46.200 ;
        RECT 25.930 45.400 29.930 45.600 ;
        RECT 25.930 44.800 26.330 45.400 ;
        RECT 25.930 44.600 29.930 44.800 ;
        RECT 25.930 44.000 26.330 44.600 ;
        RECT 25.930 43.800 29.930 44.000 ;
        RECT 25.930 43.200 26.330 43.800 ;
        RECT 25.930 43.000 29.930 43.200 ;
        RECT 25.930 42.400 26.330 43.000 ;
        RECT 25.930 42.200 29.930 42.400 ;
        RECT 30.680 42.200 30.880 49.800 ;
        RECT 31.480 42.200 31.680 49.800 ;
        RECT 32.280 42.200 32.480 49.800 ;
        RECT 33.080 42.200 33.280 49.800 ;
        RECT 33.880 42.200 34.080 49.800 ;
        RECT 35.380 50.200 35.580 57.800 ;
        RECT 36.180 50.200 36.380 57.800 ;
        RECT 36.980 50.200 37.180 57.800 ;
        RECT 37.780 50.200 37.980 57.800 ;
        RECT 38.580 50.200 38.780 57.800 ;
        RECT 39.530 57.600 43.530 57.800 ;
        RECT 43.130 57.000 43.530 57.600 ;
        RECT 39.530 56.800 43.530 57.000 ;
        RECT 43.130 56.200 43.530 56.800 ;
        RECT 39.530 56.000 43.530 56.200 ;
        RECT 43.130 55.400 43.530 56.000 ;
        RECT 39.530 55.200 43.530 55.400 ;
        RECT 43.130 54.600 43.530 55.200 ;
        RECT 39.530 54.400 43.530 54.600 ;
        RECT 43.130 53.800 43.530 54.400 ;
        RECT 39.530 53.600 43.530 53.800 ;
        RECT 43.130 53.000 43.530 53.600 ;
        RECT 39.530 52.800 43.530 53.000 ;
        RECT 43.130 52.200 43.530 52.800 ;
        RECT 39.530 52.000 43.530 52.200 ;
        RECT 43.130 51.400 43.530 52.000 ;
        RECT 39.530 51.200 43.530 51.400 ;
        RECT 43.130 50.600 43.530 51.200 ;
        RECT 39.530 50.400 43.530 50.600 ;
        RECT 43.130 50.200 43.530 50.400 ;
        RECT 35.380 49.800 43.530 50.200 ;
        RECT 35.380 42.200 35.580 49.800 ;
        RECT 36.180 42.200 36.380 49.800 ;
        RECT 36.980 42.200 37.180 49.800 ;
        RECT 37.780 42.200 37.980 49.800 ;
        RECT 38.580 42.200 38.780 49.800 ;
        RECT 43.130 49.600 43.530 49.800 ;
        RECT 39.530 49.400 43.530 49.600 ;
        RECT 43.130 48.800 43.530 49.400 ;
        RECT 39.530 48.600 43.530 48.800 ;
        RECT 43.130 48.000 43.530 48.600 ;
        RECT 39.530 47.800 43.530 48.000 ;
        RECT 43.130 47.200 43.530 47.800 ;
        RECT 39.530 47.000 43.530 47.200 ;
        RECT 43.130 46.400 43.530 47.000 ;
        RECT 39.530 46.200 43.530 46.400 ;
        RECT 43.130 45.600 43.530 46.200 ;
        RECT 39.530 45.400 43.530 45.600 ;
        RECT 43.130 44.800 43.530 45.400 ;
        RECT 39.530 44.600 43.530 44.800 ;
        RECT 43.130 44.000 43.530 44.600 ;
        RECT 39.530 43.800 43.530 44.000 ;
        RECT 43.130 43.200 43.530 43.800 ;
        RECT 39.530 43.000 43.530 43.200 ;
        RECT 43.130 42.400 43.530 43.000 ;
        RECT 39.530 42.200 43.530 42.400 ;
        RECT 45.930 57.600 49.930 57.800 ;
        RECT 45.930 57.000 46.330 57.600 ;
        RECT 45.930 56.800 49.930 57.000 ;
        RECT 45.930 56.200 46.330 56.800 ;
        RECT 45.930 56.000 49.930 56.200 ;
        RECT 45.930 55.400 46.330 56.000 ;
        RECT 45.930 55.200 49.930 55.400 ;
        RECT 45.930 54.600 46.330 55.200 ;
        RECT 45.930 54.400 49.930 54.600 ;
        RECT 45.930 53.800 46.330 54.400 ;
        RECT 45.930 53.600 49.930 53.800 ;
        RECT 45.930 53.000 46.330 53.600 ;
        RECT 45.930 52.800 49.930 53.000 ;
        RECT 45.930 52.200 46.330 52.800 ;
        RECT 45.930 52.000 49.930 52.200 ;
        RECT 45.930 51.400 46.330 52.000 ;
        RECT 45.930 51.200 49.930 51.400 ;
        RECT 45.930 50.600 46.330 51.200 ;
        RECT 45.930 50.400 49.930 50.600 ;
        RECT 45.930 50.200 46.330 50.400 ;
        RECT 50.680 50.200 50.880 57.800 ;
        RECT 51.480 50.200 51.680 57.800 ;
        RECT 52.280 50.200 52.480 57.800 ;
        RECT 53.080 50.200 53.280 57.800 ;
        RECT 53.880 50.200 54.080 57.800 ;
        RECT 45.930 49.800 54.080 50.200 ;
        RECT 45.930 49.600 46.330 49.800 ;
        RECT 45.930 49.400 49.930 49.600 ;
        RECT 45.930 48.800 46.330 49.400 ;
        RECT 45.930 48.600 49.930 48.800 ;
        RECT 45.930 48.000 46.330 48.600 ;
        RECT 45.930 47.800 49.930 48.000 ;
        RECT 45.930 47.200 46.330 47.800 ;
        RECT 45.930 47.000 49.930 47.200 ;
        RECT 45.930 46.400 46.330 47.000 ;
        RECT 45.930 46.200 49.930 46.400 ;
        RECT 45.930 45.600 46.330 46.200 ;
        RECT 45.930 45.400 49.930 45.600 ;
        RECT 45.930 44.800 46.330 45.400 ;
        RECT 45.930 44.600 49.930 44.800 ;
        RECT 45.930 44.000 46.330 44.600 ;
        RECT 45.930 43.800 49.930 44.000 ;
        RECT 45.930 43.200 46.330 43.800 ;
        RECT 45.930 43.000 49.930 43.200 ;
        RECT 45.930 42.400 46.330 43.000 ;
        RECT 45.930 42.200 49.930 42.400 ;
        RECT 50.680 42.200 50.880 49.800 ;
        RECT 51.480 42.200 51.680 49.800 ;
        RECT 52.280 42.200 52.480 49.800 ;
        RECT 53.080 42.200 53.280 49.800 ;
        RECT 53.880 42.200 54.080 49.800 ;
        RECT 55.380 50.200 55.580 57.800 ;
        RECT 56.180 50.200 56.380 57.800 ;
        RECT 56.980 50.200 57.180 57.800 ;
        RECT 57.780 50.200 57.980 57.800 ;
        RECT 58.580 50.200 58.780 57.800 ;
        RECT 59.530 57.600 63.530 57.800 ;
        RECT 63.130 57.000 63.530 57.600 ;
        RECT 59.530 56.800 63.530 57.000 ;
        RECT 63.130 56.200 63.530 56.800 ;
        RECT 59.530 56.000 63.530 56.200 ;
        RECT 63.130 55.400 63.530 56.000 ;
        RECT 59.530 55.200 63.530 55.400 ;
        RECT 63.130 54.600 63.530 55.200 ;
        RECT 59.530 54.400 63.530 54.600 ;
        RECT 63.130 53.800 63.530 54.400 ;
        RECT 59.530 53.600 63.530 53.800 ;
        RECT 63.130 53.000 63.530 53.600 ;
        RECT 59.530 52.800 63.530 53.000 ;
        RECT 63.130 52.200 63.530 52.800 ;
        RECT 59.530 52.000 63.530 52.200 ;
        RECT 63.130 51.400 63.530 52.000 ;
        RECT 59.530 51.200 63.530 51.400 ;
        RECT 63.130 50.600 63.530 51.200 ;
        RECT 59.530 50.400 63.530 50.600 ;
        RECT 63.130 50.200 63.530 50.400 ;
        RECT 55.380 49.800 63.530 50.200 ;
        RECT 55.380 42.200 55.580 49.800 ;
        RECT 56.180 42.200 56.380 49.800 ;
        RECT 56.980 42.200 57.180 49.800 ;
        RECT 57.780 42.200 57.980 49.800 ;
        RECT 58.580 42.200 58.780 49.800 ;
        RECT 63.130 49.600 63.530 49.800 ;
        RECT 59.530 49.400 63.530 49.600 ;
        RECT 63.130 48.800 63.530 49.400 ;
        RECT 59.530 48.600 63.530 48.800 ;
        RECT 63.130 48.000 63.530 48.600 ;
        RECT 59.530 47.800 63.530 48.000 ;
        RECT 63.130 47.200 63.530 47.800 ;
        RECT 59.530 47.000 63.530 47.200 ;
        RECT 63.130 46.400 63.530 47.000 ;
        RECT 59.530 46.200 63.530 46.400 ;
        RECT 63.130 45.600 63.530 46.200 ;
        RECT 59.530 45.400 63.530 45.600 ;
        RECT 63.130 44.800 63.530 45.400 ;
        RECT 59.530 44.600 63.530 44.800 ;
        RECT 63.130 44.000 63.530 44.600 ;
        RECT 59.530 43.800 63.530 44.000 ;
        RECT 63.130 43.200 63.530 43.800 ;
        RECT 59.530 43.000 63.530 43.200 ;
        RECT 63.130 42.400 63.530 43.000 ;
        RECT 59.530 42.200 63.530 42.400 ;
        RECT 65.930 57.600 69.930 57.800 ;
        RECT 65.930 57.000 66.330 57.600 ;
        RECT 65.930 56.800 69.930 57.000 ;
        RECT 65.930 56.200 66.330 56.800 ;
        RECT 65.930 56.000 69.930 56.200 ;
        RECT 65.930 55.400 66.330 56.000 ;
        RECT 65.930 55.200 69.930 55.400 ;
        RECT 65.930 54.600 66.330 55.200 ;
        RECT 65.930 54.400 69.930 54.600 ;
        RECT 65.930 53.800 66.330 54.400 ;
        RECT 65.930 53.600 69.930 53.800 ;
        RECT 65.930 53.000 66.330 53.600 ;
        RECT 65.930 52.800 69.930 53.000 ;
        RECT 65.930 52.200 66.330 52.800 ;
        RECT 65.930 52.000 69.930 52.200 ;
        RECT 65.930 51.400 66.330 52.000 ;
        RECT 65.930 51.200 69.930 51.400 ;
        RECT 65.930 50.600 66.330 51.200 ;
        RECT 65.930 50.400 69.930 50.600 ;
        RECT 65.930 50.200 66.330 50.400 ;
        RECT 70.680 50.200 70.880 57.800 ;
        RECT 71.480 50.200 71.680 57.800 ;
        RECT 72.280 50.200 72.480 57.800 ;
        RECT 73.080 50.200 73.280 57.800 ;
        RECT 73.880 50.200 74.080 57.800 ;
        RECT 65.930 49.800 74.080 50.200 ;
        RECT 65.930 49.600 66.330 49.800 ;
        RECT 65.930 49.400 69.930 49.600 ;
        RECT 65.930 48.800 66.330 49.400 ;
        RECT 65.930 48.600 69.930 48.800 ;
        RECT 65.930 48.000 66.330 48.600 ;
        RECT 65.930 47.800 69.930 48.000 ;
        RECT 65.930 47.200 66.330 47.800 ;
        RECT 65.930 47.000 69.930 47.200 ;
        RECT 65.930 46.400 66.330 47.000 ;
        RECT 65.930 46.200 69.930 46.400 ;
        RECT 65.930 45.600 66.330 46.200 ;
        RECT 65.930 45.400 69.930 45.600 ;
        RECT 65.930 44.800 66.330 45.400 ;
        RECT 65.930 44.600 69.930 44.800 ;
        RECT 65.930 44.000 66.330 44.600 ;
        RECT 65.930 43.800 69.930 44.000 ;
        RECT 65.930 43.200 66.330 43.800 ;
        RECT 65.930 43.000 69.930 43.200 ;
        RECT 65.930 42.400 66.330 43.000 ;
        RECT 65.930 42.200 69.930 42.400 ;
        RECT 70.680 42.200 70.880 49.800 ;
        RECT 71.480 42.200 71.680 49.800 ;
        RECT 72.280 42.200 72.480 49.800 ;
        RECT 73.080 42.200 73.280 49.800 ;
        RECT 73.880 42.200 74.080 49.800 ;
        RECT 75.380 50.200 75.580 57.800 ;
        RECT 76.180 50.200 76.380 57.800 ;
        RECT 76.980 50.200 77.180 57.800 ;
        RECT 77.780 50.200 77.980 57.800 ;
        RECT 78.580 50.200 78.780 57.800 ;
        RECT 79.530 57.600 83.530 57.800 ;
        RECT 83.130 57.000 83.530 57.600 ;
        RECT 79.530 56.800 83.530 57.000 ;
        RECT 83.130 56.200 83.530 56.800 ;
        RECT 79.530 56.000 83.530 56.200 ;
        RECT 83.130 55.400 83.530 56.000 ;
        RECT 79.530 55.200 83.530 55.400 ;
        RECT 83.130 54.600 83.530 55.200 ;
        RECT 79.530 54.400 83.530 54.600 ;
        RECT 83.130 53.800 83.530 54.400 ;
        RECT 79.530 53.600 83.530 53.800 ;
        RECT 83.130 53.000 83.530 53.600 ;
        RECT 79.530 52.800 83.530 53.000 ;
        RECT 83.130 52.200 83.530 52.800 ;
        RECT 79.530 52.000 83.530 52.200 ;
        RECT 83.130 51.400 83.530 52.000 ;
        RECT 79.530 51.200 83.530 51.400 ;
        RECT 83.130 50.600 83.530 51.200 ;
        RECT 79.530 50.400 83.530 50.600 ;
        RECT 83.130 50.200 83.530 50.400 ;
        RECT 75.380 49.800 83.530 50.200 ;
        RECT 75.380 42.200 75.580 49.800 ;
        RECT 76.180 42.200 76.380 49.800 ;
        RECT 76.980 42.200 77.180 49.800 ;
        RECT 77.780 42.200 77.980 49.800 ;
        RECT 78.580 42.200 78.780 49.800 ;
        RECT 83.130 49.600 83.530 49.800 ;
        RECT 79.530 49.400 83.530 49.600 ;
        RECT 83.130 48.800 83.530 49.400 ;
        RECT 79.530 48.600 83.530 48.800 ;
        RECT 83.130 48.000 83.530 48.600 ;
        RECT 79.530 47.800 83.530 48.000 ;
        RECT 83.130 47.200 83.530 47.800 ;
        RECT 79.530 47.000 83.530 47.200 ;
        RECT 83.130 46.400 83.530 47.000 ;
        RECT 79.530 46.200 83.530 46.400 ;
        RECT 83.130 45.600 83.530 46.200 ;
        RECT 79.530 45.400 83.530 45.600 ;
        RECT 83.130 44.800 83.530 45.400 ;
        RECT 79.530 44.600 83.530 44.800 ;
        RECT 83.130 44.000 83.530 44.600 ;
        RECT 79.530 43.800 83.530 44.000 ;
        RECT 83.130 43.200 83.530 43.800 ;
        RECT 79.530 43.000 83.530 43.200 ;
        RECT 83.130 42.400 83.530 43.000 ;
        RECT 79.530 42.200 83.530 42.400 ;
        RECT 85.930 57.600 89.930 57.800 ;
        RECT 85.930 57.000 86.330 57.600 ;
        RECT 85.930 56.800 89.930 57.000 ;
        RECT 85.930 56.200 86.330 56.800 ;
        RECT 85.930 56.000 89.930 56.200 ;
        RECT 85.930 55.400 86.330 56.000 ;
        RECT 85.930 55.200 89.930 55.400 ;
        RECT 85.930 54.600 86.330 55.200 ;
        RECT 85.930 54.400 89.930 54.600 ;
        RECT 85.930 53.800 86.330 54.400 ;
        RECT 85.930 53.600 89.930 53.800 ;
        RECT 85.930 53.000 86.330 53.600 ;
        RECT 85.930 52.800 89.930 53.000 ;
        RECT 85.930 52.200 86.330 52.800 ;
        RECT 85.930 52.000 89.930 52.200 ;
        RECT 85.930 51.400 86.330 52.000 ;
        RECT 85.930 51.200 89.930 51.400 ;
        RECT 85.930 50.600 86.330 51.200 ;
        RECT 85.930 50.400 89.930 50.600 ;
        RECT 85.930 50.200 86.330 50.400 ;
        RECT 90.680 50.200 90.880 57.800 ;
        RECT 91.480 50.200 91.680 57.800 ;
        RECT 92.280 50.200 92.480 57.800 ;
        RECT 93.080 50.200 93.280 57.800 ;
        RECT 93.880 50.200 94.080 57.800 ;
        RECT 85.930 49.800 94.080 50.200 ;
        RECT 85.930 49.600 86.330 49.800 ;
        RECT 85.930 49.400 89.930 49.600 ;
        RECT 85.930 48.800 86.330 49.400 ;
        RECT 85.930 48.600 89.930 48.800 ;
        RECT 85.930 48.000 86.330 48.600 ;
        RECT 85.930 47.800 89.930 48.000 ;
        RECT 85.930 47.200 86.330 47.800 ;
        RECT 85.930 47.000 89.930 47.200 ;
        RECT 85.930 46.400 86.330 47.000 ;
        RECT 85.930 46.200 89.930 46.400 ;
        RECT 85.930 45.600 86.330 46.200 ;
        RECT 85.930 45.400 89.930 45.600 ;
        RECT 85.930 44.800 86.330 45.400 ;
        RECT 85.930 44.600 89.930 44.800 ;
        RECT 85.930 44.000 86.330 44.600 ;
        RECT 85.930 43.800 89.930 44.000 ;
        RECT 85.930 43.200 86.330 43.800 ;
        RECT 85.930 43.000 89.930 43.200 ;
        RECT 85.930 42.400 86.330 43.000 ;
        RECT 85.930 42.200 89.930 42.400 ;
        RECT 90.680 42.200 90.880 49.800 ;
        RECT 91.480 42.200 91.680 49.800 ;
        RECT 92.280 42.200 92.480 49.800 ;
        RECT 93.080 42.200 93.280 49.800 ;
        RECT 93.880 42.200 94.080 49.800 ;
        RECT 95.380 50.200 95.580 57.800 ;
        RECT 96.180 50.200 96.380 57.800 ;
        RECT 96.980 50.200 97.180 57.800 ;
        RECT 97.780 50.200 97.980 57.800 ;
        RECT 98.580 50.200 98.780 57.800 ;
        RECT 99.530 57.600 103.530 57.800 ;
        RECT 103.130 57.000 103.530 57.600 ;
        RECT 99.530 56.800 103.530 57.000 ;
        RECT 103.130 56.200 103.530 56.800 ;
        RECT 99.530 56.000 103.530 56.200 ;
        RECT 103.130 55.400 103.530 56.000 ;
        RECT 99.530 55.200 103.530 55.400 ;
        RECT 103.130 54.600 103.530 55.200 ;
        RECT 99.530 54.400 103.530 54.600 ;
        RECT 103.130 53.800 103.530 54.400 ;
        RECT 99.530 53.600 103.530 53.800 ;
        RECT 103.130 53.000 103.530 53.600 ;
        RECT 99.530 52.800 103.530 53.000 ;
        RECT 103.130 52.200 103.530 52.800 ;
        RECT 99.530 52.000 103.530 52.200 ;
        RECT 103.130 51.400 103.530 52.000 ;
        RECT 99.530 51.200 103.530 51.400 ;
        RECT 103.130 50.600 103.530 51.200 ;
        RECT 99.530 50.400 103.530 50.600 ;
        RECT 103.130 50.200 103.530 50.400 ;
        RECT 95.380 49.800 103.530 50.200 ;
        RECT 95.380 42.200 95.580 49.800 ;
        RECT 96.180 42.200 96.380 49.800 ;
        RECT 96.980 42.200 97.180 49.800 ;
        RECT 97.780 42.200 97.980 49.800 ;
        RECT 98.580 42.200 98.780 49.800 ;
        RECT 103.130 49.600 103.530 49.800 ;
        RECT 99.530 49.400 103.530 49.600 ;
        RECT 103.130 48.800 103.530 49.400 ;
        RECT 99.530 48.600 103.530 48.800 ;
        RECT 103.130 48.000 103.530 48.600 ;
        RECT 99.530 47.800 103.530 48.000 ;
        RECT 103.130 47.200 103.530 47.800 ;
        RECT 99.530 47.000 103.530 47.200 ;
        RECT 103.130 46.400 103.530 47.000 ;
        RECT 99.530 46.200 103.530 46.400 ;
        RECT 103.130 45.600 103.530 46.200 ;
        RECT 99.530 45.400 103.530 45.600 ;
        RECT 103.130 44.800 103.530 45.400 ;
        RECT 99.530 44.600 103.530 44.800 ;
        RECT 103.130 44.000 103.530 44.600 ;
        RECT 99.530 43.800 103.530 44.000 ;
        RECT 103.130 43.200 103.530 43.800 ;
        RECT 99.530 43.000 103.530 43.200 ;
        RECT 103.130 42.400 103.530 43.000 ;
        RECT 99.530 42.200 103.530 42.400 ;
        RECT 105.930 57.600 109.930 57.800 ;
        RECT 105.930 57.000 106.330 57.600 ;
        RECT 105.930 56.800 109.930 57.000 ;
        RECT 105.930 56.200 106.330 56.800 ;
        RECT 105.930 56.000 109.930 56.200 ;
        RECT 105.930 55.400 106.330 56.000 ;
        RECT 105.930 55.200 109.930 55.400 ;
        RECT 105.930 54.600 106.330 55.200 ;
        RECT 105.930 54.400 109.930 54.600 ;
        RECT 105.930 53.800 106.330 54.400 ;
        RECT 105.930 53.600 109.930 53.800 ;
        RECT 105.930 53.000 106.330 53.600 ;
        RECT 105.930 52.800 109.930 53.000 ;
        RECT 105.930 52.200 106.330 52.800 ;
        RECT 105.930 52.000 109.930 52.200 ;
        RECT 105.930 51.400 106.330 52.000 ;
        RECT 105.930 51.200 109.930 51.400 ;
        RECT 105.930 50.600 106.330 51.200 ;
        RECT 105.930 50.400 109.930 50.600 ;
        RECT 105.930 50.200 106.330 50.400 ;
        RECT 110.680 50.200 110.880 57.800 ;
        RECT 111.480 50.200 111.680 57.800 ;
        RECT 112.280 50.200 112.480 57.800 ;
        RECT 113.080 50.200 113.280 57.800 ;
        RECT 113.880 50.200 114.080 57.800 ;
        RECT 105.930 49.800 114.080 50.200 ;
        RECT 105.930 49.600 106.330 49.800 ;
        RECT 105.930 49.400 109.930 49.600 ;
        RECT 105.930 48.800 106.330 49.400 ;
        RECT 105.930 48.600 109.930 48.800 ;
        RECT 105.930 48.000 106.330 48.600 ;
        RECT 105.930 47.800 109.930 48.000 ;
        RECT 105.930 47.200 106.330 47.800 ;
        RECT 105.930 47.000 109.930 47.200 ;
        RECT 105.930 46.400 106.330 47.000 ;
        RECT 105.930 46.200 109.930 46.400 ;
        RECT 105.930 45.600 106.330 46.200 ;
        RECT 105.930 45.400 109.930 45.600 ;
        RECT 105.930 44.800 106.330 45.400 ;
        RECT 105.930 44.600 109.930 44.800 ;
        RECT 105.930 44.000 106.330 44.600 ;
        RECT 105.930 43.800 109.930 44.000 ;
        RECT 105.930 43.200 106.330 43.800 ;
        RECT 105.930 43.000 109.930 43.200 ;
        RECT 105.930 42.400 106.330 43.000 ;
        RECT 105.930 42.200 109.930 42.400 ;
        RECT 110.680 42.200 110.880 49.800 ;
        RECT 111.480 42.200 111.680 49.800 ;
        RECT 112.280 42.200 112.480 49.800 ;
        RECT 113.080 42.200 113.280 49.800 ;
        RECT 113.880 42.200 114.080 49.800 ;
        RECT 115.380 50.200 115.580 57.800 ;
        RECT 116.180 50.200 116.380 57.800 ;
        RECT 116.980 50.200 117.180 57.800 ;
        RECT 117.780 50.200 117.980 57.800 ;
        RECT 118.580 50.200 118.780 57.800 ;
        RECT 119.530 57.600 123.530 57.800 ;
        RECT 123.130 57.000 123.530 57.600 ;
        RECT 119.530 56.800 123.530 57.000 ;
        RECT 123.130 56.200 123.530 56.800 ;
        RECT 119.530 56.000 123.530 56.200 ;
        RECT 123.130 55.400 123.530 56.000 ;
        RECT 119.530 55.200 123.530 55.400 ;
        RECT 123.130 54.600 123.530 55.200 ;
        RECT 119.530 54.400 123.530 54.600 ;
        RECT 123.130 53.800 123.530 54.400 ;
        RECT 119.530 53.600 123.530 53.800 ;
        RECT 123.130 53.000 123.530 53.600 ;
        RECT 119.530 52.800 123.530 53.000 ;
        RECT 123.130 52.200 123.530 52.800 ;
        RECT 119.530 52.000 123.530 52.200 ;
        RECT 123.130 51.400 123.530 52.000 ;
        RECT 119.530 51.200 123.530 51.400 ;
        RECT 123.130 50.600 123.530 51.200 ;
        RECT 130.050 50.900 130.410 51.280 ;
        RECT 130.680 50.900 131.040 51.280 ;
        RECT 131.280 50.900 131.640 51.280 ;
        RECT 119.530 50.400 123.530 50.600 ;
        RECT 123.130 50.200 123.530 50.400 ;
        RECT 130.050 50.310 130.410 50.690 ;
        RECT 130.680 50.310 131.040 50.690 ;
        RECT 131.280 50.310 131.640 50.690 ;
        RECT 115.380 49.800 123.530 50.200 ;
        RECT 115.380 42.200 115.580 49.800 ;
        RECT 116.180 42.200 116.380 49.800 ;
        RECT 116.980 42.200 117.180 49.800 ;
        RECT 117.780 42.200 117.980 49.800 ;
        RECT 118.580 42.200 118.780 49.800 ;
        RECT 123.130 49.600 123.530 49.800 ;
        RECT 119.530 49.400 123.530 49.600 ;
        RECT 123.130 48.800 123.530 49.400 ;
        RECT 119.530 48.600 123.530 48.800 ;
        RECT 123.130 48.000 123.530 48.600 ;
        RECT 119.530 47.800 123.530 48.000 ;
        RECT 123.130 47.200 123.530 47.800 ;
        RECT 119.530 47.000 123.530 47.200 ;
        RECT 123.130 46.400 123.530 47.000 ;
        RECT 119.530 46.200 123.530 46.400 ;
        RECT 123.130 45.600 123.530 46.200 ;
        RECT 119.530 45.400 123.530 45.600 ;
        RECT 123.130 44.800 123.530 45.400 ;
        RECT 119.530 44.600 123.530 44.800 ;
        RECT 123.130 44.000 123.530 44.600 ;
        RECT 119.530 43.800 123.530 44.000 ;
        RECT 123.130 43.200 123.530 43.800 ;
        RECT 119.530 43.000 123.530 43.200 ;
        RECT 123.130 42.400 123.530 43.000 ;
        RECT 119.530 42.200 123.530 42.400 ;
        RECT 5.930 37.600 9.930 37.800 ;
        RECT 5.930 37.000 6.330 37.600 ;
        RECT 5.930 36.800 9.930 37.000 ;
        RECT 5.930 36.200 6.330 36.800 ;
        RECT 5.930 36.000 9.930 36.200 ;
        RECT 5.930 35.400 6.330 36.000 ;
        RECT 5.930 35.200 9.930 35.400 ;
        RECT 5.930 34.600 6.330 35.200 ;
        RECT 5.930 34.400 9.930 34.600 ;
        RECT 5.930 33.800 6.330 34.400 ;
        RECT 5.930 33.600 9.930 33.800 ;
        RECT 5.930 33.000 6.330 33.600 ;
        RECT 5.930 32.800 9.930 33.000 ;
        RECT 5.930 32.200 6.330 32.800 ;
        RECT 5.930 32.000 9.930 32.200 ;
        RECT 5.930 31.400 6.330 32.000 ;
        RECT 5.930 31.200 9.930 31.400 ;
        RECT 5.930 30.600 6.330 31.200 ;
        RECT 5.930 30.400 9.930 30.600 ;
        RECT 5.930 30.200 6.330 30.400 ;
        RECT 10.680 30.200 10.880 37.800 ;
        RECT 11.480 30.200 11.680 37.800 ;
        RECT 12.280 30.200 12.480 37.800 ;
        RECT 13.080 30.200 13.280 37.800 ;
        RECT 13.880 30.200 14.080 37.800 ;
        RECT 5.930 29.800 14.080 30.200 ;
        RECT 5.930 29.600 6.330 29.800 ;
        RECT 5.930 29.400 9.930 29.600 ;
        RECT 5.930 28.800 6.330 29.400 ;
        RECT 5.930 28.600 9.930 28.800 ;
        RECT 5.930 28.000 6.330 28.600 ;
        RECT 5.930 27.800 9.930 28.000 ;
        RECT 5.930 27.200 6.330 27.800 ;
        RECT 5.930 27.000 9.930 27.200 ;
        RECT 5.930 26.400 6.330 27.000 ;
        RECT 5.930 26.200 9.930 26.400 ;
        RECT 5.930 25.600 6.330 26.200 ;
        RECT 5.930 25.400 9.930 25.600 ;
        RECT 5.930 24.800 6.330 25.400 ;
        RECT 5.930 24.600 9.930 24.800 ;
        RECT 5.930 24.000 6.330 24.600 ;
        RECT 5.930 23.800 9.930 24.000 ;
        RECT 5.930 23.200 6.330 23.800 ;
        RECT 5.930 23.000 9.930 23.200 ;
        RECT 5.930 22.400 6.330 23.000 ;
        RECT 5.930 22.200 9.930 22.400 ;
        RECT 10.680 22.200 10.880 29.800 ;
        RECT 11.480 22.200 11.680 29.800 ;
        RECT 12.280 22.200 12.480 29.800 ;
        RECT 13.080 22.200 13.280 29.800 ;
        RECT 13.880 22.200 14.080 29.800 ;
        RECT 15.380 30.200 15.580 37.800 ;
        RECT 16.180 30.200 16.380 37.800 ;
        RECT 16.980 30.200 17.180 37.800 ;
        RECT 17.780 30.200 17.980 37.800 ;
        RECT 18.580 30.200 18.780 37.800 ;
        RECT 19.530 37.600 23.530 37.800 ;
        RECT 23.130 37.000 23.530 37.600 ;
        RECT 19.530 36.800 23.530 37.000 ;
        RECT 23.130 36.200 23.530 36.800 ;
        RECT 19.530 36.000 23.530 36.200 ;
        RECT 23.130 35.400 23.530 36.000 ;
        RECT 19.530 35.200 23.530 35.400 ;
        RECT 23.130 34.600 23.530 35.200 ;
        RECT 19.530 34.400 23.530 34.600 ;
        RECT 23.130 33.800 23.530 34.400 ;
        RECT 19.530 33.600 23.530 33.800 ;
        RECT 23.130 33.000 23.530 33.600 ;
        RECT 19.530 32.800 23.530 33.000 ;
        RECT 23.130 32.200 23.530 32.800 ;
        RECT 19.530 32.000 23.530 32.200 ;
        RECT 23.130 31.400 23.530 32.000 ;
        RECT 19.530 31.200 23.530 31.400 ;
        RECT 23.130 30.600 23.530 31.200 ;
        RECT 19.530 30.400 23.530 30.600 ;
        RECT 23.130 30.200 23.530 30.400 ;
        RECT 15.380 29.800 23.530 30.200 ;
        RECT 15.380 22.200 15.580 29.800 ;
        RECT 16.180 22.200 16.380 29.800 ;
        RECT 16.980 22.200 17.180 29.800 ;
        RECT 17.780 22.200 17.980 29.800 ;
        RECT 18.580 22.200 18.780 29.800 ;
        RECT 23.130 29.600 23.530 29.800 ;
        RECT 19.530 29.400 23.530 29.600 ;
        RECT 23.130 28.800 23.530 29.400 ;
        RECT 19.530 28.600 23.530 28.800 ;
        RECT 23.130 28.000 23.530 28.600 ;
        RECT 19.530 27.800 23.530 28.000 ;
        RECT 23.130 27.200 23.530 27.800 ;
        RECT 19.530 27.000 23.530 27.200 ;
        RECT 23.130 26.400 23.530 27.000 ;
        RECT 19.530 26.200 23.530 26.400 ;
        RECT 23.130 25.600 23.530 26.200 ;
        RECT 19.530 25.400 23.530 25.600 ;
        RECT 23.130 24.800 23.530 25.400 ;
        RECT 19.530 24.600 23.530 24.800 ;
        RECT 23.130 24.000 23.530 24.600 ;
        RECT 19.530 23.800 23.530 24.000 ;
        RECT 23.130 23.200 23.530 23.800 ;
        RECT 19.530 23.000 23.530 23.200 ;
        RECT 23.130 22.400 23.530 23.000 ;
        RECT 19.530 22.200 23.530 22.400 ;
        RECT 25.930 37.600 29.930 37.800 ;
        RECT 25.930 37.000 26.330 37.600 ;
        RECT 25.930 36.800 29.930 37.000 ;
        RECT 25.930 36.200 26.330 36.800 ;
        RECT 25.930 36.000 29.930 36.200 ;
        RECT 25.930 35.400 26.330 36.000 ;
        RECT 25.930 35.200 29.930 35.400 ;
        RECT 25.930 34.600 26.330 35.200 ;
        RECT 25.930 34.400 29.930 34.600 ;
        RECT 25.930 33.800 26.330 34.400 ;
        RECT 25.930 33.600 29.930 33.800 ;
        RECT 25.930 33.000 26.330 33.600 ;
        RECT 25.930 32.800 29.930 33.000 ;
        RECT 25.930 32.200 26.330 32.800 ;
        RECT 25.930 32.000 29.930 32.200 ;
        RECT 25.930 31.400 26.330 32.000 ;
        RECT 25.930 31.200 29.930 31.400 ;
        RECT 25.930 30.600 26.330 31.200 ;
        RECT 25.930 30.400 29.930 30.600 ;
        RECT 25.930 30.200 26.330 30.400 ;
        RECT 30.680 30.200 30.880 37.800 ;
        RECT 31.480 30.200 31.680 37.800 ;
        RECT 32.280 30.200 32.480 37.800 ;
        RECT 33.080 30.200 33.280 37.800 ;
        RECT 33.880 30.200 34.080 37.800 ;
        RECT 25.930 29.800 34.080 30.200 ;
        RECT 25.930 29.600 26.330 29.800 ;
        RECT 25.930 29.400 29.930 29.600 ;
        RECT 25.930 28.800 26.330 29.400 ;
        RECT 25.930 28.600 29.930 28.800 ;
        RECT 25.930 28.000 26.330 28.600 ;
        RECT 25.930 27.800 29.930 28.000 ;
        RECT 25.930 27.200 26.330 27.800 ;
        RECT 25.930 27.000 29.930 27.200 ;
        RECT 25.930 26.400 26.330 27.000 ;
        RECT 25.930 26.200 29.930 26.400 ;
        RECT 25.930 25.600 26.330 26.200 ;
        RECT 25.930 25.400 29.930 25.600 ;
        RECT 25.930 24.800 26.330 25.400 ;
        RECT 25.930 24.600 29.930 24.800 ;
        RECT 25.930 24.000 26.330 24.600 ;
        RECT 25.930 23.800 29.930 24.000 ;
        RECT 25.930 23.200 26.330 23.800 ;
        RECT 25.930 23.000 29.930 23.200 ;
        RECT 25.930 22.400 26.330 23.000 ;
        RECT 25.930 22.200 29.930 22.400 ;
        RECT 30.680 22.200 30.880 29.800 ;
        RECT 31.480 22.200 31.680 29.800 ;
        RECT 32.280 22.200 32.480 29.800 ;
        RECT 33.080 22.200 33.280 29.800 ;
        RECT 33.880 22.200 34.080 29.800 ;
        RECT 35.380 30.200 35.580 37.800 ;
        RECT 36.180 30.200 36.380 37.800 ;
        RECT 36.980 30.200 37.180 37.800 ;
        RECT 37.780 30.200 37.980 37.800 ;
        RECT 38.580 30.200 38.780 37.800 ;
        RECT 39.530 37.600 43.530 37.800 ;
        RECT 43.130 37.000 43.530 37.600 ;
        RECT 39.530 36.800 43.530 37.000 ;
        RECT 43.130 36.200 43.530 36.800 ;
        RECT 39.530 36.000 43.530 36.200 ;
        RECT 43.130 35.400 43.530 36.000 ;
        RECT 39.530 35.200 43.530 35.400 ;
        RECT 43.130 34.600 43.530 35.200 ;
        RECT 39.530 34.400 43.530 34.600 ;
        RECT 43.130 33.800 43.530 34.400 ;
        RECT 39.530 33.600 43.530 33.800 ;
        RECT 43.130 33.000 43.530 33.600 ;
        RECT 39.530 32.800 43.530 33.000 ;
        RECT 43.130 32.200 43.530 32.800 ;
        RECT 39.530 32.000 43.530 32.200 ;
        RECT 43.130 31.400 43.530 32.000 ;
        RECT 39.530 31.200 43.530 31.400 ;
        RECT 43.130 30.600 43.530 31.200 ;
        RECT 39.530 30.400 43.530 30.600 ;
        RECT 43.130 30.200 43.530 30.400 ;
        RECT 35.380 29.800 43.530 30.200 ;
        RECT 35.380 22.200 35.580 29.800 ;
        RECT 36.180 22.200 36.380 29.800 ;
        RECT 36.980 22.200 37.180 29.800 ;
        RECT 37.780 22.200 37.980 29.800 ;
        RECT 38.580 22.200 38.780 29.800 ;
        RECT 43.130 29.600 43.530 29.800 ;
        RECT 39.530 29.400 43.530 29.600 ;
        RECT 43.130 28.800 43.530 29.400 ;
        RECT 39.530 28.600 43.530 28.800 ;
        RECT 43.130 28.000 43.530 28.600 ;
        RECT 39.530 27.800 43.530 28.000 ;
        RECT 43.130 27.200 43.530 27.800 ;
        RECT 39.530 27.000 43.530 27.200 ;
        RECT 43.130 26.400 43.530 27.000 ;
        RECT 39.530 26.200 43.530 26.400 ;
        RECT 43.130 25.600 43.530 26.200 ;
        RECT 39.530 25.400 43.530 25.600 ;
        RECT 43.130 24.800 43.530 25.400 ;
        RECT 39.530 24.600 43.530 24.800 ;
        RECT 43.130 24.000 43.530 24.600 ;
        RECT 39.530 23.800 43.530 24.000 ;
        RECT 43.130 23.200 43.530 23.800 ;
        RECT 39.530 23.000 43.530 23.200 ;
        RECT 43.130 22.400 43.530 23.000 ;
        RECT 39.530 22.200 43.530 22.400 ;
        RECT 45.930 37.600 49.930 37.800 ;
        RECT 45.930 37.000 46.330 37.600 ;
        RECT 45.930 36.800 49.930 37.000 ;
        RECT 45.930 36.200 46.330 36.800 ;
        RECT 45.930 36.000 49.930 36.200 ;
        RECT 45.930 35.400 46.330 36.000 ;
        RECT 45.930 35.200 49.930 35.400 ;
        RECT 45.930 34.600 46.330 35.200 ;
        RECT 45.930 34.400 49.930 34.600 ;
        RECT 45.930 33.800 46.330 34.400 ;
        RECT 45.930 33.600 49.930 33.800 ;
        RECT 45.930 33.000 46.330 33.600 ;
        RECT 45.930 32.800 49.930 33.000 ;
        RECT 45.930 32.200 46.330 32.800 ;
        RECT 45.930 32.000 49.930 32.200 ;
        RECT 45.930 31.400 46.330 32.000 ;
        RECT 45.930 31.200 49.930 31.400 ;
        RECT 45.930 30.600 46.330 31.200 ;
        RECT 45.930 30.400 49.930 30.600 ;
        RECT 45.930 30.200 46.330 30.400 ;
        RECT 50.680 30.200 50.880 37.800 ;
        RECT 51.480 30.200 51.680 37.800 ;
        RECT 52.280 30.200 52.480 37.800 ;
        RECT 53.080 30.200 53.280 37.800 ;
        RECT 53.880 30.200 54.080 37.800 ;
        RECT 45.930 29.800 54.080 30.200 ;
        RECT 45.930 29.600 46.330 29.800 ;
        RECT 45.930 29.400 49.930 29.600 ;
        RECT 45.930 28.800 46.330 29.400 ;
        RECT 45.930 28.600 49.930 28.800 ;
        RECT 45.930 28.000 46.330 28.600 ;
        RECT 45.930 27.800 49.930 28.000 ;
        RECT 45.930 27.200 46.330 27.800 ;
        RECT 45.930 27.000 49.930 27.200 ;
        RECT 45.930 26.400 46.330 27.000 ;
        RECT 45.930 26.200 49.930 26.400 ;
        RECT 45.930 25.600 46.330 26.200 ;
        RECT 45.930 25.400 49.930 25.600 ;
        RECT 45.930 24.800 46.330 25.400 ;
        RECT 45.930 24.600 49.930 24.800 ;
        RECT 45.930 24.000 46.330 24.600 ;
        RECT 45.930 23.800 49.930 24.000 ;
        RECT 45.930 23.200 46.330 23.800 ;
        RECT 45.930 23.000 49.930 23.200 ;
        RECT 45.930 22.400 46.330 23.000 ;
        RECT 45.930 22.200 49.930 22.400 ;
        RECT 50.680 22.200 50.880 29.800 ;
        RECT 51.480 22.200 51.680 29.800 ;
        RECT 52.280 22.200 52.480 29.800 ;
        RECT 53.080 22.200 53.280 29.800 ;
        RECT 53.880 22.200 54.080 29.800 ;
        RECT 55.380 30.200 55.580 37.800 ;
        RECT 56.180 30.200 56.380 37.800 ;
        RECT 56.980 30.200 57.180 37.800 ;
        RECT 57.780 30.200 57.980 37.800 ;
        RECT 58.580 30.200 58.780 37.800 ;
        RECT 59.530 37.600 63.530 37.800 ;
        RECT 63.130 37.000 63.530 37.600 ;
        RECT 59.530 36.800 63.530 37.000 ;
        RECT 63.130 36.200 63.530 36.800 ;
        RECT 59.530 36.000 63.530 36.200 ;
        RECT 63.130 35.400 63.530 36.000 ;
        RECT 59.530 35.200 63.530 35.400 ;
        RECT 63.130 34.600 63.530 35.200 ;
        RECT 59.530 34.400 63.530 34.600 ;
        RECT 63.130 33.800 63.530 34.400 ;
        RECT 59.530 33.600 63.530 33.800 ;
        RECT 63.130 33.000 63.530 33.600 ;
        RECT 59.530 32.800 63.530 33.000 ;
        RECT 63.130 32.200 63.530 32.800 ;
        RECT 59.530 32.000 63.530 32.200 ;
        RECT 63.130 31.400 63.530 32.000 ;
        RECT 59.530 31.200 63.530 31.400 ;
        RECT 63.130 30.600 63.530 31.200 ;
        RECT 59.530 30.400 63.530 30.600 ;
        RECT 63.130 30.200 63.530 30.400 ;
        RECT 55.380 29.800 63.530 30.200 ;
        RECT 55.380 22.200 55.580 29.800 ;
        RECT 56.180 22.200 56.380 29.800 ;
        RECT 56.980 22.200 57.180 29.800 ;
        RECT 57.780 22.200 57.980 29.800 ;
        RECT 58.580 22.200 58.780 29.800 ;
        RECT 63.130 29.600 63.530 29.800 ;
        RECT 59.530 29.400 63.530 29.600 ;
        RECT 63.130 28.800 63.530 29.400 ;
        RECT 59.530 28.600 63.530 28.800 ;
        RECT 63.130 28.000 63.530 28.600 ;
        RECT 59.530 27.800 63.530 28.000 ;
        RECT 63.130 27.200 63.530 27.800 ;
        RECT 59.530 27.000 63.530 27.200 ;
        RECT 63.130 26.400 63.530 27.000 ;
        RECT 59.530 26.200 63.530 26.400 ;
        RECT 63.130 25.600 63.530 26.200 ;
        RECT 59.530 25.400 63.530 25.600 ;
        RECT 63.130 24.800 63.530 25.400 ;
        RECT 59.530 24.600 63.530 24.800 ;
        RECT 63.130 24.000 63.530 24.600 ;
        RECT 59.530 23.800 63.530 24.000 ;
        RECT 63.130 23.200 63.530 23.800 ;
        RECT 59.530 23.000 63.530 23.200 ;
        RECT 63.130 22.400 63.530 23.000 ;
        RECT 59.530 22.200 63.530 22.400 ;
        RECT 65.930 37.600 69.930 37.800 ;
        RECT 65.930 37.000 66.330 37.600 ;
        RECT 65.930 36.800 69.930 37.000 ;
        RECT 65.930 36.200 66.330 36.800 ;
        RECT 65.930 36.000 69.930 36.200 ;
        RECT 65.930 35.400 66.330 36.000 ;
        RECT 65.930 35.200 69.930 35.400 ;
        RECT 65.930 34.600 66.330 35.200 ;
        RECT 65.930 34.400 69.930 34.600 ;
        RECT 65.930 33.800 66.330 34.400 ;
        RECT 65.930 33.600 69.930 33.800 ;
        RECT 65.930 33.000 66.330 33.600 ;
        RECT 65.930 32.800 69.930 33.000 ;
        RECT 65.930 32.200 66.330 32.800 ;
        RECT 65.930 32.000 69.930 32.200 ;
        RECT 65.930 31.400 66.330 32.000 ;
        RECT 65.930 31.200 69.930 31.400 ;
        RECT 65.930 30.600 66.330 31.200 ;
        RECT 65.930 30.400 69.930 30.600 ;
        RECT 65.930 30.200 66.330 30.400 ;
        RECT 70.680 30.200 70.880 37.800 ;
        RECT 71.480 30.200 71.680 37.800 ;
        RECT 72.280 30.200 72.480 37.800 ;
        RECT 73.080 30.200 73.280 37.800 ;
        RECT 73.880 30.200 74.080 37.800 ;
        RECT 65.930 29.800 74.080 30.200 ;
        RECT 65.930 29.600 66.330 29.800 ;
        RECT 65.930 29.400 69.930 29.600 ;
        RECT 65.930 28.800 66.330 29.400 ;
        RECT 65.930 28.600 69.930 28.800 ;
        RECT 65.930 28.000 66.330 28.600 ;
        RECT 65.930 27.800 69.930 28.000 ;
        RECT 65.930 27.200 66.330 27.800 ;
        RECT 65.930 27.000 69.930 27.200 ;
        RECT 65.930 26.400 66.330 27.000 ;
        RECT 65.930 26.200 69.930 26.400 ;
        RECT 65.930 25.600 66.330 26.200 ;
        RECT 65.930 25.400 69.930 25.600 ;
        RECT 65.930 24.800 66.330 25.400 ;
        RECT 65.930 24.600 69.930 24.800 ;
        RECT 65.930 24.000 66.330 24.600 ;
        RECT 65.930 23.800 69.930 24.000 ;
        RECT 65.930 23.200 66.330 23.800 ;
        RECT 65.930 23.000 69.930 23.200 ;
        RECT 65.930 22.400 66.330 23.000 ;
        RECT 65.930 22.200 69.930 22.400 ;
        RECT 70.680 22.200 70.880 29.800 ;
        RECT 71.480 22.200 71.680 29.800 ;
        RECT 72.280 22.200 72.480 29.800 ;
        RECT 73.080 22.200 73.280 29.800 ;
        RECT 73.880 22.200 74.080 29.800 ;
        RECT 75.380 30.200 75.580 37.800 ;
        RECT 76.180 30.200 76.380 37.800 ;
        RECT 76.980 30.200 77.180 37.800 ;
        RECT 77.780 30.200 77.980 37.800 ;
        RECT 78.580 30.200 78.780 37.800 ;
        RECT 79.530 37.600 83.530 37.800 ;
        RECT 83.130 37.000 83.530 37.600 ;
        RECT 79.530 36.800 83.530 37.000 ;
        RECT 83.130 36.200 83.530 36.800 ;
        RECT 79.530 36.000 83.530 36.200 ;
        RECT 83.130 35.400 83.530 36.000 ;
        RECT 79.530 35.200 83.530 35.400 ;
        RECT 83.130 34.600 83.530 35.200 ;
        RECT 79.530 34.400 83.530 34.600 ;
        RECT 83.130 33.800 83.530 34.400 ;
        RECT 79.530 33.600 83.530 33.800 ;
        RECT 83.130 33.000 83.530 33.600 ;
        RECT 79.530 32.800 83.530 33.000 ;
        RECT 83.130 32.200 83.530 32.800 ;
        RECT 79.530 32.000 83.530 32.200 ;
        RECT 83.130 31.400 83.530 32.000 ;
        RECT 79.530 31.200 83.530 31.400 ;
        RECT 83.130 30.600 83.530 31.200 ;
        RECT 79.530 30.400 83.530 30.600 ;
        RECT 83.130 30.200 83.530 30.400 ;
        RECT 75.380 29.800 83.530 30.200 ;
        RECT 75.380 22.200 75.580 29.800 ;
        RECT 76.180 22.200 76.380 29.800 ;
        RECT 76.980 22.200 77.180 29.800 ;
        RECT 77.780 22.200 77.980 29.800 ;
        RECT 78.580 22.200 78.780 29.800 ;
        RECT 83.130 29.600 83.530 29.800 ;
        RECT 79.530 29.400 83.530 29.600 ;
        RECT 83.130 28.800 83.530 29.400 ;
        RECT 79.530 28.600 83.530 28.800 ;
        RECT 83.130 28.000 83.530 28.600 ;
        RECT 79.530 27.800 83.530 28.000 ;
        RECT 83.130 27.200 83.530 27.800 ;
        RECT 79.530 27.000 83.530 27.200 ;
        RECT 83.130 26.400 83.530 27.000 ;
        RECT 79.530 26.200 83.530 26.400 ;
        RECT 83.130 25.600 83.530 26.200 ;
        RECT 79.530 25.400 83.530 25.600 ;
        RECT 83.130 24.800 83.530 25.400 ;
        RECT 79.530 24.600 83.530 24.800 ;
        RECT 83.130 24.000 83.530 24.600 ;
        RECT 79.530 23.800 83.530 24.000 ;
        RECT 83.130 23.200 83.530 23.800 ;
        RECT 79.530 23.000 83.530 23.200 ;
        RECT 83.130 22.400 83.530 23.000 ;
        RECT 79.530 22.200 83.530 22.400 ;
        RECT 85.930 37.600 89.930 37.800 ;
        RECT 85.930 37.000 86.330 37.600 ;
        RECT 85.930 36.800 89.930 37.000 ;
        RECT 85.930 36.200 86.330 36.800 ;
        RECT 85.930 36.000 89.930 36.200 ;
        RECT 85.930 35.400 86.330 36.000 ;
        RECT 85.930 35.200 89.930 35.400 ;
        RECT 85.930 34.600 86.330 35.200 ;
        RECT 85.930 34.400 89.930 34.600 ;
        RECT 85.930 33.800 86.330 34.400 ;
        RECT 85.930 33.600 89.930 33.800 ;
        RECT 85.930 33.000 86.330 33.600 ;
        RECT 85.930 32.800 89.930 33.000 ;
        RECT 85.930 32.200 86.330 32.800 ;
        RECT 85.930 32.000 89.930 32.200 ;
        RECT 85.930 31.400 86.330 32.000 ;
        RECT 85.930 31.200 89.930 31.400 ;
        RECT 85.930 30.600 86.330 31.200 ;
        RECT 85.930 30.400 89.930 30.600 ;
        RECT 85.930 30.200 86.330 30.400 ;
        RECT 90.680 30.200 90.880 37.800 ;
        RECT 91.480 30.200 91.680 37.800 ;
        RECT 92.280 30.200 92.480 37.800 ;
        RECT 93.080 30.200 93.280 37.800 ;
        RECT 93.880 30.200 94.080 37.800 ;
        RECT 85.930 29.800 94.080 30.200 ;
        RECT 85.930 29.600 86.330 29.800 ;
        RECT 85.930 29.400 89.930 29.600 ;
        RECT 85.930 28.800 86.330 29.400 ;
        RECT 85.930 28.600 89.930 28.800 ;
        RECT 85.930 28.000 86.330 28.600 ;
        RECT 85.930 27.800 89.930 28.000 ;
        RECT 85.930 27.200 86.330 27.800 ;
        RECT 85.930 27.000 89.930 27.200 ;
        RECT 85.930 26.400 86.330 27.000 ;
        RECT 85.930 26.200 89.930 26.400 ;
        RECT 85.930 25.600 86.330 26.200 ;
        RECT 85.930 25.400 89.930 25.600 ;
        RECT 85.930 24.800 86.330 25.400 ;
        RECT 85.930 24.600 89.930 24.800 ;
        RECT 85.930 24.000 86.330 24.600 ;
        RECT 85.930 23.800 89.930 24.000 ;
        RECT 85.930 23.200 86.330 23.800 ;
        RECT 85.930 23.000 89.930 23.200 ;
        RECT 85.930 22.400 86.330 23.000 ;
        RECT 85.930 22.200 89.930 22.400 ;
        RECT 90.680 22.200 90.880 29.800 ;
        RECT 91.480 22.200 91.680 29.800 ;
        RECT 92.280 22.200 92.480 29.800 ;
        RECT 93.080 22.200 93.280 29.800 ;
        RECT 93.880 22.200 94.080 29.800 ;
        RECT 95.380 30.200 95.580 37.800 ;
        RECT 96.180 30.200 96.380 37.800 ;
        RECT 96.980 30.200 97.180 37.800 ;
        RECT 97.780 30.200 97.980 37.800 ;
        RECT 98.580 30.200 98.780 37.800 ;
        RECT 99.530 37.600 103.530 37.800 ;
        RECT 103.130 37.000 103.530 37.600 ;
        RECT 99.530 36.800 103.530 37.000 ;
        RECT 103.130 36.200 103.530 36.800 ;
        RECT 99.530 36.000 103.530 36.200 ;
        RECT 103.130 35.400 103.530 36.000 ;
        RECT 99.530 35.200 103.530 35.400 ;
        RECT 103.130 34.600 103.530 35.200 ;
        RECT 99.530 34.400 103.530 34.600 ;
        RECT 103.130 33.800 103.530 34.400 ;
        RECT 99.530 33.600 103.530 33.800 ;
        RECT 103.130 33.000 103.530 33.600 ;
        RECT 99.530 32.800 103.530 33.000 ;
        RECT 103.130 32.200 103.530 32.800 ;
        RECT 99.530 32.000 103.530 32.200 ;
        RECT 103.130 31.400 103.530 32.000 ;
        RECT 99.530 31.200 103.530 31.400 ;
        RECT 103.130 30.600 103.530 31.200 ;
        RECT 99.530 30.400 103.530 30.600 ;
        RECT 103.130 30.200 103.530 30.400 ;
        RECT 95.380 29.800 103.530 30.200 ;
        RECT 95.380 22.200 95.580 29.800 ;
        RECT 96.180 22.200 96.380 29.800 ;
        RECT 96.980 22.200 97.180 29.800 ;
        RECT 97.780 22.200 97.980 29.800 ;
        RECT 98.580 22.200 98.780 29.800 ;
        RECT 103.130 29.600 103.530 29.800 ;
        RECT 99.530 29.400 103.530 29.600 ;
        RECT 103.130 28.800 103.530 29.400 ;
        RECT 99.530 28.600 103.530 28.800 ;
        RECT 103.130 28.000 103.530 28.600 ;
        RECT 99.530 27.800 103.530 28.000 ;
        RECT 103.130 27.200 103.530 27.800 ;
        RECT 99.530 27.000 103.530 27.200 ;
        RECT 103.130 26.400 103.530 27.000 ;
        RECT 99.530 26.200 103.530 26.400 ;
        RECT 103.130 25.600 103.530 26.200 ;
        RECT 99.530 25.400 103.530 25.600 ;
        RECT 103.130 24.800 103.530 25.400 ;
        RECT 99.530 24.600 103.530 24.800 ;
        RECT 103.130 24.000 103.530 24.600 ;
        RECT 99.530 23.800 103.530 24.000 ;
        RECT 103.130 23.200 103.530 23.800 ;
        RECT 99.530 23.000 103.530 23.200 ;
        RECT 103.130 22.400 103.530 23.000 ;
        RECT 99.530 22.200 103.530 22.400 ;
        RECT 105.930 37.600 109.930 37.800 ;
        RECT 105.930 37.000 106.330 37.600 ;
        RECT 105.930 36.800 109.930 37.000 ;
        RECT 105.930 36.200 106.330 36.800 ;
        RECT 105.930 36.000 109.930 36.200 ;
        RECT 105.930 35.400 106.330 36.000 ;
        RECT 105.930 35.200 109.930 35.400 ;
        RECT 105.930 34.600 106.330 35.200 ;
        RECT 105.930 34.400 109.930 34.600 ;
        RECT 105.930 33.800 106.330 34.400 ;
        RECT 105.930 33.600 109.930 33.800 ;
        RECT 105.930 33.000 106.330 33.600 ;
        RECT 105.930 32.800 109.930 33.000 ;
        RECT 105.930 32.200 106.330 32.800 ;
        RECT 105.930 32.000 109.930 32.200 ;
        RECT 105.930 31.400 106.330 32.000 ;
        RECT 105.930 31.200 109.930 31.400 ;
        RECT 105.930 30.600 106.330 31.200 ;
        RECT 105.930 30.400 109.930 30.600 ;
        RECT 105.930 30.200 106.330 30.400 ;
        RECT 110.680 30.200 110.880 37.800 ;
        RECT 111.480 30.200 111.680 37.800 ;
        RECT 112.280 30.200 112.480 37.800 ;
        RECT 113.080 30.200 113.280 37.800 ;
        RECT 113.880 30.200 114.080 37.800 ;
        RECT 105.930 29.800 114.080 30.200 ;
        RECT 105.930 29.600 106.330 29.800 ;
        RECT 105.930 29.400 109.930 29.600 ;
        RECT 105.930 28.800 106.330 29.400 ;
        RECT 105.930 28.600 109.930 28.800 ;
        RECT 105.930 28.000 106.330 28.600 ;
        RECT 105.930 27.800 109.930 28.000 ;
        RECT 105.930 27.200 106.330 27.800 ;
        RECT 105.930 27.000 109.930 27.200 ;
        RECT 105.930 26.400 106.330 27.000 ;
        RECT 105.930 26.200 109.930 26.400 ;
        RECT 105.930 25.600 106.330 26.200 ;
        RECT 105.930 25.400 109.930 25.600 ;
        RECT 105.930 24.800 106.330 25.400 ;
        RECT 105.930 24.600 109.930 24.800 ;
        RECT 105.930 24.000 106.330 24.600 ;
        RECT 105.930 23.800 109.930 24.000 ;
        RECT 105.930 23.200 106.330 23.800 ;
        RECT 105.930 23.000 109.930 23.200 ;
        RECT 105.930 22.400 106.330 23.000 ;
        RECT 105.930 22.200 109.930 22.400 ;
        RECT 110.680 22.200 110.880 29.800 ;
        RECT 111.480 22.200 111.680 29.800 ;
        RECT 112.280 22.200 112.480 29.800 ;
        RECT 113.080 22.200 113.280 29.800 ;
        RECT 113.880 22.200 114.080 29.800 ;
        RECT 115.380 30.200 115.580 37.800 ;
        RECT 116.180 30.200 116.380 37.800 ;
        RECT 116.980 30.200 117.180 37.800 ;
        RECT 117.780 30.200 117.980 37.800 ;
        RECT 118.580 30.200 118.780 37.800 ;
        RECT 119.530 37.600 123.530 37.800 ;
        RECT 123.130 37.000 123.530 37.600 ;
        RECT 119.530 36.800 123.530 37.000 ;
        RECT 123.130 36.200 123.530 36.800 ;
        RECT 119.530 36.000 123.530 36.200 ;
        RECT 123.130 35.400 123.530 36.000 ;
        RECT 119.530 35.200 123.530 35.400 ;
        RECT 123.130 34.600 123.530 35.200 ;
        RECT 119.530 34.400 123.530 34.600 ;
        RECT 123.130 33.800 123.530 34.400 ;
        RECT 119.530 33.600 123.530 33.800 ;
        RECT 123.130 33.000 123.530 33.600 ;
        RECT 119.530 32.800 123.530 33.000 ;
        RECT 123.130 32.200 123.530 32.800 ;
        RECT 119.530 32.000 123.530 32.200 ;
        RECT 123.130 31.400 123.530 32.000 ;
        RECT 119.530 31.200 123.530 31.400 ;
        RECT 123.130 30.600 123.530 31.200 ;
        RECT 130.050 31.080 130.410 31.460 ;
        RECT 130.680 31.080 131.040 31.460 ;
        RECT 131.280 31.080 131.640 31.460 ;
        RECT 119.530 30.400 123.530 30.600 ;
        RECT 130.050 30.490 130.410 30.870 ;
        RECT 130.680 30.490 131.040 30.870 ;
        RECT 131.280 30.490 131.640 30.870 ;
        RECT 123.130 30.200 123.530 30.400 ;
        RECT 115.380 29.800 123.530 30.200 ;
        RECT 115.380 22.200 115.580 29.800 ;
        RECT 116.180 22.200 116.380 29.800 ;
        RECT 116.980 22.200 117.180 29.800 ;
        RECT 117.780 22.200 117.980 29.800 ;
        RECT 118.580 22.200 118.780 29.800 ;
        RECT 123.130 29.600 123.530 29.800 ;
        RECT 119.530 29.400 123.530 29.600 ;
        RECT 123.130 28.800 123.530 29.400 ;
        RECT 119.530 28.600 123.530 28.800 ;
        RECT 123.130 28.000 123.530 28.600 ;
        RECT 119.530 27.800 123.530 28.000 ;
        RECT 123.130 27.200 123.530 27.800 ;
        RECT 119.530 27.000 123.530 27.200 ;
        RECT 123.130 26.400 123.530 27.000 ;
        RECT 119.530 26.200 123.530 26.400 ;
        RECT 123.130 25.600 123.530 26.200 ;
        RECT 119.530 25.400 123.530 25.600 ;
        RECT 123.130 24.800 123.530 25.400 ;
        RECT 119.530 24.600 123.530 24.800 ;
        RECT 123.130 24.000 123.530 24.600 ;
        RECT 119.530 23.800 123.530 24.000 ;
        RECT 123.130 23.200 123.530 23.800 ;
        RECT 119.530 23.000 123.530 23.200 ;
        RECT 123.130 22.400 123.530 23.000 ;
        RECT 119.530 22.200 123.530 22.400 ;
        RECT 5.930 17.600 9.930 17.800 ;
        RECT 5.930 17.000 6.330 17.600 ;
        RECT 5.930 16.800 9.930 17.000 ;
        RECT 5.930 16.200 6.330 16.800 ;
        RECT 5.930 16.000 9.930 16.200 ;
        RECT 5.930 15.400 6.330 16.000 ;
        RECT 5.930 15.200 9.930 15.400 ;
        RECT 5.930 14.600 6.330 15.200 ;
        RECT 5.930 14.400 9.930 14.600 ;
        RECT 5.930 13.800 6.330 14.400 ;
        RECT 5.930 13.600 9.930 13.800 ;
        RECT 5.930 13.000 6.330 13.600 ;
        RECT 5.930 12.800 9.930 13.000 ;
        RECT 5.930 12.200 6.330 12.800 ;
        RECT 5.930 12.000 9.930 12.200 ;
        RECT 5.930 11.400 6.330 12.000 ;
        RECT 5.930 11.200 9.930 11.400 ;
        RECT 5.930 10.600 6.330 11.200 ;
        RECT 5.930 10.400 9.930 10.600 ;
        RECT 5.930 10.200 6.330 10.400 ;
        RECT 10.680 10.200 10.880 17.800 ;
        RECT 11.480 10.200 11.680 17.800 ;
        RECT 12.280 10.200 12.480 17.800 ;
        RECT 13.080 10.200 13.280 17.800 ;
        RECT 13.880 10.200 14.080 17.800 ;
        RECT 5.930 9.800 14.080 10.200 ;
        RECT 5.930 9.600 6.330 9.800 ;
        RECT 5.930 9.400 9.930 9.600 ;
        RECT 5.930 8.800 6.330 9.400 ;
        RECT 5.930 8.600 9.930 8.800 ;
        RECT 5.930 8.000 6.330 8.600 ;
        RECT 5.930 7.800 9.930 8.000 ;
        RECT 5.930 7.200 6.330 7.800 ;
        RECT 5.930 7.000 9.930 7.200 ;
        RECT 5.930 6.400 6.330 7.000 ;
        RECT 5.930 6.200 9.930 6.400 ;
        RECT 5.930 5.600 6.330 6.200 ;
        RECT 5.930 5.400 9.930 5.600 ;
        RECT 5.930 4.800 6.330 5.400 ;
        RECT 5.930 4.600 9.930 4.800 ;
        RECT 5.930 4.000 6.330 4.600 ;
        RECT 5.930 3.800 9.930 4.000 ;
        RECT 5.930 3.200 6.330 3.800 ;
        RECT 5.930 3.000 9.930 3.200 ;
        RECT 5.930 2.400 6.330 3.000 ;
        RECT 5.930 2.200 9.930 2.400 ;
        RECT 10.680 2.200 10.880 9.800 ;
        RECT 11.480 2.200 11.680 9.800 ;
        RECT 12.280 2.200 12.480 9.800 ;
        RECT 13.080 2.200 13.280 9.800 ;
        RECT 13.880 2.200 14.080 9.800 ;
        RECT 15.380 10.200 15.580 17.800 ;
        RECT 16.180 10.200 16.380 17.800 ;
        RECT 16.980 10.200 17.180 17.800 ;
        RECT 17.780 10.200 17.980 17.800 ;
        RECT 18.580 10.200 18.780 17.800 ;
        RECT 19.530 17.600 23.530 17.800 ;
        RECT 23.130 17.000 23.530 17.600 ;
        RECT 19.530 16.800 23.530 17.000 ;
        RECT 23.130 16.200 23.530 16.800 ;
        RECT 19.530 16.000 23.530 16.200 ;
        RECT 23.130 15.400 23.530 16.000 ;
        RECT 19.530 15.200 23.530 15.400 ;
        RECT 23.130 14.600 23.530 15.200 ;
        RECT 19.530 14.400 23.530 14.600 ;
        RECT 23.130 13.800 23.530 14.400 ;
        RECT 19.530 13.600 23.530 13.800 ;
        RECT 23.130 13.000 23.530 13.600 ;
        RECT 19.530 12.800 23.530 13.000 ;
        RECT 23.130 12.200 23.530 12.800 ;
        RECT 19.530 12.000 23.530 12.200 ;
        RECT 23.130 11.400 23.530 12.000 ;
        RECT 19.530 11.200 23.530 11.400 ;
        RECT 23.130 10.600 23.530 11.200 ;
        RECT 19.530 10.400 23.530 10.600 ;
        RECT 23.130 10.200 23.530 10.400 ;
        RECT 15.380 9.800 23.530 10.200 ;
        RECT 15.380 2.200 15.580 9.800 ;
        RECT 16.180 2.200 16.380 9.800 ;
        RECT 16.980 2.200 17.180 9.800 ;
        RECT 17.780 2.200 17.980 9.800 ;
        RECT 18.580 2.200 18.780 9.800 ;
        RECT 23.130 9.600 23.530 9.800 ;
        RECT 19.530 9.400 23.530 9.600 ;
        RECT 23.130 8.800 23.530 9.400 ;
        RECT 19.530 8.600 23.530 8.800 ;
        RECT 23.130 8.000 23.530 8.600 ;
        RECT 19.530 7.800 23.530 8.000 ;
        RECT 23.130 7.200 23.530 7.800 ;
        RECT 19.530 7.000 23.530 7.200 ;
        RECT 23.130 6.400 23.530 7.000 ;
        RECT 19.530 6.200 23.530 6.400 ;
        RECT 23.130 5.600 23.530 6.200 ;
        RECT 19.530 5.400 23.530 5.600 ;
        RECT 23.130 4.800 23.530 5.400 ;
        RECT 19.530 4.600 23.530 4.800 ;
        RECT 23.130 4.000 23.530 4.600 ;
        RECT 19.530 3.800 23.530 4.000 ;
        RECT 23.130 3.200 23.530 3.800 ;
        RECT 19.530 3.000 23.530 3.200 ;
        RECT 23.130 2.400 23.530 3.000 ;
        RECT 19.530 2.200 23.530 2.400 ;
        RECT 25.930 17.600 29.930 17.800 ;
        RECT 25.930 17.000 26.330 17.600 ;
        RECT 25.930 16.800 29.930 17.000 ;
        RECT 25.930 16.200 26.330 16.800 ;
        RECT 25.930 16.000 29.930 16.200 ;
        RECT 25.930 15.400 26.330 16.000 ;
        RECT 25.930 15.200 29.930 15.400 ;
        RECT 25.930 14.600 26.330 15.200 ;
        RECT 25.930 14.400 29.930 14.600 ;
        RECT 25.930 13.800 26.330 14.400 ;
        RECT 25.930 13.600 29.930 13.800 ;
        RECT 25.930 13.000 26.330 13.600 ;
        RECT 25.930 12.800 29.930 13.000 ;
        RECT 25.930 12.200 26.330 12.800 ;
        RECT 25.930 12.000 29.930 12.200 ;
        RECT 25.930 11.400 26.330 12.000 ;
        RECT 25.930 11.200 29.930 11.400 ;
        RECT 25.930 10.600 26.330 11.200 ;
        RECT 25.930 10.400 29.930 10.600 ;
        RECT 25.930 10.200 26.330 10.400 ;
        RECT 30.680 10.200 30.880 17.800 ;
        RECT 31.480 10.200 31.680 17.800 ;
        RECT 32.280 10.200 32.480 17.800 ;
        RECT 33.080 10.200 33.280 17.800 ;
        RECT 33.880 10.200 34.080 17.800 ;
        RECT 25.930 9.800 34.080 10.200 ;
        RECT 25.930 9.600 26.330 9.800 ;
        RECT 25.930 9.400 29.930 9.600 ;
        RECT 25.930 8.800 26.330 9.400 ;
        RECT 25.930 8.600 29.930 8.800 ;
        RECT 25.930 8.000 26.330 8.600 ;
        RECT 25.930 7.800 29.930 8.000 ;
        RECT 25.930 7.200 26.330 7.800 ;
        RECT 25.930 7.000 29.930 7.200 ;
        RECT 25.930 6.400 26.330 7.000 ;
        RECT 25.930 6.200 29.930 6.400 ;
        RECT 25.930 5.600 26.330 6.200 ;
        RECT 25.930 5.400 29.930 5.600 ;
        RECT 25.930 4.800 26.330 5.400 ;
        RECT 25.930 4.600 29.930 4.800 ;
        RECT 25.930 4.000 26.330 4.600 ;
        RECT 25.930 3.800 29.930 4.000 ;
        RECT 25.930 3.200 26.330 3.800 ;
        RECT 25.930 3.000 29.930 3.200 ;
        RECT 25.930 2.400 26.330 3.000 ;
        RECT 25.930 2.200 29.930 2.400 ;
        RECT 30.680 2.200 30.880 9.800 ;
        RECT 31.480 2.200 31.680 9.800 ;
        RECT 32.280 2.200 32.480 9.800 ;
        RECT 33.080 2.200 33.280 9.800 ;
        RECT 33.880 2.200 34.080 9.800 ;
        RECT 35.380 10.200 35.580 17.800 ;
        RECT 36.180 10.200 36.380 17.800 ;
        RECT 36.980 10.200 37.180 17.800 ;
        RECT 37.780 10.200 37.980 17.800 ;
        RECT 38.580 10.200 38.780 17.800 ;
        RECT 39.530 17.600 43.530 17.800 ;
        RECT 43.130 17.000 43.530 17.600 ;
        RECT 39.530 16.800 43.530 17.000 ;
        RECT 43.130 16.200 43.530 16.800 ;
        RECT 39.530 16.000 43.530 16.200 ;
        RECT 43.130 15.400 43.530 16.000 ;
        RECT 39.530 15.200 43.530 15.400 ;
        RECT 43.130 14.600 43.530 15.200 ;
        RECT 39.530 14.400 43.530 14.600 ;
        RECT 43.130 13.800 43.530 14.400 ;
        RECT 39.530 13.600 43.530 13.800 ;
        RECT 43.130 13.000 43.530 13.600 ;
        RECT 39.530 12.800 43.530 13.000 ;
        RECT 43.130 12.200 43.530 12.800 ;
        RECT 39.530 12.000 43.530 12.200 ;
        RECT 43.130 11.400 43.530 12.000 ;
        RECT 39.530 11.200 43.530 11.400 ;
        RECT 43.130 10.600 43.530 11.200 ;
        RECT 39.530 10.400 43.530 10.600 ;
        RECT 43.130 10.200 43.530 10.400 ;
        RECT 35.380 9.800 43.530 10.200 ;
        RECT 35.380 2.200 35.580 9.800 ;
        RECT 36.180 2.200 36.380 9.800 ;
        RECT 36.980 2.200 37.180 9.800 ;
        RECT 37.780 2.200 37.980 9.800 ;
        RECT 38.580 2.200 38.780 9.800 ;
        RECT 43.130 9.600 43.530 9.800 ;
        RECT 39.530 9.400 43.530 9.600 ;
        RECT 43.130 8.800 43.530 9.400 ;
        RECT 39.530 8.600 43.530 8.800 ;
        RECT 43.130 8.000 43.530 8.600 ;
        RECT 39.530 7.800 43.530 8.000 ;
        RECT 43.130 7.200 43.530 7.800 ;
        RECT 39.530 7.000 43.530 7.200 ;
        RECT 43.130 6.400 43.530 7.000 ;
        RECT 39.530 6.200 43.530 6.400 ;
        RECT 43.130 5.600 43.530 6.200 ;
        RECT 39.530 5.400 43.530 5.600 ;
        RECT 43.130 4.800 43.530 5.400 ;
        RECT 39.530 4.600 43.530 4.800 ;
        RECT 43.130 4.000 43.530 4.600 ;
        RECT 39.530 3.800 43.530 4.000 ;
        RECT 43.130 3.200 43.530 3.800 ;
        RECT 39.530 3.000 43.530 3.200 ;
        RECT 43.130 2.400 43.530 3.000 ;
        RECT 39.530 2.200 43.530 2.400 ;
        RECT 45.930 17.600 49.930 17.800 ;
        RECT 45.930 17.000 46.330 17.600 ;
        RECT 45.930 16.800 49.930 17.000 ;
        RECT 45.930 16.200 46.330 16.800 ;
        RECT 45.930 16.000 49.930 16.200 ;
        RECT 45.930 15.400 46.330 16.000 ;
        RECT 45.930 15.200 49.930 15.400 ;
        RECT 45.930 14.600 46.330 15.200 ;
        RECT 45.930 14.400 49.930 14.600 ;
        RECT 45.930 13.800 46.330 14.400 ;
        RECT 45.930 13.600 49.930 13.800 ;
        RECT 45.930 13.000 46.330 13.600 ;
        RECT 45.930 12.800 49.930 13.000 ;
        RECT 45.930 12.200 46.330 12.800 ;
        RECT 45.930 12.000 49.930 12.200 ;
        RECT 45.930 11.400 46.330 12.000 ;
        RECT 45.930 11.200 49.930 11.400 ;
        RECT 45.930 10.600 46.330 11.200 ;
        RECT 45.930 10.400 49.930 10.600 ;
        RECT 45.930 10.200 46.330 10.400 ;
        RECT 50.680 10.200 50.880 17.800 ;
        RECT 51.480 10.200 51.680 17.800 ;
        RECT 52.280 10.200 52.480 17.800 ;
        RECT 53.080 10.200 53.280 17.800 ;
        RECT 53.880 10.200 54.080 17.800 ;
        RECT 45.930 9.800 54.080 10.200 ;
        RECT 45.930 9.600 46.330 9.800 ;
        RECT 45.930 9.400 49.930 9.600 ;
        RECT 45.930 8.800 46.330 9.400 ;
        RECT 45.930 8.600 49.930 8.800 ;
        RECT 45.930 8.000 46.330 8.600 ;
        RECT 45.930 7.800 49.930 8.000 ;
        RECT 45.930 7.200 46.330 7.800 ;
        RECT 45.930 7.000 49.930 7.200 ;
        RECT 45.930 6.400 46.330 7.000 ;
        RECT 45.930 6.200 49.930 6.400 ;
        RECT 45.930 5.600 46.330 6.200 ;
        RECT 45.930 5.400 49.930 5.600 ;
        RECT 45.930 4.800 46.330 5.400 ;
        RECT 45.930 4.600 49.930 4.800 ;
        RECT 45.930 4.000 46.330 4.600 ;
        RECT 45.930 3.800 49.930 4.000 ;
        RECT 45.930 3.200 46.330 3.800 ;
        RECT 45.930 3.000 49.930 3.200 ;
        RECT 45.930 2.400 46.330 3.000 ;
        RECT 45.930 2.200 49.930 2.400 ;
        RECT 50.680 2.200 50.880 9.800 ;
        RECT 51.480 2.200 51.680 9.800 ;
        RECT 52.280 2.200 52.480 9.800 ;
        RECT 53.080 2.200 53.280 9.800 ;
        RECT 53.880 2.200 54.080 9.800 ;
        RECT 55.380 10.200 55.580 17.800 ;
        RECT 56.180 10.200 56.380 17.800 ;
        RECT 56.980 10.200 57.180 17.800 ;
        RECT 57.780 10.200 57.980 17.800 ;
        RECT 58.580 10.200 58.780 17.800 ;
        RECT 59.530 17.600 63.530 17.800 ;
        RECT 63.130 17.000 63.530 17.600 ;
        RECT 59.530 16.800 63.530 17.000 ;
        RECT 63.130 16.200 63.530 16.800 ;
        RECT 59.530 16.000 63.530 16.200 ;
        RECT 63.130 15.400 63.530 16.000 ;
        RECT 59.530 15.200 63.530 15.400 ;
        RECT 63.130 14.600 63.530 15.200 ;
        RECT 59.530 14.400 63.530 14.600 ;
        RECT 63.130 13.800 63.530 14.400 ;
        RECT 59.530 13.600 63.530 13.800 ;
        RECT 63.130 13.000 63.530 13.600 ;
        RECT 59.530 12.800 63.530 13.000 ;
        RECT 63.130 12.200 63.530 12.800 ;
        RECT 59.530 12.000 63.530 12.200 ;
        RECT 63.130 11.400 63.530 12.000 ;
        RECT 59.530 11.200 63.530 11.400 ;
        RECT 63.130 10.600 63.530 11.200 ;
        RECT 59.530 10.400 63.530 10.600 ;
        RECT 63.130 10.200 63.530 10.400 ;
        RECT 55.380 9.800 63.530 10.200 ;
        RECT 55.380 2.200 55.580 9.800 ;
        RECT 56.180 2.200 56.380 9.800 ;
        RECT 56.980 2.200 57.180 9.800 ;
        RECT 57.780 2.200 57.980 9.800 ;
        RECT 58.580 2.200 58.780 9.800 ;
        RECT 63.130 9.600 63.530 9.800 ;
        RECT 59.530 9.400 63.530 9.600 ;
        RECT 63.130 8.800 63.530 9.400 ;
        RECT 59.530 8.600 63.530 8.800 ;
        RECT 63.130 8.000 63.530 8.600 ;
        RECT 59.530 7.800 63.530 8.000 ;
        RECT 63.130 7.200 63.530 7.800 ;
        RECT 59.530 7.000 63.530 7.200 ;
        RECT 63.130 6.400 63.530 7.000 ;
        RECT 59.530 6.200 63.530 6.400 ;
        RECT 63.130 5.600 63.530 6.200 ;
        RECT 59.530 5.400 63.530 5.600 ;
        RECT 63.130 4.800 63.530 5.400 ;
        RECT 59.530 4.600 63.530 4.800 ;
        RECT 63.130 4.000 63.530 4.600 ;
        RECT 59.530 3.800 63.530 4.000 ;
        RECT 63.130 3.200 63.530 3.800 ;
        RECT 59.530 3.000 63.530 3.200 ;
        RECT 63.130 2.400 63.530 3.000 ;
        RECT 59.530 2.200 63.530 2.400 ;
        RECT 65.930 17.600 69.930 17.800 ;
        RECT 65.930 17.000 66.330 17.600 ;
        RECT 65.930 16.800 69.930 17.000 ;
        RECT 65.930 16.200 66.330 16.800 ;
        RECT 65.930 16.000 69.930 16.200 ;
        RECT 65.930 15.400 66.330 16.000 ;
        RECT 65.930 15.200 69.930 15.400 ;
        RECT 65.930 14.600 66.330 15.200 ;
        RECT 65.930 14.400 69.930 14.600 ;
        RECT 65.930 13.800 66.330 14.400 ;
        RECT 65.930 13.600 69.930 13.800 ;
        RECT 65.930 13.000 66.330 13.600 ;
        RECT 65.930 12.800 69.930 13.000 ;
        RECT 65.930 12.200 66.330 12.800 ;
        RECT 65.930 12.000 69.930 12.200 ;
        RECT 65.930 11.400 66.330 12.000 ;
        RECT 65.930 11.200 69.930 11.400 ;
        RECT 65.930 10.600 66.330 11.200 ;
        RECT 65.930 10.400 69.930 10.600 ;
        RECT 65.930 10.200 66.330 10.400 ;
        RECT 70.680 10.200 70.880 17.800 ;
        RECT 71.480 10.200 71.680 17.800 ;
        RECT 72.280 10.200 72.480 17.800 ;
        RECT 73.080 10.200 73.280 17.800 ;
        RECT 73.880 10.200 74.080 17.800 ;
        RECT 65.930 9.800 74.080 10.200 ;
        RECT 65.930 9.600 66.330 9.800 ;
        RECT 65.930 9.400 69.930 9.600 ;
        RECT 65.930 8.800 66.330 9.400 ;
        RECT 65.930 8.600 69.930 8.800 ;
        RECT 65.930 8.000 66.330 8.600 ;
        RECT 65.930 7.800 69.930 8.000 ;
        RECT 65.930 7.200 66.330 7.800 ;
        RECT 65.930 7.000 69.930 7.200 ;
        RECT 65.930 6.400 66.330 7.000 ;
        RECT 65.930 6.200 69.930 6.400 ;
        RECT 65.930 5.600 66.330 6.200 ;
        RECT 65.930 5.400 69.930 5.600 ;
        RECT 65.930 4.800 66.330 5.400 ;
        RECT 65.930 4.600 69.930 4.800 ;
        RECT 65.930 4.000 66.330 4.600 ;
        RECT 65.930 3.800 69.930 4.000 ;
        RECT 65.930 3.200 66.330 3.800 ;
        RECT 65.930 3.000 69.930 3.200 ;
        RECT 65.930 2.400 66.330 3.000 ;
        RECT 65.930 2.200 69.930 2.400 ;
        RECT 70.680 2.200 70.880 9.800 ;
        RECT 71.480 2.200 71.680 9.800 ;
        RECT 72.280 2.200 72.480 9.800 ;
        RECT 73.080 2.200 73.280 9.800 ;
        RECT 73.880 2.200 74.080 9.800 ;
        RECT 75.380 10.200 75.580 17.800 ;
        RECT 76.180 10.200 76.380 17.800 ;
        RECT 76.980 10.200 77.180 17.800 ;
        RECT 77.780 10.200 77.980 17.800 ;
        RECT 78.580 10.200 78.780 17.800 ;
        RECT 79.530 17.600 83.530 17.800 ;
        RECT 83.130 17.000 83.530 17.600 ;
        RECT 79.530 16.800 83.530 17.000 ;
        RECT 83.130 16.200 83.530 16.800 ;
        RECT 79.530 16.000 83.530 16.200 ;
        RECT 83.130 15.400 83.530 16.000 ;
        RECT 79.530 15.200 83.530 15.400 ;
        RECT 83.130 14.600 83.530 15.200 ;
        RECT 79.530 14.400 83.530 14.600 ;
        RECT 83.130 13.800 83.530 14.400 ;
        RECT 79.530 13.600 83.530 13.800 ;
        RECT 83.130 13.000 83.530 13.600 ;
        RECT 79.530 12.800 83.530 13.000 ;
        RECT 83.130 12.200 83.530 12.800 ;
        RECT 79.530 12.000 83.530 12.200 ;
        RECT 83.130 11.400 83.530 12.000 ;
        RECT 79.530 11.200 83.530 11.400 ;
        RECT 83.130 10.600 83.530 11.200 ;
        RECT 79.530 10.400 83.530 10.600 ;
        RECT 83.130 10.200 83.530 10.400 ;
        RECT 75.380 9.800 83.530 10.200 ;
        RECT 75.380 2.200 75.580 9.800 ;
        RECT 76.180 2.200 76.380 9.800 ;
        RECT 76.980 2.200 77.180 9.800 ;
        RECT 77.780 2.200 77.980 9.800 ;
        RECT 78.580 2.200 78.780 9.800 ;
        RECT 83.130 9.600 83.530 9.800 ;
        RECT 79.530 9.400 83.530 9.600 ;
        RECT 83.130 8.800 83.530 9.400 ;
        RECT 79.530 8.600 83.530 8.800 ;
        RECT 83.130 8.000 83.530 8.600 ;
        RECT 79.530 7.800 83.530 8.000 ;
        RECT 83.130 7.200 83.530 7.800 ;
        RECT 79.530 7.000 83.530 7.200 ;
        RECT 83.130 6.400 83.530 7.000 ;
        RECT 79.530 6.200 83.530 6.400 ;
        RECT 83.130 5.600 83.530 6.200 ;
        RECT 79.530 5.400 83.530 5.600 ;
        RECT 83.130 4.800 83.530 5.400 ;
        RECT 79.530 4.600 83.530 4.800 ;
        RECT 83.130 4.000 83.530 4.600 ;
        RECT 79.530 3.800 83.530 4.000 ;
        RECT 83.130 3.200 83.530 3.800 ;
        RECT 79.530 3.000 83.530 3.200 ;
        RECT 83.130 2.400 83.530 3.000 ;
        RECT 79.530 2.200 83.530 2.400 ;
        RECT 85.930 17.600 89.930 17.800 ;
        RECT 85.930 17.000 86.330 17.600 ;
        RECT 85.930 16.800 89.930 17.000 ;
        RECT 85.930 16.200 86.330 16.800 ;
        RECT 85.930 16.000 89.930 16.200 ;
        RECT 85.930 15.400 86.330 16.000 ;
        RECT 85.930 15.200 89.930 15.400 ;
        RECT 85.930 14.600 86.330 15.200 ;
        RECT 85.930 14.400 89.930 14.600 ;
        RECT 85.930 13.800 86.330 14.400 ;
        RECT 85.930 13.600 89.930 13.800 ;
        RECT 85.930 13.000 86.330 13.600 ;
        RECT 85.930 12.800 89.930 13.000 ;
        RECT 85.930 12.200 86.330 12.800 ;
        RECT 85.930 12.000 89.930 12.200 ;
        RECT 85.930 11.400 86.330 12.000 ;
        RECT 85.930 11.200 89.930 11.400 ;
        RECT 85.930 10.600 86.330 11.200 ;
        RECT 85.930 10.400 89.930 10.600 ;
        RECT 85.930 10.200 86.330 10.400 ;
        RECT 90.680 10.200 90.880 17.800 ;
        RECT 91.480 10.200 91.680 17.800 ;
        RECT 92.280 10.200 92.480 17.800 ;
        RECT 93.080 10.200 93.280 17.800 ;
        RECT 93.880 10.200 94.080 17.800 ;
        RECT 85.930 9.800 94.080 10.200 ;
        RECT 85.930 9.600 86.330 9.800 ;
        RECT 85.930 9.400 89.930 9.600 ;
        RECT 85.930 8.800 86.330 9.400 ;
        RECT 85.930 8.600 89.930 8.800 ;
        RECT 85.930 8.000 86.330 8.600 ;
        RECT 85.930 7.800 89.930 8.000 ;
        RECT 85.930 7.200 86.330 7.800 ;
        RECT 85.930 7.000 89.930 7.200 ;
        RECT 85.930 6.400 86.330 7.000 ;
        RECT 85.930 6.200 89.930 6.400 ;
        RECT 85.930 5.600 86.330 6.200 ;
        RECT 85.930 5.400 89.930 5.600 ;
        RECT 85.930 4.800 86.330 5.400 ;
        RECT 85.930 4.600 89.930 4.800 ;
        RECT 85.930 4.000 86.330 4.600 ;
        RECT 85.930 3.800 89.930 4.000 ;
        RECT 85.930 3.200 86.330 3.800 ;
        RECT 85.930 3.000 89.930 3.200 ;
        RECT 85.930 2.400 86.330 3.000 ;
        RECT 85.930 2.200 89.930 2.400 ;
        RECT 90.680 2.200 90.880 9.800 ;
        RECT 91.480 2.200 91.680 9.800 ;
        RECT 92.280 2.200 92.480 9.800 ;
        RECT 93.080 2.200 93.280 9.800 ;
        RECT 93.880 2.200 94.080 9.800 ;
        RECT 95.380 10.200 95.580 17.800 ;
        RECT 96.180 10.200 96.380 17.800 ;
        RECT 96.980 10.200 97.180 17.800 ;
        RECT 97.780 10.200 97.980 17.800 ;
        RECT 98.580 10.200 98.780 17.800 ;
        RECT 99.530 17.600 103.530 17.800 ;
        RECT 103.130 17.000 103.530 17.600 ;
        RECT 99.530 16.800 103.530 17.000 ;
        RECT 103.130 16.200 103.530 16.800 ;
        RECT 99.530 16.000 103.530 16.200 ;
        RECT 103.130 15.400 103.530 16.000 ;
        RECT 99.530 15.200 103.530 15.400 ;
        RECT 103.130 14.600 103.530 15.200 ;
        RECT 99.530 14.400 103.530 14.600 ;
        RECT 103.130 13.800 103.530 14.400 ;
        RECT 99.530 13.600 103.530 13.800 ;
        RECT 103.130 13.000 103.530 13.600 ;
        RECT 99.530 12.800 103.530 13.000 ;
        RECT 103.130 12.200 103.530 12.800 ;
        RECT 99.530 12.000 103.530 12.200 ;
        RECT 103.130 11.400 103.530 12.000 ;
        RECT 99.530 11.200 103.530 11.400 ;
        RECT 103.130 10.600 103.530 11.200 ;
        RECT 99.530 10.400 103.530 10.600 ;
        RECT 103.130 10.200 103.530 10.400 ;
        RECT 95.380 9.800 103.530 10.200 ;
        RECT 95.380 2.200 95.580 9.800 ;
        RECT 96.180 2.200 96.380 9.800 ;
        RECT 96.980 2.200 97.180 9.800 ;
        RECT 97.780 2.200 97.980 9.800 ;
        RECT 98.580 2.200 98.780 9.800 ;
        RECT 103.130 9.600 103.530 9.800 ;
        RECT 99.530 9.400 103.530 9.600 ;
        RECT 103.130 8.800 103.530 9.400 ;
        RECT 99.530 8.600 103.530 8.800 ;
        RECT 103.130 8.000 103.530 8.600 ;
        RECT 99.530 7.800 103.530 8.000 ;
        RECT 103.130 7.200 103.530 7.800 ;
        RECT 99.530 7.000 103.530 7.200 ;
        RECT 103.130 6.400 103.530 7.000 ;
        RECT 99.530 6.200 103.530 6.400 ;
        RECT 103.130 5.600 103.530 6.200 ;
        RECT 99.530 5.400 103.530 5.600 ;
        RECT 103.130 4.800 103.530 5.400 ;
        RECT 99.530 4.600 103.530 4.800 ;
        RECT 103.130 4.000 103.530 4.600 ;
        RECT 99.530 3.800 103.530 4.000 ;
        RECT 103.130 3.200 103.530 3.800 ;
        RECT 99.530 3.000 103.530 3.200 ;
        RECT 103.130 2.400 103.530 3.000 ;
        RECT 99.530 2.200 103.530 2.400 ;
        RECT 105.930 17.600 109.930 17.800 ;
        RECT 105.930 17.000 106.330 17.600 ;
        RECT 105.930 16.800 109.930 17.000 ;
        RECT 105.930 16.200 106.330 16.800 ;
        RECT 105.930 16.000 109.930 16.200 ;
        RECT 105.930 15.400 106.330 16.000 ;
        RECT 105.930 15.200 109.930 15.400 ;
        RECT 105.930 14.600 106.330 15.200 ;
        RECT 105.930 14.400 109.930 14.600 ;
        RECT 105.930 13.800 106.330 14.400 ;
        RECT 105.930 13.600 109.930 13.800 ;
        RECT 105.930 13.000 106.330 13.600 ;
        RECT 105.930 12.800 109.930 13.000 ;
        RECT 105.930 12.200 106.330 12.800 ;
        RECT 105.930 12.000 109.930 12.200 ;
        RECT 105.930 11.400 106.330 12.000 ;
        RECT 105.930 11.200 109.930 11.400 ;
        RECT 105.930 10.600 106.330 11.200 ;
        RECT 105.930 10.400 109.930 10.600 ;
        RECT 105.930 10.200 106.330 10.400 ;
        RECT 110.680 10.200 110.880 17.800 ;
        RECT 111.480 10.200 111.680 17.800 ;
        RECT 112.280 10.200 112.480 17.800 ;
        RECT 113.080 10.200 113.280 17.800 ;
        RECT 113.880 10.200 114.080 17.800 ;
        RECT 105.930 9.800 114.080 10.200 ;
        RECT 105.930 9.600 106.330 9.800 ;
        RECT 105.930 9.400 109.930 9.600 ;
        RECT 105.930 8.800 106.330 9.400 ;
        RECT 105.930 8.600 109.930 8.800 ;
        RECT 105.930 8.000 106.330 8.600 ;
        RECT 105.930 7.800 109.930 8.000 ;
        RECT 105.930 7.200 106.330 7.800 ;
        RECT 105.930 7.000 109.930 7.200 ;
        RECT 105.930 6.400 106.330 7.000 ;
        RECT 105.930 6.200 109.930 6.400 ;
        RECT 105.930 5.600 106.330 6.200 ;
        RECT 105.930 5.400 109.930 5.600 ;
        RECT 105.930 4.800 106.330 5.400 ;
        RECT 105.930 4.600 109.930 4.800 ;
        RECT 105.930 4.000 106.330 4.600 ;
        RECT 105.930 3.800 109.930 4.000 ;
        RECT 105.930 3.200 106.330 3.800 ;
        RECT 105.930 3.000 109.930 3.200 ;
        RECT 105.930 2.400 106.330 3.000 ;
        RECT 105.930 2.200 109.930 2.400 ;
        RECT 110.680 2.200 110.880 9.800 ;
        RECT 111.480 2.200 111.680 9.800 ;
        RECT 112.280 2.200 112.480 9.800 ;
        RECT 113.080 2.200 113.280 9.800 ;
        RECT 113.880 2.200 114.080 9.800 ;
        RECT 115.380 10.200 115.580 17.800 ;
        RECT 116.180 10.200 116.380 17.800 ;
        RECT 116.980 10.200 117.180 17.800 ;
        RECT 117.780 10.200 117.980 17.800 ;
        RECT 118.580 10.200 118.780 17.800 ;
        RECT 119.530 17.600 123.530 17.800 ;
        RECT 123.130 17.000 123.530 17.600 ;
        RECT 119.530 16.800 123.530 17.000 ;
        RECT 123.130 16.200 123.530 16.800 ;
        RECT 119.530 16.000 123.530 16.200 ;
        RECT 123.130 15.400 123.530 16.000 ;
        RECT 119.530 15.200 123.530 15.400 ;
        RECT 123.130 14.600 123.530 15.200 ;
        RECT 119.530 14.400 123.530 14.600 ;
        RECT 123.130 13.800 123.530 14.400 ;
        RECT 119.530 13.600 123.530 13.800 ;
        RECT 123.130 13.000 123.530 13.600 ;
        RECT 119.530 12.800 123.530 13.000 ;
        RECT 123.130 12.200 123.530 12.800 ;
        RECT 119.530 12.000 123.530 12.200 ;
        RECT 123.130 11.400 123.530 12.000 ;
        RECT 119.530 11.200 123.530 11.400 ;
        RECT 123.130 10.600 123.530 11.200 ;
        RECT 130.050 11.020 130.410 11.400 ;
        RECT 130.680 11.020 131.040 11.400 ;
        RECT 131.280 11.020 131.640 11.400 ;
        RECT 119.530 10.400 123.530 10.600 ;
        RECT 130.050 10.430 130.410 10.810 ;
        RECT 130.680 10.430 131.040 10.810 ;
        RECT 131.280 10.430 131.640 10.810 ;
        RECT 123.130 10.200 123.530 10.400 ;
        RECT 115.380 9.800 123.530 10.200 ;
        RECT 115.380 2.200 115.580 9.800 ;
        RECT 116.180 2.200 116.380 9.800 ;
        RECT 116.980 2.200 117.180 9.800 ;
        RECT 117.780 2.200 117.980 9.800 ;
        RECT 118.580 2.200 118.780 9.800 ;
        RECT 123.130 9.600 123.530 9.800 ;
        RECT 119.530 9.400 123.530 9.600 ;
        RECT 123.130 8.800 123.530 9.400 ;
        RECT 119.530 8.600 123.530 8.800 ;
        RECT 123.130 8.000 123.530 8.600 ;
        RECT 119.530 7.800 123.530 8.000 ;
        RECT 123.130 7.200 123.530 7.800 ;
        RECT 119.530 7.000 123.530 7.200 ;
        RECT 123.130 6.400 123.530 7.000 ;
        RECT 119.530 6.200 123.530 6.400 ;
        RECT 123.130 5.600 123.530 6.200 ;
        RECT 119.530 5.400 123.530 5.600 ;
        RECT 123.130 4.800 123.530 5.400 ;
        RECT 119.530 4.600 123.530 4.800 ;
        RECT 123.130 4.000 123.530 4.600 ;
        RECT 119.530 3.800 123.530 4.000 ;
        RECT 123.130 3.200 123.530 3.800 ;
        RECT 119.530 3.000 123.530 3.200 ;
        RECT 123.130 2.400 123.530 3.000 ;
        RECT 119.530 2.200 123.530 2.400 ;
      LAYER mcon ;
        RECT 5.980 334.300 6.280 334.750 ;
        RECT 5.980 333.550 6.280 334.000 ;
        RECT 5.980 332.800 6.280 333.250 ;
        RECT 5.980 332.050 6.280 332.500 ;
        RECT 5.980 331.300 6.280 331.750 ;
        RECT 5.980 330.550 6.280 331.000 ;
        RECT 5.980 329.800 6.280 330.250 ;
        RECT 5.980 329.050 6.280 329.500 ;
        RECT 5.980 328.300 6.280 328.750 ;
        RECT 5.980 327.550 6.280 328.000 ;
        RECT 5.980 326.800 6.280 327.250 ;
        RECT 5.980 326.050 6.280 326.500 ;
        RECT 5.980 325.300 6.280 325.750 ;
        RECT 23.180 334.300 23.480 334.750 ;
        RECT 23.180 333.550 23.480 334.000 ;
        RECT 23.180 332.800 23.480 333.250 ;
        RECT 23.180 332.050 23.480 332.500 ;
        RECT 23.180 331.300 23.480 331.750 ;
        RECT 23.180 330.550 23.480 331.000 ;
        RECT 23.180 329.800 23.480 330.250 ;
        RECT 23.180 329.050 23.480 329.500 ;
        RECT 23.180 328.300 23.480 328.750 ;
        RECT 23.180 327.550 23.480 328.000 ;
        RECT 23.180 326.800 23.480 327.250 ;
        RECT 23.180 326.050 23.480 326.500 ;
        RECT 23.180 325.300 23.480 325.750 ;
        RECT 25.980 334.300 26.280 334.750 ;
        RECT 25.980 333.550 26.280 334.000 ;
        RECT 25.980 332.800 26.280 333.250 ;
        RECT 25.980 332.050 26.280 332.500 ;
        RECT 25.980 331.300 26.280 331.750 ;
        RECT 25.980 330.550 26.280 331.000 ;
        RECT 25.980 329.800 26.280 330.250 ;
        RECT 25.980 329.050 26.280 329.500 ;
        RECT 25.980 328.300 26.280 328.750 ;
        RECT 25.980 327.550 26.280 328.000 ;
        RECT 25.980 326.800 26.280 327.250 ;
        RECT 25.980 326.050 26.280 326.500 ;
        RECT 25.980 325.300 26.280 325.750 ;
        RECT 43.180 334.300 43.480 334.750 ;
        RECT 43.180 333.550 43.480 334.000 ;
        RECT 43.180 332.800 43.480 333.250 ;
        RECT 43.180 332.050 43.480 332.500 ;
        RECT 43.180 331.300 43.480 331.750 ;
        RECT 43.180 330.550 43.480 331.000 ;
        RECT 43.180 329.800 43.480 330.250 ;
        RECT 43.180 329.050 43.480 329.500 ;
        RECT 43.180 328.300 43.480 328.750 ;
        RECT 43.180 327.550 43.480 328.000 ;
        RECT 43.180 326.800 43.480 327.250 ;
        RECT 43.180 326.050 43.480 326.500 ;
        RECT 43.180 325.300 43.480 325.750 ;
        RECT 45.980 334.300 46.280 334.750 ;
        RECT 45.980 333.550 46.280 334.000 ;
        RECT 45.980 332.800 46.280 333.250 ;
        RECT 45.980 332.050 46.280 332.500 ;
        RECT 45.980 331.300 46.280 331.750 ;
        RECT 45.980 330.550 46.280 331.000 ;
        RECT 45.980 329.800 46.280 330.250 ;
        RECT 45.980 329.050 46.280 329.500 ;
        RECT 45.980 328.300 46.280 328.750 ;
        RECT 45.980 327.550 46.280 328.000 ;
        RECT 45.980 326.800 46.280 327.250 ;
        RECT 45.980 326.050 46.280 326.500 ;
        RECT 45.980 325.300 46.280 325.750 ;
        RECT 63.180 334.300 63.480 334.750 ;
        RECT 63.180 333.550 63.480 334.000 ;
        RECT 63.180 332.800 63.480 333.250 ;
        RECT 63.180 332.050 63.480 332.500 ;
        RECT 63.180 331.300 63.480 331.750 ;
        RECT 63.180 330.550 63.480 331.000 ;
        RECT 63.180 329.800 63.480 330.250 ;
        RECT 63.180 329.050 63.480 329.500 ;
        RECT 63.180 328.300 63.480 328.750 ;
        RECT 63.180 327.550 63.480 328.000 ;
        RECT 63.180 326.800 63.480 327.250 ;
        RECT 63.180 326.050 63.480 326.500 ;
        RECT 63.180 325.300 63.480 325.750 ;
        RECT 65.980 334.300 66.280 334.750 ;
        RECT 65.980 333.550 66.280 334.000 ;
        RECT 65.980 332.800 66.280 333.250 ;
        RECT 65.980 332.050 66.280 332.500 ;
        RECT 65.980 331.300 66.280 331.750 ;
        RECT 65.980 330.550 66.280 331.000 ;
        RECT 65.980 329.800 66.280 330.250 ;
        RECT 65.980 329.050 66.280 329.500 ;
        RECT 65.980 328.300 66.280 328.750 ;
        RECT 65.980 327.550 66.280 328.000 ;
        RECT 65.980 326.800 66.280 327.250 ;
        RECT 65.980 326.050 66.280 326.500 ;
        RECT 65.980 325.300 66.280 325.750 ;
        RECT 83.180 334.300 83.480 334.750 ;
        RECT 83.180 333.550 83.480 334.000 ;
        RECT 83.180 332.800 83.480 333.250 ;
        RECT 83.180 332.050 83.480 332.500 ;
        RECT 83.180 331.300 83.480 331.750 ;
        RECT 83.180 330.550 83.480 331.000 ;
        RECT 83.180 329.800 83.480 330.250 ;
        RECT 83.180 329.050 83.480 329.500 ;
        RECT 83.180 328.300 83.480 328.750 ;
        RECT 83.180 327.550 83.480 328.000 ;
        RECT 83.180 326.800 83.480 327.250 ;
        RECT 83.180 326.050 83.480 326.500 ;
        RECT 83.180 325.300 83.480 325.750 ;
        RECT 85.980 334.300 86.280 334.750 ;
        RECT 85.980 333.550 86.280 334.000 ;
        RECT 85.980 332.800 86.280 333.250 ;
        RECT 85.980 332.050 86.280 332.500 ;
        RECT 85.980 331.300 86.280 331.750 ;
        RECT 85.980 330.550 86.280 331.000 ;
        RECT 85.980 329.800 86.280 330.250 ;
        RECT 85.980 329.050 86.280 329.500 ;
        RECT 85.980 328.300 86.280 328.750 ;
        RECT 85.980 327.550 86.280 328.000 ;
        RECT 85.980 326.800 86.280 327.250 ;
        RECT 85.980 326.050 86.280 326.500 ;
        RECT 85.980 325.300 86.280 325.750 ;
        RECT 103.180 334.300 103.480 334.750 ;
        RECT 103.180 333.550 103.480 334.000 ;
        RECT 103.180 332.800 103.480 333.250 ;
        RECT 103.180 332.050 103.480 332.500 ;
        RECT 103.180 331.300 103.480 331.750 ;
        RECT 103.180 330.550 103.480 331.000 ;
        RECT 103.180 329.800 103.480 330.250 ;
        RECT 103.180 329.050 103.480 329.500 ;
        RECT 103.180 328.300 103.480 328.750 ;
        RECT 103.180 327.550 103.480 328.000 ;
        RECT 103.180 326.800 103.480 327.250 ;
        RECT 103.180 326.050 103.480 326.500 ;
        RECT 103.180 325.300 103.480 325.750 ;
        RECT 105.980 334.300 106.280 334.750 ;
        RECT 105.980 333.550 106.280 334.000 ;
        RECT 105.980 332.800 106.280 333.250 ;
        RECT 105.980 332.050 106.280 332.500 ;
        RECT 105.980 331.300 106.280 331.750 ;
        RECT 105.980 330.550 106.280 331.000 ;
        RECT 105.980 329.800 106.280 330.250 ;
        RECT 105.980 329.050 106.280 329.500 ;
        RECT 105.980 328.300 106.280 328.750 ;
        RECT 105.980 327.550 106.280 328.000 ;
        RECT 105.980 326.800 106.280 327.250 ;
        RECT 105.980 326.050 106.280 326.500 ;
        RECT 105.980 325.300 106.280 325.750 ;
        RECT 123.180 334.300 123.480 334.750 ;
        RECT 123.180 333.550 123.480 334.000 ;
        RECT 123.180 332.800 123.480 333.250 ;
        RECT 123.180 332.050 123.480 332.500 ;
        RECT 123.180 331.300 123.480 331.750 ;
        RECT 123.180 330.550 123.480 331.000 ;
        RECT 123.180 329.800 123.480 330.250 ;
        RECT 123.180 329.050 123.480 329.500 ;
        RECT 123.180 328.300 123.480 328.750 ;
        RECT 123.180 327.550 123.480 328.000 ;
        RECT 123.180 326.800 123.480 327.250 ;
        RECT 123.180 326.050 123.480 326.500 ;
        RECT 123.180 325.300 123.480 325.750 ;
        RECT 5.980 314.300 6.280 314.750 ;
        RECT 5.980 313.550 6.280 314.000 ;
        RECT 5.980 312.800 6.280 313.250 ;
        RECT 5.980 312.050 6.280 312.500 ;
        RECT 5.980 311.300 6.280 311.750 ;
        RECT 5.980 310.550 6.280 311.000 ;
        RECT 5.980 309.800 6.280 310.250 ;
        RECT 5.980 309.050 6.280 309.500 ;
        RECT 5.980 308.300 6.280 308.750 ;
        RECT 5.980 307.550 6.280 308.000 ;
        RECT 5.980 306.800 6.280 307.250 ;
        RECT 5.980 306.050 6.280 306.500 ;
        RECT 5.980 305.300 6.280 305.750 ;
        RECT 23.180 314.300 23.480 314.750 ;
        RECT 23.180 313.550 23.480 314.000 ;
        RECT 23.180 312.800 23.480 313.250 ;
        RECT 23.180 312.050 23.480 312.500 ;
        RECT 23.180 311.300 23.480 311.750 ;
        RECT 23.180 310.550 23.480 311.000 ;
        RECT 23.180 309.800 23.480 310.250 ;
        RECT 23.180 309.050 23.480 309.500 ;
        RECT 23.180 308.300 23.480 308.750 ;
        RECT 23.180 307.550 23.480 308.000 ;
        RECT 23.180 306.800 23.480 307.250 ;
        RECT 23.180 306.050 23.480 306.500 ;
        RECT 23.180 305.300 23.480 305.750 ;
        RECT 25.980 314.300 26.280 314.750 ;
        RECT 25.980 313.550 26.280 314.000 ;
        RECT 25.980 312.800 26.280 313.250 ;
        RECT 25.980 312.050 26.280 312.500 ;
        RECT 25.980 311.300 26.280 311.750 ;
        RECT 25.980 310.550 26.280 311.000 ;
        RECT 25.980 309.800 26.280 310.250 ;
        RECT 25.980 309.050 26.280 309.500 ;
        RECT 25.980 308.300 26.280 308.750 ;
        RECT 25.980 307.550 26.280 308.000 ;
        RECT 25.980 306.800 26.280 307.250 ;
        RECT 25.980 306.050 26.280 306.500 ;
        RECT 25.980 305.300 26.280 305.750 ;
        RECT 43.180 314.300 43.480 314.750 ;
        RECT 43.180 313.550 43.480 314.000 ;
        RECT 43.180 312.800 43.480 313.250 ;
        RECT 43.180 312.050 43.480 312.500 ;
        RECT 43.180 311.300 43.480 311.750 ;
        RECT 43.180 310.550 43.480 311.000 ;
        RECT 43.180 309.800 43.480 310.250 ;
        RECT 43.180 309.050 43.480 309.500 ;
        RECT 43.180 308.300 43.480 308.750 ;
        RECT 43.180 307.550 43.480 308.000 ;
        RECT 43.180 306.800 43.480 307.250 ;
        RECT 43.180 306.050 43.480 306.500 ;
        RECT 43.180 305.300 43.480 305.750 ;
        RECT 45.980 314.300 46.280 314.750 ;
        RECT 45.980 313.550 46.280 314.000 ;
        RECT 45.980 312.800 46.280 313.250 ;
        RECT 45.980 312.050 46.280 312.500 ;
        RECT 45.980 311.300 46.280 311.750 ;
        RECT 45.980 310.550 46.280 311.000 ;
        RECT 45.980 309.800 46.280 310.250 ;
        RECT 45.980 309.050 46.280 309.500 ;
        RECT 45.980 308.300 46.280 308.750 ;
        RECT 45.980 307.550 46.280 308.000 ;
        RECT 45.980 306.800 46.280 307.250 ;
        RECT 45.980 306.050 46.280 306.500 ;
        RECT 45.980 305.300 46.280 305.750 ;
        RECT 63.180 314.300 63.480 314.750 ;
        RECT 63.180 313.550 63.480 314.000 ;
        RECT 63.180 312.800 63.480 313.250 ;
        RECT 63.180 312.050 63.480 312.500 ;
        RECT 63.180 311.300 63.480 311.750 ;
        RECT 63.180 310.550 63.480 311.000 ;
        RECT 63.180 309.800 63.480 310.250 ;
        RECT 63.180 309.050 63.480 309.500 ;
        RECT 63.180 308.300 63.480 308.750 ;
        RECT 63.180 307.550 63.480 308.000 ;
        RECT 63.180 306.800 63.480 307.250 ;
        RECT 63.180 306.050 63.480 306.500 ;
        RECT 63.180 305.300 63.480 305.750 ;
        RECT 65.980 314.300 66.280 314.750 ;
        RECT 65.980 313.550 66.280 314.000 ;
        RECT 65.980 312.800 66.280 313.250 ;
        RECT 65.980 312.050 66.280 312.500 ;
        RECT 65.980 311.300 66.280 311.750 ;
        RECT 65.980 310.550 66.280 311.000 ;
        RECT 65.980 309.800 66.280 310.250 ;
        RECT 65.980 309.050 66.280 309.500 ;
        RECT 65.980 308.300 66.280 308.750 ;
        RECT 65.980 307.550 66.280 308.000 ;
        RECT 65.980 306.800 66.280 307.250 ;
        RECT 65.980 306.050 66.280 306.500 ;
        RECT 65.980 305.300 66.280 305.750 ;
        RECT 83.180 314.300 83.480 314.750 ;
        RECT 83.180 313.550 83.480 314.000 ;
        RECT 83.180 312.800 83.480 313.250 ;
        RECT 83.180 312.050 83.480 312.500 ;
        RECT 83.180 311.300 83.480 311.750 ;
        RECT 83.180 310.550 83.480 311.000 ;
        RECT 83.180 309.800 83.480 310.250 ;
        RECT 83.180 309.050 83.480 309.500 ;
        RECT 83.180 308.300 83.480 308.750 ;
        RECT 83.180 307.550 83.480 308.000 ;
        RECT 83.180 306.800 83.480 307.250 ;
        RECT 83.180 306.050 83.480 306.500 ;
        RECT 83.180 305.300 83.480 305.750 ;
        RECT 85.980 314.300 86.280 314.750 ;
        RECT 85.980 313.550 86.280 314.000 ;
        RECT 85.980 312.800 86.280 313.250 ;
        RECT 85.980 312.050 86.280 312.500 ;
        RECT 85.980 311.300 86.280 311.750 ;
        RECT 85.980 310.550 86.280 311.000 ;
        RECT 85.980 309.800 86.280 310.250 ;
        RECT 85.980 309.050 86.280 309.500 ;
        RECT 85.980 308.300 86.280 308.750 ;
        RECT 85.980 307.550 86.280 308.000 ;
        RECT 85.980 306.800 86.280 307.250 ;
        RECT 85.980 306.050 86.280 306.500 ;
        RECT 85.980 305.300 86.280 305.750 ;
        RECT 103.180 314.300 103.480 314.750 ;
        RECT 103.180 313.550 103.480 314.000 ;
        RECT 103.180 312.800 103.480 313.250 ;
        RECT 103.180 312.050 103.480 312.500 ;
        RECT 103.180 311.300 103.480 311.750 ;
        RECT 103.180 310.550 103.480 311.000 ;
        RECT 103.180 309.800 103.480 310.250 ;
        RECT 103.180 309.050 103.480 309.500 ;
        RECT 103.180 308.300 103.480 308.750 ;
        RECT 103.180 307.550 103.480 308.000 ;
        RECT 103.180 306.800 103.480 307.250 ;
        RECT 103.180 306.050 103.480 306.500 ;
        RECT 103.180 305.300 103.480 305.750 ;
        RECT 105.980 314.300 106.280 314.750 ;
        RECT 105.980 313.550 106.280 314.000 ;
        RECT 105.980 312.800 106.280 313.250 ;
        RECT 105.980 312.050 106.280 312.500 ;
        RECT 105.980 311.300 106.280 311.750 ;
        RECT 105.980 310.550 106.280 311.000 ;
        RECT 105.980 309.800 106.280 310.250 ;
        RECT 105.980 309.050 106.280 309.500 ;
        RECT 105.980 308.300 106.280 308.750 ;
        RECT 105.980 307.550 106.280 308.000 ;
        RECT 105.980 306.800 106.280 307.250 ;
        RECT 105.980 306.050 106.280 306.500 ;
        RECT 105.980 305.300 106.280 305.750 ;
        RECT 123.180 314.300 123.480 314.750 ;
        RECT 123.180 313.550 123.480 314.000 ;
        RECT 123.180 312.800 123.480 313.250 ;
        RECT 123.180 312.050 123.480 312.500 ;
        RECT 123.180 311.300 123.480 311.750 ;
        RECT 123.180 310.550 123.480 311.000 ;
        RECT 123.180 309.800 123.480 310.250 ;
        RECT 123.180 309.050 123.480 309.500 ;
        RECT 123.180 308.300 123.480 308.750 ;
        RECT 123.180 307.550 123.480 308.000 ;
        RECT 123.180 306.800 123.480 307.250 ;
        RECT 123.180 306.050 123.480 306.500 ;
        RECT 123.180 305.300 123.480 305.750 ;
        RECT 5.980 294.300 6.280 294.750 ;
        RECT 5.980 293.550 6.280 294.000 ;
        RECT 5.980 292.800 6.280 293.250 ;
        RECT 5.980 292.050 6.280 292.500 ;
        RECT 5.980 291.300 6.280 291.750 ;
        RECT 5.980 290.550 6.280 291.000 ;
        RECT 5.980 289.800 6.280 290.250 ;
        RECT 5.980 289.050 6.280 289.500 ;
        RECT 5.980 288.300 6.280 288.750 ;
        RECT 5.980 287.550 6.280 288.000 ;
        RECT 5.980 286.800 6.280 287.250 ;
        RECT 5.980 286.050 6.280 286.500 ;
        RECT 5.980 285.300 6.280 285.750 ;
        RECT 23.180 294.300 23.480 294.750 ;
        RECT 23.180 293.550 23.480 294.000 ;
        RECT 23.180 292.800 23.480 293.250 ;
        RECT 23.180 292.050 23.480 292.500 ;
        RECT 23.180 291.300 23.480 291.750 ;
        RECT 23.180 290.550 23.480 291.000 ;
        RECT 23.180 289.800 23.480 290.250 ;
        RECT 23.180 289.050 23.480 289.500 ;
        RECT 23.180 288.300 23.480 288.750 ;
        RECT 23.180 287.550 23.480 288.000 ;
        RECT 23.180 286.800 23.480 287.250 ;
        RECT 23.180 286.050 23.480 286.500 ;
        RECT 23.180 285.300 23.480 285.750 ;
        RECT 25.980 294.300 26.280 294.750 ;
        RECT 25.980 293.550 26.280 294.000 ;
        RECT 25.980 292.800 26.280 293.250 ;
        RECT 25.980 292.050 26.280 292.500 ;
        RECT 25.980 291.300 26.280 291.750 ;
        RECT 25.980 290.550 26.280 291.000 ;
        RECT 25.980 289.800 26.280 290.250 ;
        RECT 25.980 289.050 26.280 289.500 ;
        RECT 25.980 288.300 26.280 288.750 ;
        RECT 25.980 287.550 26.280 288.000 ;
        RECT 25.980 286.800 26.280 287.250 ;
        RECT 25.980 286.050 26.280 286.500 ;
        RECT 25.980 285.300 26.280 285.750 ;
        RECT 43.180 294.300 43.480 294.750 ;
        RECT 43.180 293.550 43.480 294.000 ;
        RECT 43.180 292.800 43.480 293.250 ;
        RECT 43.180 292.050 43.480 292.500 ;
        RECT 43.180 291.300 43.480 291.750 ;
        RECT 43.180 290.550 43.480 291.000 ;
        RECT 43.180 289.800 43.480 290.250 ;
        RECT 43.180 289.050 43.480 289.500 ;
        RECT 43.180 288.300 43.480 288.750 ;
        RECT 43.180 287.550 43.480 288.000 ;
        RECT 43.180 286.800 43.480 287.250 ;
        RECT 43.180 286.050 43.480 286.500 ;
        RECT 43.180 285.300 43.480 285.750 ;
        RECT 45.980 294.300 46.280 294.750 ;
        RECT 45.980 293.550 46.280 294.000 ;
        RECT 45.980 292.800 46.280 293.250 ;
        RECT 45.980 292.050 46.280 292.500 ;
        RECT 45.980 291.300 46.280 291.750 ;
        RECT 45.980 290.550 46.280 291.000 ;
        RECT 45.980 289.800 46.280 290.250 ;
        RECT 45.980 289.050 46.280 289.500 ;
        RECT 45.980 288.300 46.280 288.750 ;
        RECT 45.980 287.550 46.280 288.000 ;
        RECT 45.980 286.800 46.280 287.250 ;
        RECT 45.980 286.050 46.280 286.500 ;
        RECT 45.980 285.300 46.280 285.750 ;
        RECT 63.180 294.300 63.480 294.750 ;
        RECT 63.180 293.550 63.480 294.000 ;
        RECT 63.180 292.800 63.480 293.250 ;
        RECT 63.180 292.050 63.480 292.500 ;
        RECT 63.180 291.300 63.480 291.750 ;
        RECT 63.180 290.550 63.480 291.000 ;
        RECT 63.180 289.800 63.480 290.250 ;
        RECT 63.180 289.050 63.480 289.500 ;
        RECT 63.180 288.300 63.480 288.750 ;
        RECT 63.180 287.550 63.480 288.000 ;
        RECT 63.180 286.800 63.480 287.250 ;
        RECT 63.180 286.050 63.480 286.500 ;
        RECT 63.180 285.300 63.480 285.750 ;
        RECT 65.980 294.300 66.280 294.750 ;
        RECT 65.980 293.550 66.280 294.000 ;
        RECT 65.980 292.800 66.280 293.250 ;
        RECT 65.980 292.050 66.280 292.500 ;
        RECT 65.980 291.300 66.280 291.750 ;
        RECT 65.980 290.550 66.280 291.000 ;
        RECT 65.980 289.800 66.280 290.250 ;
        RECT 65.980 289.050 66.280 289.500 ;
        RECT 65.980 288.300 66.280 288.750 ;
        RECT 65.980 287.550 66.280 288.000 ;
        RECT 65.980 286.800 66.280 287.250 ;
        RECT 65.980 286.050 66.280 286.500 ;
        RECT 65.980 285.300 66.280 285.750 ;
        RECT 83.180 294.300 83.480 294.750 ;
        RECT 83.180 293.550 83.480 294.000 ;
        RECT 83.180 292.800 83.480 293.250 ;
        RECT 83.180 292.050 83.480 292.500 ;
        RECT 83.180 291.300 83.480 291.750 ;
        RECT 83.180 290.550 83.480 291.000 ;
        RECT 83.180 289.800 83.480 290.250 ;
        RECT 83.180 289.050 83.480 289.500 ;
        RECT 83.180 288.300 83.480 288.750 ;
        RECT 83.180 287.550 83.480 288.000 ;
        RECT 83.180 286.800 83.480 287.250 ;
        RECT 83.180 286.050 83.480 286.500 ;
        RECT 83.180 285.300 83.480 285.750 ;
        RECT 85.980 294.300 86.280 294.750 ;
        RECT 85.980 293.550 86.280 294.000 ;
        RECT 85.980 292.800 86.280 293.250 ;
        RECT 85.980 292.050 86.280 292.500 ;
        RECT 85.980 291.300 86.280 291.750 ;
        RECT 85.980 290.550 86.280 291.000 ;
        RECT 85.980 289.800 86.280 290.250 ;
        RECT 85.980 289.050 86.280 289.500 ;
        RECT 85.980 288.300 86.280 288.750 ;
        RECT 85.980 287.550 86.280 288.000 ;
        RECT 85.980 286.800 86.280 287.250 ;
        RECT 85.980 286.050 86.280 286.500 ;
        RECT 85.980 285.300 86.280 285.750 ;
        RECT 103.180 294.300 103.480 294.750 ;
        RECT 103.180 293.550 103.480 294.000 ;
        RECT 103.180 292.800 103.480 293.250 ;
        RECT 103.180 292.050 103.480 292.500 ;
        RECT 103.180 291.300 103.480 291.750 ;
        RECT 103.180 290.550 103.480 291.000 ;
        RECT 103.180 289.800 103.480 290.250 ;
        RECT 103.180 289.050 103.480 289.500 ;
        RECT 103.180 288.300 103.480 288.750 ;
        RECT 103.180 287.550 103.480 288.000 ;
        RECT 103.180 286.800 103.480 287.250 ;
        RECT 103.180 286.050 103.480 286.500 ;
        RECT 103.180 285.300 103.480 285.750 ;
        RECT 105.980 294.300 106.280 294.750 ;
        RECT 105.980 293.550 106.280 294.000 ;
        RECT 105.980 292.800 106.280 293.250 ;
        RECT 105.980 292.050 106.280 292.500 ;
        RECT 105.980 291.300 106.280 291.750 ;
        RECT 105.980 290.550 106.280 291.000 ;
        RECT 105.980 289.800 106.280 290.250 ;
        RECT 105.980 289.050 106.280 289.500 ;
        RECT 105.980 288.300 106.280 288.750 ;
        RECT 105.980 287.550 106.280 288.000 ;
        RECT 105.980 286.800 106.280 287.250 ;
        RECT 105.980 286.050 106.280 286.500 ;
        RECT 105.980 285.300 106.280 285.750 ;
        RECT 123.180 294.300 123.480 294.750 ;
        RECT 123.180 293.550 123.480 294.000 ;
        RECT 123.180 292.800 123.480 293.250 ;
        RECT 123.180 292.050 123.480 292.500 ;
        RECT 123.180 291.300 123.480 291.750 ;
        RECT 123.180 290.550 123.480 291.000 ;
        RECT 123.180 289.800 123.480 290.250 ;
        RECT 123.180 289.050 123.480 289.500 ;
        RECT 123.180 288.300 123.480 288.750 ;
        RECT 123.180 287.550 123.480 288.000 ;
        RECT 123.180 286.800 123.480 287.250 ;
        RECT 123.180 286.050 123.480 286.500 ;
        RECT 123.180 285.300 123.480 285.750 ;
        RECT 5.980 274.300 6.280 274.750 ;
        RECT 5.980 273.550 6.280 274.000 ;
        RECT 5.980 272.800 6.280 273.250 ;
        RECT 5.980 272.050 6.280 272.500 ;
        RECT 5.980 271.300 6.280 271.750 ;
        RECT 5.980 270.550 6.280 271.000 ;
        RECT 5.980 269.800 6.280 270.250 ;
        RECT 5.980 269.050 6.280 269.500 ;
        RECT 5.980 268.300 6.280 268.750 ;
        RECT 5.980 267.550 6.280 268.000 ;
        RECT 5.980 266.800 6.280 267.250 ;
        RECT 5.980 266.050 6.280 266.500 ;
        RECT 5.980 265.300 6.280 265.750 ;
        RECT 23.180 274.300 23.480 274.750 ;
        RECT 23.180 273.550 23.480 274.000 ;
        RECT 23.180 272.800 23.480 273.250 ;
        RECT 23.180 272.050 23.480 272.500 ;
        RECT 23.180 271.300 23.480 271.750 ;
        RECT 23.180 270.550 23.480 271.000 ;
        RECT 23.180 269.800 23.480 270.250 ;
        RECT 23.180 269.050 23.480 269.500 ;
        RECT 23.180 268.300 23.480 268.750 ;
        RECT 23.180 267.550 23.480 268.000 ;
        RECT 23.180 266.800 23.480 267.250 ;
        RECT 23.180 266.050 23.480 266.500 ;
        RECT 23.180 265.300 23.480 265.750 ;
        RECT 25.980 274.300 26.280 274.750 ;
        RECT 25.980 273.550 26.280 274.000 ;
        RECT 25.980 272.800 26.280 273.250 ;
        RECT 25.980 272.050 26.280 272.500 ;
        RECT 25.980 271.300 26.280 271.750 ;
        RECT 25.980 270.550 26.280 271.000 ;
        RECT 25.980 269.800 26.280 270.250 ;
        RECT 25.980 269.050 26.280 269.500 ;
        RECT 25.980 268.300 26.280 268.750 ;
        RECT 25.980 267.550 26.280 268.000 ;
        RECT 25.980 266.800 26.280 267.250 ;
        RECT 25.980 266.050 26.280 266.500 ;
        RECT 25.980 265.300 26.280 265.750 ;
        RECT 43.180 274.300 43.480 274.750 ;
        RECT 43.180 273.550 43.480 274.000 ;
        RECT 43.180 272.800 43.480 273.250 ;
        RECT 43.180 272.050 43.480 272.500 ;
        RECT 43.180 271.300 43.480 271.750 ;
        RECT 43.180 270.550 43.480 271.000 ;
        RECT 43.180 269.800 43.480 270.250 ;
        RECT 43.180 269.050 43.480 269.500 ;
        RECT 43.180 268.300 43.480 268.750 ;
        RECT 43.180 267.550 43.480 268.000 ;
        RECT 43.180 266.800 43.480 267.250 ;
        RECT 43.180 266.050 43.480 266.500 ;
        RECT 43.180 265.300 43.480 265.750 ;
        RECT 45.980 274.300 46.280 274.750 ;
        RECT 45.980 273.550 46.280 274.000 ;
        RECT 45.980 272.800 46.280 273.250 ;
        RECT 45.980 272.050 46.280 272.500 ;
        RECT 45.980 271.300 46.280 271.750 ;
        RECT 45.980 270.550 46.280 271.000 ;
        RECT 45.980 269.800 46.280 270.250 ;
        RECT 45.980 269.050 46.280 269.500 ;
        RECT 45.980 268.300 46.280 268.750 ;
        RECT 45.980 267.550 46.280 268.000 ;
        RECT 45.980 266.800 46.280 267.250 ;
        RECT 45.980 266.050 46.280 266.500 ;
        RECT 45.980 265.300 46.280 265.750 ;
        RECT 63.180 274.300 63.480 274.750 ;
        RECT 63.180 273.550 63.480 274.000 ;
        RECT 63.180 272.800 63.480 273.250 ;
        RECT 63.180 272.050 63.480 272.500 ;
        RECT 63.180 271.300 63.480 271.750 ;
        RECT 63.180 270.550 63.480 271.000 ;
        RECT 63.180 269.800 63.480 270.250 ;
        RECT 63.180 269.050 63.480 269.500 ;
        RECT 63.180 268.300 63.480 268.750 ;
        RECT 63.180 267.550 63.480 268.000 ;
        RECT 63.180 266.800 63.480 267.250 ;
        RECT 63.180 266.050 63.480 266.500 ;
        RECT 63.180 265.300 63.480 265.750 ;
        RECT 65.980 274.300 66.280 274.750 ;
        RECT 65.980 273.550 66.280 274.000 ;
        RECT 65.980 272.800 66.280 273.250 ;
        RECT 65.980 272.050 66.280 272.500 ;
        RECT 65.980 271.300 66.280 271.750 ;
        RECT 65.980 270.550 66.280 271.000 ;
        RECT 65.980 269.800 66.280 270.250 ;
        RECT 65.980 269.050 66.280 269.500 ;
        RECT 65.980 268.300 66.280 268.750 ;
        RECT 65.980 267.550 66.280 268.000 ;
        RECT 65.980 266.800 66.280 267.250 ;
        RECT 65.980 266.050 66.280 266.500 ;
        RECT 65.980 265.300 66.280 265.750 ;
        RECT 83.180 274.300 83.480 274.750 ;
        RECT 83.180 273.550 83.480 274.000 ;
        RECT 83.180 272.800 83.480 273.250 ;
        RECT 83.180 272.050 83.480 272.500 ;
        RECT 83.180 271.300 83.480 271.750 ;
        RECT 83.180 270.550 83.480 271.000 ;
        RECT 83.180 269.800 83.480 270.250 ;
        RECT 83.180 269.050 83.480 269.500 ;
        RECT 83.180 268.300 83.480 268.750 ;
        RECT 83.180 267.550 83.480 268.000 ;
        RECT 83.180 266.800 83.480 267.250 ;
        RECT 83.180 266.050 83.480 266.500 ;
        RECT 83.180 265.300 83.480 265.750 ;
        RECT 85.980 274.300 86.280 274.750 ;
        RECT 85.980 273.550 86.280 274.000 ;
        RECT 85.980 272.800 86.280 273.250 ;
        RECT 85.980 272.050 86.280 272.500 ;
        RECT 85.980 271.300 86.280 271.750 ;
        RECT 85.980 270.550 86.280 271.000 ;
        RECT 85.980 269.800 86.280 270.250 ;
        RECT 85.980 269.050 86.280 269.500 ;
        RECT 85.980 268.300 86.280 268.750 ;
        RECT 85.980 267.550 86.280 268.000 ;
        RECT 85.980 266.800 86.280 267.250 ;
        RECT 85.980 266.050 86.280 266.500 ;
        RECT 85.980 265.300 86.280 265.750 ;
        RECT 103.180 274.300 103.480 274.750 ;
        RECT 103.180 273.550 103.480 274.000 ;
        RECT 103.180 272.800 103.480 273.250 ;
        RECT 103.180 272.050 103.480 272.500 ;
        RECT 103.180 271.300 103.480 271.750 ;
        RECT 103.180 270.550 103.480 271.000 ;
        RECT 103.180 269.800 103.480 270.250 ;
        RECT 103.180 269.050 103.480 269.500 ;
        RECT 103.180 268.300 103.480 268.750 ;
        RECT 103.180 267.550 103.480 268.000 ;
        RECT 103.180 266.800 103.480 267.250 ;
        RECT 103.180 266.050 103.480 266.500 ;
        RECT 103.180 265.300 103.480 265.750 ;
        RECT 105.980 274.300 106.280 274.750 ;
        RECT 105.980 273.550 106.280 274.000 ;
        RECT 105.980 272.800 106.280 273.250 ;
        RECT 105.980 272.050 106.280 272.500 ;
        RECT 105.980 271.300 106.280 271.750 ;
        RECT 105.980 270.550 106.280 271.000 ;
        RECT 105.980 269.800 106.280 270.250 ;
        RECT 105.980 269.050 106.280 269.500 ;
        RECT 105.980 268.300 106.280 268.750 ;
        RECT 105.980 267.550 106.280 268.000 ;
        RECT 105.980 266.800 106.280 267.250 ;
        RECT 105.980 266.050 106.280 266.500 ;
        RECT 105.980 265.300 106.280 265.750 ;
        RECT 123.180 274.300 123.480 274.750 ;
        RECT 123.180 273.550 123.480 274.000 ;
        RECT 123.180 272.800 123.480 273.250 ;
        RECT 123.180 272.050 123.480 272.500 ;
        RECT 123.180 271.300 123.480 271.750 ;
        RECT 123.180 270.550 123.480 271.000 ;
        RECT 123.180 269.800 123.480 270.250 ;
        RECT 123.180 269.050 123.480 269.500 ;
        RECT 123.180 268.300 123.480 268.750 ;
        RECT 123.180 267.550 123.480 268.000 ;
        RECT 123.180 266.800 123.480 267.250 ;
        RECT 123.180 266.050 123.480 266.500 ;
        RECT 123.180 265.300 123.480 265.750 ;
        RECT 5.980 254.300 6.280 254.750 ;
        RECT 5.980 253.550 6.280 254.000 ;
        RECT 5.980 252.800 6.280 253.250 ;
        RECT 5.980 252.050 6.280 252.500 ;
        RECT 5.980 251.300 6.280 251.750 ;
        RECT 5.980 250.550 6.280 251.000 ;
        RECT 5.980 249.800 6.280 250.250 ;
        RECT 5.980 249.050 6.280 249.500 ;
        RECT 5.980 248.300 6.280 248.750 ;
        RECT 5.980 247.550 6.280 248.000 ;
        RECT 5.980 246.800 6.280 247.250 ;
        RECT 5.980 246.050 6.280 246.500 ;
        RECT 5.980 245.300 6.280 245.750 ;
        RECT 23.180 254.300 23.480 254.750 ;
        RECT 23.180 253.550 23.480 254.000 ;
        RECT 23.180 252.800 23.480 253.250 ;
        RECT 23.180 252.050 23.480 252.500 ;
        RECT 23.180 251.300 23.480 251.750 ;
        RECT 23.180 250.550 23.480 251.000 ;
        RECT 23.180 249.800 23.480 250.250 ;
        RECT 23.180 249.050 23.480 249.500 ;
        RECT 23.180 248.300 23.480 248.750 ;
        RECT 23.180 247.550 23.480 248.000 ;
        RECT 23.180 246.800 23.480 247.250 ;
        RECT 23.180 246.050 23.480 246.500 ;
        RECT 23.180 245.300 23.480 245.750 ;
        RECT 25.980 254.300 26.280 254.750 ;
        RECT 25.980 253.550 26.280 254.000 ;
        RECT 25.980 252.800 26.280 253.250 ;
        RECT 25.980 252.050 26.280 252.500 ;
        RECT 25.980 251.300 26.280 251.750 ;
        RECT 25.980 250.550 26.280 251.000 ;
        RECT 25.980 249.800 26.280 250.250 ;
        RECT 25.980 249.050 26.280 249.500 ;
        RECT 25.980 248.300 26.280 248.750 ;
        RECT 25.980 247.550 26.280 248.000 ;
        RECT 25.980 246.800 26.280 247.250 ;
        RECT 25.980 246.050 26.280 246.500 ;
        RECT 25.980 245.300 26.280 245.750 ;
        RECT 43.180 254.300 43.480 254.750 ;
        RECT 43.180 253.550 43.480 254.000 ;
        RECT 43.180 252.800 43.480 253.250 ;
        RECT 43.180 252.050 43.480 252.500 ;
        RECT 43.180 251.300 43.480 251.750 ;
        RECT 43.180 250.550 43.480 251.000 ;
        RECT 43.180 249.800 43.480 250.250 ;
        RECT 43.180 249.050 43.480 249.500 ;
        RECT 43.180 248.300 43.480 248.750 ;
        RECT 43.180 247.550 43.480 248.000 ;
        RECT 43.180 246.800 43.480 247.250 ;
        RECT 43.180 246.050 43.480 246.500 ;
        RECT 43.180 245.300 43.480 245.750 ;
        RECT 45.980 254.300 46.280 254.750 ;
        RECT 45.980 253.550 46.280 254.000 ;
        RECT 45.980 252.800 46.280 253.250 ;
        RECT 45.980 252.050 46.280 252.500 ;
        RECT 45.980 251.300 46.280 251.750 ;
        RECT 45.980 250.550 46.280 251.000 ;
        RECT 45.980 249.800 46.280 250.250 ;
        RECT 45.980 249.050 46.280 249.500 ;
        RECT 45.980 248.300 46.280 248.750 ;
        RECT 45.980 247.550 46.280 248.000 ;
        RECT 45.980 246.800 46.280 247.250 ;
        RECT 45.980 246.050 46.280 246.500 ;
        RECT 45.980 245.300 46.280 245.750 ;
        RECT 63.180 254.300 63.480 254.750 ;
        RECT 63.180 253.550 63.480 254.000 ;
        RECT 63.180 252.800 63.480 253.250 ;
        RECT 63.180 252.050 63.480 252.500 ;
        RECT 63.180 251.300 63.480 251.750 ;
        RECT 63.180 250.550 63.480 251.000 ;
        RECT 63.180 249.800 63.480 250.250 ;
        RECT 63.180 249.050 63.480 249.500 ;
        RECT 63.180 248.300 63.480 248.750 ;
        RECT 63.180 247.550 63.480 248.000 ;
        RECT 63.180 246.800 63.480 247.250 ;
        RECT 63.180 246.050 63.480 246.500 ;
        RECT 63.180 245.300 63.480 245.750 ;
        RECT 65.980 254.300 66.280 254.750 ;
        RECT 65.980 253.550 66.280 254.000 ;
        RECT 65.980 252.800 66.280 253.250 ;
        RECT 65.980 252.050 66.280 252.500 ;
        RECT 65.980 251.300 66.280 251.750 ;
        RECT 65.980 250.550 66.280 251.000 ;
        RECT 65.980 249.800 66.280 250.250 ;
        RECT 65.980 249.050 66.280 249.500 ;
        RECT 65.980 248.300 66.280 248.750 ;
        RECT 65.980 247.550 66.280 248.000 ;
        RECT 65.980 246.800 66.280 247.250 ;
        RECT 65.980 246.050 66.280 246.500 ;
        RECT 65.980 245.300 66.280 245.750 ;
        RECT 83.180 254.300 83.480 254.750 ;
        RECT 83.180 253.550 83.480 254.000 ;
        RECT 83.180 252.800 83.480 253.250 ;
        RECT 83.180 252.050 83.480 252.500 ;
        RECT 83.180 251.300 83.480 251.750 ;
        RECT 83.180 250.550 83.480 251.000 ;
        RECT 83.180 249.800 83.480 250.250 ;
        RECT 83.180 249.050 83.480 249.500 ;
        RECT 83.180 248.300 83.480 248.750 ;
        RECT 83.180 247.550 83.480 248.000 ;
        RECT 83.180 246.800 83.480 247.250 ;
        RECT 83.180 246.050 83.480 246.500 ;
        RECT 83.180 245.300 83.480 245.750 ;
        RECT 85.980 254.300 86.280 254.750 ;
        RECT 85.980 253.550 86.280 254.000 ;
        RECT 85.980 252.800 86.280 253.250 ;
        RECT 85.980 252.050 86.280 252.500 ;
        RECT 85.980 251.300 86.280 251.750 ;
        RECT 85.980 250.550 86.280 251.000 ;
        RECT 85.980 249.800 86.280 250.250 ;
        RECT 85.980 249.050 86.280 249.500 ;
        RECT 85.980 248.300 86.280 248.750 ;
        RECT 85.980 247.550 86.280 248.000 ;
        RECT 85.980 246.800 86.280 247.250 ;
        RECT 85.980 246.050 86.280 246.500 ;
        RECT 85.980 245.300 86.280 245.750 ;
        RECT 103.180 254.300 103.480 254.750 ;
        RECT 103.180 253.550 103.480 254.000 ;
        RECT 103.180 252.800 103.480 253.250 ;
        RECT 103.180 252.050 103.480 252.500 ;
        RECT 103.180 251.300 103.480 251.750 ;
        RECT 103.180 250.550 103.480 251.000 ;
        RECT 103.180 249.800 103.480 250.250 ;
        RECT 103.180 249.050 103.480 249.500 ;
        RECT 103.180 248.300 103.480 248.750 ;
        RECT 103.180 247.550 103.480 248.000 ;
        RECT 103.180 246.800 103.480 247.250 ;
        RECT 103.180 246.050 103.480 246.500 ;
        RECT 103.180 245.300 103.480 245.750 ;
        RECT 105.980 254.300 106.280 254.750 ;
        RECT 105.980 253.550 106.280 254.000 ;
        RECT 105.980 252.800 106.280 253.250 ;
        RECT 105.980 252.050 106.280 252.500 ;
        RECT 105.980 251.300 106.280 251.750 ;
        RECT 105.980 250.550 106.280 251.000 ;
        RECT 105.980 249.800 106.280 250.250 ;
        RECT 105.980 249.050 106.280 249.500 ;
        RECT 105.980 248.300 106.280 248.750 ;
        RECT 105.980 247.550 106.280 248.000 ;
        RECT 105.980 246.800 106.280 247.250 ;
        RECT 105.980 246.050 106.280 246.500 ;
        RECT 105.980 245.300 106.280 245.750 ;
        RECT 123.180 254.300 123.480 254.750 ;
        RECT 123.180 253.550 123.480 254.000 ;
        RECT 123.180 252.800 123.480 253.250 ;
        RECT 123.180 252.050 123.480 252.500 ;
        RECT 123.180 251.300 123.480 251.750 ;
        RECT 123.180 250.550 123.480 251.000 ;
        RECT 123.180 249.800 123.480 250.250 ;
        RECT 123.180 249.050 123.480 249.500 ;
        RECT 123.180 248.300 123.480 248.750 ;
        RECT 123.180 247.550 123.480 248.000 ;
        RECT 123.180 246.800 123.480 247.250 ;
        RECT 123.180 246.050 123.480 246.500 ;
        RECT 123.180 245.300 123.480 245.750 ;
        RECT 5.980 234.300 6.280 234.750 ;
        RECT 5.980 233.550 6.280 234.000 ;
        RECT 5.980 232.800 6.280 233.250 ;
        RECT 5.980 232.050 6.280 232.500 ;
        RECT 5.980 231.300 6.280 231.750 ;
        RECT 5.980 230.550 6.280 231.000 ;
        RECT 5.980 229.800 6.280 230.250 ;
        RECT 5.980 229.050 6.280 229.500 ;
        RECT 5.980 228.300 6.280 228.750 ;
        RECT 5.980 227.550 6.280 228.000 ;
        RECT 5.980 226.800 6.280 227.250 ;
        RECT 5.980 226.050 6.280 226.500 ;
        RECT 5.980 225.300 6.280 225.750 ;
        RECT 23.180 234.300 23.480 234.750 ;
        RECT 23.180 233.550 23.480 234.000 ;
        RECT 23.180 232.800 23.480 233.250 ;
        RECT 23.180 232.050 23.480 232.500 ;
        RECT 23.180 231.300 23.480 231.750 ;
        RECT 23.180 230.550 23.480 231.000 ;
        RECT 23.180 229.800 23.480 230.250 ;
        RECT 23.180 229.050 23.480 229.500 ;
        RECT 23.180 228.300 23.480 228.750 ;
        RECT 23.180 227.550 23.480 228.000 ;
        RECT 23.180 226.800 23.480 227.250 ;
        RECT 23.180 226.050 23.480 226.500 ;
        RECT 23.180 225.300 23.480 225.750 ;
        RECT 25.980 234.300 26.280 234.750 ;
        RECT 25.980 233.550 26.280 234.000 ;
        RECT 25.980 232.800 26.280 233.250 ;
        RECT 25.980 232.050 26.280 232.500 ;
        RECT 25.980 231.300 26.280 231.750 ;
        RECT 25.980 230.550 26.280 231.000 ;
        RECT 25.980 229.800 26.280 230.250 ;
        RECT 25.980 229.050 26.280 229.500 ;
        RECT 25.980 228.300 26.280 228.750 ;
        RECT 25.980 227.550 26.280 228.000 ;
        RECT 25.980 226.800 26.280 227.250 ;
        RECT 25.980 226.050 26.280 226.500 ;
        RECT 25.980 225.300 26.280 225.750 ;
        RECT 43.180 234.300 43.480 234.750 ;
        RECT 43.180 233.550 43.480 234.000 ;
        RECT 43.180 232.800 43.480 233.250 ;
        RECT 43.180 232.050 43.480 232.500 ;
        RECT 43.180 231.300 43.480 231.750 ;
        RECT 43.180 230.550 43.480 231.000 ;
        RECT 43.180 229.800 43.480 230.250 ;
        RECT 43.180 229.050 43.480 229.500 ;
        RECT 43.180 228.300 43.480 228.750 ;
        RECT 43.180 227.550 43.480 228.000 ;
        RECT 43.180 226.800 43.480 227.250 ;
        RECT 43.180 226.050 43.480 226.500 ;
        RECT 43.180 225.300 43.480 225.750 ;
        RECT 45.980 234.300 46.280 234.750 ;
        RECT 45.980 233.550 46.280 234.000 ;
        RECT 45.980 232.800 46.280 233.250 ;
        RECT 45.980 232.050 46.280 232.500 ;
        RECT 45.980 231.300 46.280 231.750 ;
        RECT 45.980 230.550 46.280 231.000 ;
        RECT 45.980 229.800 46.280 230.250 ;
        RECT 45.980 229.050 46.280 229.500 ;
        RECT 45.980 228.300 46.280 228.750 ;
        RECT 45.980 227.550 46.280 228.000 ;
        RECT 45.980 226.800 46.280 227.250 ;
        RECT 45.980 226.050 46.280 226.500 ;
        RECT 45.980 225.300 46.280 225.750 ;
        RECT 63.180 234.300 63.480 234.750 ;
        RECT 63.180 233.550 63.480 234.000 ;
        RECT 63.180 232.800 63.480 233.250 ;
        RECT 63.180 232.050 63.480 232.500 ;
        RECT 63.180 231.300 63.480 231.750 ;
        RECT 63.180 230.550 63.480 231.000 ;
        RECT 63.180 229.800 63.480 230.250 ;
        RECT 63.180 229.050 63.480 229.500 ;
        RECT 63.180 228.300 63.480 228.750 ;
        RECT 63.180 227.550 63.480 228.000 ;
        RECT 63.180 226.800 63.480 227.250 ;
        RECT 63.180 226.050 63.480 226.500 ;
        RECT 63.180 225.300 63.480 225.750 ;
        RECT 65.980 234.300 66.280 234.750 ;
        RECT 65.980 233.550 66.280 234.000 ;
        RECT 65.980 232.800 66.280 233.250 ;
        RECT 65.980 232.050 66.280 232.500 ;
        RECT 65.980 231.300 66.280 231.750 ;
        RECT 65.980 230.550 66.280 231.000 ;
        RECT 65.980 229.800 66.280 230.250 ;
        RECT 65.980 229.050 66.280 229.500 ;
        RECT 65.980 228.300 66.280 228.750 ;
        RECT 65.980 227.550 66.280 228.000 ;
        RECT 65.980 226.800 66.280 227.250 ;
        RECT 65.980 226.050 66.280 226.500 ;
        RECT 65.980 225.300 66.280 225.750 ;
        RECT 83.180 234.300 83.480 234.750 ;
        RECT 83.180 233.550 83.480 234.000 ;
        RECT 83.180 232.800 83.480 233.250 ;
        RECT 83.180 232.050 83.480 232.500 ;
        RECT 83.180 231.300 83.480 231.750 ;
        RECT 83.180 230.550 83.480 231.000 ;
        RECT 83.180 229.800 83.480 230.250 ;
        RECT 83.180 229.050 83.480 229.500 ;
        RECT 83.180 228.300 83.480 228.750 ;
        RECT 83.180 227.550 83.480 228.000 ;
        RECT 83.180 226.800 83.480 227.250 ;
        RECT 83.180 226.050 83.480 226.500 ;
        RECT 83.180 225.300 83.480 225.750 ;
        RECT 85.980 234.300 86.280 234.750 ;
        RECT 85.980 233.550 86.280 234.000 ;
        RECT 85.980 232.800 86.280 233.250 ;
        RECT 85.980 232.050 86.280 232.500 ;
        RECT 85.980 231.300 86.280 231.750 ;
        RECT 85.980 230.550 86.280 231.000 ;
        RECT 85.980 229.800 86.280 230.250 ;
        RECT 85.980 229.050 86.280 229.500 ;
        RECT 85.980 228.300 86.280 228.750 ;
        RECT 85.980 227.550 86.280 228.000 ;
        RECT 85.980 226.800 86.280 227.250 ;
        RECT 85.980 226.050 86.280 226.500 ;
        RECT 85.980 225.300 86.280 225.750 ;
        RECT 103.180 234.300 103.480 234.750 ;
        RECT 103.180 233.550 103.480 234.000 ;
        RECT 103.180 232.800 103.480 233.250 ;
        RECT 103.180 232.050 103.480 232.500 ;
        RECT 103.180 231.300 103.480 231.750 ;
        RECT 103.180 230.550 103.480 231.000 ;
        RECT 103.180 229.800 103.480 230.250 ;
        RECT 103.180 229.050 103.480 229.500 ;
        RECT 103.180 228.300 103.480 228.750 ;
        RECT 103.180 227.550 103.480 228.000 ;
        RECT 103.180 226.800 103.480 227.250 ;
        RECT 103.180 226.050 103.480 226.500 ;
        RECT 103.180 225.300 103.480 225.750 ;
        RECT 105.980 234.300 106.280 234.750 ;
        RECT 105.980 233.550 106.280 234.000 ;
        RECT 105.980 232.800 106.280 233.250 ;
        RECT 105.980 232.050 106.280 232.500 ;
        RECT 105.980 231.300 106.280 231.750 ;
        RECT 105.980 230.550 106.280 231.000 ;
        RECT 105.980 229.800 106.280 230.250 ;
        RECT 105.980 229.050 106.280 229.500 ;
        RECT 105.980 228.300 106.280 228.750 ;
        RECT 105.980 227.550 106.280 228.000 ;
        RECT 105.980 226.800 106.280 227.250 ;
        RECT 105.980 226.050 106.280 226.500 ;
        RECT 105.980 225.300 106.280 225.750 ;
        RECT 123.180 234.300 123.480 234.750 ;
        RECT 123.180 233.550 123.480 234.000 ;
        RECT 123.180 232.800 123.480 233.250 ;
        RECT 123.180 232.050 123.480 232.500 ;
        RECT 123.180 231.300 123.480 231.750 ;
        RECT 123.180 230.550 123.480 231.000 ;
        RECT 123.180 229.800 123.480 230.250 ;
        RECT 123.180 229.050 123.480 229.500 ;
        RECT 123.180 228.300 123.480 228.750 ;
        RECT 123.180 227.550 123.480 228.000 ;
        RECT 123.180 226.800 123.480 227.250 ;
        RECT 123.180 226.050 123.480 226.500 ;
        RECT 123.180 225.300 123.480 225.750 ;
        RECT 5.980 214.300 6.280 214.750 ;
        RECT 5.980 213.550 6.280 214.000 ;
        RECT 5.980 212.800 6.280 213.250 ;
        RECT 5.980 212.050 6.280 212.500 ;
        RECT 5.980 211.300 6.280 211.750 ;
        RECT 5.980 210.550 6.280 211.000 ;
        RECT 5.980 209.800 6.280 210.250 ;
        RECT 5.980 209.050 6.280 209.500 ;
        RECT 5.980 208.300 6.280 208.750 ;
        RECT 5.980 207.550 6.280 208.000 ;
        RECT 5.980 206.800 6.280 207.250 ;
        RECT 5.980 206.050 6.280 206.500 ;
        RECT 5.980 205.300 6.280 205.750 ;
        RECT 23.180 214.300 23.480 214.750 ;
        RECT 23.180 213.550 23.480 214.000 ;
        RECT 23.180 212.800 23.480 213.250 ;
        RECT 23.180 212.050 23.480 212.500 ;
        RECT 23.180 211.300 23.480 211.750 ;
        RECT 23.180 210.550 23.480 211.000 ;
        RECT 23.180 209.800 23.480 210.250 ;
        RECT 23.180 209.050 23.480 209.500 ;
        RECT 23.180 208.300 23.480 208.750 ;
        RECT 23.180 207.550 23.480 208.000 ;
        RECT 23.180 206.800 23.480 207.250 ;
        RECT 23.180 206.050 23.480 206.500 ;
        RECT 23.180 205.300 23.480 205.750 ;
        RECT 25.980 214.300 26.280 214.750 ;
        RECT 25.980 213.550 26.280 214.000 ;
        RECT 25.980 212.800 26.280 213.250 ;
        RECT 25.980 212.050 26.280 212.500 ;
        RECT 25.980 211.300 26.280 211.750 ;
        RECT 25.980 210.550 26.280 211.000 ;
        RECT 25.980 209.800 26.280 210.250 ;
        RECT 25.980 209.050 26.280 209.500 ;
        RECT 25.980 208.300 26.280 208.750 ;
        RECT 25.980 207.550 26.280 208.000 ;
        RECT 25.980 206.800 26.280 207.250 ;
        RECT 25.980 206.050 26.280 206.500 ;
        RECT 25.980 205.300 26.280 205.750 ;
        RECT 43.180 214.300 43.480 214.750 ;
        RECT 43.180 213.550 43.480 214.000 ;
        RECT 43.180 212.800 43.480 213.250 ;
        RECT 43.180 212.050 43.480 212.500 ;
        RECT 43.180 211.300 43.480 211.750 ;
        RECT 43.180 210.550 43.480 211.000 ;
        RECT 43.180 209.800 43.480 210.250 ;
        RECT 43.180 209.050 43.480 209.500 ;
        RECT 43.180 208.300 43.480 208.750 ;
        RECT 43.180 207.550 43.480 208.000 ;
        RECT 43.180 206.800 43.480 207.250 ;
        RECT 43.180 206.050 43.480 206.500 ;
        RECT 43.180 205.300 43.480 205.750 ;
        RECT 45.980 214.300 46.280 214.750 ;
        RECT 45.980 213.550 46.280 214.000 ;
        RECT 45.980 212.800 46.280 213.250 ;
        RECT 45.980 212.050 46.280 212.500 ;
        RECT 45.980 211.300 46.280 211.750 ;
        RECT 45.980 210.550 46.280 211.000 ;
        RECT 45.980 209.800 46.280 210.250 ;
        RECT 45.980 209.050 46.280 209.500 ;
        RECT 45.980 208.300 46.280 208.750 ;
        RECT 45.980 207.550 46.280 208.000 ;
        RECT 45.980 206.800 46.280 207.250 ;
        RECT 45.980 206.050 46.280 206.500 ;
        RECT 45.980 205.300 46.280 205.750 ;
        RECT 63.180 214.300 63.480 214.750 ;
        RECT 63.180 213.550 63.480 214.000 ;
        RECT 63.180 212.800 63.480 213.250 ;
        RECT 63.180 212.050 63.480 212.500 ;
        RECT 63.180 211.300 63.480 211.750 ;
        RECT 63.180 210.550 63.480 211.000 ;
        RECT 63.180 209.800 63.480 210.250 ;
        RECT 63.180 209.050 63.480 209.500 ;
        RECT 63.180 208.300 63.480 208.750 ;
        RECT 63.180 207.550 63.480 208.000 ;
        RECT 63.180 206.800 63.480 207.250 ;
        RECT 63.180 206.050 63.480 206.500 ;
        RECT 63.180 205.300 63.480 205.750 ;
        RECT 65.980 214.300 66.280 214.750 ;
        RECT 65.980 213.550 66.280 214.000 ;
        RECT 65.980 212.800 66.280 213.250 ;
        RECT 65.980 212.050 66.280 212.500 ;
        RECT 65.980 211.300 66.280 211.750 ;
        RECT 65.980 210.550 66.280 211.000 ;
        RECT 65.980 209.800 66.280 210.250 ;
        RECT 65.980 209.050 66.280 209.500 ;
        RECT 65.980 208.300 66.280 208.750 ;
        RECT 65.980 207.550 66.280 208.000 ;
        RECT 65.980 206.800 66.280 207.250 ;
        RECT 65.980 206.050 66.280 206.500 ;
        RECT 65.980 205.300 66.280 205.750 ;
        RECT 83.180 214.300 83.480 214.750 ;
        RECT 83.180 213.550 83.480 214.000 ;
        RECT 83.180 212.800 83.480 213.250 ;
        RECT 83.180 212.050 83.480 212.500 ;
        RECT 83.180 211.300 83.480 211.750 ;
        RECT 83.180 210.550 83.480 211.000 ;
        RECT 83.180 209.800 83.480 210.250 ;
        RECT 83.180 209.050 83.480 209.500 ;
        RECT 83.180 208.300 83.480 208.750 ;
        RECT 83.180 207.550 83.480 208.000 ;
        RECT 83.180 206.800 83.480 207.250 ;
        RECT 83.180 206.050 83.480 206.500 ;
        RECT 83.180 205.300 83.480 205.750 ;
        RECT 85.980 214.300 86.280 214.750 ;
        RECT 85.980 213.550 86.280 214.000 ;
        RECT 85.980 212.800 86.280 213.250 ;
        RECT 85.980 212.050 86.280 212.500 ;
        RECT 85.980 211.300 86.280 211.750 ;
        RECT 85.980 210.550 86.280 211.000 ;
        RECT 85.980 209.800 86.280 210.250 ;
        RECT 85.980 209.050 86.280 209.500 ;
        RECT 85.980 208.300 86.280 208.750 ;
        RECT 85.980 207.550 86.280 208.000 ;
        RECT 85.980 206.800 86.280 207.250 ;
        RECT 85.980 206.050 86.280 206.500 ;
        RECT 85.980 205.300 86.280 205.750 ;
        RECT 103.180 214.300 103.480 214.750 ;
        RECT 103.180 213.550 103.480 214.000 ;
        RECT 103.180 212.800 103.480 213.250 ;
        RECT 103.180 212.050 103.480 212.500 ;
        RECT 103.180 211.300 103.480 211.750 ;
        RECT 103.180 210.550 103.480 211.000 ;
        RECT 103.180 209.800 103.480 210.250 ;
        RECT 103.180 209.050 103.480 209.500 ;
        RECT 103.180 208.300 103.480 208.750 ;
        RECT 103.180 207.550 103.480 208.000 ;
        RECT 103.180 206.800 103.480 207.250 ;
        RECT 103.180 206.050 103.480 206.500 ;
        RECT 103.180 205.300 103.480 205.750 ;
        RECT 105.980 214.300 106.280 214.750 ;
        RECT 105.980 213.550 106.280 214.000 ;
        RECT 105.980 212.800 106.280 213.250 ;
        RECT 105.980 212.050 106.280 212.500 ;
        RECT 105.980 211.300 106.280 211.750 ;
        RECT 105.980 210.550 106.280 211.000 ;
        RECT 105.980 209.800 106.280 210.250 ;
        RECT 105.980 209.050 106.280 209.500 ;
        RECT 105.980 208.300 106.280 208.750 ;
        RECT 105.980 207.550 106.280 208.000 ;
        RECT 105.980 206.800 106.280 207.250 ;
        RECT 105.980 206.050 106.280 206.500 ;
        RECT 105.980 205.300 106.280 205.750 ;
        RECT 123.180 214.300 123.480 214.750 ;
        RECT 123.180 213.550 123.480 214.000 ;
        RECT 123.180 212.800 123.480 213.250 ;
        RECT 123.180 212.050 123.480 212.500 ;
        RECT 123.180 211.300 123.480 211.750 ;
        RECT 123.180 210.550 123.480 211.000 ;
        RECT 123.180 209.800 123.480 210.250 ;
        RECT 123.180 209.050 123.480 209.500 ;
        RECT 123.180 208.300 123.480 208.750 ;
        RECT 123.180 207.550 123.480 208.000 ;
        RECT 123.180 206.800 123.480 207.250 ;
        RECT 123.180 206.050 123.480 206.500 ;
        RECT 123.180 205.300 123.480 205.750 ;
        RECT 9.425 176.405 10.015 176.975 ;
        RECT 10.205 176.405 10.795 176.975 ;
        RECT 10.985 176.405 11.575 176.975 ;
        RECT 10.175 174.445 10.345 174.720 ;
        RECT 11.755 174.445 11.925 174.720 ;
        RECT 12.395 174.445 12.570 174.745 ;
        RECT 13.985 174.450 14.155 174.745 ;
        RECT 5.980 134.300 6.280 134.750 ;
        RECT 5.980 133.550 6.280 134.000 ;
        RECT 5.980 132.800 6.280 133.250 ;
        RECT 5.980 132.050 6.280 132.500 ;
        RECT 5.980 131.300 6.280 131.750 ;
        RECT 5.980 130.550 6.280 131.000 ;
        RECT 5.980 129.800 6.280 130.250 ;
        RECT 5.980 129.050 6.280 129.500 ;
        RECT 5.980 128.300 6.280 128.750 ;
        RECT 5.980 127.550 6.280 128.000 ;
        RECT 5.980 126.800 6.280 127.250 ;
        RECT 5.980 126.050 6.280 126.500 ;
        RECT 5.980 125.300 6.280 125.750 ;
        RECT 23.180 134.300 23.480 134.750 ;
        RECT 23.180 133.550 23.480 134.000 ;
        RECT 23.180 132.800 23.480 133.250 ;
        RECT 23.180 132.050 23.480 132.500 ;
        RECT 23.180 131.300 23.480 131.750 ;
        RECT 23.180 130.550 23.480 131.000 ;
        RECT 23.180 129.800 23.480 130.250 ;
        RECT 23.180 129.050 23.480 129.500 ;
        RECT 23.180 128.300 23.480 128.750 ;
        RECT 23.180 127.550 23.480 128.000 ;
        RECT 23.180 126.800 23.480 127.250 ;
        RECT 23.180 126.050 23.480 126.500 ;
        RECT 23.180 125.300 23.480 125.750 ;
        RECT 25.980 134.300 26.280 134.750 ;
        RECT 25.980 133.550 26.280 134.000 ;
        RECT 25.980 132.800 26.280 133.250 ;
        RECT 25.980 132.050 26.280 132.500 ;
        RECT 25.980 131.300 26.280 131.750 ;
        RECT 25.980 130.550 26.280 131.000 ;
        RECT 25.980 129.800 26.280 130.250 ;
        RECT 25.980 129.050 26.280 129.500 ;
        RECT 25.980 128.300 26.280 128.750 ;
        RECT 25.980 127.550 26.280 128.000 ;
        RECT 25.980 126.800 26.280 127.250 ;
        RECT 25.980 126.050 26.280 126.500 ;
        RECT 25.980 125.300 26.280 125.750 ;
        RECT 43.180 134.300 43.480 134.750 ;
        RECT 43.180 133.550 43.480 134.000 ;
        RECT 43.180 132.800 43.480 133.250 ;
        RECT 43.180 132.050 43.480 132.500 ;
        RECT 43.180 131.300 43.480 131.750 ;
        RECT 43.180 130.550 43.480 131.000 ;
        RECT 43.180 129.800 43.480 130.250 ;
        RECT 43.180 129.050 43.480 129.500 ;
        RECT 43.180 128.300 43.480 128.750 ;
        RECT 43.180 127.550 43.480 128.000 ;
        RECT 43.180 126.800 43.480 127.250 ;
        RECT 43.180 126.050 43.480 126.500 ;
        RECT 43.180 125.300 43.480 125.750 ;
        RECT 45.980 134.300 46.280 134.750 ;
        RECT 45.980 133.550 46.280 134.000 ;
        RECT 45.980 132.800 46.280 133.250 ;
        RECT 45.980 132.050 46.280 132.500 ;
        RECT 45.980 131.300 46.280 131.750 ;
        RECT 45.980 130.550 46.280 131.000 ;
        RECT 45.980 129.800 46.280 130.250 ;
        RECT 45.980 129.050 46.280 129.500 ;
        RECT 45.980 128.300 46.280 128.750 ;
        RECT 45.980 127.550 46.280 128.000 ;
        RECT 45.980 126.800 46.280 127.250 ;
        RECT 45.980 126.050 46.280 126.500 ;
        RECT 45.980 125.300 46.280 125.750 ;
        RECT 63.180 134.300 63.480 134.750 ;
        RECT 63.180 133.550 63.480 134.000 ;
        RECT 63.180 132.800 63.480 133.250 ;
        RECT 63.180 132.050 63.480 132.500 ;
        RECT 63.180 131.300 63.480 131.750 ;
        RECT 63.180 130.550 63.480 131.000 ;
        RECT 63.180 129.800 63.480 130.250 ;
        RECT 63.180 129.050 63.480 129.500 ;
        RECT 63.180 128.300 63.480 128.750 ;
        RECT 63.180 127.550 63.480 128.000 ;
        RECT 63.180 126.800 63.480 127.250 ;
        RECT 63.180 126.050 63.480 126.500 ;
        RECT 63.180 125.300 63.480 125.750 ;
        RECT 65.980 134.300 66.280 134.750 ;
        RECT 65.980 133.550 66.280 134.000 ;
        RECT 65.980 132.800 66.280 133.250 ;
        RECT 65.980 132.050 66.280 132.500 ;
        RECT 65.980 131.300 66.280 131.750 ;
        RECT 65.980 130.550 66.280 131.000 ;
        RECT 65.980 129.800 66.280 130.250 ;
        RECT 65.980 129.050 66.280 129.500 ;
        RECT 65.980 128.300 66.280 128.750 ;
        RECT 65.980 127.550 66.280 128.000 ;
        RECT 65.980 126.800 66.280 127.250 ;
        RECT 65.980 126.050 66.280 126.500 ;
        RECT 65.980 125.300 66.280 125.750 ;
        RECT 83.180 134.300 83.480 134.750 ;
        RECT 83.180 133.550 83.480 134.000 ;
        RECT 83.180 132.800 83.480 133.250 ;
        RECT 83.180 132.050 83.480 132.500 ;
        RECT 83.180 131.300 83.480 131.750 ;
        RECT 83.180 130.550 83.480 131.000 ;
        RECT 83.180 129.800 83.480 130.250 ;
        RECT 83.180 129.050 83.480 129.500 ;
        RECT 83.180 128.300 83.480 128.750 ;
        RECT 83.180 127.550 83.480 128.000 ;
        RECT 83.180 126.800 83.480 127.250 ;
        RECT 83.180 126.050 83.480 126.500 ;
        RECT 83.180 125.300 83.480 125.750 ;
        RECT 85.980 134.300 86.280 134.750 ;
        RECT 85.980 133.550 86.280 134.000 ;
        RECT 85.980 132.800 86.280 133.250 ;
        RECT 85.980 132.050 86.280 132.500 ;
        RECT 85.980 131.300 86.280 131.750 ;
        RECT 85.980 130.550 86.280 131.000 ;
        RECT 85.980 129.800 86.280 130.250 ;
        RECT 85.980 129.050 86.280 129.500 ;
        RECT 85.980 128.300 86.280 128.750 ;
        RECT 85.980 127.550 86.280 128.000 ;
        RECT 85.980 126.800 86.280 127.250 ;
        RECT 85.980 126.050 86.280 126.500 ;
        RECT 85.980 125.300 86.280 125.750 ;
        RECT 103.180 134.300 103.480 134.750 ;
        RECT 103.180 133.550 103.480 134.000 ;
        RECT 103.180 132.800 103.480 133.250 ;
        RECT 103.180 132.050 103.480 132.500 ;
        RECT 103.180 131.300 103.480 131.750 ;
        RECT 103.180 130.550 103.480 131.000 ;
        RECT 103.180 129.800 103.480 130.250 ;
        RECT 103.180 129.050 103.480 129.500 ;
        RECT 103.180 128.300 103.480 128.750 ;
        RECT 103.180 127.550 103.480 128.000 ;
        RECT 103.180 126.800 103.480 127.250 ;
        RECT 103.180 126.050 103.480 126.500 ;
        RECT 103.180 125.300 103.480 125.750 ;
        RECT 105.980 134.300 106.280 134.750 ;
        RECT 105.980 133.550 106.280 134.000 ;
        RECT 105.980 132.800 106.280 133.250 ;
        RECT 105.980 132.050 106.280 132.500 ;
        RECT 105.980 131.300 106.280 131.750 ;
        RECT 105.980 130.550 106.280 131.000 ;
        RECT 105.980 129.800 106.280 130.250 ;
        RECT 105.980 129.050 106.280 129.500 ;
        RECT 105.980 128.300 106.280 128.750 ;
        RECT 105.980 127.550 106.280 128.000 ;
        RECT 105.980 126.800 106.280 127.250 ;
        RECT 105.980 126.050 106.280 126.500 ;
        RECT 105.980 125.300 106.280 125.750 ;
        RECT 123.180 134.300 123.480 134.750 ;
        RECT 123.180 133.550 123.480 134.000 ;
        RECT 123.180 132.800 123.480 133.250 ;
        RECT 123.180 132.050 123.480 132.500 ;
        RECT 123.180 131.300 123.480 131.750 ;
        RECT 123.180 130.550 123.480 131.000 ;
        RECT 123.180 129.800 123.480 130.250 ;
        RECT 123.180 129.050 123.480 129.500 ;
        RECT 123.180 128.300 123.480 128.750 ;
        RECT 123.180 127.550 123.480 128.000 ;
        RECT 123.180 126.800 123.480 127.250 ;
        RECT 123.180 126.050 123.480 126.500 ;
        RECT 123.180 125.300 123.480 125.750 ;
        RECT 5.980 114.300 6.280 114.750 ;
        RECT 5.980 113.550 6.280 114.000 ;
        RECT 5.980 112.800 6.280 113.250 ;
        RECT 5.980 112.050 6.280 112.500 ;
        RECT 5.980 111.300 6.280 111.750 ;
        RECT 5.980 110.550 6.280 111.000 ;
        RECT 5.980 109.800 6.280 110.250 ;
        RECT 5.980 109.050 6.280 109.500 ;
        RECT 5.980 108.300 6.280 108.750 ;
        RECT 5.980 107.550 6.280 108.000 ;
        RECT 5.980 106.800 6.280 107.250 ;
        RECT 5.980 106.050 6.280 106.500 ;
        RECT 5.980 105.300 6.280 105.750 ;
        RECT 23.180 114.300 23.480 114.750 ;
        RECT 23.180 113.550 23.480 114.000 ;
        RECT 23.180 112.800 23.480 113.250 ;
        RECT 23.180 112.050 23.480 112.500 ;
        RECT 23.180 111.300 23.480 111.750 ;
        RECT 23.180 110.550 23.480 111.000 ;
        RECT 23.180 109.800 23.480 110.250 ;
        RECT 23.180 109.050 23.480 109.500 ;
        RECT 23.180 108.300 23.480 108.750 ;
        RECT 23.180 107.550 23.480 108.000 ;
        RECT 23.180 106.800 23.480 107.250 ;
        RECT 23.180 106.050 23.480 106.500 ;
        RECT 23.180 105.300 23.480 105.750 ;
        RECT 25.980 114.300 26.280 114.750 ;
        RECT 25.980 113.550 26.280 114.000 ;
        RECT 25.980 112.800 26.280 113.250 ;
        RECT 25.980 112.050 26.280 112.500 ;
        RECT 25.980 111.300 26.280 111.750 ;
        RECT 25.980 110.550 26.280 111.000 ;
        RECT 25.980 109.800 26.280 110.250 ;
        RECT 25.980 109.050 26.280 109.500 ;
        RECT 25.980 108.300 26.280 108.750 ;
        RECT 25.980 107.550 26.280 108.000 ;
        RECT 25.980 106.800 26.280 107.250 ;
        RECT 25.980 106.050 26.280 106.500 ;
        RECT 25.980 105.300 26.280 105.750 ;
        RECT 43.180 114.300 43.480 114.750 ;
        RECT 43.180 113.550 43.480 114.000 ;
        RECT 43.180 112.800 43.480 113.250 ;
        RECT 43.180 112.050 43.480 112.500 ;
        RECT 43.180 111.300 43.480 111.750 ;
        RECT 43.180 110.550 43.480 111.000 ;
        RECT 43.180 109.800 43.480 110.250 ;
        RECT 43.180 109.050 43.480 109.500 ;
        RECT 43.180 108.300 43.480 108.750 ;
        RECT 43.180 107.550 43.480 108.000 ;
        RECT 43.180 106.800 43.480 107.250 ;
        RECT 43.180 106.050 43.480 106.500 ;
        RECT 43.180 105.300 43.480 105.750 ;
        RECT 45.980 114.300 46.280 114.750 ;
        RECT 45.980 113.550 46.280 114.000 ;
        RECT 45.980 112.800 46.280 113.250 ;
        RECT 45.980 112.050 46.280 112.500 ;
        RECT 45.980 111.300 46.280 111.750 ;
        RECT 45.980 110.550 46.280 111.000 ;
        RECT 45.980 109.800 46.280 110.250 ;
        RECT 45.980 109.050 46.280 109.500 ;
        RECT 45.980 108.300 46.280 108.750 ;
        RECT 45.980 107.550 46.280 108.000 ;
        RECT 45.980 106.800 46.280 107.250 ;
        RECT 45.980 106.050 46.280 106.500 ;
        RECT 45.980 105.300 46.280 105.750 ;
        RECT 63.180 114.300 63.480 114.750 ;
        RECT 63.180 113.550 63.480 114.000 ;
        RECT 63.180 112.800 63.480 113.250 ;
        RECT 63.180 112.050 63.480 112.500 ;
        RECT 63.180 111.300 63.480 111.750 ;
        RECT 63.180 110.550 63.480 111.000 ;
        RECT 63.180 109.800 63.480 110.250 ;
        RECT 63.180 109.050 63.480 109.500 ;
        RECT 63.180 108.300 63.480 108.750 ;
        RECT 63.180 107.550 63.480 108.000 ;
        RECT 63.180 106.800 63.480 107.250 ;
        RECT 63.180 106.050 63.480 106.500 ;
        RECT 63.180 105.300 63.480 105.750 ;
        RECT 65.980 114.300 66.280 114.750 ;
        RECT 65.980 113.550 66.280 114.000 ;
        RECT 65.980 112.800 66.280 113.250 ;
        RECT 65.980 112.050 66.280 112.500 ;
        RECT 65.980 111.300 66.280 111.750 ;
        RECT 65.980 110.550 66.280 111.000 ;
        RECT 65.980 109.800 66.280 110.250 ;
        RECT 65.980 109.050 66.280 109.500 ;
        RECT 65.980 108.300 66.280 108.750 ;
        RECT 65.980 107.550 66.280 108.000 ;
        RECT 65.980 106.800 66.280 107.250 ;
        RECT 65.980 106.050 66.280 106.500 ;
        RECT 65.980 105.300 66.280 105.750 ;
        RECT 83.180 114.300 83.480 114.750 ;
        RECT 83.180 113.550 83.480 114.000 ;
        RECT 83.180 112.800 83.480 113.250 ;
        RECT 83.180 112.050 83.480 112.500 ;
        RECT 83.180 111.300 83.480 111.750 ;
        RECT 83.180 110.550 83.480 111.000 ;
        RECT 83.180 109.800 83.480 110.250 ;
        RECT 83.180 109.050 83.480 109.500 ;
        RECT 83.180 108.300 83.480 108.750 ;
        RECT 83.180 107.550 83.480 108.000 ;
        RECT 83.180 106.800 83.480 107.250 ;
        RECT 83.180 106.050 83.480 106.500 ;
        RECT 83.180 105.300 83.480 105.750 ;
        RECT 85.980 114.300 86.280 114.750 ;
        RECT 85.980 113.550 86.280 114.000 ;
        RECT 85.980 112.800 86.280 113.250 ;
        RECT 85.980 112.050 86.280 112.500 ;
        RECT 85.980 111.300 86.280 111.750 ;
        RECT 85.980 110.550 86.280 111.000 ;
        RECT 85.980 109.800 86.280 110.250 ;
        RECT 85.980 109.050 86.280 109.500 ;
        RECT 85.980 108.300 86.280 108.750 ;
        RECT 85.980 107.550 86.280 108.000 ;
        RECT 85.980 106.800 86.280 107.250 ;
        RECT 85.980 106.050 86.280 106.500 ;
        RECT 85.980 105.300 86.280 105.750 ;
        RECT 103.180 114.300 103.480 114.750 ;
        RECT 103.180 113.550 103.480 114.000 ;
        RECT 103.180 112.800 103.480 113.250 ;
        RECT 103.180 112.050 103.480 112.500 ;
        RECT 103.180 111.300 103.480 111.750 ;
        RECT 103.180 110.550 103.480 111.000 ;
        RECT 103.180 109.800 103.480 110.250 ;
        RECT 103.180 109.050 103.480 109.500 ;
        RECT 103.180 108.300 103.480 108.750 ;
        RECT 103.180 107.550 103.480 108.000 ;
        RECT 103.180 106.800 103.480 107.250 ;
        RECT 103.180 106.050 103.480 106.500 ;
        RECT 103.180 105.300 103.480 105.750 ;
        RECT 105.980 114.300 106.280 114.750 ;
        RECT 105.980 113.550 106.280 114.000 ;
        RECT 105.980 112.800 106.280 113.250 ;
        RECT 105.980 112.050 106.280 112.500 ;
        RECT 105.980 111.300 106.280 111.750 ;
        RECT 105.980 110.550 106.280 111.000 ;
        RECT 105.980 109.800 106.280 110.250 ;
        RECT 105.980 109.050 106.280 109.500 ;
        RECT 105.980 108.300 106.280 108.750 ;
        RECT 105.980 107.550 106.280 108.000 ;
        RECT 105.980 106.800 106.280 107.250 ;
        RECT 105.980 106.050 106.280 106.500 ;
        RECT 105.980 105.300 106.280 105.750 ;
        RECT 123.180 114.300 123.480 114.750 ;
        RECT 123.180 113.550 123.480 114.000 ;
        RECT 123.180 112.800 123.480 113.250 ;
        RECT 123.180 112.050 123.480 112.500 ;
        RECT 123.180 111.300 123.480 111.750 ;
        RECT 123.180 110.550 123.480 111.000 ;
        RECT 123.180 109.800 123.480 110.250 ;
        RECT 123.180 109.050 123.480 109.500 ;
        RECT 123.180 108.300 123.480 108.750 ;
        RECT 123.180 107.550 123.480 108.000 ;
        RECT 123.180 106.800 123.480 107.250 ;
        RECT 123.180 106.050 123.480 106.500 ;
        RECT 123.180 105.300 123.480 105.750 ;
        RECT 5.980 94.300 6.280 94.750 ;
        RECT 5.980 93.550 6.280 94.000 ;
        RECT 5.980 92.800 6.280 93.250 ;
        RECT 5.980 92.050 6.280 92.500 ;
        RECT 5.980 91.300 6.280 91.750 ;
        RECT 5.980 90.550 6.280 91.000 ;
        RECT 5.980 89.800 6.280 90.250 ;
        RECT 5.980 89.050 6.280 89.500 ;
        RECT 5.980 88.300 6.280 88.750 ;
        RECT 5.980 87.550 6.280 88.000 ;
        RECT 5.980 86.800 6.280 87.250 ;
        RECT 5.980 86.050 6.280 86.500 ;
        RECT 5.980 85.300 6.280 85.750 ;
        RECT 23.180 94.300 23.480 94.750 ;
        RECT 23.180 93.550 23.480 94.000 ;
        RECT 23.180 92.800 23.480 93.250 ;
        RECT 23.180 92.050 23.480 92.500 ;
        RECT 23.180 91.300 23.480 91.750 ;
        RECT 23.180 90.550 23.480 91.000 ;
        RECT 23.180 89.800 23.480 90.250 ;
        RECT 23.180 89.050 23.480 89.500 ;
        RECT 23.180 88.300 23.480 88.750 ;
        RECT 23.180 87.550 23.480 88.000 ;
        RECT 23.180 86.800 23.480 87.250 ;
        RECT 23.180 86.050 23.480 86.500 ;
        RECT 23.180 85.300 23.480 85.750 ;
        RECT 25.980 94.300 26.280 94.750 ;
        RECT 25.980 93.550 26.280 94.000 ;
        RECT 25.980 92.800 26.280 93.250 ;
        RECT 25.980 92.050 26.280 92.500 ;
        RECT 25.980 91.300 26.280 91.750 ;
        RECT 25.980 90.550 26.280 91.000 ;
        RECT 25.980 89.800 26.280 90.250 ;
        RECT 25.980 89.050 26.280 89.500 ;
        RECT 25.980 88.300 26.280 88.750 ;
        RECT 25.980 87.550 26.280 88.000 ;
        RECT 25.980 86.800 26.280 87.250 ;
        RECT 25.980 86.050 26.280 86.500 ;
        RECT 25.980 85.300 26.280 85.750 ;
        RECT 43.180 94.300 43.480 94.750 ;
        RECT 43.180 93.550 43.480 94.000 ;
        RECT 43.180 92.800 43.480 93.250 ;
        RECT 43.180 92.050 43.480 92.500 ;
        RECT 43.180 91.300 43.480 91.750 ;
        RECT 43.180 90.550 43.480 91.000 ;
        RECT 43.180 89.800 43.480 90.250 ;
        RECT 43.180 89.050 43.480 89.500 ;
        RECT 43.180 88.300 43.480 88.750 ;
        RECT 43.180 87.550 43.480 88.000 ;
        RECT 43.180 86.800 43.480 87.250 ;
        RECT 43.180 86.050 43.480 86.500 ;
        RECT 43.180 85.300 43.480 85.750 ;
        RECT 45.980 94.300 46.280 94.750 ;
        RECT 45.980 93.550 46.280 94.000 ;
        RECT 45.980 92.800 46.280 93.250 ;
        RECT 45.980 92.050 46.280 92.500 ;
        RECT 45.980 91.300 46.280 91.750 ;
        RECT 45.980 90.550 46.280 91.000 ;
        RECT 45.980 89.800 46.280 90.250 ;
        RECT 45.980 89.050 46.280 89.500 ;
        RECT 45.980 88.300 46.280 88.750 ;
        RECT 45.980 87.550 46.280 88.000 ;
        RECT 45.980 86.800 46.280 87.250 ;
        RECT 45.980 86.050 46.280 86.500 ;
        RECT 45.980 85.300 46.280 85.750 ;
        RECT 63.180 94.300 63.480 94.750 ;
        RECT 63.180 93.550 63.480 94.000 ;
        RECT 63.180 92.800 63.480 93.250 ;
        RECT 63.180 92.050 63.480 92.500 ;
        RECT 63.180 91.300 63.480 91.750 ;
        RECT 63.180 90.550 63.480 91.000 ;
        RECT 63.180 89.800 63.480 90.250 ;
        RECT 63.180 89.050 63.480 89.500 ;
        RECT 63.180 88.300 63.480 88.750 ;
        RECT 63.180 87.550 63.480 88.000 ;
        RECT 63.180 86.800 63.480 87.250 ;
        RECT 63.180 86.050 63.480 86.500 ;
        RECT 63.180 85.300 63.480 85.750 ;
        RECT 65.980 94.300 66.280 94.750 ;
        RECT 65.980 93.550 66.280 94.000 ;
        RECT 65.980 92.800 66.280 93.250 ;
        RECT 65.980 92.050 66.280 92.500 ;
        RECT 65.980 91.300 66.280 91.750 ;
        RECT 65.980 90.550 66.280 91.000 ;
        RECT 65.980 89.800 66.280 90.250 ;
        RECT 65.980 89.050 66.280 89.500 ;
        RECT 65.980 88.300 66.280 88.750 ;
        RECT 65.980 87.550 66.280 88.000 ;
        RECT 65.980 86.800 66.280 87.250 ;
        RECT 65.980 86.050 66.280 86.500 ;
        RECT 65.980 85.300 66.280 85.750 ;
        RECT 83.180 94.300 83.480 94.750 ;
        RECT 83.180 93.550 83.480 94.000 ;
        RECT 83.180 92.800 83.480 93.250 ;
        RECT 83.180 92.050 83.480 92.500 ;
        RECT 83.180 91.300 83.480 91.750 ;
        RECT 83.180 90.550 83.480 91.000 ;
        RECT 83.180 89.800 83.480 90.250 ;
        RECT 83.180 89.050 83.480 89.500 ;
        RECT 83.180 88.300 83.480 88.750 ;
        RECT 83.180 87.550 83.480 88.000 ;
        RECT 83.180 86.800 83.480 87.250 ;
        RECT 83.180 86.050 83.480 86.500 ;
        RECT 83.180 85.300 83.480 85.750 ;
        RECT 85.980 94.300 86.280 94.750 ;
        RECT 85.980 93.550 86.280 94.000 ;
        RECT 85.980 92.800 86.280 93.250 ;
        RECT 85.980 92.050 86.280 92.500 ;
        RECT 85.980 91.300 86.280 91.750 ;
        RECT 85.980 90.550 86.280 91.000 ;
        RECT 85.980 89.800 86.280 90.250 ;
        RECT 85.980 89.050 86.280 89.500 ;
        RECT 85.980 88.300 86.280 88.750 ;
        RECT 85.980 87.550 86.280 88.000 ;
        RECT 85.980 86.800 86.280 87.250 ;
        RECT 85.980 86.050 86.280 86.500 ;
        RECT 85.980 85.300 86.280 85.750 ;
        RECT 103.180 94.300 103.480 94.750 ;
        RECT 103.180 93.550 103.480 94.000 ;
        RECT 103.180 92.800 103.480 93.250 ;
        RECT 103.180 92.050 103.480 92.500 ;
        RECT 103.180 91.300 103.480 91.750 ;
        RECT 103.180 90.550 103.480 91.000 ;
        RECT 103.180 89.800 103.480 90.250 ;
        RECT 103.180 89.050 103.480 89.500 ;
        RECT 103.180 88.300 103.480 88.750 ;
        RECT 103.180 87.550 103.480 88.000 ;
        RECT 103.180 86.800 103.480 87.250 ;
        RECT 103.180 86.050 103.480 86.500 ;
        RECT 103.180 85.300 103.480 85.750 ;
        RECT 105.980 94.300 106.280 94.750 ;
        RECT 105.980 93.550 106.280 94.000 ;
        RECT 105.980 92.800 106.280 93.250 ;
        RECT 105.980 92.050 106.280 92.500 ;
        RECT 105.980 91.300 106.280 91.750 ;
        RECT 105.980 90.550 106.280 91.000 ;
        RECT 105.980 89.800 106.280 90.250 ;
        RECT 105.980 89.050 106.280 89.500 ;
        RECT 105.980 88.300 106.280 88.750 ;
        RECT 105.980 87.550 106.280 88.000 ;
        RECT 105.980 86.800 106.280 87.250 ;
        RECT 105.980 86.050 106.280 86.500 ;
        RECT 105.980 85.300 106.280 85.750 ;
        RECT 123.180 94.300 123.480 94.750 ;
        RECT 123.180 93.550 123.480 94.000 ;
        RECT 123.180 92.800 123.480 93.250 ;
        RECT 123.180 92.050 123.480 92.500 ;
        RECT 123.180 91.300 123.480 91.750 ;
        RECT 123.180 90.550 123.480 91.000 ;
        RECT 123.180 89.800 123.480 90.250 ;
        RECT 123.180 89.050 123.480 89.500 ;
        RECT 123.180 88.300 123.480 88.750 ;
        RECT 123.180 87.550 123.480 88.000 ;
        RECT 123.180 86.800 123.480 87.250 ;
        RECT 123.180 86.050 123.480 86.500 ;
        RECT 123.180 85.300 123.480 85.750 ;
        RECT 5.980 74.300 6.280 74.750 ;
        RECT 5.980 73.550 6.280 74.000 ;
        RECT 5.980 72.800 6.280 73.250 ;
        RECT 5.980 72.050 6.280 72.500 ;
        RECT 5.980 71.300 6.280 71.750 ;
        RECT 5.980 70.550 6.280 71.000 ;
        RECT 5.980 69.800 6.280 70.250 ;
        RECT 5.980 69.050 6.280 69.500 ;
        RECT 5.980 68.300 6.280 68.750 ;
        RECT 5.980 67.550 6.280 68.000 ;
        RECT 5.980 66.800 6.280 67.250 ;
        RECT 5.980 66.050 6.280 66.500 ;
        RECT 5.980 65.300 6.280 65.750 ;
        RECT 23.180 74.300 23.480 74.750 ;
        RECT 23.180 73.550 23.480 74.000 ;
        RECT 23.180 72.800 23.480 73.250 ;
        RECT 23.180 72.050 23.480 72.500 ;
        RECT 23.180 71.300 23.480 71.750 ;
        RECT 23.180 70.550 23.480 71.000 ;
        RECT 23.180 69.800 23.480 70.250 ;
        RECT 23.180 69.050 23.480 69.500 ;
        RECT 23.180 68.300 23.480 68.750 ;
        RECT 23.180 67.550 23.480 68.000 ;
        RECT 23.180 66.800 23.480 67.250 ;
        RECT 23.180 66.050 23.480 66.500 ;
        RECT 23.180 65.300 23.480 65.750 ;
        RECT 25.980 74.300 26.280 74.750 ;
        RECT 25.980 73.550 26.280 74.000 ;
        RECT 25.980 72.800 26.280 73.250 ;
        RECT 25.980 72.050 26.280 72.500 ;
        RECT 25.980 71.300 26.280 71.750 ;
        RECT 25.980 70.550 26.280 71.000 ;
        RECT 25.980 69.800 26.280 70.250 ;
        RECT 25.980 69.050 26.280 69.500 ;
        RECT 25.980 68.300 26.280 68.750 ;
        RECT 25.980 67.550 26.280 68.000 ;
        RECT 25.980 66.800 26.280 67.250 ;
        RECT 25.980 66.050 26.280 66.500 ;
        RECT 25.980 65.300 26.280 65.750 ;
        RECT 43.180 74.300 43.480 74.750 ;
        RECT 43.180 73.550 43.480 74.000 ;
        RECT 43.180 72.800 43.480 73.250 ;
        RECT 43.180 72.050 43.480 72.500 ;
        RECT 43.180 71.300 43.480 71.750 ;
        RECT 43.180 70.550 43.480 71.000 ;
        RECT 43.180 69.800 43.480 70.250 ;
        RECT 43.180 69.050 43.480 69.500 ;
        RECT 43.180 68.300 43.480 68.750 ;
        RECT 43.180 67.550 43.480 68.000 ;
        RECT 43.180 66.800 43.480 67.250 ;
        RECT 43.180 66.050 43.480 66.500 ;
        RECT 43.180 65.300 43.480 65.750 ;
        RECT 45.980 74.300 46.280 74.750 ;
        RECT 45.980 73.550 46.280 74.000 ;
        RECT 45.980 72.800 46.280 73.250 ;
        RECT 45.980 72.050 46.280 72.500 ;
        RECT 45.980 71.300 46.280 71.750 ;
        RECT 45.980 70.550 46.280 71.000 ;
        RECT 45.980 69.800 46.280 70.250 ;
        RECT 45.980 69.050 46.280 69.500 ;
        RECT 45.980 68.300 46.280 68.750 ;
        RECT 45.980 67.550 46.280 68.000 ;
        RECT 45.980 66.800 46.280 67.250 ;
        RECT 45.980 66.050 46.280 66.500 ;
        RECT 45.980 65.300 46.280 65.750 ;
        RECT 63.180 74.300 63.480 74.750 ;
        RECT 63.180 73.550 63.480 74.000 ;
        RECT 63.180 72.800 63.480 73.250 ;
        RECT 63.180 72.050 63.480 72.500 ;
        RECT 63.180 71.300 63.480 71.750 ;
        RECT 63.180 70.550 63.480 71.000 ;
        RECT 63.180 69.800 63.480 70.250 ;
        RECT 63.180 69.050 63.480 69.500 ;
        RECT 63.180 68.300 63.480 68.750 ;
        RECT 63.180 67.550 63.480 68.000 ;
        RECT 63.180 66.800 63.480 67.250 ;
        RECT 63.180 66.050 63.480 66.500 ;
        RECT 63.180 65.300 63.480 65.750 ;
        RECT 65.980 74.300 66.280 74.750 ;
        RECT 65.980 73.550 66.280 74.000 ;
        RECT 65.980 72.800 66.280 73.250 ;
        RECT 65.980 72.050 66.280 72.500 ;
        RECT 65.980 71.300 66.280 71.750 ;
        RECT 65.980 70.550 66.280 71.000 ;
        RECT 65.980 69.800 66.280 70.250 ;
        RECT 65.980 69.050 66.280 69.500 ;
        RECT 65.980 68.300 66.280 68.750 ;
        RECT 65.980 67.550 66.280 68.000 ;
        RECT 65.980 66.800 66.280 67.250 ;
        RECT 65.980 66.050 66.280 66.500 ;
        RECT 65.980 65.300 66.280 65.750 ;
        RECT 83.180 74.300 83.480 74.750 ;
        RECT 83.180 73.550 83.480 74.000 ;
        RECT 83.180 72.800 83.480 73.250 ;
        RECT 83.180 72.050 83.480 72.500 ;
        RECT 83.180 71.300 83.480 71.750 ;
        RECT 83.180 70.550 83.480 71.000 ;
        RECT 83.180 69.800 83.480 70.250 ;
        RECT 83.180 69.050 83.480 69.500 ;
        RECT 83.180 68.300 83.480 68.750 ;
        RECT 83.180 67.550 83.480 68.000 ;
        RECT 83.180 66.800 83.480 67.250 ;
        RECT 83.180 66.050 83.480 66.500 ;
        RECT 83.180 65.300 83.480 65.750 ;
        RECT 85.980 74.300 86.280 74.750 ;
        RECT 85.980 73.550 86.280 74.000 ;
        RECT 85.980 72.800 86.280 73.250 ;
        RECT 85.980 72.050 86.280 72.500 ;
        RECT 85.980 71.300 86.280 71.750 ;
        RECT 85.980 70.550 86.280 71.000 ;
        RECT 85.980 69.800 86.280 70.250 ;
        RECT 85.980 69.050 86.280 69.500 ;
        RECT 85.980 68.300 86.280 68.750 ;
        RECT 85.980 67.550 86.280 68.000 ;
        RECT 85.980 66.800 86.280 67.250 ;
        RECT 85.980 66.050 86.280 66.500 ;
        RECT 85.980 65.300 86.280 65.750 ;
        RECT 103.180 74.300 103.480 74.750 ;
        RECT 103.180 73.550 103.480 74.000 ;
        RECT 103.180 72.800 103.480 73.250 ;
        RECT 103.180 72.050 103.480 72.500 ;
        RECT 103.180 71.300 103.480 71.750 ;
        RECT 103.180 70.550 103.480 71.000 ;
        RECT 103.180 69.800 103.480 70.250 ;
        RECT 103.180 69.050 103.480 69.500 ;
        RECT 103.180 68.300 103.480 68.750 ;
        RECT 103.180 67.550 103.480 68.000 ;
        RECT 103.180 66.800 103.480 67.250 ;
        RECT 103.180 66.050 103.480 66.500 ;
        RECT 103.180 65.300 103.480 65.750 ;
        RECT 105.980 74.300 106.280 74.750 ;
        RECT 105.980 73.550 106.280 74.000 ;
        RECT 105.980 72.800 106.280 73.250 ;
        RECT 105.980 72.050 106.280 72.500 ;
        RECT 105.980 71.300 106.280 71.750 ;
        RECT 105.980 70.550 106.280 71.000 ;
        RECT 105.980 69.800 106.280 70.250 ;
        RECT 105.980 69.050 106.280 69.500 ;
        RECT 105.980 68.300 106.280 68.750 ;
        RECT 105.980 67.550 106.280 68.000 ;
        RECT 105.980 66.800 106.280 67.250 ;
        RECT 105.980 66.050 106.280 66.500 ;
        RECT 105.980 65.300 106.280 65.750 ;
        RECT 123.180 74.300 123.480 74.750 ;
        RECT 123.180 73.550 123.480 74.000 ;
        RECT 123.180 72.800 123.480 73.250 ;
        RECT 123.180 72.050 123.480 72.500 ;
        RECT 123.180 71.300 123.480 71.750 ;
        RECT 123.180 70.550 123.480 71.000 ;
        RECT 123.180 69.800 123.480 70.250 ;
        RECT 123.180 69.050 123.480 69.500 ;
        RECT 123.180 68.300 123.480 68.750 ;
        RECT 123.180 67.550 123.480 68.000 ;
        RECT 123.180 66.800 123.480 67.250 ;
        RECT 123.180 66.050 123.480 66.500 ;
        RECT 123.180 65.300 123.480 65.750 ;
        RECT 5.980 54.300 6.280 54.750 ;
        RECT 5.980 53.550 6.280 54.000 ;
        RECT 5.980 52.800 6.280 53.250 ;
        RECT 5.980 52.050 6.280 52.500 ;
        RECT 5.980 51.300 6.280 51.750 ;
        RECT 5.980 50.550 6.280 51.000 ;
        RECT 5.980 49.800 6.280 50.250 ;
        RECT 5.980 49.050 6.280 49.500 ;
        RECT 5.980 48.300 6.280 48.750 ;
        RECT 5.980 47.550 6.280 48.000 ;
        RECT 5.980 46.800 6.280 47.250 ;
        RECT 5.980 46.050 6.280 46.500 ;
        RECT 5.980 45.300 6.280 45.750 ;
        RECT 23.180 54.300 23.480 54.750 ;
        RECT 23.180 53.550 23.480 54.000 ;
        RECT 23.180 52.800 23.480 53.250 ;
        RECT 23.180 52.050 23.480 52.500 ;
        RECT 23.180 51.300 23.480 51.750 ;
        RECT 23.180 50.550 23.480 51.000 ;
        RECT 23.180 49.800 23.480 50.250 ;
        RECT 23.180 49.050 23.480 49.500 ;
        RECT 23.180 48.300 23.480 48.750 ;
        RECT 23.180 47.550 23.480 48.000 ;
        RECT 23.180 46.800 23.480 47.250 ;
        RECT 23.180 46.050 23.480 46.500 ;
        RECT 23.180 45.300 23.480 45.750 ;
        RECT 25.980 54.300 26.280 54.750 ;
        RECT 25.980 53.550 26.280 54.000 ;
        RECT 25.980 52.800 26.280 53.250 ;
        RECT 25.980 52.050 26.280 52.500 ;
        RECT 25.980 51.300 26.280 51.750 ;
        RECT 25.980 50.550 26.280 51.000 ;
        RECT 25.980 49.800 26.280 50.250 ;
        RECT 25.980 49.050 26.280 49.500 ;
        RECT 25.980 48.300 26.280 48.750 ;
        RECT 25.980 47.550 26.280 48.000 ;
        RECT 25.980 46.800 26.280 47.250 ;
        RECT 25.980 46.050 26.280 46.500 ;
        RECT 25.980 45.300 26.280 45.750 ;
        RECT 43.180 54.300 43.480 54.750 ;
        RECT 43.180 53.550 43.480 54.000 ;
        RECT 43.180 52.800 43.480 53.250 ;
        RECT 43.180 52.050 43.480 52.500 ;
        RECT 43.180 51.300 43.480 51.750 ;
        RECT 43.180 50.550 43.480 51.000 ;
        RECT 43.180 49.800 43.480 50.250 ;
        RECT 43.180 49.050 43.480 49.500 ;
        RECT 43.180 48.300 43.480 48.750 ;
        RECT 43.180 47.550 43.480 48.000 ;
        RECT 43.180 46.800 43.480 47.250 ;
        RECT 43.180 46.050 43.480 46.500 ;
        RECT 43.180 45.300 43.480 45.750 ;
        RECT 45.980 54.300 46.280 54.750 ;
        RECT 45.980 53.550 46.280 54.000 ;
        RECT 45.980 52.800 46.280 53.250 ;
        RECT 45.980 52.050 46.280 52.500 ;
        RECT 45.980 51.300 46.280 51.750 ;
        RECT 45.980 50.550 46.280 51.000 ;
        RECT 45.980 49.800 46.280 50.250 ;
        RECT 45.980 49.050 46.280 49.500 ;
        RECT 45.980 48.300 46.280 48.750 ;
        RECT 45.980 47.550 46.280 48.000 ;
        RECT 45.980 46.800 46.280 47.250 ;
        RECT 45.980 46.050 46.280 46.500 ;
        RECT 45.980 45.300 46.280 45.750 ;
        RECT 63.180 54.300 63.480 54.750 ;
        RECT 63.180 53.550 63.480 54.000 ;
        RECT 63.180 52.800 63.480 53.250 ;
        RECT 63.180 52.050 63.480 52.500 ;
        RECT 63.180 51.300 63.480 51.750 ;
        RECT 63.180 50.550 63.480 51.000 ;
        RECT 63.180 49.800 63.480 50.250 ;
        RECT 63.180 49.050 63.480 49.500 ;
        RECT 63.180 48.300 63.480 48.750 ;
        RECT 63.180 47.550 63.480 48.000 ;
        RECT 63.180 46.800 63.480 47.250 ;
        RECT 63.180 46.050 63.480 46.500 ;
        RECT 63.180 45.300 63.480 45.750 ;
        RECT 65.980 54.300 66.280 54.750 ;
        RECT 65.980 53.550 66.280 54.000 ;
        RECT 65.980 52.800 66.280 53.250 ;
        RECT 65.980 52.050 66.280 52.500 ;
        RECT 65.980 51.300 66.280 51.750 ;
        RECT 65.980 50.550 66.280 51.000 ;
        RECT 65.980 49.800 66.280 50.250 ;
        RECT 65.980 49.050 66.280 49.500 ;
        RECT 65.980 48.300 66.280 48.750 ;
        RECT 65.980 47.550 66.280 48.000 ;
        RECT 65.980 46.800 66.280 47.250 ;
        RECT 65.980 46.050 66.280 46.500 ;
        RECT 65.980 45.300 66.280 45.750 ;
        RECT 83.180 54.300 83.480 54.750 ;
        RECT 83.180 53.550 83.480 54.000 ;
        RECT 83.180 52.800 83.480 53.250 ;
        RECT 83.180 52.050 83.480 52.500 ;
        RECT 83.180 51.300 83.480 51.750 ;
        RECT 83.180 50.550 83.480 51.000 ;
        RECT 83.180 49.800 83.480 50.250 ;
        RECT 83.180 49.050 83.480 49.500 ;
        RECT 83.180 48.300 83.480 48.750 ;
        RECT 83.180 47.550 83.480 48.000 ;
        RECT 83.180 46.800 83.480 47.250 ;
        RECT 83.180 46.050 83.480 46.500 ;
        RECT 83.180 45.300 83.480 45.750 ;
        RECT 85.980 54.300 86.280 54.750 ;
        RECT 85.980 53.550 86.280 54.000 ;
        RECT 85.980 52.800 86.280 53.250 ;
        RECT 85.980 52.050 86.280 52.500 ;
        RECT 85.980 51.300 86.280 51.750 ;
        RECT 85.980 50.550 86.280 51.000 ;
        RECT 85.980 49.800 86.280 50.250 ;
        RECT 85.980 49.050 86.280 49.500 ;
        RECT 85.980 48.300 86.280 48.750 ;
        RECT 85.980 47.550 86.280 48.000 ;
        RECT 85.980 46.800 86.280 47.250 ;
        RECT 85.980 46.050 86.280 46.500 ;
        RECT 85.980 45.300 86.280 45.750 ;
        RECT 103.180 54.300 103.480 54.750 ;
        RECT 103.180 53.550 103.480 54.000 ;
        RECT 103.180 52.800 103.480 53.250 ;
        RECT 103.180 52.050 103.480 52.500 ;
        RECT 103.180 51.300 103.480 51.750 ;
        RECT 103.180 50.550 103.480 51.000 ;
        RECT 103.180 49.800 103.480 50.250 ;
        RECT 103.180 49.050 103.480 49.500 ;
        RECT 103.180 48.300 103.480 48.750 ;
        RECT 103.180 47.550 103.480 48.000 ;
        RECT 103.180 46.800 103.480 47.250 ;
        RECT 103.180 46.050 103.480 46.500 ;
        RECT 103.180 45.300 103.480 45.750 ;
        RECT 105.980 54.300 106.280 54.750 ;
        RECT 105.980 53.550 106.280 54.000 ;
        RECT 105.980 52.800 106.280 53.250 ;
        RECT 105.980 52.050 106.280 52.500 ;
        RECT 105.980 51.300 106.280 51.750 ;
        RECT 105.980 50.550 106.280 51.000 ;
        RECT 105.980 49.800 106.280 50.250 ;
        RECT 105.980 49.050 106.280 49.500 ;
        RECT 105.980 48.300 106.280 48.750 ;
        RECT 105.980 47.550 106.280 48.000 ;
        RECT 105.980 46.800 106.280 47.250 ;
        RECT 105.980 46.050 106.280 46.500 ;
        RECT 105.980 45.300 106.280 45.750 ;
        RECT 123.180 54.300 123.480 54.750 ;
        RECT 123.180 53.550 123.480 54.000 ;
        RECT 123.180 52.800 123.480 53.250 ;
        RECT 123.180 52.050 123.480 52.500 ;
        RECT 123.180 51.300 123.480 51.750 ;
        RECT 123.180 50.550 123.480 51.000 ;
        RECT 123.180 49.800 123.480 50.250 ;
        RECT 123.180 49.050 123.480 49.500 ;
        RECT 123.180 48.300 123.480 48.750 ;
        RECT 123.180 47.550 123.480 48.000 ;
        RECT 123.180 46.800 123.480 47.250 ;
        RECT 123.180 46.050 123.480 46.500 ;
        RECT 123.180 45.300 123.480 45.750 ;
        RECT 5.980 34.300 6.280 34.750 ;
        RECT 5.980 33.550 6.280 34.000 ;
        RECT 5.980 32.800 6.280 33.250 ;
        RECT 5.980 32.050 6.280 32.500 ;
        RECT 5.980 31.300 6.280 31.750 ;
        RECT 5.980 30.550 6.280 31.000 ;
        RECT 5.980 29.800 6.280 30.250 ;
        RECT 5.980 29.050 6.280 29.500 ;
        RECT 5.980 28.300 6.280 28.750 ;
        RECT 5.980 27.550 6.280 28.000 ;
        RECT 5.980 26.800 6.280 27.250 ;
        RECT 5.980 26.050 6.280 26.500 ;
        RECT 5.980 25.300 6.280 25.750 ;
        RECT 23.180 34.300 23.480 34.750 ;
        RECT 23.180 33.550 23.480 34.000 ;
        RECT 23.180 32.800 23.480 33.250 ;
        RECT 23.180 32.050 23.480 32.500 ;
        RECT 23.180 31.300 23.480 31.750 ;
        RECT 23.180 30.550 23.480 31.000 ;
        RECT 23.180 29.800 23.480 30.250 ;
        RECT 23.180 29.050 23.480 29.500 ;
        RECT 23.180 28.300 23.480 28.750 ;
        RECT 23.180 27.550 23.480 28.000 ;
        RECT 23.180 26.800 23.480 27.250 ;
        RECT 23.180 26.050 23.480 26.500 ;
        RECT 23.180 25.300 23.480 25.750 ;
        RECT 25.980 34.300 26.280 34.750 ;
        RECT 25.980 33.550 26.280 34.000 ;
        RECT 25.980 32.800 26.280 33.250 ;
        RECT 25.980 32.050 26.280 32.500 ;
        RECT 25.980 31.300 26.280 31.750 ;
        RECT 25.980 30.550 26.280 31.000 ;
        RECT 25.980 29.800 26.280 30.250 ;
        RECT 25.980 29.050 26.280 29.500 ;
        RECT 25.980 28.300 26.280 28.750 ;
        RECT 25.980 27.550 26.280 28.000 ;
        RECT 25.980 26.800 26.280 27.250 ;
        RECT 25.980 26.050 26.280 26.500 ;
        RECT 25.980 25.300 26.280 25.750 ;
        RECT 43.180 34.300 43.480 34.750 ;
        RECT 43.180 33.550 43.480 34.000 ;
        RECT 43.180 32.800 43.480 33.250 ;
        RECT 43.180 32.050 43.480 32.500 ;
        RECT 43.180 31.300 43.480 31.750 ;
        RECT 43.180 30.550 43.480 31.000 ;
        RECT 43.180 29.800 43.480 30.250 ;
        RECT 43.180 29.050 43.480 29.500 ;
        RECT 43.180 28.300 43.480 28.750 ;
        RECT 43.180 27.550 43.480 28.000 ;
        RECT 43.180 26.800 43.480 27.250 ;
        RECT 43.180 26.050 43.480 26.500 ;
        RECT 43.180 25.300 43.480 25.750 ;
        RECT 45.980 34.300 46.280 34.750 ;
        RECT 45.980 33.550 46.280 34.000 ;
        RECT 45.980 32.800 46.280 33.250 ;
        RECT 45.980 32.050 46.280 32.500 ;
        RECT 45.980 31.300 46.280 31.750 ;
        RECT 45.980 30.550 46.280 31.000 ;
        RECT 45.980 29.800 46.280 30.250 ;
        RECT 45.980 29.050 46.280 29.500 ;
        RECT 45.980 28.300 46.280 28.750 ;
        RECT 45.980 27.550 46.280 28.000 ;
        RECT 45.980 26.800 46.280 27.250 ;
        RECT 45.980 26.050 46.280 26.500 ;
        RECT 45.980 25.300 46.280 25.750 ;
        RECT 63.180 34.300 63.480 34.750 ;
        RECT 63.180 33.550 63.480 34.000 ;
        RECT 63.180 32.800 63.480 33.250 ;
        RECT 63.180 32.050 63.480 32.500 ;
        RECT 63.180 31.300 63.480 31.750 ;
        RECT 63.180 30.550 63.480 31.000 ;
        RECT 63.180 29.800 63.480 30.250 ;
        RECT 63.180 29.050 63.480 29.500 ;
        RECT 63.180 28.300 63.480 28.750 ;
        RECT 63.180 27.550 63.480 28.000 ;
        RECT 63.180 26.800 63.480 27.250 ;
        RECT 63.180 26.050 63.480 26.500 ;
        RECT 63.180 25.300 63.480 25.750 ;
        RECT 65.980 34.300 66.280 34.750 ;
        RECT 65.980 33.550 66.280 34.000 ;
        RECT 65.980 32.800 66.280 33.250 ;
        RECT 65.980 32.050 66.280 32.500 ;
        RECT 65.980 31.300 66.280 31.750 ;
        RECT 65.980 30.550 66.280 31.000 ;
        RECT 65.980 29.800 66.280 30.250 ;
        RECT 65.980 29.050 66.280 29.500 ;
        RECT 65.980 28.300 66.280 28.750 ;
        RECT 65.980 27.550 66.280 28.000 ;
        RECT 65.980 26.800 66.280 27.250 ;
        RECT 65.980 26.050 66.280 26.500 ;
        RECT 65.980 25.300 66.280 25.750 ;
        RECT 83.180 34.300 83.480 34.750 ;
        RECT 83.180 33.550 83.480 34.000 ;
        RECT 83.180 32.800 83.480 33.250 ;
        RECT 83.180 32.050 83.480 32.500 ;
        RECT 83.180 31.300 83.480 31.750 ;
        RECT 83.180 30.550 83.480 31.000 ;
        RECT 83.180 29.800 83.480 30.250 ;
        RECT 83.180 29.050 83.480 29.500 ;
        RECT 83.180 28.300 83.480 28.750 ;
        RECT 83.180 27.550 83.480 28.000 ;
        RECT 83.180 26.800 83.480 27.250 ;
        RECT 83.180 26.050 83.480 26.500 ;
        RECT 83.180 25.300 83.480 25.750 ;
        RECT 85.980 34.300 86.280 34.750 ;
        RECT 85.980 33.550 86.280 34.000 ;
        RECT 85.980 32.800 86.280 33.250 ;
        RECT 85.980 32.050 86.280 32.500 ;
        RECT 85.980 31.300 86.280 31.750 ;
        RECT 85.980 30.550 86.280 31.000 ;
        RECT 85.980 29.800 86.280 30.250 ;
        RECT 85.980 29.050 86.280 29.500 ;
        RECT 85.980 28.300 86.280 28.750 ;
        RECT 85.980 27.550 86.280 28.000 ;
        RECT 85.980 26.800 86.280 27.250 ;
        RECT 85.980 26.050 86.280 26.500 ;
        RECT 85.980 25.300 86.280 25.750 ;
        RECT 103.180 34.300 103.480 34.750 ;
        RECT 103.180 33.550 103.480 34.000 ;
        RECT 103.180 32.800 103.480 33.250 ;
        RECT 103.180 32.050 103.480 32.500 ;
        RECT 103.180 31.300 103.480 31.750 ;
        RECT 103.180 30.550 103.480 31.000 ;
        RECT 103.180 29.800 103.480 30.250 ;
        RECT 103.180 29.050 103.480 29.500 ;
        RECT 103.180 28.300 103.480 28.750 ;
        RECT 103.180 27.550 103.480 28.000 ;
        RECT 103.180 26.800 103.480 27.250 ;
        RECT 103.180 26.050 103.480 26.500 ;
        RECT 103.180 25.300 103.480 25.750 ;
        RECT 105.980 34.300 106.280 34.750 ;
        RECT 105.980 33.550 106.280 34.000 ;
        RECT 105.980 32.800 106.280 33.250 ;
        RECT 105.980 32.050 106.280 32.500 ;
        RECT 105.980 31.300 106.280 31.750 ;
        RECT 105.980 30.550 106.280 31.000 ;
        RECT 105.980 29.800 106.280 30.250 ;
        RECT 105.980 29.050 106.280 29.500 ;
        RECT 105.980 28.300 106.280 28.750 ;
        RECT 105.980 27.550 106.280 28.000 ;
        RECT 105.980 26.800 106.280 27.250 ;
        RECT 105.980 26.050 106.280 26.500 ;
        RECT 105.980 25.300 106.280 25.750 ;
        RECT 123.180 34.300 123.480 34.750 ;
        RECT 123.180 33.550 123.480 34.000 ;
        RECT 123.180 32.800 123.480 33.250 ;
        RECT 123.180 32.050 123.480 32.500 ;
        RECT 123.180 31.300 123.480 31.750 ;
        RECT 123.180 30.550 123.480 31.000 ;
        RECT 123.180 29.800 123.480 30.250 ;
        RECT 123.180 29.050 123.480 29.500 ;
        RECT 123.180 28.300 123.480 28.750 ;
        RECT 123.180 27.550 123.480 28.000 ;
        RECT 123.180 26.800 123.480 27.250 ;
        RECT 123.180 26.050 123.480 26.500 ;
        RECT 123.180 25.300 123.480 25.750 ;
        RECT 5.980 14.300 6.280 14.750 ;
        RECT 5.980 13.550 6.280 14.000 ;
        RECT 5.980 12.800 6.280 13.250 ;
        RECT 5.980 12.050 6.280 12.500 ;
        RECT 5.980 11.300 6.280 11.750 ;
        RECT 5.980 10.550 6.280 11.000 ;
        RECT 5.980 9.800 6.280 10.250 ;
        RECT 5.980 9.050 6.280 9.500 ;
        RECT 5.980 8.300 6.280 8.750 ;
        RECT 5.980 7.550 6.280 8.000 ;
        RECT 5.980 6.800 6.280 7.250 ;
        RECT 5.980 6.050 6.280 6.500 ;
        RECT 5.980 5.300 6.280 5.750 ;
        RECT 23.180 14.300 23.480 14.750 ;
        RECT 23.180 13.550 23.480 14.000 ;
        RECT 23.180 12.800 23.480 13.250 ;
        RECT 23.180 12.050 23.480 12.500 ;
        RECT 23.180 11.300 23.480 11.750 ;
        RECT 23.180 10.550 23.480 11.000 ;
        RECT 23.180 9.800 23.480 10.250 ;
        RECT 23.180 9.050 23.480 9.500 ;
        RECT 23.180 8.300 23.480 8.750 ;
        RECT 23.180 7.550 23.480 8.000 ;
        RECT 23.180 6.800 23.480 7.250 ;
        RECT 23.180 6.050 23.480 6.500 ;
        RECT 23.180 5.300 23.480 5.750 ;
        RECT 25.980 14.300 26.280 14.750 ;
        RECT 25.980 13.550 26.280 14.000 ;
        RECT 25.980 12.800 26.280 13.250 ;
        RECT 25.980 12.050 26.280 12.500 ;
        RECT 25.980 11.300 26.280 11.750 ;
        RECT 25.980 10.550 26.280 11.000 ;
        RECT 25.980 9.800 26.280 10.250 ;
        RECT 25.980 9.050 26.280 9.500 ;
        RECT 25.980 8.300 26.280 8.750 ;
        RECT 25.980 7.550 26.280 8.000 ;
        RECT 25.980 6.800 26.280 7.250 ;
        RECT 25.980 6.050 26.280 6.500 ;
        RECT 25.980 5.300 26.280 5.750 ;
        RECT 43.180 14.300 43.480 14.750 ;
        RECT 43.180 13.550 43.480 14.000 ;
        RECT 43.180 12.800 43.480 13.250 ;
        RECT 43.180 12.050 43.480 12.500 ;
        RECT 43.180 11.300 43.480 11.750 ;
        RECT 43.180 10.550 43.480 11.000 ;
        RECT 43.180 9.800 43.480 10.250 ;
        RECT 43.180 9.050 43.480 9.500 ;
        RECT 43.180 8.300 43.480 8.750 ;
        RECT 43.180 7.550 43.480 8.000 ;
        RECT 43.180 6.800 43.480 7.250 ;
        RECT 43.180 6.050 43.480 6.500 ;
        RECT 43.180 5.300 43.480 5.750 ;
        RECT 45.980 14.300 46.280 14.750 ;
        RECT 45.980 13.550 46.280 14.000 ;
        RECT 45.980 12.800 46.280 13.250 ;
        RECT 45.980 12.050 46.280 12.500 ;
        RECT 45.980 11.300 46.280 11.750 ;
        RECT 45.980 10.550 46.280 11.000 ;
        RECT 45.980 9.800 46.280 10.250 ;
        RECT 45.980 9.050 46.280 9.500 ;
        RECT 45.980 8.300 46.280 8.750 ;
        RECT 45.980 7.550 46.280 8.000 ;
        RECT 45.980 6.800 46.280 7.250 ;
        RECT 45.980 6.050 46.280 6.500 ;
        RECT 45.980 5.300 46.280 5.750 ;
        RECT 63.180 14.300 63.480 14.750 ;
        RECT 63.180 13.550 63.480 14.000 ;
        RECT 63.180 12.800 63.480 13.250 ;
        RECT 63.180 12.050 63.480 12.500 ;
        RECT 63.180 11.300 63.480 11.750 ;
        RECT 63.180 10.550 63.480 11.000 ;
        RECT 63.180 9.800 63.480 10.250 ;
        RECT 63.180 9.050 63.480 9.500 ;
        RECT 63.180 8.300 63.480 8.750 ;
        RECT 63.180 7.550 63.480 8.000 ;
        RECT 63.180 6.800 63.480 7.250 ;
        RECT 63.180 6.050 63.480 6.500 ;
        RECT 63.180 5.300 63.480 5.750 ;
        RECT 65.980 14.300 66.280 14.750 ;
        RECT 65.980 13.550 66.280 14.000 ;
        RECT 65.980 12.800 66.280 13.250 ;
        RECT 65.980 12.050 66.280 12.500 ;
        RECT 65.980 11.300 66.280 11.750 ;
        RECT 65.980 10.550 66.280 11.000 ;
        RECT 65.980 9.800 66.280 10.250 ;
        RECT 65.980 9.050 66.280 9.500 ;
        RECT 65.980 8.300 66.280 8.750 ;
        RECT 65.980 7.550 66.280 8.000 ;
        RECT 65.980 6.800 66.280 7.250 ;
        RECT 65.980 6.050 66.280 6.500 ;
        RECT 65.980 5.300 66.280 5.750 ;
        RECT 83.180 14.300 83.480 14.750 ;
        RECT 83.180 13.550 83.480 14.000 ;
        RECT 83.180 12.800 83.480 13.250 ;
        RECT 83.180 12.050 83.480 12.500 ;
        RECT 83.180 11.300 83.480 11.750 ;
        RECT 83.180 10.550 83.480 11.000 ;
        RECT 83.180 9.800 83.480 10.250 ;
        RECT 83.180 9.050 83.480 9.500 ;
        RECT 83.180 8.300 83.480 8.750 ;
        RECT 83.180 7.550 83.480 8.000 ;
        RECT 83.180 6.800 83.480 7.250 ;
        RECT 83.180 6.050 83.480 6.500 ;
        RECT 83.180 5.300 83.480 5.750 ;
        RECT 85.980 14.300 86.280 14.750 ;
        RECT 85.980 13.550 86.280 14.000 ;
        RECT 85.980 12.800 86.280 13.250 ;
        RECT 85.980 12.050 86.280 12.500 ;
        RECT 85.980 11.300 86.280 11.750 ;
        RECT 85.980 10.550 86.280 11.000 ;
        RECT 85.980 9.800 86.280 10.250 ;
        RECT 85.980 9.050 86.280 9.500 ;
        RECT 85.980 8.300 86.280 8.750 ;
        RECT 85.980 7.550 86.280 8.000 ;
        RECT 85.980 6.800 86.280 7.250 ;
        RECT 85.980 6.050 86.280 6.500 ;
        RECT 85.980 5.300 86.280 5.750 ;
        RECT 103.180 14.300 103.480 14.750 ;
        RECT 103.180 13.550 103.480 14.000 ;
        RECT 103.180 12.800 103.480 13.250 ;
        RECT 103.180 12.050 103.480 12.500 ;
        RECT 103.180 11.300 103.480 11.750 ;
        RECT 103.180 10.550 103.480 11.000 ;
        RECT 103.180 9.800 103.480 10.250 ;
        RECT 103.180 9.050 103.480 9.500 ;
        RECT 103.180 8.300 103.480 8.750 ;
        RECT 103.180 7.550 103.480 8.000 ;
        RECT 103.180 6.800 103.480 7.250 ;
        RECT 103.180 6.050 103.480 6.500 ;
        RECT 103.180 5.300 103.480 5.750 ;
        RECT 105.980 14.300 106.280 14.750 ;
        RECT 105.980 13.550 106.280 14.000 ;
        RECT 105.980 12.800 106.280 13.250 ;
        RECT 105.980 12.050 106.280 12.500 ;
        RECT 105.980 11.300 106.280 11.750 ;
        RECT 105.980 10.550 106.280 11.000 ;
        RECT 105.980 9.800 106.280 10.250 ;
        RECT 105.980 9.050 106.280 9.500 ;
        RECT 105.980 8.300 106.280 8.750 ;
        RECT 105.980 7.550 106.280 8.000 ;
        RECT 105.980 6.800 106.280 7.250 ;
        RECT 105.980 6.050 106.280 6.500 ;
        RECT 105.980 5.300 106.280 5.750 ;
        RECT 123.180 14.300 123.480 14.750 ;
        RECT 123.180 13.550 123.480 14.000 ;
        RECT 123.180 12.800 123.480 13.250 ;
        RECT 123.180 12.050 123.480 12.500 ;
        RECT 123.180 11.300 123.480 11.750 ;
        RECT 123.180 10.550 123.480 11.000 ;
        RECT 123.180 9.800 123.480 10.250 ;
        RECT 123.180 9.050 123.480 9.500 ;
        RECT 123.180 8.300 123.480 8.750 ;
        RECT 123.180 7.550 123.480 8.000 ;
        RECT 123.180 6.800 123.480 7.250 ;
        RECT 123.180 6.050 123.480 6.500 ;
        RECT 123.180 5.300 123.480 5.750 ;
      LAYER met1 ;
        RECT 11.530 338.800 17.930 340.000 ;
        RECT 31.530 338.800 37.930 340.000 ;
        RECT 51.530 338.800 57.930 340.000 ;
        RECT 71.530 338.800 77.930 340.000 ;
        RECT 91.530 338.800 97.930 340.000 ;
        RECT 111.530 338.800 117.930 340.000 ;
        RECT 14.230 338.150 15.230 338.800 ;
        RECT 34.230 338.150 35.230 338.800 ;
        RECT 54.230 338.150 55.230 338.800 ;
        RECT 74.230 338.150 75.230 338.800 ;
        RECT 94.230 338.150 95.230 338.800 ;
        RECT 114.230 338.150 115.230 338.800 ;
        RECT 10.880 338.000 18.580 338.150 ;
        RECT 30.880 338.000 38.580 338.150 ;
        RECT 50.880 338.000 58.580 338.150 ;
        RECT 70.880 338.000 78.580 338.150 ;
        RECT 90.880 338.000 98.580 338.150 ;
        RECT 110.880 338.000 118.580 338.150 ;
        RECT 5.930 333.200 6.680 335.000 ;
        RECT 4.730 330.450 6.680 333.200 ;
        RECT 4.730 329.550 4.880 330.450 ;
        RECT 5.530 330.300 6.680 330.450 ;
        RECT 6.830 330.300 6.980 337.850 ;
        RECT 7.430 330.300 7.580 337.850 ;
        RECT 8.030 330.300 8.180 337.850 ;
        RECT 8.630 330.300 8.780 337.850 ;
        RECT 9.230 330.300 9.380 337.850 ;
        RECT 9.830 330.300 9.980 337.850 ;
        RECT 14.230 337.550 15.230 338.000 ;
        RECT 10.880 337.400 18.580 337.550 ;
        RECT 14.230 336.950 15.230 337.400 ;
        RECT 10.880 336.800 18.580 336.950 ;
        RECT 14.230 336.350 15.230 336.800 ;
        RECT 10.880 336.200 18.580 336.350 ;
        RECT 14.230 335.750 15.230 336.200 ;
        RECT 10.880 335.600 18.580 335.750 ;
        RECT 14.230 335.150 15.230 335.600 ;
        RECT 10.880 335.000 18.580 335.150 ;
        RECT 14.230 334.550 15.230 335.000 ;
        RECT 10.880 334.400 18.580 334.550 ;
        RECT 14.230 333.950 15.230 334.400 ;
        RECT 10.880 333.800 18.580 333.950 ;
        RECT 14.230 333.350 15.230 333.800 ;
        RECT 10.880 333.200 18.580 333.350 ;
        RECT 14.230 332.750 15.230 333.200 ;
        RECT 10.880 332.600 18.580 332.750 ;
        RECT 14.230 332.150 15.230 332.600 ;
        RECT 10.880 332.000 18.580 332.150 ;
        RECT 14.230 331.550 15.230 332.000 ;
        RECT 10.880 331.400 18.580 331.550 ;
        RECT 14.230 330.950 15.230 331.400 ;
        RECT 10.880 330.800 18.580 330.950 ;
        RECT 14.230 330.300 15.230 330.800 ;
        RECT 19.480 330.300 19.630 337.850 ;
        RECT 20.080 330.300 20.230 337.850 ;
        RECT 20.680 330.300 20.830 337.850 ;
        RECT 21.280 330.300 21.430 337.850 ;
        RECT 21.880 330.300 22.030 337.850 ;
        RECT 22.480 330.300 22.630 337.850 ;
        RECT 22.780 333.200 23.530 335.000 ;
        RECT 25.930 333.200 26.680 335.000 ;
        RECT 22.780 330.450 26.680 333.200 ;
        RECT 22.780 330.300 23.930 330.450 ;
        RECT 5.530 329.700 23.930 330.300 ;
        RECT 5.530 329.550 6.680 329.700 ;
        RECT 4.730 326.800 6.680 329.550 ;
        RECT 5.930 325.050 6.680 326.800 ;
        RECT 6.830 322.150 6.980 329.700 ;
        RECT 7.430 322.150 7.580 329.700 ;
        RECT 8.030 322.150 8.180 329.700 ;
        RECT 8.630 322.150 8.780 329.700 ;
        RECT 9.230 322.150 9.380 329.700 ;
        RECT 9.830 322.150 9.980 329.700 ;
        RECT 14.230 329.200 15.230 329.700 ;
        RECT 10.880 329.050 18.580 329.200 ;
        RECT 14.230 328.600 15.230 329.050 ;
        RECT 10.880 328.450 18.580 328.600 ;
        RECT 14.230 328.000 15.230 328.450 ;
        RECT 10.880 327.850 18.580 328.000 ;
        RECT 14.230 327.400 15.230 327.850 ;
        RECT 10.880 327.250 18.580 327.400 ;
        RECT 14.230 326.800 15.230 327.250 ;
        RECT 10.880 326.650 18.580 326.800 ;
        RECT 14.230 326.200 15.230 326.650 ;
        RECT 10.880 326.050 18.580 326.200 ;
        RECT 14.230 325.600 15.230 326.050 ;
        RECT 10.880 325.450 18.580 325.600 ;
        RECT 14.230 325.000 15.230 325.450 ;
        RECT 10.880 324.850 18.580 325.000 ;
        RECT 14.230 324.400 15.230 324.850 ;
        RECT 10.880 324.250 18.580 324.400 ;
        RECT 14.230 323.800 15.230 324.250 ;
        RECT 10.880 323.650 18.580 323.800 ;
        RECT 14.230 323.200 15.230 323.650 ;
        RECT 10.880 323.050 18.580 323.200 ;
        RECT 14.230 322.600 15.230 323.050 ;
        RECT 10.880 322.450 18.580 322.600 ;
        RECT 14.230 322.000 15.230 322.450 ;
        RECT 19.480 322.150 19.630 329.700 ;
        RECT 20.080 322.150 20.230 329.700 ;
        RECT 20.680 322.150 20.830 329.700 ;
        RECT 21.280 322.150 21.430 329.700 ;
        RECT 21.880 322.150 22.030 329.700 ;
        RECT 22.480 322.150 22.630 329.700 ;
        RECT 22.780 329.550 23.930 329.700 ;
        RECT 24.580 329.550 24.880 330.450 ;
        RECT 25.530 330.300 26.680 330.450 ;
        RECT 26.830 330.300 26.980 337.850 ;
        RECT 27.430 330.300 27.580 337.850 ;
        RECT 28.030 330.300 28.180 337.850 ;
        RECT 28.630 330.300 28.780 337.850 ;
        RECT 29.230 330.300 29.380 337.850 ;
        RECT 29.830 330.300 29.980 337.850 ;
        RECT 34.230 337.550 35.230 338.000 ;
        RECT 30.880 337.400 38.580 337.550 ;
        RECT 34.230 336.950 35.230 337.400 ;
        RECT 30.880 336.800 38.580 336.950 ;
        RECT 34.230 336.350 35.230 336.800 ;
        RECT 30.880 336.200 38.580 336.350 ;
        RECT 34.230 335.750 35.230 336.200 ;
        RECT 30.880 335.600 38.580 335.750 ;
        RECT 34.230 335.150 35.230 335.600 ;
        RECT 30.880 335.000 38.580 335.150 ;
        RECT 34.230 334.550 35.230 335.000 ;
        RECT 30.880 334.400 38.580 334.550 ;
        RECT 34.230 333.950 35.230 334.400 ;
        RECT 30.880 333.800 38.580 333.950 ;
        RECT 34.230 333.350 35.230 333.800 ;
        RECT 30.880 333.200 38.580 333.350 ;
        RECT 34.230 332.750 35.230 333.200 ;
        RECT 30.880 332.600 38.580 332.750 ;
        RECT 34.230 332.150 35.230 332.600 ;
        RECT 30.880 332.000 38.580 332.150 ;
        RECT 34.230 331.550 35.230 332.000 ;
        RECT 30.880 331.400 38.580 331.550 ;
        RECT 34.230 330.950 35.230 331.400 ;
        RECT 30.880 330.800 38.580 330.950 ;
        RECT 34.230 330.300 35.230 330.800 ;
        RECT 39.480 330.300 39.630 337.850 ;
        RECT 40.080 330.300 40.230 337.850 ;
        RECT 40.680 330.300 40.830 337.850 ;
        RECT 41.280 330.300 41.430 337.850 ;
        RECT 41.880 330.300 42.030 337.850 ;
        RECT 42.480 330.300 42.630 337.850 ;
        RECT 42.780 333.200 43.530 335.000 ;
        RECT 45.930 333.200 46.680 335.000 ;
        RECT 42.780 330.450 46.680 333.200 ;
        RECT 42.780 330.300 43.930 330.450 ;
        RECT 25.530 329.700 43.930 330.300 ;
        RECT 25.530 329.550 26.680 329.700 ;
        RECT 22.780 326.800 26.680 329.550 ;
        RECT 22.780 325.050 23.530 326.800 ;
        RECT 25.930 325.050 26.680 326.800 ;
        RECT 26.830 322.150 26.980 329.700 ;
        RECT 27.430 322.150 27.580 329.700 ;
        RECT 28.030 322.150 28.180 329.700 ;
        RECT 28.630 322.150 28.780 329.700 ;
        RECT 29.230 322.150 29.380 329.700 ;
        RECT 29.830 322.150 29.980 329.700 ;
        RECT 34.230 329.200 35.230 329.700 ;
        RECT 30.880 329.050 38.580 329.200 ;
        RECT 34.230 328.600 35.230 329.050 ;
        RECT 30.880 328.450 38.580 328.600 ;
        RECT 34.230 328.000 35.230 328.450 ;
        RECT 30.880 327.850 38.580 328.000 ;
        RECT 34.230 327.400 35.230 327.850 ;
        RECT 30.880 327.250 38.580 327.400 ;
        RECT 34.230 326.800 35.230 327.250 ;
        RECT 30.880 326.650 38.580 326.800 ;
        RECT 34.230 326.200 35.230 326.650 ;
        RECT 30.880 326.050 38.580 326.200 ;
        RECT 34.230 325.600 35.230 326.050 ;
        RECT 30.880 325.450 38.580 325.600 ;
        RECT 34.230 325.000 35.230 325.450 ;
        RECT 30.880 324.850 38.580 325.000 ;
        RECT 34.230 324.400 35.230 324.850 ;
        RECT 30.880 324.250 38.580 324.400 ;
        RECT 34.230 323.800 35.230 324.250 ;
        RECT 30.880 323.650 38.580 323.800 ;
        RECT 34.230 323.200 35.230 323.650 ;
        RECT 30.880 323.050 38.580 323.200 ;
        RECT 34.230 322.600 35.230 323.050 ;
        RECT 30.880 322.450 38.580 322.600 ;
        RECT 34.230 322.000 35.230 322.450 ;
        RECT 39.480 322.150 39.630 329.700 ;
        RECT 40.080 322.150 40.230 329.700 ;
        RECT 40.680 322.150 40.830 329.700 ;
        RECT 41.280 322.150 41.430 329.700 ;
        RECT 41.880 322.150 42.030 329.700 ;
        RECT 42.480 322.150 42.630 329.700 ;
        RECT 42.780 329.550 43.930 329.700 ;
        RECT 44.580 329.550 44.880 330.450 ;
        RECT 45.530 330.300 46.680 330.450 ;
        RECT 46.830 330.300 46.980 337.850 ;
        RECT 47.430 330.300 47.580 337.850 ;
        RECT 48.030 330.300 48.180 337.850 ;
        RECT 48.630 330.300 48.780 337.850 ;
        RECT 49.230 330.300 49.380 337.850 ;
        RECT 49.830 330.300 49.980 337.850 ;
        RECT 54.230 337.550 55.230 338.000 ;
        RECT 50.880 337.400 58.580 337.550 ;
        RECT 54.230 336.950 55.230 337.400 ;
        RECT 50.880 336.800 58.580 336.950 ;
        RECT 54.230 336.350 55.230 336.800 ;
        RECT 50.880 336.200 58.580 336.350 ;
        RECT 54.230 335.750 55.230 336.200 ;
        RECT 50.880 335.600 58.580 335.750 ;
        RECT 54.230 335.150 55.230 335.600 ;
        RECT 50.880 335.000 58.580 335.150 ;
        RECT 54.230 334.550 55.230 335.000 ;
        RECT 50.880 334.400 58.580 334.550 ;
        RECT 54.230 333.950 55.230 334.400 ;
        RECT 50.880 333.800 58.580 333.950 ;
        RECT 54.230 333.350 55.230 333.800 ;
        RECT 50.880 333.200 58.580 333.350 ;
        RECT 54.230 332.750 55.230 333.200 ;
        RECT 50.880 332.600 58.580 332.750 ;
        RECT 54.230 332.150 55.230 332.600 ;
        RECT 50.880 332.000 58.580 332.150 ;
        RECT 54.230 331.550 55.230 332.000 ;
        RECT 50.880 331.400 58.580 331.550 ;
        RECT 54.230 330.950 55.230 331.400 ;
        RECT 50.880 330.800 58.580 330.950 ;
        RECT 54.230 330.300 55.230 330.800 ;
        RECT 59.480 330.300 59.630 337.850 ;
        RECT 60.080 330.300 60.230 337.850 ;
        RECT 60.680 330.300 60.830 337.850 ;
        RECT 61.280 330.300 61.430 337.850 ;
        RECT 61.880 330.300 62.030 337.850 ;
        RECT 62.480 330.300 62.630 337.850 ;
        RECT 62.780 333.200 63.530 335.000 ;
        RECT 65.930 333.200 66.680 335.000 ;
        RECT 62.780 330.450 66.680 333.200 ;
        RECT 62.780 330.300 63.930 330.450 ;
        RECT 45.530 329.700 63.930 330.300 ;
        RECT 45.530 329.550 46.680 329.700 ;
        RECT 42.780 326.800 46.680 329.550 ;
        RECT 42.780 325.050 43.530 326.800 ;
        RECT 45.930 325.050 46.680 326.800 ;
        RECT 46.830 322.150 46.980 329.700 ;
        RECT 47.430 322.150 47.580 329.700 ;
        RECT 48.030 322.150 48.180 329.700 ;
        RECT 48.630 322.150 48.780 329.700 ;
        RECT 49.230 322.150 49.380 329.700 ;
        RECT 49.830 322.150 49.980 329.700 ;
        RECT 54.230 329.200 55.230 329.700 ;
        RECT 50.880 329.050 58.580 329.200 ;
        RECT 54.230 328.600 55.230 329.050 ;
        RECT 50.880 328.450 58.580 328.600 ;
        RECT 54.230 328.000 55.230 328.450 ;
        RECT 50.880 327.850 58.580 328.000 ;
        RECT 54.230 327.400 55.230 327.850 ;
        RECT 50.880 327.250 58.580 327.400 ;
        RECT 54.230 326.800 55.230 327.250 ;
        RECT 50.880 326.650 58.580 326.800 ;
        RECT 54.230 326.200 55.230 326.650 ;
        RECT 50.880 326.050 58.580 326.200 ;
        RECT 54.230 325.600 55.230 326.050 ;
        RECT 50.880 325.450 58.580 325.600 ;
        RECT 54.230 325.000 55.230 325.450 ;
        RECT 50.880 324.850 58.580 325.000 ;
        RECT 54.230 324.400 55.230 324.850 ;
        RECT 50.880 324.250 58.580 324.400 ;
        RECT 54.230 323.800 55.230 324.250 ;
        RECT 50.880 323.650 58.580 323.800 ;
        RECT 54.230 323.200 55.230 323.650 ;
        RECT 50.880 323.050 58.580 323.200 ;
        RECT 54.230 322.600 55.230 323.050 ;
        RECT 50.880 322.450 58.580 322.600 ;
        RECT 54.230 322.000 55.230 322.450 ;
        RECT 59.480 322.150 59.630 329.700 ;
        RECT 60.080 322.150 60.230 329.700 ;
        RECT 60.680 322.150 60.830 329.700 ;
        RECT 61.280 322.150 61.430 329.700 ;
        RECT 61.880 322.150 62.030 329.700 ;
        RECT 62.480 322.150 62.630 329.700 ;
        RECT 62.780 329.550 63.930 329.700 ;
        RECT 64.580 329.550 64.880 330.450 ;
        RECT 65.530 330.300 66.680 330.450 ;
        RECT 66.830 330.300 66.980 337.850 ;
        RECT 67.430 330.300 67.580 337.850 ;
        RECT 68.030 330.300 68.180 337.850 ;
        RECT 68.630 330.300 68.780 337.850 ;
        RECT 69.230 330.300 69.380 337.850 ;
        RECT 69.830 330.300 69.980 337.850 ;
        RECT 74.230 337.550 75.230 338.000 ;
        RECT 70.880 337.400 78.580 337.550 ;
        RECT 74.230 336.950 75.230 337.400 ;
        RECT 70.880 336.800 78.580 336.950 ;
        RECT 74.230 336.350 75.230 336.800 ;
        RECT 70.880 336.200 78.580 336.350 ;
        RECT 74.230 335.750 75.230 336.200 ;
        RECT 70.880 335.600 78.580 335.750 ;
        RECT 74.230 335.150 75.230 335.600 ;
        RECT 70.880 335.000 78.580 335.150 ;
        RECT 74.230 334.550 75.230 335.000 ;
        RECT 70.880 334.400 78.580 334.550 ;
        RECT 74.230 333.950 75.230 334.400 ;
        RECT 70.880 333.800 78.580 333.950 ;
        RECT 74.230 333.350 75.230 333.800 ;
        RECT 70.880 333.200 78.580 333.350 ;
        RECT 74.230 332.750 75.230 333.200 ;
        RECT 70.880 332.600 78.580 332.750 ;
        RECT 74.230 332.150 75.230 332.600 ;
        RECT 70.880 332.000 78.580 332.150 ;
        RECT 74.230 331.550 75.230 332.000 ;
        RECT 70.880 331.400 78.580 331.550 ;
        RECT 74.230 330.950 75.230 331.400 ;
        RECT 70.880 330.800 78.580 330.950 ;
        RECT 74.230 330.300 75.230 330.800 ;
        RECT 79.480 330.300 79.630 337.850 ;
        RECT 80.080 330.300 80.230 337.850 ;
        RECT 80.680 330.300 80.830 337.850 ;
        RECT 81.280 330.300 81.430 337.850 ;
        RECT 81.880 330.300 82.030 337.850 ;
        RECT 82.480 330.300 82.630 337.850 ;
        RECT 82.780 333.200 83.530 335.000 ;
        RECT 85.930 333.200 86.680 335.000 ;
        RECT 82.780 330.450 86.680 333.200 ;
        RECT 82.780 330.300 83.930 330.450 ;
        RECT 65.530 329.700 83.930 330.300 ;
        RECT 65.530 329.550 66.680 329.700 ;
        RECT 62.780 326.800 66.680 329.550 ;
        RECT 62.780 325.050 63.530 326.800 ;
        RECT 65.930 325.050 66.680 326.800 ;
        RECT 66.830 322.150 66.980 329.700 ;
        RECT 67.430 322.150 67.580 329.700 ;
        RECT 68.030 322.150 68.180 329.700 ;
        RECT 68.630 322.150 68.780 329.700 ;
        RECT 69.230 322.150 69.380 329.700 ;
        RECT 69.830 322.150 69.980 329.700 ;
        RECT 74.230 329.200 75.230 329.700 ;
        RECT 70.880 329.050 78.580 329.200 ;
        RECT 74.230 328.600 75.230 329.050 ;
        RECT 70.880 328.450 78.580 328.600 ;
        RECT 74.230 328.000 75.230 328.450 ;
        RECT 70.880 327.850 78.580 328.000 ;
        RECT 74.230 327.400 75.230 327.850 ;
        RECT 70.880 327.250 78.580 327.400 ;
        RECT 74.230 326.800 75.230 327.250 ;
        RECT 70.880 326.650 78.580 326.800 ;
        RECT 74.230 326.200 75.230 326.650 ;
        RECT 70.880 326.050 78.580 326.200 ;
        RECT 74.230 325.600 75.230 326.050 ;
        RECT 70.880 325.450 78.580 325.600 ;
        RECT 74.230 325.000 75.230 325.450 ;
        RECT 70.880 324.850 78.580 325.000 ;
        RECT 74.230 324.400 75.230 324.850 ;
        RECT 70.880 324.250 78.580 324.400 ;
        RECT 74.230 323.800 75.230 324.250 ;
        RECT 70.880 323.650 78.580 323.800 ;
        RECT 74.230 323.200 75.230 323.650 ;
        RECT 70.880 323.050 78.580 323.200 ;
        RECT 74.230 322.600 75.230 323.050 ;
        RECT 70.880 322.450 78.580 322.600 ;
        RECT 74.230 322.000 75.230 322.450 ;
        RECT 79.480 322.150 79.630 329.700 ;
        RECT 80.080 322.150 80.230 329.700 ;
        RECT 80.680 322.150 80.830 329.700 ;
        RECT 81.280 322.150 81.430 329.700 ;
        RECT 81.880 322.150 82.030 329.700 ;
        RECT 82.480 322.150 82.630 329.700 ;
        RECT 82.780 329.550 83.930 329.700 ;
        RECT 84.580 329.550 84.880 330.450 ;
        RECT 85.530 330.300 86.680 330.450 ;
        RECT 86.830 330.300 86.980 337.850 ;
        RECT 87.430 330.300 87.580 337.850 ;
        RECT 88.030 330.300 88.180 337.850 ;
        RECT 88.630 330.300 88.780 337.850 ;
        RECT 89.230 330.300 89.380 337.850 ;
        RECT 89.830 330.300 89.980 337.850 ;
        RECT 94.230 337.550 95.230 338.000 ;
        RECT 90.880 337.400 98.580 337.550 ;
        RECT 94.230 336.950 95.230 337.400 ;
        RECT 90.880 336.800 98.580 336.950 ;
        RECT 94.230 336.350 95.230 336.800 ;
        RECT 90.880 336.200 98.580 336.350 ;
        RECT 94.230 335.750 95.230 336.200 ;
        RECT 90.880 335.600 98.580 335.750 ;
        RECT 94.230 335.150 95.230 335.600 ;
        RECT 90.880 335.000 98.580 335.150 ;
        RECT 94.230 334.550 95.230 335.000 ;
        RECT 90.880 334.400 98.580 334.550 ;
        RECT 94.230 333.950 95.230 334.400 ;
        RECT 90.880 333.800 98.580 333.950 ;
        RECT 94.230 333.350 95.230 333.800 ;
        RECT 90.880 333.200 98.580 333.350 ;
        RECT 94.230 332.750 95.230 333.200 ;
        RECT 90.880 332.600 98.580 332.750 ;
        RECT 94.230 332.150 95.230 332.600 ;
        RECT 90.880 332.000 98.580 332.150 ;
        RECT 94.230 331.550 95.230 332.000 ;
        RECT 90.880 331.400 98.580 331.550 ;
        RECT 94.230 330.950 95.230 331.400 ;
        RECT 90.880 330.800 98.580 330.950 ;
        RECT 94.230 330.300 95.230 330.800 ;
        RECT 99.480 330.300 99.630 337.850 ;
        RECT 100.080 330.300 100.230 337.850 ;
        RECT 100.680 330.300 100.830 337.850 ;
        RECT 101.280 330.300 101.430 337.850 ;
        RECT 101.880 330.300 102.030 337.850 ;
        RECT 102.480 330.300 102.630 337.850 ;
        RECT 102.780 333.200 103.530 335.000 ;
        RECT 105.930 333.200 106.680 335.000 ;
        RECT 102.780 330.450 106.680 333.200 ;
        RECT 102.780 330.300 103.930 330.450 ;
        RECT 85.530 329.700 103.930 330.300 ;
        RECT 85.530 329.550 86.680 329.700 ;
        RECT 82.780 326.800 86.680 329.550 ;
        RECT 82.780 325.050 83.530 326.800 ;
        RECT 85.930 325.050 86.680 326.800 ;
        RECT 86.830 322.150 86.980 329.700 ;
        RECT 87.430 322.150 87.580 329.700 ;
        RECT 88.030 322.150 88.180 329.700 ;
        RECT 88.630 322.150 88.780 329.700 ;
        RECT 89.230 322.150 89.380 329.700 ;
        RECT 89.830 322.150 89.980 329.700 ;
        RECT 94.230 329.200 95.230 329.700 ;
        RECT 90.880 329.050 98.580 329.200 ;
        RECT 94.230 328.600 95.230 329.050 ;
        RECT 90.880 328.450 98.580 328.600 ;
        RECT 94.230 328.000 95.230 328.450 ;
        RECT 90.880 327.850 98.580 328.000 ;
        RECT 94.230 327.400 95.230 327.850 ;
        RECT 90.880 327.250 98.580 327.400 ;
        RECT 94.230 326.800 95.230 327.250 ;
        RECT 90.880 326.650 98.580 326.800 ;
        RECT 94.230 326.200 95.230 326.650 ;
        RECT 90.880 326.050 98.580 326.200 ;
        RECT 94.230 325.600 95.230 326.050 ;
        RECT 90.880 325.450 98.580 325.600 ;
        RECT 94.230 325.000 95.230 325.450 ;
        RECT 90.880 324.850 98.580 325.000 ;
        RECT 94.230 324.400 95.230 324.850 ;
        RECT 90.880 324.250 98.580 324.400 ;
        RECT 94.230 323.800 95.230 324.250 ;
        RECT 90.880 323.650 98.580 323.800 ;
        RECT 94.230 323.200 95.230 323.650 ;
        RECT 90.880 323.050 98.580 323.200 ;
        RECT 94.230 322.600 95.230 323.050 ;
        RECT 90.880 322.450 98.580 322.600 ;
        RECT 94.230 322.000 95.230 322.450 ;
        RECT 99.480 322.150 99.630 329.700 ;
        RECT 100.080 322.150 100.230 329.700 ;
        RECT 100.680 322.150 100.830 329.700 ;
        RECT 101.280 322.150 101.430 329.700 ;
        RECT 101.880 322.150 102.030 329.700 ;
        RECT 102.480 322.150 102.630 329.700 ;
        RECT 102.780 329.550 103.930 329.700 ;
        RECT 104.580 329.550 104.880 330.450 ;
        RECT 105.530 330.300 106.680 330.450 ;
        RECT 106.830 330.300 106.980 337.850 ;
        RECT 107.430 330.300 107.580 337.850 ;
        RECT 108.030 330.300 108.180 337.850 ;
        RECT 108.630 330.300 108.780 337.850 ;
        RECT 109.230 330.300 109.380 337.850 ;
        RECT 109.830 330.300 109.980 337.850 ;
        RECT 114.230 337.550 115.230 338.000 ;
        RECT 110.880 337.400 118.580 337.550 ;
        RECT 114.230 336.950 115.230 337.400 ;
        RECT 110.880 336.800 118.580 336.950 ;
        RECT 114.230 336.350 115.230 336.800 ;
        RECT 110.880 336.200 118.580 336.350 ;
        RECT 114.230 335.750 115.230 336.200 ;
        RECT 110.880 335.600 118.580 335.750 ;
        RECT 114.230 335.150 115.230 335.600 ;
        RECT 110.880 335.000 118.580 335.150 ;
        RECT 114.230 334.550 115.230 335.000 ;
        RECT 110.880 334.400 118.580 334.550 ;
        RECT 114.230 333.950 115.230 334.400 ;
        RECT 110.880 333.800 118.580 333.950 ;
        RECT 114.230 333.350 115.230 333.800 ;
        RECT 110.880 333.200 118.580 333.350 ;
        RECT 114.230 332.750 115.230 333.200 ;
        RECT 110.880 332.600 118.580 332.750 ;
        RECT 114.230 332.150 115.230 332.600 ;
        RECT 110.880 332.000 118.580 332.150 ;
        RECT 114.230 331.550 115.230 332.000 ;
        RECT 110.880 331.400 118.580 331.550 ;
        RECT 114.230 330.950 115.230 331.400 ;
        RECT 110.880 330.800 118.580 330.950 ;
        RECT 114.230 330.300 115.230 330.800 ;
        RECT 119.480 330.300 119.630 337.850 ;
        RECT 120.080 330.300 120.230 337.850 ;
        RECT 120.680 330.300 120.830 337.850 ;
        RECT 121.280 330.300 121.430 337.850 ;
        RECT 121.880 330.300 122.030 337.850 ;
        RECT 122.480 330.300 122.630 337.850 ;
        RECT 122.780 333.200 123.530 335.000 ;
        RECT 122.780 330.480 124.730 333.200 ;
        RECT 122.780 330.450 131.850 330.480 ;
        RECT 122.780 330.300 123.930 330.450 ;
        RECT 105.530 329.700 123.930 330.300 ;
        RECT 105.530 329.550 106.680 329.700 ;
        RECT 102.780 326.800 106.680 329.550 ;
        RECT 102.780 325.050 103.530 326.800 ;
        RECT 105.930 325.050 106.680 326.800 ;
        RECT 106.830 322.150 106.980 329.700 ;
        RECT 107.430 322.150 107.580 329.700 ;
        RECT 108.030 322.150 108.180 329.700 ;
        RECT 108.630 322.150 108.780 329.700 ;
        RECT 109.230 322.150 109.380 329.700 ;
        RECT 109.830 322.150 109.980 329.700 ;
        RECT 114.230 329.200 115.230 329.700 ;
        RECT 110.880 329.050 118.580 329.200 ;
        RECT 114.230 328.600 115.230 329.050 ;
        RECT 110.880 328.450 118.580 328.600 ;
        RECT 114.230 328.000 115.230 328.450 ;
        RECT 110.880 327.850 118.580 328.000 ;
        RECT 114.230 327.400 115.230 327.850 ;
        RECT 110.880 327.250 118.580 327.400 ;
        RECT 114.230 326.800 115.230 327.250 ;
        RECT 110.880 326.650 118.580 326.800 ;
        RECT 114.230 326.200 115.230 326.650 ;
        RECT 110.880 326.050 118.580 326.200 ;
        RECT 114.230 325.600 115.230 326.050 ;
        RECT 110.880 325.450 118.580 325.600 ;
        RECT 114.230 325.000 115.230 325.450 ;
        RECT 110.880 324.850 118.580 325.000 ;
        RECT 114.230 324.400 115.230 324.850 ;
        RECT 110.880 324.250 118.580 324.400 ;
        RECT 114.230 323.800 115.230 324.250 ;
        RECT 110.880 323.650 118.580 323.800 ;
        RECT 114.230 323.200 115.230 323.650 ;
        RECT 110.880 323.050 118.580 323.200 ;
        RECT 114.230 322.600 115.230 323.050 ;
        RECT 110.880 322.450 118.580 322.600 ;
        RECT 114.230 322.000 115.230 322.450 ;
        RECT 119.480 322.150 119.630 329.700 ;
        RECT 120.080 322.150 120.230 329.700 ;
        RECT 120.680 322.150 120.830 329.700 ;
        RECT 121.280 322.150 121.430 329.700 ;
        RECT 121.880 322.150 122.030 329.700 ;
        RECT 122.480 322.150 122.630 329.700 ;
        RECT 122.780 329.550 123.930 329.700 ;
        RECT 124.580 329.550 131.850 330.450 ;
        RECT 122.780 329.205 131.850 329.550 ;
        RECT 122.780 326.800 124.730 329.205 ;
        RECT 122.780 325.050 123.530 326.800 ;
        RECT 10.880 321.850 18.580 322.000 ;
        RECT 30.880 321.850 38.580 322.000 ;
        RECT 50.880 321.850 58.580 322.000 ;
        RECT 70.880 321.850 78.580 322.000 ;
        RECT 90.880 321.850 98.580 322.000 ;
        RECT 110.880 321.850 118.580 322.000 ;
        RECT 14.230 321.200 15.230 321.850 ;
        RECT 34.230 321.200 35.230 321.850 ;
        RECT 54.230 321.200 55.230 321.850 ;
        RECT 74.230 321.200 75.230 321.850 ;
        RECT 94.230 321.200 95.230 321.850 ;
        RECT 114.230 321.200 115.230 321.850 ;
        RECT 11.530 318.800 17.930 321.200 ;
        RECT 31.530 318.800 37.930 321.200 ;
        RECT 51.530 318.800 57.930 321.200 ;
        RECT 71.530 318.800 77.930 321.200 ;
        RECT 91.530 318.800 97.930 321.200 ;
        RECT 111.530 318.800 117.930 321.200 ;
        RECT 14.230 318.150 15.230 318.800 ;
        RECT 34.230 318.150 35.230 318.800 ;
        RECT 54.230 318.150 55.230 318.800 ;
        RECT 74.230 318.150 75.230 318.800 ;
        RECT 94.230 318.150 95.230 318.800 ;
        RECT 114.230 318.150 115.230 318.800 ;
        RECT 10.880 318.000 18.580 318.150 ;
        RECT 30.880 318.000 38.580 318.150 ;
        RECT 50.880 318.000 58.580 318.150 ;
        RECT 70.880 318.000 78.580 318.150 ;
        RECT 90.880 318.000 98.580 318.150 ;
        RECT 110.880 318.000 118.580 318.150 ;
        RECT 5.930 313.200 6.680 315.000 ;
        RECT 4.730 310.450 6.680 313.200 ;
        RECT 4.730 309.550 4.880 310.450 ;
        RECT 5.530 310.300 6.680 310.450 ;
        RECT 6.830 310.300 6.980 317.850 ;
        RECT 7.430 310.300 7.580 317.850 ;
        RECT 8.030 310.300 8.180 317.850 ;
        RECT 8.630 310.300 8.780 317.850 ;
        RECT 9.230 310.300 9.380 317.850 ;
        RECT 9.830 310.300 9.980 317.850 ;
        RECT 14.230 317.550 15.230 318.000 ;
        RECT 10.880 317.400 18.580 317.550 ;
        RECT 14.230 316.950 15.230 317.400 ;
        RECT 10.880 316.800 18.580 316.950 ;
        RECT 14.230 316.350 15.230 316.800 ;
        RECT 10.880 316.200 18.580 316.350 ;
        RECT 14.230 315.750 15.230 316.200 ;
        RECT 10.880 315.600 18.580 315.750 ;
        RECT 14.230 315.150 15.230 315.600 ;
        RECT 10.880 315.000 18.580 315.150 ;
        RECT 14.230 314.550 15.230 315.000 ;
        RECT 10.880 314.400 18.580 314.550 ;
        RECT 14.230 313.950 15.230 314.400 ;
        RECT 10.880 313.800 18.580 313.950 ;
        RECT 14.230 313.350 15.230 313.800 ;
        RECT 10.880 313.200 18.580 313.350 ;
        RECT 14.230 312.750 15.230 313.200 ;
        RECT 10.880 312.600 18.580 312.750 ;
        RECT 14.230 312.150 15.230 312.600 ;
        RECT 10.880 312.000 18.580 312.150 ;
        RECT 14.230 311.550 15.230 312.000 ;
        RECT 10.880 311.400 18.580 311.550 ;
        RECT 14.230 310.950 15.230 311.400 ;
        RECT 10.880 310.800 18.580 310.950 ;
        RECT 14.230 310.300 15.230 310.800 ;
        RECT 19.480 310.300 19.630 317.850 ;
        RECT 20.080 310.300 20.230 317.850 ;
        RECT 20.680 310.300 20.830 317.850 ;
        RECT 21.280 310.300 21.430 317.850 ;
        RECT 21.880 310.300 22.030 317.850 ;
        RECT 22.480 310.300 22.630 317.850 ;
        RECT 22.780 313.200 23.530 315.000 ;
        RECT 25.930 313.200 26.680 315.000 ;
        RECT 22.780 310.450 26.680 313.200 ;
        RECT 22.780 310.300 23.930 310.450 ;
        RECT 5.530 309.700 23.930 310.300 ;
        RECT 5.530 309.550 6.680 309.700 ;
        RECT 4.730 306.800 6.680 309.550 ;
        RECT 5.930 305.050 6.680 306.800 ;
        RECT 6.830 302.150 6.980 309.700 ;
        RECT 7.430 302.150 7.580 309.700 ;
        RECT 8.030 302.150 8.180 309.700 ;
        RECT 8.630 302.150 8.780 309.700 ;
        RECT 9.230 302.150 9.380 309.700 ;
        RECT 9.830 302.150 9.980 309.700 ;
        RECT 14.230 309.200 15.230 309.700 ;
        RECT 10.880 309.050 18.580 309.200 ;
        RECT 14.230 308.600 15.230 309.050 ;
        RECT 10.880 308.450 18.580 308.600 ;
        RECT 14.230 308.000 15.230 308.450 ;
        RECT 10.880 307.850 18.580 308.000 ;
        RECT 14.230 307.400 15.230 307.850 ;
        RECT 10.880 307.250 18.580 307.400 ;
        RECT 14.230 306.800 15.230 307.250 ;
        RECT 10.880 306.650 18.580 306.800 ;
        RECT 14.230 306.200 15.230 306.650 ;
        RECT 10.880 306.050 18.580 306.200 ;
        RECT 14.230 305.600 15.230 306.050 ;
        RECT 10.880 305.450 18.580 305.600 ;
        RECT 14.230 305.000 15.230 305.450 ;
        RECT 10.880 304.850 18.580 305.000 ;
        RECT 14.230 304.400 15.230 304.850 ;
        RECT 10.880 304.250 18.580 304.400 ;
        RECT 14.230 303.800 15.230 304.250 ;
        RECT 10.880 303.650 18.580 303.800 ;
        RECT 14.230 303.200 15.230 303.650 ;
        RECT 10.880 303.050 18.580 303.200 ;
        RECT 14.230 302.600 15.230 303.050 ;
        RECT 10.880 302.450 18.580 302.600 ;
        RECT 14.230 302.000 15.230 302.450 ;
        RECT 19.480 302.150 19.630 309.700 ;
        RECT 20.080 302.150 20.230 309.700 ;
        RECT 20.680 302.150 20.830 309.700 ;
        RECT 21.280 302.150 21.430 309.700 ;
        RECT 21.880 302.150 22.030 309.700 ;
        RECT 22.480 302.150 22.630 309.700 ;
        RECT 22.780 309.550 23.930 309.700 ;
        RECT 24.580 309.550 24.880 310.450 ;
        RECT 25.530 310.300 26.680 310.450 ;
        RECT 26.830 310.300 26.980 317.850 ;
        RECT 27.430 310.300 27.580 317.850 ;
        RECT 28.030 310.300 28.180 317.850 ;
        RECT 28.630 310.300 28.780 317.850 ;
        RECT 29.230 310.300 29.380 317.850 ;
        RECT 29.830 310.300 29.980 317.850 ;
        RECT 34.230 317.550 35.230 318.000 ;
        RECT 30.880 317.400 38.580 317.550 ;
        RECT 34.230 316.950 35.230 317.400 ;
        RECT 30.880 316.800 38.580 316.950 ;
        RECT 34.230 316.350 35.230 316.800 ;
        RECT 30.880 316.200 38.580 316.350 ;
        RECT 34.230 315.750 35.230 316.200 ;
        RECT 30.880 315.600 38.580 315.750 ;
        RECT 34.230 315.150 35.230 315.600 ;
        RECT 30.880 315.000 38.580 315.150 ;
        RECT 34.230 314.550 35.230 315.000 ;
        RECT 30.880 314.400 38.580 314.550 ;
        RECT 34.230 313.950 35.230 314.400 ;
        RECT 30.880 313.800 38.580 313.950 ;
        RECT 34.230 313.350 35.230 313.800 ;
        RECT 30.880 313.200 38.580 313.350 ;
        RECT 34.230 312.750 35.230 313.200 ;
        RECT 30.880 312.600 38.580 312.750 ;
        RECT 34.230 312.150 35.230 312.600 ;
        RECT 30.880 312.000 38.580 312.150 ;
        RECT 34.230 311.550 35.230 312.000 ;
        RECT 30.880 311.400 38.580 311.550 ;
        RECT 34.230 310.950 35.230 311.400 ;
        RECT 30.880 310.800 38.580 310.950 ;
        RECT 34.230 310.300 35.230 310.800 ;
        RECT 39.480 310.300 39.630 317.850 ;
        RECT 40.080 310.300 40.230 317.850 ;
        RECT 40.680 310.300 40.830 317.850 ;
        RECT 41.280 310.300 41.430 317.850 ;
        RECT 41.880 310.300 42.030 317.850 ;
        RECT 42.480 310.300 42.630 317.850 ;
        RECT 42.780 313.200 43.530 315.000 ;
        RECT 45.930 313.200 46.680 315.000 ;
        RECT 42.780 310.450 46.680 313.200 ;
        RECT 42.780 310.300 43.930 310.450 ;
        RECT 25.530 309.700 43.930 310.300 ;
        RECT 25.530 309.550 26.680 309.700 ;
        RECT 22.780 306.800 26.680 309.550 ;
        RECT 22.780 305.050 23.530 306.800 ;
        RECT 25.930 305.050 26.680 306.800 ;
        RECT 26.830 302.150 26.980 309.700 ;
        RECT 27.430 302.150 27.580 309.700 ;
        RECT 28.030 302.150 28.180 309.700 ;
        RECT 28.630 302.150 28.780 309.700 ;
        RECT 29.230 302.150 29.380 309.700 ;
        RECT 29.830 302.150 29.980 309.700 ;
        RECT 34.230 309.200 35.230 309.700 ;
        RECT 30.880 309.050 38.580 309.200 ;
        RECT 34.230 308.600 35.230 309.050 ;
        RECT 30.880 308.450 38.580 308.600 ;
        RECT 34.230 308.000 35.230 308.450 ;
        RECT 30.880 307.850 38.580 308.000 ;
        RECT 34.230 307.400 35.230 307.850 ;
        RECT 30.880 307.250 38.580 307.400 ;
        RECT 34.230 306.800 35.230 307.250 ;
        RECT 30.880 306.650 38.580 306.800 ;
        RECT 34.230 306.200 35.230 306.650 ;
        RECT 30.880 306.050 38.580 306.200 ;
        RECT 34.230 305.600 35.230 306.050 ;
        RECT 30.880 305.450 38.580 305.600 ;
        RECT 34.230 305.000 35.230 305.450 ;
        RECT 30.880 304.850 38.580 305.000 ;
        RECT 34.230 304.400 35.230 304.850 ;
        RECT 30.880 304.250 38.580 304.400 ;
        RECT 34.230 303.800 35.230 304.250 ;
        RECT 30.880 303.650 38.580 303.800 ;
        RECT 34.230 303.200 35.230 303.650 ;
        RECT 30.880 303.050 38.580 303.200 ;
        RECT 34.230 302.600 35.230 303.050 ;
        RECT 30.880 302.450 38.580 302.600 ;
        RECT 34.230 302.000 35.230 302.450 ;
        RECT 39.480 302.150 39.630 309.700 ;
        RECT 40.080 302.150 40.230 309.700 ;
        RECT 40.680 302.150 40.830 309.700 ;
        RECT 41.280 302.150 41.430 309.700 ;
        RECT 41.880 302.150 42.030 309.700 ;
        RECT 42.480 302.150 42.630 309.700 ;
        RECT 42.780 309.550 43.930 309.700 ;
        RECT 44.580 309.550 44.880 310.450 ;
        RECT 45.530 310.300 46.680 310.450 ;
        RECT 46.830 310.300 46.980 317.850 ;
        RECT 47.430 310.300 47.580 317.850 ;
        RECT 48.030 310.300 48.180 317.850 ;
        RECT 48.630 310.300 48.780 317.850 ;
        RECT 49.230 310.300 49.380 317.850 ;
        RECT 49.830 310.300 49.980 317.850 ;
        RECT 54.230 317.550 55.230 318.000 ;
        RECT 50.880 317.400 58.580 317.550 ;
        RECT 54.230 316.950 55.230 317.400 ;
        RECT 50.880 316.800 58.580 316.950 ;
        RECT 54.230 316.350 55.230 316.800 ;
        RECT 50.880 316.200 58.580 316.350 ;
        RECT 54.230 315.750 55.230 316.200 ;
        RECT 50.880 315.600 58.580 315.750 ;
        RECT 54.230 315.150 55.230 315.600 ;
        RECT 50.880 315.000 58.580 315.150 ;
        RECT 54.230 314.550 55.230 315.000 ;
        RECT 50.880 314.400 58.580 314.550 ;
        RECT 54.230 313.950 55.230 314.400 ;
        RECT 50.880 313.800 58.580 313.950 ;
        RECT 54.230 313.350 55.230 313.800 ;
        RECT 50.880 313.200 58.580 313.350 ;
        RECT 54.230 312.750 55.230 313.200 ;
        RECT 50.880 312.600 58.580 312.750 ;
        RECT 54.230 312.150 55.230 312.600 ;
        RECT 50.880 312.000 58.580 312.150 ;
        RECT 54.230 311.550 55.230 312.000 ;
        RECT 50.880 311.400 58.580 311.550 ;
        RECT 54.230 310.950 55.230 311.400 ;
        RECT 50.880 310.800 58.580 310.950 ;
        RECT 54.230 310.300 55.230 310.800 ;
        RECT 59.480 310.300 59.630 317.850 ;
        RECT 60.080 310.300 60.230 317.850 ;
        RECT 60.680 310.300 60.830 317.850 ;
        RECT 61.280 310.300 61.430 317.850 ;
        RECT 61.880 310.300 62.030 317.850 ;
        RECT 62.480 310.300 62.630 317.850 ;
        RECT 62.780 313.200 63.530 315.000 ;
        RECT 65.930 313.200 66.680 315.000 ;
        RECT 62.780 310.450 66.680 313.200 ;
        RECT 62.780 310.300 63.930 310.450 ;
        RECT 45.530 309.700 63.930 310.300 ;
        RECT 45.530 309.550 46.680 309.700 ;
        RECT 42.780 306.800 46.680 309.550 ;
        RECT 42.780 305.050 43.530 306.800 ;
        RECT 45.930 305.050 46.680 306.800 ;
        RECT 46.830 302.150 46.980 309.700 ;
        RECT 47.430 302.150 47.580 309.700 ;
        RECT 48.030 302.150 48.180 309.700 ;
        RECT 48.630 302.150 48.780 309.700 ;
        RECT 49.230 302.150 49.380 309.700 ;
        RECT 49.830 302.150 49.980 309.700 ;
        RECT 54.230 309.200 55.230 309.700 ;
        RECT 50.880 309.050 58.580 309.200 ;
        RECT 54.230 308.600 55.230 309.050 ;
        RECT 50.880 308.450 58.580 308.600 ;
        RECT 54.230 308.000 55.230 308.450 ;
        RECT 50.880 307.850 58.580 308.000 ;
        RECT 54.230 307.400 55.230 307.850 ;
        RECT 50.880 307.250 58.580 307.400 ;
        RECT 54.230 306.800 55.230 307.250 ;
        RECT 50.880 306.650 58.580 306.800 ;
        RECT 54.230 306.200 55.230 306.650 ;
        RECT 50.880 306.050 58.580 306.200 ;
        RECT 54.230 305.600 55.230 306.050 ;
        RECT 50.880 305.450 58.580 305.600 ;
        RECT 54.230 305.000 55.230 305.450 ;
        RECT 50.880 304.850 58.580 305.000 ;
        RECT 54.230 304.400 55.230 304.850 ;
        RECT 50.880 304.250 58.580 304.400 ;
        RECT 54.230 303.800 55.230 304.250 ;
        RECT 50.880 303.650 58.580 303.800 ;
        RECT 54.230 303.200 55.230 303.650 ;
        RECT 50.880 303.050 58.580 303.200 ;
        RECT 54.230 302.600 55.230 303.050 ;
        RECT 50.880 302.450 58.580 302.600 ;
        RECT 54.230 302.000 55.230 302.450 ;
        RECT 59.480 302.150 59.630 309.700 ;
        RECT 60.080 302.150 60.230 309.700 ;
        RECT 60.680 302.150 60.830 309.700 ;
        RECT 61.280 302.150 61.430 309.700 ;
        RECT 61.880 302.150 62.030 309.700 ;
        RECT 62.480 302.150 62.630 309.700 ;
        RECT 62.780 309.550 63.930 309.700 ;
        RECT 64.580 309.550 64.880 310.450 ;
        RECT 65.530 310.300 66.680 310.450 ;
        RECT 66.830 310.300 66.980 317.850 ;
        RECT 67.430 310.300 67.580 317.850 ;
        RECT 68.030 310.300 68.180 317.850 ;
        RECT 68.630 310.300 68.780 317.850 ;
        RECT 69.230 310.300 69.380 317.850 ;
        RECT 69.830 310.300 69.980 317.850 ;
        RECT 74.230 317.550 75.230 318.000 ;
        RECT 70.880 317.400 78.580 317.550 ;
        RECT 74.230 316.950 75.230 317.400 ;
        RECT 70.880 316.800 78.580 316.950 ;
        RECT 74.230 316.350 75.230 316.800 ;
        RECT 70.880 316.200 78.580 316.350 ;
        RECT 74.230 315.750 75.230 316.200 ;
        RECT 70.880 315.600 78.580 315.750 ;
        RECT 74.230 315.150 75.230 315.600 ;
        RECT 70.880 315.000 78.580 315.150 ;
        RECT 74.230 314.550 75.230 315.000 ;
        RECT 70.880 314.400 78.580 314.550 ;
        RECT 74.230 313.950 75.230 314.400 ;
        RECT 70.880 313.800 78.580 313.950 ;
        RECT 74.230 313.350 75.230 313.800 ;
        RECT 70.880 313.200 78.580 313.350 ;
        RECT 74.230 312.750 75.230 313.200 ;
        RECT 70.880 312.600 78.580 312.750 ;
        RECT 74.230 312.150 75.230 312.600 ;
        RECT 70.880 312.000 78.580 312.150 ;
        RECT 74.230 311.550 75.230 312.000 ;
        RECT 70.880 311.400 78.580 311.550 ;
        RECT 74.230 310.950 75.230 311.400 ;
        RECT 70.880 310.800 78.580 310.950 ;
        RECT 74.230 310.300 75.230 310.800 ;
        RECT 79.480 310.300 79.630 317.850 ;
        RECT 80.080 310.300 80.230 317.850 ;
        RECT 80.680 310.300 80.830 317.850 ;
        RECT 81.280 310.300 81.430 317.850 ;
        RECT 81.880 310.300 82.030 317.850 ;
        RECT 82.480 310.300 82.630 317.850 ;
        RECT 82.780 313.200 83.530 315.000 ;
        RECT 85.930 313.200 86.680 315.000 ;
        RECT 82.780 310.450 86.680 313.200 ;
        RECT 82.780 310.300 83.930 310.450 ;
        RECT 65.530 309.700 83.930 310.300 ;
        RECT 65.530 309.550 66.680 309.700 ;
        RECT 62.780 306.800 66.680 309.550 ;
        RECT 62.780 305.050 63.530 306.800 ;
        RECT 65.930 305.050 66.680 306.800 ;
        RECT 66.830 302.150 66.980 309.700 ;
        RECT 67.430 302.150 67.580 309.700 ;
        RECT 68.030 302.150 68.180 309.700 ;
        RECT 68.630 302.150 68.780 309.700 ;
        RECT 69.230 302.150 69.380 309.700 ;
        RECT 69.830 302.150 69.980 309.700 ;
        RECT 74.230 309.200 75.230 309.700 ;
        RECT 70.880 309.050 78.580 309.200 ;
        RECT 74.230 308.600 75.230 309.050 ;
        RECT 70.880 308.450 78.580 308.600 ;
        RECT 74.230 308.000 75.230 308.450 ;
        RECT 70.880 307.850 78.580 308.000 ;
        RECT 74.230 307.400 75.230 307.850 ;
        RECT 70.880 307.250 78.580 307.400 ;
        RECT 74.230 306.800 75.230 307.250 ;
        RECT 70.880 306.650 78.580 306.800 ;
        RECT 74.230 306.200 75.230 306.650 ;
        RECT 70.880 306.050 78.580 306.200 ;
        RECT 74.230 305.600 75.230 306.050 ;
        RECT 70.880 305.450 78.580 305.600 ;
        RECT 74.230 305.000 75.230 305.450 ;
        RECT 70.880 304.850 78.580 305.000 ;
        RECT 74.230 304.400 75.230 304.850 ;
        RECT 70.880 304.250 78.580 304.400 ;
        RECT 74.230 303.800 75.230 304.250 ;
        RECT 70.880 303.650 78.580 303.800 ;
        RECT 74.230 303.200 75.230 303.650 ;
        RECT 70.880 303.050 78.580 303.200 ;
        RECT 74.230 302.600 75.230 303.050 ;
        RECT 70.880 302.450 78.580 302.600 ;
        RECT 74.230 302.000 75.230 302.450 ;
        RECT 79.480 302.150 79.630 309.700 ;
        RECT 80.080 302.150 80.230 309.700 ;
        RECT 80.680 302.150 80.830 309.700 ;
        RECT 81.280 302.150 81.430 309.700 ;
        RECT 81.880 302.150 82.030 309.700 ;
        RECT 82.480 302.150 82.630 309.700 ;
        RECT 82.780 309.550 83.930 309.700 ;
        RECT 84.580 309.550 84.880 310.450 ;
        RECT 85.530 310.300 86.680 310.450 ;
        RECT 86.830 310.300 86.980 317.850 ;
        RECT 87.430 310.300 87.580 317.850 ;
        RECT 88.030 310.300 88.180 317.850 ;
        RECT 88.630 310.300 88.780 317.850 ;
        RECT 89.230 310.300 89.380 317.850 ;
        RECT 89.830 310.300 89.980 317.850 ;
        RECT 94.230 317.550 95.230 318.000 ;
        RECT 90.880 317.400 98.580 317.550 ;
        RECT 94.230 316.950 95.230 317.400 ;
        RECT 90.880 316.800 98.580 316.950 ;
        RECT 94.230 316.350 95.230 316.800 ;
        RECT 90.880 316.200 98.580 316.350 ;
        RECT 94.230 315.750 95.230 316.200 ;
        RECT 90.880 315.600 98.580 315.750 ;
        RECT 94.230 315.150 95.230 315.600 ;
        RECT 90.880 315.000 98.580 315.150 ;
        RECT 94.230 314.550 95.230 315.000 ;
        RECT 90.880 314.400 98.580 314.550 ;
        RECT 94.230 313.950 95.230 314.400 ;
        RECT 90.880 313.800 98.580 313.950 ;
        RECT 94.230 313.350 95.230 313.800 ;
        RECT 90.880 313.200 98.580 313.350 ;
        RECT 94.230 312.750 95.230 313.200 ;
        RECT 90.880 312.600 98.580 312.750 ;
        RECT 94.230 312.150 95.230 312.600 ;
        RECT 90.880 312.000 98.580 312.150 ;
        RECT 94.230 311.550 95.230 312.000 ;
        RECT 90.880 311.400 98.580 311.550 ;
        RECT 94.230 310.950 95.230 311.400 ;
        RECT 90.880 310.800 98.580 310.950 ;
        RECT 94.230 310.300 95.230 310.800 ;
        RECT 99.480 310.300 99.630 317.850 ;
        RECT 100.080 310.300 100.230 317.850 ;
        RECT 100.680 310.300 100.830 317.850 ;
        RECT 101.280 310.300 101.430 317.850 ;
        RECT 101.880 310.300 102.030 317.850 ;
        RECT 102.480 310.300 102.630 317.850 ;
        RECT 102.780 313.200 103.530 315.000 ;
        RECT 105.930 313.200 106.680 315.000 ;
        RECT 102.780 310.450 106.680 313.200 ;
        RECT 102.780 310.300 103.930 310.450 ;
        RECT 85.530 309.700 103.930 310.300 ;
        RECT 85.530 309.550 86.680 309.700 ;
        RECT 82.780 306.800 86.680 309.550 ;
        RECT 82.780 305.050 83.530 306.800 ;
        RECT 85.930 305.050 86.680 306.800 ;
        RECT 86.830 302.150 86.980 309.700 ;
        RECT 87.430 302.150 87.580 309.700 ;
        RECT 88.030 302.150 88.180 309.700 ;
        RECT 88.630 302.150 88.780 309.700 ;
        RECT 89.230 302.150 89.380 309.700 ;
        RECT 89.830 302.150 89.980 309.700 ;
        RECT 94.230 309.200 95.230 309.700 ;
        RECT 90.880 309.050 98.580 309.200 ;
        RECT 94.230 308.600 95.230 309.050 ;
        RECT 90.880 308.450 98.580 308.600 ;
        RECT 94.230 308.000 95.230 308.450 ;
        RECT 90.880 307.850 98.580 308.000 ;
        RECT 94.230 307.400 95.230 307.850 ;
        RECT 90.880 307.250 98.580 307.400 ;
        RECT 94.230 306.800 95.230 307.250 ;
        RECT 90.880 306.650 98.580 306.800 ;
        RECT 94.230 306.200 95.230 306.650 ;
        RECT 90.880 306.050 98.580 306.200 ;
        RECT 94.230 305.600 95.230 306.050 ;
        RECT 90.880 305.450 98.580 305.600 ;
        RECT 94.230 305.000 95.230 305.450 ;
        RECT 90.880 304.850 98.580 305.000 ;
        RECT 94.230 304.400 95.230 304.850 ;
        RECT 90.880 304.250 98.580 304.400 ;
        RECT 94.230 303.800 95.230 304.250 ;
        RECT 90.880 303.650 98.580 303.800 ;
        RECT 94.230 303.200 95.230 303.650 ;
        RECT 90.880 303.050 98.580 303.200 ;
        RECT 94.230 302.600 95.230 303.050 ;
        RECT 90.880 302.450 98.580 302.600 ;
        RECT 94.230 302.000 95.230 302.450 ;
        RECT 99.480 302.150 99.630 309.700 ;
        RECT 100.080 302.150 100.230 309.700 ;
        RECT 100.680 302.150 100.830 309.700 ;
        RECT 101.280 302.150 101.430 309.700 ;
        RECT 101.880 302.150 102.030 309.700 ;
        RECT 102.480 302.150 102.630 309.700 ;
        RECT 102.780 309.550 103.930 309.700 ;
        RECT 104.580 309.550 104.880 310.450 ;
        RECT 105.530 310.300 106.680 310.450 ;
        RECT 106.830 310.300 106.980 317.850 ;
        RECT 107.430 310.300 107.580 317.850 ;
        RECT 108.030 310.300 108.180 317.850 ;
        RECT 108.630 310.300 108.780 317.850 ;
        RECT 109.230 310.300 109.380 317.850 ;
        RECT 109.830 310.300 109.980 317.850 ;
        RECT 114.230 317.550 115.230 318.000 ;
        RECT 110.880 317.400 118.580 317.550 ;
        RECT 114.230 316.950 115.230 317.400 ;
        RECT 110.880 316.800 118.580 316.950 ;
        RECT 114.230 316.350 115.230 316.800 ;
        RECT 110.880 316.200 118.580 316.350 ;
        RECT 114.230 315.750 115.230 316.200 ;
        RECT 110.880 315.600 118.580 315.750 ;
        RECT 114.230 315.150 115.230 315.600 ;
        RECT 110.880 315.000 118.580 315.150 ;
        RECT 114.230 314.550 115.230 315.000 ;
        RECT 110.880 314.400 118.580 314.550 ;
        RECT 114.230 313.950 115.230 314.400 ;
        RECT 110.880 313.800 118.580 313.950 ;
        RECT 114.230 313.350 115.230 313.800 ;
        RECT 110.880 313.200 118.580 313.350 ;
        RECT 114.230 312.750 115.230 313.200 ;
        RECT 110.880 312.600 118.580 312.750 ;
        RECT 114.230 312.150 115.230 312.600 ;
        RECT 110.880 312.000 118.580 312.150 ;
        RECT 114.230 311.550 115.230 312.000 ;
        RECT 110.880 311.400 118.580 311.550 ;
        RECT 114.230 310.950 115.230 311.400 ;
        RECT 110.880 310.800 118.580 310.950 ;
        RECT 114.230 310.300 115.230 310.800 ;
        RECT 119.480 310.300 119.630 317.850 ;
        RECT 120.080 310.300 120.230 317.850 ;
        RECT 120.680 310.300 120.830 317.850 ;
        RECT 121.280 310.300 121.430 317.850 ;
        RECT 121.880 310.300 122.030 317.850 ;
        RECT 122.480 310.300 122.630 317.850 ;
        RECT 122.780 313.200 123.530 315.000 ;
        RECT 122.780 310.450 124.730 313.200 ;
        RECT 122.780 310.300 123.930 310.450 ;
        RECT 105.530 309.700 123.930 310.300 ;
        RECT 105.530 309.550 106.680 309.700 ;
        RECT 102.780 306.800 106.680 309.550 ;
        RECT 102.780 305.050 103.530 306.800 ;
        RECT 105.930 305.050 106.680 306.800 ;
        RECT 106.830 302.150 106.980 309.700 ;
        RECT 107.430 302.150 107.580 309.700 ;
        RECT 108.030 302.150 108.180 309.700 ;
        RECT 108.630 302.150 108.780 309.700 ;
        RECT 109.230 302.150 109.380 309.700 ;
        RECT 109.830 302.150 109.980 309.700 ;
        RECT 114.230 309.200 115.230 309.700 ;
        RECT 110.880 309.050 118.580 309.200 ;
        RECT 114.230 308.600 115.230 309.050 ;
        RECT 110.880 308.450 118.580 308.600 ;
        RECT 114.230 308.000 115.230 308.450 ;
        RECT 110.880 307.850 118.580 308.000 ;
        RECT 114.230 307.400 115.230 307.850 ;
        RECT 110.880 307.250 118.580 307.400 ;
        RECT 114.230 306.800 115.230 307.250 ;
        RECT 110.880 306.650 118.580 306.800 ;
        RECT 114.230 306.200 115.230 306.650 ;
        RECT 110.880 306.050 118.580 306.200 ;
        RECT 114.230 305.600 115.230 306.050 ;
        RECT 110.880 305.450 118.580 305.600 ;
        RECT 114.230 305.000 115.230 305.450 ;
        RECT 110.880 304.850 118.580 305.000 ;
        RECT 114.230 304.400 115.230 304.850 ;
        RECT 110.880 304.250 118.580 304.400 ;
        RECT 114.230 303.800 115.230 304.250 ;
        RECT 110.880 303.650 118.580 303.800 ;
        RECT 114.230 303.200 115.230 303.650 ;
        RECT 110.880 303.050 118.580 303.200 ;
        RECT 114.230 302.600 115.230 303.050 ;
        RECT 110.880 302.450 118.580 302.600 ;
        RECT 114.230 302.000 115.230 302.450 ;
        RECT 119.480 302.150 119.630 309.700 ;
        RECT 120.080 302.150 120.230 309.700 ;
        RECT 120.680 302.150 120.830 309.700 ;
        RECT 121.280 302.150 121.430 309.700 ;
        RECT 121.880 302.150 122.030 309.700 ;
        RECT 122.480 302.150 122.630 309.700 ;
        RECT 122.780 309.550 123.930 309.700 ;
        RECT 124.580 310.415 124.730 310.450 ;
        RECT 124.580 309.550 131.850 310.415 ;
        RECT 122.780 309.140 131.850 309.550 ;
        RECT 122.780 306.800 124.730 309.140 ;
        RECT 122.780 305.050 123.530 306.800 ;
        RECT 10.880 301.850 18.580 302.000 ;
        RECT 30.880 301.850 38.580 302.000 ;
        RECT 50.880 301.850 58.580 302.000 ;
        RECT 70.880 301.850 78.580 302.000 ;
        RECT 90.880 301.850 98.580 302.000 ;
        RECT 110.880 301.850 118.580 302.000 ;
        RECT 14.230 301.200 15.230 301.850 ;
        RECT 34.230 301.200 35.230 301.850 ;
        RECT 54.230 301.200 55.230 301.850 ;
        RECT 74.230 301.200 75.230 301.850 ;
        RECT 94.230 301.200 95.230 301.850 ;
        RECT 114.230 301.200 115.230 301.850 ;
        RECT 11.530 298.800 17.930 301.200 ;
        RECT 31.530 298.800 37.930 301.200 ;
        RECT 51.530 298.800 57.930 301.200 ;
        RECT 71.530 298.800 77.930 301.200 ;
        RECT 91.530 298.800 97.930 301.200 ;
        RECT 111.530 298.800 117.930 301.200 ;
        RECT 14.230 298.150 15.230 298.800 ;
        RECT 34.230 298.150 35.230 298.800 ;
        RECT 54.230 298.150 55.230 298.800 ;
        RECT 74.230 298.150 75.230 298.800 ;
        RECT 94.230 298.150 95.230 298.800 ;
        RECT 114.230 298.150 115.230 298.800 ;
        RECT 10.880 298.000 18.580 298.150 ;
        RECT 30.880 298.000 38.580 298.150 ;
        RECT 50.880 298.000 58.580 298.150 ;
        RECT 70.880 298.000 78.580 298.150 ;
        RECT 90.880 298.000 98.580 298.150 ;
        RECT 110.880 298.000 118.580 298.150 ;
        RECT 5.930 293.200 6.680 295.000 ;
        RECT 4.730 290.450 6.680 293.200 ;
        RECT 4.730 289.550 4.880 290.450 ;
        RECT 5.530 290.300 6.680 290.450 ;
        RECT 6.830 290.300 6.980 297.850 ;
        RECT 7.430 290.300 7.580 297.850 ;
        RECT 8.030 290.300 8.180 297.850 ;
        RECT 8.630 290.300 8.780 297.850 ;
        RECT 9.230 290.300 9.380 297.850 ;
        RECT 9.830 290.300 9.980 297.850 ;
        RECT 14.230 297.550 15.230 298.000 ;
        RECT 10.880 297.400 18.580 297.550 ;
        RECT 14.230 296.950 15.230 297.400 ;
        RECT 10.880 296.800 18.580 296.950 ;
        RECT 14.230 296.350 15.230 296.800 ;
        RECT 10.880 296.200 18.580 296.350 ;
        RECT 14.230 295.750 15.230 296.200 ;
        RECT 10.880 295.600 18.580 295.750 ;
        RECT 14.230 295.150 15.230 295.600 ;
        RECT 10.880 295.000 18.580 295.150 ;
        RECT 14.230 294.550 15.230 295.000 ;
        RECT 10.880 294.400 18.580 294.550 ;
        RECT 14.230 293.950 15.230 294.400 ;
        RECT 10.880 293.800 18.580 293.950 ;
        RECT 14.230 293.350 15.230 293.800 ;
        RECT 10.880 293.200 18.580 293.350 ;
        RECT 14.230 292.750 15.230 293.200 ;
        RECT 10.880 292.600 18.580 292.750 ;
        RECT 14.230 292.150 15.230 292.600 ;
        RECT 10.880 292.000 18.580 292.150 ;
        RECT 14.230 291.550 15.230 292.000 ;
        RECT 10.880 291.400 18.580 291.550 ;
        RECT 14.230 290.950 15.230 291.400 ;
        RECT 10.880 290.800 18.580 290.950 ;
        RECT 14.230 290.300 15.230 290.800 ;
        RECT 19.480 290.300 19.630 297.850 ;
        RECT 20.080 290.300 20.230 297.850 ;
        RECT 20.680 290.300 20.830 297.850 ;
        RECT 21.280 290.300 21.430 297.850 ;
        RECT 21.880 290.300 22.030 297.850 ;
        RECT 22.480 290.300 22.630 297.850 ;
        RECT 22.780 293.200 23.530 295.000 ;
        RECT 25.930 293.200 26.680 295.000 ;
        RECT 22.780 290.450 26.680 293.200 ;
        RECT 22.780 290.300 23.930 290.450 ;
        RECT 5.530 289.700 23.930 290.300 ;
        RECT 5.530 289.550 6.680 289.700 ;
        RECT 4.730 286.800 6.680 289.550 ;
        RECT 5.930 285.050 6.680 286.800 ;
        RECT 6.830 282.150 6.980 289.700 ;
        RECT 7.430 282.150 7.580 289.700 ;
        RECT 8.030 282.150 8.180 289.700 ;
        RECT 8.630 282.150 8.780 289.700 ;
        RECT 9.230 282.150 9.380 289.700 ;
        RECT 9.830 282.150 9.980 289.700 ;
        RECT 14.230 289.200 15.230 289.700 ;
        RECT 10.880 289.050 18.580 289.200 ;
        RECT 14.230 288.600 15.230 289.050 ;
        RECT 10.880 288.450 18.580 288.600 ;
        RECT 14.230 288.000 15.230 288.450 ;
        RECT 10.880 287.850 18.580 288.000 ;
        RECT 14.230 287.400 15.230 287.850 ;
        RECT 10.880 287.250 18.580 287.400 ;
        RECT 14.230 286.800 15.230 287.250 ;
        RECT 10.880 286.650 18.580 286.800 ;
        RECT 14.230 286.200 15.230 286.650 ;
        RECT 10.880 286.050 18.580 286.200 ;
        RECT 14.230 285.600 15.230 286.050 ;
        RECT 10.880 285.450 18.580 285.600 ;
        RECT 14.230 285.000 15.230 285.450 ;
        RECT 10.880 284.850 18.580 285.000 ;
        RECT 14.230 284.400 15.230 284.850 ;
        RECT 10.880 284.250 18.580 284.400 ;
        RECT 14.230 283.800 15.230 284.250 ;
        RECT 10.880 283.650 18.580 283.800 ;
        RECT 14.230 283.200 15.230 283.650 ;
        RECT 10.880 283.050 18.580 283.200 ;
        RECT 14.230 282.600 15.230 283.050 ;
        RECT 10.880 282.450 18.580 282.600 ;
        RECT 14.230 282.000 15.230 282.450 ;
        RECT 19.480 282.150 19.630 289.700 ;
        RECT 20.080 282.150 20.230 289.700 ;
        RECT 20.680 282.150 20.830 289.700 ;
        RECT 21.280 282.150 21.430 289.700 ;
        RECT 21.880 282.150 22.030 289.700 ;
        RECT 22.480 282.150 22.630 289.700 ;
        RECT 22.780 289.550 23.930 289.700 ;
        RECT 24.580 289.550 24.880 290.450 ;
        RECT 25.530 290.300 26.680 290.450 ;
        RECT 26.830 290.300 26.980 297.850 ;
        RECT 27.430 290.300 27.580 297.850 ;
        RECT 28.030 290.300 28.180 297.850 ;
        RECT 28.630 290.300 28.780 297.850 ;
        RECT 29.230 290.300 29.380 297.850 ;
        RECT 29.830 290.300 29.980 297.850 ;
        RECT 34.230 297.550 35.230 298.000 ;
        RECT 30.880 297.400 38.580 297.550 ;
        RECT 34.230 296.950 35.230 297.400 ;
        RECT 30.880 296.800 38.580 296.950 ;
        RECT 34.230 296.350 35.230 296.800 ;
        RECT 30.880 296.200 38.580 296.350 ;
        RECT 34.230 295.750 35.230 296.200 ;
        RECT 30.880 295.600 38.580 295.750 ;
        RECT 34.230 295.150 35.230 295.600 ;
        RECT 30.880 295.000 38.580 295.150 ;
        RECT 34.230 294.550 35.230 295.000 ;
        RECT 30.880 294.400 38.580 294.550 ;
        RECT 34.230 293.950 35.230 294.400 ;
        RECT 30.880 293.800 38.580 293.950 ;
        RECT 34.230 293.350 35.230 293.800 ;
        RECT 30.880 293.200 38.580 293.350 ;
        RECT 34.230 292.750 35.230 293.200 ;
        RECT 30.880 292.600 38.580 292.750 ;
        RECT 34.230 292.150 35.230 292.600 ;
        RECT 30.880 292.000 38.580 292.150 ;
        RECT 34.230 291.550 35.230 292.000 ;
        RECT 30.880 291.400 38.580 291.550 ;
        RECT 34.230 290.950 35.230 291.400 ;
        RECT 30.880 290.800 38.580 290.950 ;
        RECT 34.230 290.300 35.230 290.800 ;
        RECT 39.480 290.300 39.630 297.850 ;
        RECT 40.080 290.300 40.230 297.850 ;
        RECT 40.680 290.300 40.830 297.850 ;
        RECT 41.280 290.300 41.430 297.850 ;
        RECT 41.880 290.300 42.030 297.850 ;
        RECT 42.480 290.300 42.630 297.850 ;
        RECT 42.780 293.200 43.530 295.000 ;
        RECT 45.930 293.200 46.680 295.000 ;
        RECT 42.780 290.450 46.680 293.200 ;
        RECT 42.780 290.300 43.930 290.450 ;
        RECT 25.530 289.700 43.930 290.300 ;
        RECT 25.530 289.550 26.680 289.700 ;
        RECT 22.780 286.800 26.680 289.550 ;
        RECT 22.780 285.050 23.530 286.800 ;
        RECT 25.930 285.050 26.680 286.800 ;
        RECT 26.830 282.150 26.980 289.700 ;
        RECT 27.430 282.150 27.580 289.700 ;
        RECT 28.030 282.150 28.180 289.700 ;
        RECT 28.630 282.150 28.780 289.700 ;
        RECT 29.230 282.150 29.380 289.700 ;
        RECT 29.830 282.150 29.980 289.700 ;
        RECT 34.230 289.200 35.230 289.700 ;
        RECT 30.880 289.050 38.580 289.200 ;
        RECT 34.230 288.600 35.230 289.050 ;
        RECT 30.880 288.450 38.580 288.600 ;
        RECT 34.230 288.000 35.230 288.450 ;
        RECT 30.880 287.850 38.580 288.000 ;
        RECT 34.230 287.400 35.230 287.850 ;
        RECT 30.880 287.250 38.580 287.400 ;
        RECT 34.230 286.800 35.230 287.250 ;
        RECT 30.880 286.650 38.580 286.800 ;
        RECT 34.230 286.200 35.230 286.650 ;
        RECT 30.880 286.050 38.580 286.200 ;
        RECT 34.230 285.600 35.230 286.050 ;
        RECT 30.880 285.450 38.580 285.600 ;
        RECT 34.230 285.000 35.230 285.450 ;
        RECT 30.880 284.850 38.580 285.000 ;
        RECT 34.230 284.400 35.230 284.850 ;
        RECT 30.880 284.250 38.580 284.400 ;
        RECT 34.230 283.800 35.230 284.250 ;
        RECT 30.880 283.650 38.580 283.800 ;
        RECT 34.230 283.200 35.230 283.650 ;
        RECT 30.880 283.050 38.580 283.200 ;
        RECT 34.230 282.600 35.230 283.050 ;
        RECT 30.880 282.450 38.580 282.600 ;
        RECT 34.230 282.000 35.230 282.450 ;
        RECT 39.480 282.150 39.630 289.700 ;
        RECT 40.080 282.150 40.230 289.700 ;
        RECT 40.680 282.150 40.830 289.700 ;
        RECT 41.280 282.150 41.430 289.700 ;
        RECT 41.880 282.150 42.030 289.700 ;
        RECT 42.480 282.150 42.630 289.700 ;
        RECT 42.780 289.550 43.930 289.700 ;
        RECT 44.580 289.550 44.880 290.450 ;
        RECT 45.530 290.300 46.680 290.450 ;
        RECT 46.830 290.300 46.980 297.850 ;
        RECT 47.430 290.300 47.580 297.850 ;
        RECT 48.030 290.300 48.180 297.850 ;
        RECT 48.630 290.300 48.780 297.850 ;
        RECT 49.230 290.300 49.380 297.850 ;
        RECT 49.830 290.300 49.980 297.850 ;
        RECT 54.230 297.550 55.230 298.000 ;
        RECT 50.880 297.400 58.580 297.550 ;
        RECT 54.230 296.950 55.230 297.400 ;
        RECT 50.880 296.800 58.580 296.950 ;
        RECT 54.230 296.350 55.230 296.800 ;
        RECT 50.880 296.200 58.580 296.350 ;
        RECT 54.230 295.750 55.230 296.200 ;
        RECT 50.880 295.600 58.580 295.750 ;
        RECT 54.230 295.150 55.230 295.600 ;
        RECT 50.880 295.000 58.580 295.150 ;
        RECT 54.230 294.550 55.230 295.000 ;
        RECT 50.880 294.400 58.580 294.550 ;
        RECT 54.230 293.950 55.230 294.400 ;
        RECT 50.880 293.800 58.580 293.950 ;
        RECT 54.230 293.350 55.230 293.800 ;
        RECT 50.880 293.200 58.580 293.350 ;
        RECT 54.230 292.750 55.230 293.200 ;
        RECT 50.880 292.600 58.580 292.750 ;
        RECT 54.230 292.150 55.230 292.600 ;
        RECT 50.880 292.000 58.580 292.150 ;
        RECT 54.230 291.550 55.230 292.000 ;
        RECT 50.880 291.400 58.580 291.550 ;
        RECT 54.230 290.950 55.230 291.400 ;
        RECT 50.880 290.800 58.580 290.950 ;
        RECT 54.230 290.300 55.230 290.800 ;
        RECT 59.480 290.300 59.630 297.850 ;
        RECT 60.080 290.300 60.230 297.850 ;
        RECT 60.680 290.300 60.830 297.850 ;
        RECT 61.280 290.300 61.430 297.850 ;
        RECT 61.880 290.300 62.030 297.850 ;
        RECT 62.480 290.300 62.630 297.850 ;
        RECT 62.780 293.200 63.530 295.000 ;
        RECT 65.930 293.200 66.680 295.000 ;
        RECT 62.780 290.450 66.680 293.200 ;
        RECT 62.780 290.300 63.930 290.450 ;
        RECT 45.530 289.700 63.930 290.300 ;
        RECT 45.530 289.550 46.680 289.700 ;
        RECT 42.780 286.800 46.680 289.550 ;
        RECT 42.780 285.050 43.530 286.800 ;
        RECT 45.930 285.050 46.680 286.800 ;
        RECT 46.830 282.150 46.980 289.700 ;
        RECT 47.430 282.150 47.580 289.700 ;
        RECT 48.030 282.150 48.180 289.700 ;
        RECT 48.630 282.150 48.780 289.700 ;
        RECT 49.230 282.150 49.380 289.700 ;
        RECT 49.830 282.150 49.980 289.700 ;
        RECT 54.230 289.200 55.230 289.700 ;
        RECT 50.880 289.050 58.580 289.200 ;
        RECT 54.230 288.600 55.230 289.050 ;
        RECT 50.880 288.450 58.580 288.600 ;
        RECT 54.230 288.000 55.230 288.450 ;
        RECT 50.880 287.850 58.580 288.000 ;
        RECT 54.230 287.400 55.230 287.850 ;
        RECT 50.880 287.250 58.580 287.400 ;
        RECT 54.230 286.800 55.230 287.250 ;
        RECT 50.880 286.650 58.580 286.800 ;
        RECT 54.230 286.200 55.230 286.650 ;
        RECT 50.880 286.050 58.580 286.200 ;
        RECT 54.230 285.600 55.230 286.050 ;
        RECT 50.880 285.450 58.580 285.600 ;
        RECT 54.230 285.000 55.230 285.450 ;
        RECT 50.880 284.850 58.580 285.000 ;
        RECT 54.230 284.400 55.230 284.850 ;
        RECT 50.880 284.250 58.580 284.400 ;
        RECT 54.230 283.800 55.230 284.250 ;
        RECT 50.880 283.650 58.580 283.800 ;
        RECT 54.230 283.200 55.230 283.650 ;
        RECT 50.880 283.050 58.580 283.200 ;
        RECT 54.230 282.600 55.230 283.050 ;
        RECT 50.880 282.450 58.580 282.600 ;
        RECT 54.230 282.000 55.230 282.450 ;
        RECT 59.480 282.150 59.630 289.700 ;
        RECT 60.080 282.150 60.230 289.700 ;
        RECT 60.680 282.150 60.830 289.700 ;
        RECT 61.280 282.150 61.430 289.700 ;
        RECT 61.880 282.150 62.030 289.700 ;
        RECT 62.480 282.150 62.630 289.700 ;
        RECT 62.780 289.550 63.930 289.700 ;
        RECT 64.580 289.550 64.880 290.450 ;
        RECT 65.530 290.300 66.680 290.450 ;
        RECT 66.830 290.300 66.980 297.850 ;
        RECT 67.430 290.300 67.580 297.850 ;
        RECT 68.030 290.300 68.180 297.850 ;
        RECT 68.630 290.300 68.780 297.850 ;
        RECT 69.230 290.300 69.380 297.850 ;
        RECT 69.830 290.300 69.980 297.850 ;
        RECT 74.230 297.550 75.230 298.000 ;
        RECT 70.880 297.400 78.580 297.550 ;
        RECT 74.230 296.950 75.230 297.400 ;
        RECT 70.880 296.800 78.580 296.950 ;
        RECT 74.230 296.350 75.230 296.800 ;
        RECT 70.880 296.200 78.580 296.350 ;
        RECT 74.230 295.750 75.230 296.200 ;
        RECT 70.880 295.600 78.580 295.750 ;
        RECT 74.230 295.150 75.230 295.600 ;
        RECT 70.880 295.000 78.580 295.150 ;
        RECT 74.230 294.550 75.230 295.000 ;
        RECT 70.880 294.400 78.580 294.550 ;
        RECT 74.230 293.950 75.230 294.400 ;
        RECT 70.880 293.800 78.580 293.950 ;
        RECT 74.230 293.350 75.230 293.800 ;
        RECT 70.880 293.200 78.580 293.350 ;
        RECT 74.230 292.750 75.230 293.200 ;
        RECT 70.880 292.600 78.580 292.750 ;
        RECT 74.230 292.150 75.230 292.600 ;
        RECT 70.880 292.000 78.580 292.150 ;
        RECT 74.230 291.550 75.230 292.000 ;
        RECT 70.880 291.400 78.580 291.550 ;
        RECT 74.230 290.950 75.230 291.400 ;
        RECT 70.880 290.800 78.580 290.950 ;
        RECT 74.230 290.300 75.230 290.800 ;
        RECT 79.480 290.300 79.630 297.850 ;
        RECT 80.080 290.300 80.230 297.850 ;
        RECT 80.680 290.300 80.830 297.850 ;
        RECT 81.280 290.300 81.430 297.850 ;
        RECT 81.880 290.300 82.030 297.850 ;
        RECT 82.480 290.300 82.630 297.850 ;
        RECT 82.780 293.200 83.530 295.000 ;
        RECT 85.930 293.200 86.680 295.000 ;
        RECT 82.780 290.450 86.680 293.200 ;
        RECT 82.780 290.300 83.930 290.450 ;
        RECT 65.530 289.700 83.930 290.300 ;
        RECT 65.530 289.550 66.680 289.700 ;
        RECT 62.780 286.800 66.680 289.550 ;
        RECT 62.780 285.050 63.530 286.800 ;
        RECT 65.930 285.050 66.680 286.800 ;
        RECT 66.830 282.150 66.980 289.700 ;
        RECT 67.430 282.150 67.580 289.700 ;
        RECT 68.030 282.150 68.180 289.700 ;
        RECT 68.630 282.150 68.780 289.700 ;
        RECT 69.230 282.150 69.380 289.700 ;
        RECT 69.830 282.150 69.980 289.700 ;
        RECT 74.230 289.200 75.230 289.700 ;
        RECT 70.880 289.050 78.580 289.200 ;
        RECT 74.230 288.600 75.230 289.050 ;
        RECT 70.880 288.450 78.580 288.600 ;
        RECT 74.230 288.000 75.230 288.450 ;
        RECT 70.880 287.850 78.580 288.000 ;
        RECT 74.230 287.400 75.230 287.850 ;
        RECT 70.880 287.250 78.580 287.400 ;
        RECT 74.230 286.800 75.230 287.250 ;
        RECT 70.880 286.650 78.580 286.800 ;
        RECT 74.230 286.200 75.230 286.650 ;
        RECT 70.880 286.050 78.580 286.200 ;
        RECT 74.230 285.600 75.230 286.050 ;
        RECT 70.880 285.450 78.580 285.600 ;
        RECT 74.230 285.000 75.230 285.450 ;
        RECT 70.880 284.850 78.580 285.000 ;
        RECT 74.230 284.400 75.230 284.850 ;
        RECT 70.880 284.250 78.580 284.400 ;
        RECT 74.230 283.800 75.230 284.250 ;
        RECT 70.880 283.650 78.580 283.800 ;
        RECT 74.230 283.200 75.230 283.650 ;
        RECT 70.880 283.050 78.580 283.200 ;
        RECT 74.230 282.600 75.230 283.050 ;
        RECT 70.880 282.450 78.580 282.600 ;
        RECT 74.230 282.000 75.230 282.450 ;
        RECT 79.480 282.150 79.630 289.700 ;
        RECT 80.080 282.150 80.230 289.700 ;
        RECT 80.680 282.150 80.830 289.700 ;
        RECT 81.280 282.150 81.430 289.700 ;
        RECT 81.880 282.150 82.030 289.700 ;
        RECT 82.480 282.150 82.630 289.700 ;
        RECT 82.780 289.550 83.930 289.700 ;
        RECT 84.580 289.550 84.880 290.450 ;
        RECT 85.530 290.300 86.680 290.450 ;
        RECT 86.830 290.300 86.980 297.850 ;
        RECT 87.430 290.300 87.580 297.850 ;
        RECT 88.030 290.300 88.180 297.850 ;
        RECT 88.630 290.300 88.780 297.850 ;
        RECT 89.230 290.300 89.380 297.850 ;
        RECT 89.830 290.300 89.980 297.850 ;
        RECT 94.230 297.550 95.230 298.000 ;
        RECT 90.880 297.400 98.580 297.550 ;
        RECT 94.230 296.950 95.230 297.400 ;
        RECT 90.880 296.800 98.580 296.950 ;
        RECT 94.230 296.350 95.230 296.800 ;
        RECT 90.880 296.200 98.580 296.350 ;
        RECT 94.230 295.750 95.230 296.200 ;
        RECT 90.880 295.600 98.580 295.750 ;
        RECT 94.230 295.150 95.230 295.600 ;
        RECT 90.880 295.000 98.580 295.150 ;
        RECT 94.230 294.550 95.230 295.000 ;
        RECT 90.880 294.400 98.580 294.550 ;
        RECT 94.230 293.950 95.230 294.400 ;
        RECT 90.880 293.800 98.580 293.950 ;
        RECT 94.230 293.350 95.230 293.800 ;
        RECT 90.880 293.200 98.580 293.350 ;
        RECT 94.230 292.750 95.230 293.200 ;
        RECT 90.880 292.600 98.580 292.750 ;
        RECT 94.230 292.150 95.230 292.600 ;
        RECT 90.880 292.000 98.580 292.150 ;
        RECT 94.230 291.550 95.230 292.000 ;
        RECT 90.880 291.400 98.580 291.550 ;
        RECT 94.230 290.950 95.230 291.400 ;
        RECT 90.880 290.800 98.580 290.950 ;
        RECT 94.230 290.300 95.230 290.800 ;
        RECT 99.480 290.300 99.630 297.850 ;
        RECT 100.080 290.300 100.230 297.850 ;
        RECT 100.680 290.300 100.830 297.850 ;
        RECT 101.280 290.300 101.430 297.850 ;
        RECT 101.880 290.300 102.030 297.850 ;
        RECT 102.480 290.300 102.630 297.850 ;
        RECT 102.780 293.200 103.530 295.000 ;
        RECT 105.930 293.200 106.680 295.000 ;
        RECT 102.780 290.450 106.680 293.200 ;
        RECT 102.780 290.300 103.930 290.450 ;
        RECT 85.530 289.700 103.930 290.300 ;
        RECT 85.530 289.550 86.680 289.700 ;
        RECT 82.780 286.800 86.680 289.550 ;
        RECT 82.780 285.050 83.530 286.800 ;
        RECT 85.930 285.050 86.680 286.800 ;
        RECT 86.830 282.150 86.980 289.700 ;
        RECT 87.430 282.150 87.580 289.700 ;
        RECT 88.030 282.150 88.180 289.700 ;
        RECT 88.630 282.150 88.780 289.700 ;
        RECT 89.230 282.150 89.380 289.700 ;
        RECT 89.830 282.150 89.980 289.700 ;
        RECT 94.230 289.200 95.230 289.700 ;
        RECT 90.880 289.050 98.580 289.200 ;
        RECT 94.230 288.600 95.230 289.050 ;
        RECT 90.880 288.450 98.580 288.600 ;
        RECT 94.230 288.000 95.230 288.450 ;
        RECT 90.880 287.850 98.580 288.000 ;
        RECT 94.230 287.400 95.230 287.850 ;
        RECT 90.880 287.250 98.580 287.400 ;
        RECT 94.230 286.800 95.230 287.250 ;
        RECT 90.880 286.650 98.580 286.800 ;
        RECT 94.230 286.200 95.230 286.650 ;
        RECT 90.880 286.050 98.580 286.200 ;
        RECT 94.230 285.600 95.230 286.050 ;
        RECT 90.880 285.450 98.580 285.600 ;
        RECT 94.230 285.000 95.230 285.450 ;
        RECT 90.880 284.850 98.580 285.000 ;
        RECT 94.230 284.400 95.230 284.850 ;
        RECT 90.880 284.250 98.580 284.400 ;
        RECT 94.230 283.800 95.230 284.250 ;
        RECT 90.880 283.650 98.580 283.800 ;
        RECT 94.230 283.200 95.230 283.650 ;
        RECT 90.880 283.050 98.580 283.200 ;
        RECT 94.230 282.600 95.230 283.050 ;
        RECT 90.880 282.450 98.580 282.600 ;
        RECT 94.230 282.000 95.230 282.450 ;
        RECT 99.480 282.150 99.630 289.700 ;
        RECT 100.080 282.150 100.230 289.700 ;
        RECT 100.680 282.150 100.830 289.700 ;
        RECT 101.280 282.150 101.430 289.700 ;
        RECT 101.880 282.150 102.030 289.700 ;
        RECT 102.480 282.150 102.630 289.700 ;
        RECT 102.780 289.550 103.930 289.700 ;
        RECT 104.580 289.550 104.880 290.450 ;
        RECT 105.530 290.300 106.680 290.450 ;
        RECT 106.830 290.300 106.980 297.850 ;
        RECT 107.430 290.300 107.580 297.850 ;
        RECT 108.030 290.300 108.180 297.850 ;
        RECT 108.630 290.300 108.780 297.850 ;
        RECT 109.230 290.300 109.380 297.850 ;
        RECT 109.830 290.300 109.980 297.850 ;
        RECT 114.230 297.550 115.230 298.000 ;
        RECT 110.880 297.400 118.580 297.550 ;
        RECT 114.230 296.950 115.230 297.400 ;
        RECT 110.880 296.800 118.580 296.950 ;
        RECT 114.230 296.350 115.230 296.800 ;
        RECT 110.880 296.200 118.580 296.350 ;
        RECT 114.230 295.750 115.230 296.200 ;
        RECT 110.880 295.600 118.580 295.750 ;
        RECT 114.230 295.150 115.230 295.600 ;
        RECT 110.880 295.000 118.580 295.150 ;
        RECT 114.230 294.550 115.230 295.000 ;
        RECT 110.880 294.400 118.580 294.550 ;
        RECT 114.230 293.950 115.230 294.400 ;
        RECT 110.880 293.800 118.580 293.950 ;
        RECT 114.230 293.350 115.230 293.800 ;
        RECT 110.880 293.200 118.580 293.350 ;
        RECT 114.230 292.750 115.230 293.200 ;
        RECT 110.880 292.600 118.580 292.750 ;
        RECT 114.230 292.150 115.230 292.600 ;
        RECT 110.880 292.000 118.580 292.150 ;
        RECT 114.230 291.550 115.230 292.000 ;
        RECT 110.880 291.400 118.580 291.550 ;
        RECT 114.230 290.950 115.230 291.400 ;
        RECT 110.880 290.800 118.580 290.950 ;
        RECT 114.230 290.300 115.230 290.800 ;
        RECT 119.480 290.300 119.630 297.850 ;
        RECT 120.080 290.300 120.230 297.850 ;
        RECT 120.680 290.300 120.830 297.850 ;
        RECT 121.280 290.300 121.430 297.850 ;
        RECT 121.880 290.300 122.030 297.850 ;
        RECT 122.480 290.300 122.630 297.850 ;
        RECT 122.780 293.200 123.530 295.000 ;
        RECT 122.780 290.450 124.730 293.200 ;
        RECT 122.780 290.300 123.930 290.450 ;
        RECT 105.530 289.700 123.930 290.300 ;
        RECT 105.530 289.550 106.680 289.700 ;
        RECT 102.780 286.800 106.680 289.550 ;
        RECT 102.780 285.050 103.530 286.800 ;
        RECT 105.930 285.050 106.680 286.800 ;
        RECT 106.830 282.150 106.980 289.700 ;
        RECT 107.430 282.150 107.580 289.700 ;
        RECT 108.030 282.150 108.180 289.700 ;
        RECT 108.630 282.150 108.780 289.700 ;
        RECT 109.230 282.150 109.380 289.700 ;
        RECT 109.830 282.150 109.980 289.700 ;
        RECT 114.230 289.200 115.230 289.700 ;
        RECT 110.880 289.050 118.580 289.200 ;
        RECT 114.230 288.600 115.230 289.050 ;
        RECT 110.880 288.450 118.580 288.600 ;
        RECT 114.230 288.000 115.230 288.450 ;
        RECT 110.880 287.850 118.580 288.000 ;
        RECT 114.230 287.400 115.230 287.850 ;
        RECT 110.880 287.250 118.580 287.400 ;
        RECT 114.230 286.800 115.230 287.250 ;
        RECT 110.880 286.650 118.580 286.800 ;
        RECT 114.230 286.200 115.230 286.650 ;
        RECT 110.880 286.050 118.580 286.200 ;
        RECT 114.230 285.600 115.230 286.050 ;
        RECT 110.880 285.450 118.580 285.600 ;
        RECT 114.230 285.000 115.230 285.450 ;
        RECT 110.880 284.850 118.580 285.000 ;
        RECT 114.230 284.400 115.230 284.850 ;
        RECT 110.880 284.250 118.580 284.400 ;
        RECT 114.230 283.800 115.230 284.250 ;
        RECT 110.880 283.650 118.580 283.800 ;
        RECT 114.230 283.200 115.230 283.650 ;
        RECT 110.880 283.050 118.580 283.200 ;
        RECT 114.230 282.600 115.230 283.050 ;
        RECT 110.880 282.450 118.580 282.600 ;
        RECT 114.230 282.000 115.230 282.450 ;
        RECT 119.480 282.150 119.630 289.700 ;
        RECT 120.080 282.150 120.230 289.700 ;
        RECT 120.680 282.150 120.830 289.700 ;
        RECT 121.280 282.150 121.430 289.700 ;
        RECT 121.880 282.150 122.030 289.700 ;
        RECT 122.480 282.150 122.630 289.700 ;
        RECT 122.780 289.550 123.930 289.700 ;
        RECT 124.580 290.410 124.730 290.450 ;
        RECT 124.580 289.550 131.850 290.410 ;
        RECT 122.780 289.135 131.850 289.550 ;
        RECT 122.780 286.800 124.730 289.135 ;
        RECT 122.780 285.050 123.530 286.800 ;
        RECT 10.880 281.850 18.580 282.000 ;
        RECT 30.880 281.850 38.580 282.000 ;
        RECT 50.880 281.850 58.580 282.000 ;
        RECT 70.880 281.850 78.580 282.000 ;
        RECT 90.880 281.850 98.580 282.000 ;
        RECT 110.880 281.850 118.580 282.000 ;
        RECT 14.230 281.200 15.230 281.850 ;
        RECT 34.230 281.200 35.230 281.850 ;
        RECT 54.230 281.200 55.230 281.850 ;
        RECT 74.230 281.200 75.230 281.850 ;
        RECT 94.230 281.200 95.230 281.850 ;
        RECT 114.230 281.200 115.230 281.850 ;
        RECT 11.530 278.800 17.930 281.200 ;
        RECT 31.530 278.800 37.930 281.200 ;
        RECT 51.530 278.800 57.930 281.200 ;
        RECT 71.530 278.800 77.930 281.200 ;
        RECT 91.530 278.800 97.930 281.200 ;
        RECT 111.530 278.800 117.930 281.200 ;
        RECT 14.230 278.150 15.230 278.800 ;
        RECT 34.230 278.150 35.230 278.800 ;
        RECT 54.230 278.150 55.230 278.800 ;
        RECT 74.230 278.150 75.230 278.800 ;
        RECT 94.230 278.150 95.230 278.800 ;
        RECT 114.230 278.150 115.230 278.800 ;
        RECT 10.880 278.000 18.580 278.150 ;
        RECT 30.880 278.000 38.580 278.150 ;
        RECT 50.880 278.000 58.580 278.150 ;
        RECT 70.880 278.000 78.580 278.150 ;
        RECT 90.880 278.000 98.580 278.150 ;
        RECT 110.880 278.000 118.580 278.150 ;
        RECT 5.930 273.200 6.680 275.000 ;
        RECT 4.730 270.450 6.680 273.200 ;
        RECT 4.730 269.550 4.880 270.450 ;
        RECT 5.530 270.300 6.680 270.450 ;
        RECT 6.830 270.300 6.980 277.850 ;
        RECT 7.430 270.300 7.580 277.850 ;
        RECT 8.030 270.300 8.180 277.850 ;
        RECT 8.630 270.300 8.780 277.850 ;
        RECT 9.230 270.300 9.380 277.850 ;
        RECT 9.830 270.300 9.980 277.850 ;
        RECT 14.230 277.550 15.230 278.000 ;
        RECT 10.880 277.400 18.580 277.550 ;
        RECT 14.230 276.950 15.230 277.400 ;
        RECT 10.880 276.800 18.580 276.950 ;
        RECT 14.230 276.350 15.230 276.800 ;
        RECT 10.880 276.200 18.580 276.350 ;
        RECT 14.230 275.750 15.230 276.200 ;
        RECT 10.880 275.600 18.580 275.750 ;
        RECT 14.230 275.150 15.230 275.600 ;
        RECT 10.880 275.000 18.580 275.150 ;
        RECT 14.230 274.550 15.230 275.000 ;
        RECT 10.880 274.400 18.580 274.550 ;
        RECT 14.230 273.950 15.230 274.400 ;
        RECT 10.880 273.800 18.580 273.950 ;
        RECT 14.230 273.350 15.230 273.800 ;
        RECT 10.880 273.200 18.580 273.350 ;
        RECT 14.230 272.750 15.230 273.200 ;
        RECT 10.880 272.600 18.580 272.750 ;
        RECT 14.230 272.150 15.230 272.600 ;
        RECT 10.880 272.000 18.580 272.150 ;
        RECT 14.230 271.550 15.230 272.000 ;
        RECT 10.880 271.400 18.580 271.550 ;
        RECT 14.230 270.950 15.230 271.400 ;
        RECT 10.880 270.800 18.580 270.950 ;
        RECT 14.230 270.300 15.230 270.800 ;
        RECT 19.480 270.300 19.630 277.850 ;
        RECT 20.080 270.300 20.230 277.850 ;
        RECT 20.680 270.300 20.830 277.850 ;
        RECT 21.280 270.300 21.430 277.850 ;
        RECT 21.880 270.300 22.030 277.850 ;
        RECT 22.480 270.300 22.630 277.850 ;
        RECT 22.780 273.200 23.530 275.000 ;
        RECT 25.930 273.200 26.680 275.000 ;
        RECT 22.780 270.450 26.680 273.200 ;
        RECT 22.780 270.300 23.930 270.450 ;
        RECT 5.530 269.700 23.930 270.300 ;
        RECT 5.530 269.550 6.680 269.700 ;
        RECT 4.730 266.800 6.680 269.550 ;
        RECT 5.930 265.050 6.680 266.800 ;
        RECT 6.830 262.150 6.980 269.700 ;
        RECT 7.430 262.150 7.580 269.700 ;
        RECT 8.030 262.150 8.180 269.700 ;
        RECT 8.630 262.150 8.780 269.700 ;
        RECT 9.230 262.150 9.380 269.700 ;
        RECT 9.830 262.150 9.980 269.700 ;
        RECT 14.230 269.200 15.230 269.700 ;
        RECT 10.880 269.050 18.580 269.200 ;
        RECT 14.230 268.600 15.230 269.050 ;
        RECT 10.880 268.450 18.580 268.600 ;
        RECT 14.230 268.000 15.230 268.450 ;
        RECT 10.880 267.850 18.580 268.000 ;
        RECT 14.230 267.400 15.230 267.850 ;
        RECT 10.880 267.250 18.580 267.400 ;
        RECT 14.230 266.800 15.230 267.250 ;
        RECT 10.880 266.650 18.580 266.800 ;
        RECT 14.230 266.200 15.230 266.650 ;
        RECT 10.880 266.050 18.580 266.200 ;
        RECT 14.230 265.600 15.230 266.050 ;
        RECT 10.880 265.450 18.580 265.600 ;
        RECT 14.230 265.000 15.230 265.450 ;
        RECT 10.880 264.850 18.580 265.000 ;
        RECT 14.230 264.400 15.230 264.850 ;
        RECT 10.880 264.250 18.580 264.400 ;
        RECT 14.230 263.800 15.230 264.250 ;
        RECT 10.880 263.650 18.580 263.800 ;
        RECT 14.230 263.200 15.230 263.650 ;
        RECT 10.880 263.050 18.580 263.200 ;
        RECT 14.230 262.600 15.230 263.050 ;
        RECT 10.880 262.450 18.580 262.600 ;
        RECT 14.230 262.000 15.230 262.450 ;
        RECT 19.480 262.150 19.630 269.700 ;
        RECT 20.080 262.150 20.230 269.700 ;
        RECT 20.680 262.150 20.830 269.700 ;
        RECT 21.280 262.150 21.430 269.700 ;
        RECT 21.880 262.150 22.030 269.700 ;
        RECT 22.480 262.150 22.630 269.700 ;
        RECT 22.780 269.550 23.930 269.700 ;
        RECT 24.580 269.550 24.880 270.450 ;
        RECT 25.530 270.300 26.680 270.450 ;
        RECT 26.830 270.300 26.980 277.850 ;
        RECT 27.430 270.300 27.580 277.850 ;
        RECT 28.030 270.300 28.180 277.850 ;
        RECT 28.630 270.300 28.780 277.850 ;
        RECT 29.230 270.300 29.380 277.850 ;
        RECT 29.830 270.300 29.980 277.850 ;
        RECT 34.230 277.550 35.230 278.000 ;
        RECT 30.880 277.400 38.580 277.550 ;
        RECT 34.230 276.950 35.230 277.400 ;
        RECT 30.880 276.800 38.580 276.950 ;
        RECT 34.230 276.350 35.230 276.800 ;
        RECT 30.880 276.200 38.580 276.350 ;
        RECT 34.230 275.750 35.230 276.200 ;
        RECT 30.880 275.600 38.580 275.750 ;
        RECT 34.230 275.150 35.230 275.600 ;
        RECT 30.880 275.000 38.580 275.150 ;
        RECT 34.230 274.550 35.230 275.000 ;
        RECT 30.880 274.400 38.580 274.550 ;
        RECT 34.230 273.950 35.230 274.400 ;
        RECT 30.880 273.800 38.580 273.950 ;
        RECT 34.230 273.350 35.230 273.800 ;
        RECT 30.880 273.200 38.580 273.350 ;
        RECT 34.230 272.750 35.230 273.200 ;
        RECT 30.880 272.600 38.580 272.750 ;
        RECT 34.230 272.150 35.230 272.600 ;
        RECT 30.880 272.000 38.580 272.150 ;
        RECT 34.230 271.550 35.230 272.000 ;
        RECT 30.880 271.400 38.580 271.550 ;
        RECT 34.230 270.950 35.230 271.400 ;
        RECT 30.880 270.800 38.580 270.950 ;
        RECT 34.230 270.300 35.230 270.800 ;
        RECT 39.480 270.300 39.630 277.850 ;
        RECT 40.080 270.300 40.230 277.850 ;
        RECT 40.680 270.300 40.830 277.850 ;
        RECT 41.280 270.300 41.430 277.850 ;
        RECT 41.880 270.300 42.030 277.850 ;
        RECT 42.480 270.300 42.630 277.850 ;
        RECT 42.780 273.200 43.530 275.000 ;
        RECT 45.930 273.200 46.680 275.000 ;
        RECT 42.780 270.450 46.680 273.200 ;
        RECT 42.780 270.300 43.930 270.450 ;
        RECT 25.530 269.700 43.930 270.300 ;
        RECT 25.530 269.550 26.680 269.700 ;
        RECT 22.780 266.800 26.680 269.550 ;
        RECT 22.780 265.050 23.530 266.800 ;
        RECT 25.930 265.050 26.680 266.800 ;
        RECT 26.830 262.150 26.980 269.700 ;
        RECT 27.430 262.150 27.580 269.700 ;
        RECT 28.030 262.150 28.180 269.700 ;
        RECT 28.630 262.150 28.780 269.700 ;
        RECT 29.230 262.150 29.380 269.700 ;
        RECT 29.830 262.150 29.980 269.700 ;
        RECT 34.230 269.200 35.230 269.700 ;
        RECT 30.880 269.050 38.580 269.200 ;
        RECT 34.230 268.600 35.230 269.050 ;
        RECT 30.880 268.450 38.580 268.600 ;
        RECT 34.230 268.000 35.230 268.450 ;
        RECT 30.880 267.850 38.580 268.000 ;
        RECT 34.230 267.400 35.230 267.850 ;
        RECT 30.880 267.250 38.580 267.400 ;
        RECT 34.230 266.800 35.230 267.250 ;
        RECT 30.880 266.650 38.580 266.800 ;
        RECT 34.230 266.200 35.230 266.650 ;
        RECT 30.880 266.050 38.580 266.200 ;
        RECT 34.230 265.600 35.230 266.050 ;
        RECT 30.880 265.450 38.580 265.600 ;
        RECT 34.230 265.000 35.230 265.450 ;
        RECT 30.880 264.850 38.580 265.000 ;
        RECT 34.230 264.400 35.230 264.850 ;
        RECT 30.880 264.250 38.580 264.400 ;
        RECT 34.230 263.800 35.230 264.250 ;
        RECT 30.880 263.650 38.580 263.800 ;
        RECT 34.230 263.200 35.230 263.650 ;
        RECT 30.880 263.050 38.580 263.200 ;
        RECT 34.230 262.600 35.230 263.050 ;
        RECT 30.880 262.450 38.580 262.600 ;
        RECT 34.230 262.000 35.230 262.450 ;
        RECT 39.480 262.150 39.630 269.700 ;
        RECT 40.080 262.150 40.230 269.700 ;
        RECT 40.680 262.150 40.830 269.700 ;
        RECT 41.280 262.150 41.430 269.700 ;
        RECT 41.880 262.150 42.030 269.700 ;
        RECT 42.480 262.150 42.630 269.700 ;
        RECT 42.780 269.550 43.930 269.700 ;
        RECT 44.580 269.550 44.880 270.450 ;
        RECT 45.530 270.300 46.680 270.450 ;
        RECT 46.830 270.300 46.980 277.850 ;
        RECT 47.430 270.300 47.580 277.850 ;
        RECT 48.030 270.300 48.180 277.850 ;
        RECT 48.630 270.300 48.780 277.850 ;
        RECT 49.230 270.300 49.380 277.850 ;
        RECT 49.830 270.300 49.980 277.850 ;
        RECT 54.230 277.550 55.230 278.000 ;
        RECT 50.880 277.400 58.580 277.550 ;
        RECT 54.230 276.950 55.230 277.400 ;
        RECT 50.880 276.800 58.580 276.950 ;
        RECT 54.230 276.350 55.230 276.800 ;
        RECT 50.880 276.200 58.580 276.350 ;
        RECT 54.230 275.750 55.230 276.200 ;
        RECT 50.880 275.600 58.580 275.750 ;
        RECT 54.230 275.150 55.230 275.600 ;
        RECT 50.880 275.000 58.580 275.150 ;
        RECT 54.230 274.550 55.230 275.000 ;
        RECT 50.880 274.400 58.580 274.550 ;
        RECT 54.230 273.950 55.230 274.400 ;
        RECT 50.880 273.800 58.580 273.950 ;
        RECT 54.230 273.350 55.230 273.800 ;
        RECT 50.880 273.200 58.580 273.350 ;
        RECT 54.230 272.750 55.230 273.200 ;
        RECT 50.880 272.600 58.580 272.750 ;
        RECT 54.230 272.150 55.230 272.600 ;
        RECT 50.880 272.000 58.580 272.150 ;
        RECT 54.230 271.550 55.230 272.000 ;
        RECT 50.880 271.400 58.580 271.550 ;
        RECT 54.230 270.950 55.230 271.400 ;
        RECT 50.880 270.800 58.580 270.950 ;
        RECT 54.230 270.300 55.230 270.800 ;
        RECT 59.480 270.300 59.630 277.850 ;
        RECT 60.080 270.300 60.230 277.850 ;
        RECT 60.680 270.300 60.830 277.850 ;
        RECT 61.280 270.300 61.430 277.850 ;
        RECT 61.880 270.300 62.030 277.850 ;
        RECT 62.480 270.300 62.630 277.850 ;
        RECT 62.780 273.200 63.530 275.000 ;
        RECT 65.930 273.200 66.680 275.000 ;
        RECT 62.780 270.450 66.680 273.200 ;
        RECT 62.780 270.300 63.930 270.450 ;
        RECT 45.530 269.700 63.930 270.300 ;
        RECT 45.530 269.550 46.680 269.700 ;
        RECT 42.780 266.800 46.680 269.550 ;
        RECT 42.780 265.050 43.530 266.800 ;
        RECT 45.930 265.050 46.680 266.800 ;
        RECT 46.830 262.150 46.980 269.700 ;
        RECT 47.430 262.150 47.580 269.700 ;
        RECT 48.030 262.150 48.180 269.700 ;
        RECT 48.630 262.150 48.780 269.700 ;
        RECT 49.230 262.150 49.380 269.700 ;
        RECT 49.830 262.150 49.980 269.700 ;
        RECT 54.230 269.200 55.230 269.700 ;
        RECT 50.880 269.050 58.580 269.200 ;
        RECT 54.230 268.600 55.230 269.050 ;
        RECT 50.880 268.450 58.580 268.600 ;
        RECT 54.230 268.000 55.230 268.450 ;
        RECT 50.880 267.850 58.580 268.000 ;
        RECT 54.230 267.400 55.230 267.850 ;
        RECT 50.880 267.250 58.580 267.400 ;
        RECT 54.230 266.800 55.230 267.250 ;
        RECT 50.880 266.650 58.580 266.800 ;
        RECT 54.230 266.200 55.230 266.650 ;
        RECT 50.880 266.050 58.580 266.200 ;
        RECT 54.230 265.600 55.230 266.050 ;
        RECT 50.880 265.450 58.580 265.600 ;
        RECT 54.230 265.000 55.230 265.450 ;
        RECT 50.880 264.850 58.580 265.000 ;
        RECT 54.230 264.400 55.230 264.850 ;
        RECT 50.880 264.250 58.580 264.400 ;
        RECT 54.230 263.800 55.230 264.250 ;
        RECT 50.880 263.650 58.580 263.800 ;
        RECT 54.230 263.200 55.230 263.650 ;
        RECT 50.880 263.050 58.580 263.200 ;
        RECT 54.230 262.600 55.230 263.050 ;
        RECT 50.880 262.450 58.580 262.600 ;
        RECT 54.230 262.000 55.230 262.450 ;
        RECT 59.480 262.150 59.630 269.700 ;
        RECT 60.080 262.150 60.230 269.700 ;
        RECT 60.680 262.150 60.830 269.700 ;
        RECT 61.280 262.150 61.430 269.700 ;
        RECT 61.880 262.150 62.030 269.700 ;
        RECT 62.480 262.150 62.630 269.700 ;
        RECT 62.780 269.550 63.930 269.700 ;
        RECT 64.580 269.550 64.880 270.450 ;
        RECT 65.530 270.300 66.680 270.450 ;
        RECT 66.830 270.300 66.980 277.850 ;
        RECT 67.430 270.300 67.580 277.850 ;
        RECT 68.030 270.300 68.180 277.850 ;
        RECT 68.630 270.300 68.780 277.850 ;
        RECT 69.230 270.300 69.380 277.850 ;
        RECT 69.830 270.300 69.980 277.850 ;
        RECT 74.230 277.550 75.230 278.000 ;
        RECT 70.880 277.400 78.580 277.550 ;
        RECT 74.230 276.950 75.230 277.400 ;
        RECT 70.880 276.800 78.580 276.950 ;
        RECT 74.230 276.350 75.230 276.800 ;
        RECT 70.880 276.200 78.580 276.350 ;
        RECT 74.230 275.750 75.230 276.200 ;
        RECT 70.880 275.600 78.580 275.750 ;
        RECT 74.230 275.150 75.230 275.600 ;
        RECT 70.880 275.000 78.580 275.150 ;
        RECT 74.230 274.550 75.230 275.000 ;
        RECT 70.880 274.400 78.580 274.550 ;
        RECT 74.230 273.950 75.230 274.400 ;
        RECT 70.880 273.800 78.580 273.950 ;
        RECT 74.230 273.350 75.230 273.800 ;
        RECT 70.880 273.200 78.580 273.350 ;
        RECT 74.230 272.750 75.230 273.200 ;
        RECT 70.880 272.600 78.580 272.750 ;
        RECT 74.230 272.150 75.230 272.600 ;
        RECT 70.880 272.000 78.580 272.150 ;
        RECT 74.230 271.550 75.230 272.000 ;
        RECT 70.880 271.400 78.580 271.550 ;
        RECT 74.230 270.950 75.230 271.400 ;
        RECT 70.880 270.800 78.580 270.950 ;
        RECT 74.230 270.300 75.230 270.800 ;
        RECT 79.480 270.300 79.630 277.850 ;
        RECT 80.080 270.300 80.230 277.850 ;
        RECT 80.680 270.300 80.830 277.850 ;
        RECT 81.280 270.300 81.430 277.850 ;
        RECT 81.880 270.300 82.030 277.850 ;
        RECT 82.480 270.300 82.630 277.850 ;
        RECT 82.780 273.200 83.530 275.000 ;
        RECT 85.930 273.200 86.680 275.000 ;
        RECT 82.780 270.450 86.680 273.200 ;
        RECT 82.780 270.300 83.930 270.450 ;
        RECT 65.530 269.700 83.930 270.300 ;
        RECT 65.530 269.550 66.680 269.700 ;
        RECT 62.780 266.800 66.680 269.550 ;
        RECT 62.780 265.050 63.530 266.800 ;
        RECT 65.930 265.050 66.680 266.800 ;
        RECT 66.830 262.150 66.980 269.700 ;
        RECT 67.430 262.150 67.580 269.700 ;
        RECT 68.030 262.150 68.180 269.700 ;
        RECT 68.630 262.150 68.780 269.700 ;
        RECT 69.230 262.150 69.380 269.700 ;
        RECT 69.830 262.150 69.980 269.700 ;
        RECT 74.230 269.200 75.230 269.700 ;
        RECT 70.880 269.050 78.580 269.200 ;
        RECT 74.230 268.600 75.230 269.050 ;
        RECT 70.880 268.450 78.580 268.600 ;
        RECT 74.230 268.000 75.230 268.450 ;
        RECT 70.880 267.850 78.580 268.000 ;
        RECT 74.230 267.400 75.230 267.850 ;
        RECT 70.880 267.250 78.580 267.400 ;
        RECT 74.230 266.800 75.230 267.250 ;
        RECT 70.880 266.650 78.580 266.800 ;
        RECT 74.230 266.200 75.230 266.650 ;
        RECT 70.880 266.050 78.580 266.200 ;
        RECT 74.230 265.600 75.230 266.050 ;
        RECT 70.880 265.450 78.580 265.600 ;
        RECT 74.230 265.000 75.230 265.450 ;
        RECT 70.880 264.850 78.580 265.000 ;
        RECT 74.230 264.400 75.230 264.850 ;
        RECT 70.880 264.250 78.580 264.400 ;
        RECT 74.230 263.800 75.230 264.250 ;
        RECT 70.880 263.650 78.580 263.800 ;
        RECT 74.230 263.200 75.230 263.650 ;
        RECT 70.880 263.050 78.580 263.200 ;
        RECT 74.230 262.600 75.230 263.050 ;
        RECT 70.880 262.450 78.580 262.600 ;
        RECT 74.230 262.000 75.230 262.450 ;
        RECT 79.480 262.150 79.630 269.700 ;
        RECT 80.080 262.150 80.230 269.700 ;
        RECT 80.680 262.150 80.830 269.700 ;
        RECT 81.280 262.150 81.430 269.700 ;
        RECT 81.880 262.150 82.030 269.700 ;
        RECT 82.480 262.150 82.630 269.700 ;
        RECT 82.780 269.550 83.930 269.700 ;
        RECT 84.580 269.550 84.880 270.450 ;
        RECT 85.530 270.300 86.680 270.450 ;
        RECT 86.830 270.300 86.980 277.850 ;
        RECT 87.430 270.300 87.580 277.850 ;
        RECT 88.030 270.300 88.180 277.850 ;
        RECT 88.630 270.300 88.780 277.850 ;
        RECT 89.230 270.300 89.380 277.850 ;
        RECT 89.830 270.300 89.980 277.850 ;
        RECT 94.230 277.550 95.230 278.000 ;
        RECT 90.880 277.400 98.580 277.550 ;
        RECT 94.230 276.950 95.230 277.400 ;
        RECT 90.880 276.800 98.580 276.950 ;
        RECT 94.230 276.350 95.230 276.800 ;
        RECT 90.880 276.200 98.580 276.350 ;
        RECT 94.230 275.750 95.230 276.200 ;
        RECT 90.880 275.600 98.580 275.750 ;
        RECT 94.230 275.150 95.230 275.600 ;
        RECT 90.880 275.000 98.580 275.150 ;
        RECT 94.230 274.550 95.230 275.000 ;
        RECT 90.880 274.400 98.580 274.550 ;
        RECT 94.230 273.950 95.230 274.400 ;
        RECT 90.880 273.800 98.580 273.950 ;
        RECT 94.230 273.350 95.230 273.800 ;
        RECT 90.880 273.200 98.580 273.350 ;
        RECT 94.230 272.750 95.230 273.200 ;
        RECT 90.880 272.600 98.580 272.750 ;
        RECT 94.230 272.150 95.230 272.600 ;
        RECT 90.880 272.000 98.580 272.150 ;
        RECT 94.230 271.550 95.230 272.000 ;
        RECT 90.880 271.400 98.580 271.550 ;
        RECT 94.230 270.950 95.230 271.400 ;
        RECT 90.880 270.800 98.580 270.950 ;
        RECT 94.230 270.300 95.230 270.800 ;
        RECT 99.480 270.300 99.630 277.850 ;
        RECT 100.080 270.300 100.230 277.850 ;
        RECT 100.680 270.300 100.830 277.850 ;
        RECT 101.280 270.300 101.430 277.850 ;
        RECT 101.880 270.300 102.030 277.850 ;
        RECT 102.480 270.300 102.630 277.850 ;
        RECT 102.780 273.200 103.530 275.000 ;
        RECT 105.930 273.200 106.680 275.000 ;
        RECT 102.780 270.450 106.680 273.200 ;
        RECT 102.780 270.300 103.930 270.450 ;
        RECT 85.530 269.700 103.930 270.300 ;
        RECT 85.530 269.550 86.680 269.700 ;
        RECT 82.780 266.800 86.680 269.550 ;
        RECT 82.780 265.050 83.530 266.800 ;
        RECT 85.930 265.050 86.680 266.800 ;
        RECT 86.830 262.150 86.980 269.700 ;
        RECT 87.430 262.150 87.580 269.700 ;
        RECT 88.030 262.150 88.180 269.700 ;
        RECT 88.630 262.150 88.780 269.700 ;
        RECT 89.230 262.150 89.380 269.700 ;
        RECT 89.830 262.150 89.980 269.700 ;
        RECT 94.230 269.200 95.230 269.700 ;
        RECT 90.880 269.050 98.580 269.200 ;
        RECT 94.230 268.600 95.230 269.050 ;
        RECT 90.880 268.450 98.580 268.600 ;
        RECT 94.230 268.000 95.230 268.450 ;
        RECT 90.880 267.850 98.580 268.000 ;
        RECT 94.230 267.400 95.230 267.850 ;
        RECT 90.880 267.250 98.580 267.400 ;
        RECT 94.230 266.800 95.230 267.250 ;
        RECT 90.880 266.650 98.580 266.800 ;
        RECT 94.230 266.200 95.230 266.650 ;
        RECT 90.880 266.050 98.580 266.200 ;
        RECT 94.230 265.600 95.230 266.050 ;
        RECT 90.880 265.450 98.580 265.600 ;
        RECT 94.230 265.000 95.230 265.450 ;
        RECT 90.880 264.850 98.580 265.000 ;
        RECT 94.230 264.400 95.230 264.850 ;
        RECT 90.880 264.250 98.580 264.400 ;
        RECT 94.230 263.800 95.230 264.250 ;
        RECT 90.880 263.650 98.580 263.800 ;
        RECT 94.230 263.200 95.230 263.650 ;
        RECT 90.880 263.050 98.580 263.200 ;
        RECT 94.230 262.600 95.230 263.050 ;
        RECT 90.880 262.450 98.580 262.600 ;
        RECT 94.230 262.000 95.230 262.450 ;
        RECT 99.480 262.150 99.630 269.700 ;
        RECT 100.080 262.150 100.230 269.700 ;
        RECT 100.680 262.150 100.830 269.700 ;
        RECT 101.280 262.150 101.430 269.700 ;
        RECT 101.880 262.150 102.030 269.700 ;
        RECT 102.480 262.150 102.630 269.700 ;
        RECT 102.780 269.550 103.930 269.700 ;
        RECT 104.580 269.550 104.880 270.450 ;
        RECT 105.530 270.300 106.680 270.450 ;
        RECT 106.830 270.300 106.980 277.850 ;
        RECT 107.430 270.300 107.580 277.850 ;
        RECT 108.030 270.300 108.180 277.850 ;
        RECT 108.630 270.300 108.780 277.850 ;
        RECT 109.230 270.300 109.380 277.850 ;
        RECT 109.830 270.300 109.980 277.850 ;
        RECT 114.230 277.550 115.230 278.000 ;
        RECT 110.880 277.400 118.580 277.550 ;
        RECT 114.230 276.950 115.230 277.400 ;
        RECT 110.880 276.800 118.580 276.950 ;
        RECT 114.230 276.350 115.230 276.800 ;
        RECT 110.880 276.200 118.580 276.350 ;
        RECT 114.230 275.750 115.230 276.200 ;
        RECT 110.880 275.600 118.580 275.750 ;
        RECT 114.230 275.150 115.230 275.600 ;
        RECT 110.880 275.000 118.580 275.150 ;
        RECT 114.230 274.550 115.230 275.000 ;
        RECT 110.880 274.400 118.580 274.550 ;
        RECT 114.230 273.950 115.230 274.400 ;
        RECT 110.880 273.800 118.580 273.950 ;
        RECT 114.230 273.350 115.230 273.800 ;
        RECT 110.880 273.200 118.580 273.350 ;
        RECT 114.230 272.750 115.230 273.200 ;
        RECT 110.880 272.600 118.580 272.750 ;
        RECT 114.230 272.150 115.230 272.600 ;
        RECT 110.880 272.000 118.580 272.150 ;
        RECT 114.230 271.550 115.230 272.000 ;
        RECT 110.880 271.400 118.580 271.550 ;
        RECT 114.230 270.950 115.230 271.400 ;
        RECT 110.880 270.800 118.580 270.950 ;
        RECT 114.230 270.300 115.230 270.800 ;
        RECT 119.480 270.300 119.630 277.850 ;
        RECT 120.080 270.300 120.230 277.850 ;
        RECT 120.680 270.300 120.830 277.850 ;
        RECT 121.280 270.300 121.430 277.850 ;
        RECT 121.880 270.300 122.030 277.850 ;
        RECT 122.480 270.300 122.630 277.850 ;
        RECT 122.780 273.200 123.530 275.000 ;
        RECT 122.780 270.605 124.730 273.200 ;
        RECT 122.780 270.450 131.850 270.605 ;
        RECT 122.780 270.300 123.930 270.450 ;
        RECT 105.530 269.700 123.930 270.300 ;
        RECT 105.530 269.550 106.680 269.700 ;
        RECT 102.780 266.800 106.680 269.550 ;
        RECT 102.780 265.050 103.530 266.800 ;
        RECT 105.930 265.050 106.680 266.800 ;
        RECT 106.830 262.150 106.980 269.700 ;
        RECT 107.430 262.150 107.580 269.700 ;
        RECT 108.030 262.150 108.180 269.700 ;
        RECT 108.630 262.150 108.780 269.700 ;
        RECT 109.230 262.150 109.380 269.700 ;
        RECT 109.830 262.150 109.980 269.700 ;
        RECT 114.230 269.200 115.230 269.700 ;
        RECT 110.880 269.050 118.580 269.200 ;
        RECT 114.230 268.600 115.230 269.050 ;
        RECT 110.880 268.450 118.580 268.600 ;
        RECT 114.230 268.000 115.230 268.450 ;
        RECT 110.880 267.850 118.580 268.000 ;
        RECT 114.230 267.400 115.230 267.850 ;
        RECT 110.880 267.250 118.580 267.400 ;
        RECT 114.230 266.800 115.230 267.250 ;
        RECT 110.880 266.650 118.580 266.800 ;
        RECT 114.230 266.200 115.230 266.650 ;
        RECT 110.880 266.050 118.580 266.200 ;
        RECT 114.230 265.600 115.230 266.050 ;
        RECT 110.880 265.450 118.580 265.600 ;
        RECT 114.230 265.000 115.230 265.450 ;
        RECT 110.880 264.850 118.580 265.000 ;
        RECT 114.230 264.400 115.230 264.850 ;
        RECT 110.880 264.250 118.580 264.400 ;
        RECT 114.230 263.800 115.230 264.250 ;
        RECT 110.880 263.650 118.580 263.800 ;
        RECT 114.230 263.200 115.230 263.650 ;
        RECT 110.880 263.050 118.580 263.200 ;
        RECT 114.230 262.600 115.230 263.050 ;
        RECT 110.880 262.450 118.580 262.600 ;
        RECT 114.230 262.000 115.230 262.450 ;
        RECT 119.480 262.150 119.630 269.700 ;
        RECT 120.080 262.150 120.230 269.700 ;
        RECT 120.680 262.150 120.830 269.700 ;
        RECT 121.280 262.150 121.430 269.700 ;
        RECT 121.880 262.150 122.030 269.700 ;
        RECT 122.480 262.150 122.630 269.700 ;
        RECT 122.780 269.550 123.930 269.700 ;
        RECT 124.580 269.550 131.850 270.450 ;
        RECT 122.780 269.330 131.850 269.550 ;
        RECT 122.780 266.800 124.730 269.330 ;
        RECT 122.780 265.050 123.530 266.800 ;
        RECT 10.880 261.850 18.580 262.000 ;
        RECT 30.880 261.850 38.580 262.000 ;
        RECT 50.880 261.850 58.580 262.000 ;
        RECT 70.880 261.850 78.580 262.000 ;
        RECT 90.880 261.850 98.580 262.000 ;
        RECT 110.880 261.850 118.580 262.000 ;
        RECT 14.230 261.200 15.230 261.850 ;
        RECT 34.230 261.200 35.230 261.850 ;
        RECT 54.230 261.200 55.230 261.850 ;
        RECT 74.230 261.200 75.230 261.850 ;
        RECT 94.230 261.200 95.230 261.850 ;
        RECT 114.230 261.200 115.230 261.850 ;
        RECT 11.530 258.800 17.930 261.200 ;
        RECT 31.530 258.800 37.930 261.200 ;
        RECT 51.530 258.800 57.930 261.200 ;
        RECT 71.530 258.800 77.930 261.200 ;
        RECT 91.530 258.800 97.930 261.200 ;
        RECT 111.530 258.800 117.930 261.200 ;
        RECT 14.230 258.150 15.230 258.800 ;
        RECT 34.230 258.150 35.230 258.800 ;
        RECT 54.230 258.150 55.230 258.800 ;
        RECT 74.230 258.150 75.230 258.800 ;
        RECT 94.230 258.150 95.230 258.800 ;
        RECT 114.230 258.150 115.230 258.800 ;
        RECT 10.880 258.000 18.580 258.150 ;
        RECT 30.880 258.000 38.580 258.150 ;
        RECT 50.880 258.000 58.580 258.150 ;
        RECT 70.880 258.000 78.580 258.150 ;
        RECT 90.880 258.000 98.580 258.150 ;
        RECT 110.880 258.000 118.580 258.150 ;
        RECT 5.930 253.200 6.680 255.000 ;
        RECT 4.730 250.450 6.680 253.200 ;
        RECT 4.730 249.550 4.880 250.450 ;
        RECT 5.530 250.300 6.680 250.450 ;
        RECT 6.830 250.300 6.980 257.850 ;
        RECT 7.430 250.300 7.580 257.850 ;
        RECT 8.030 250.300 8.180 257.850 ;
        RECT 8.630 250.300 8.780 257.850 ;
        RECT 9.230 250.300 9.380 257.850 ;
        RECT 9.830 250.300 9.980 257.850 ;
        RECT 14.230 257.550 15.230 258.000 ;
        RECT 10.880 257.400 18.580 257.550 ;
        RECT 14.230 256.950 15.230 257.400 ;
        RECT 10.880 256.800 18.580 256.950 ;
        RECT 14.230 256.350 15.230 256.800 ;
        RECT 10.880 256.200 18.580 256.350 ;
        RECT 14.230 255.750 15.230 256.200 ;
        RECT 10.880 255.600 18.580 255.750 ;
        RECT 14.230 255.150 15.230 255.600 ;
        RECT 10.880 255.000 18.580 255.150 ;
        RECT 14.230 254.550 15.230 255.000 ;
        RECT 10.880 254.400 18.580 254.550 ;
        RECT 14.230 253.950 15.230 254.400 ;
        RECT 10.880 253.800 18.580 253.950 ;
        RECT 14.230 253.350 15.230 253.800 ;
        RECT 10.880 253.200 18.580 253.350 ;
        RECT 14.230 252.750 15.230 253.200 ;
        RECT 10.880 252.600 18.580 252.750 ;
        RECT 14.230 252.150 15.230 252.600 ;
        RECT 10.880 252.000 18.580 252.150 ;
        RECT 14.230 251.550 15.230 252.000 ;
        RECT 10.880 251.400 18.580 251.550 ;
        RECT 14.230 250.950 15.230 251.400 ;
        RECT 10.880 250.800 18.580 250.950 ;
        RECT 14.230 250.300 15.230 250.800 ;
        RECT 19.480 250.300 19.630 257.850 ;
        RECT 20.080 250.300 20.230 257.850 ;
        RECT 20.680 250.300 20.830 257.850 ;
        RECT 21.280 250.300 21.430 257.850 ;
        RECT 21.880 250.300 22.030 257.850 ;
        RECT 22.480 250.300 22.630 257.850 ;
        RECT 22.780 253.200 23.530 255.000 ;
        RECT 25.930 253.200 26.680 255.000 ;
        RECT 22.780 250.450 26.680 253.200 ;
        RECT 22.780 250.300 23.930 250.450 ;
        RECT 5.530 249.700 23.930 250.300 ;
        RECT 5.530 249.550 6.680 249.700 ;
        RECT 4.730 246.800 6.680 249.550 ;
        RECT 5.930 245.050 6.680 246.800 ;
        RECT 6.830 242.150 6.980 249.700 ;
        RECT 7.430 242.150 7.580 249.700 ;
        RECT 8.030 242.150 8.180 249.700 ;
        RECT 8.630 242.150 8.780 249.700 ;
        RECT 9.230 242.150 9.380 249.700 ;
        RECT 9.830 242.150 9.980 249.700 ;
        RECT 14.230 249.200 15.230 249.700 ;
        RECT 10.880 249.050 18.580 249.200 ;
        RECT 14.230 248.600 15.230 249.050 ;
        RECT 10.880 248.450 18.580 248.600 ;
        RECT 14.230 248.000 15.230 248.450 ;
        RECT 10.880 247.850 18.580 248.000 ;
        RECT 14.230 247.400 15.230 247.850 ;
        RECT 10.880 247.250 18.580 247.400 ;
        RECT 14.230 246.800 15.230 247.250 ;
        RECT 10.880 246.650 18.580 246.800 ;
        RECT 14.230 246.200 15.230 246.650 ;
        RECT 10.880 246.050 18.580 246.200 ;
        RECT 14.230 245.600 15.230 246.050 ;
        RECT 10.880 245.450 18.580 245.600 ;
        RECT 14.230 245.000 15.230 245.450 ;
        RECT 10.880 244.850 18.580 245.000 ;
        RECT 14.230 244.400 15.230 244.850 ;
        RECT 10.880 244.250 18.580 244.400 ;
        RECT 14.230 243.800 15.230 244.250 ;
        RECT 10.880 243.650 18.580 243.800 ;
        RECT 14.230 243.200 15.230 243.650 ;
        RECT 10.880 243.050 18.580 243.200 ;
        RECT 14.230 242.600 15.230 243.050 ;
        RECT 10.880 242.450 18.580 242.600 ;
        RECT 14.230 242.000 15.230 242.450 ;
        RECT 19.480 242.150 19.630 249.700 ;
        RECT 20.080 242.150 20.230 249.700 ;
        RECT 20.680 242.150 20.830 249.700 ;
        RECT 21.280 242.150 21.430 249.700 ;
        RECT 21.880 242.150 22.030 249.700 ;
        RECT 22.480 242.150 22.630 249.700 ;
        RECT 22.780 249.550 23.930 249.700 ;
        RECT 24.580 249.550 24.880 250.450 ;
        RECT 25.530 250.300 26.680 250.450 ;
        RECT 26.830 250.300 26.980 257.850 ;
        RECT 27.430 250.300 27.580 257.850 ;
        RECT 28.030 250.300 28.180 257.850 ;
        RECT 28.630 250.300 28.780 257.850 ;
        RECT 29.230 250.300 29.380 257.850 ;
        RECT 29.830 250.300 29.980 257.850 ;
        RECT 34.230 257.550 35.230 258.000 ;
        RECT 30.880 257.400 38.580 257.550 ;
        RECT 34.230 256.950 35.230 257.400 ;
        RECT 30.880 256.800 38.580 256.950 ;
        RECT 34.230 256.350 35.230 256.800 ;
        RECT 30.880 256.200 38.580 256.350 ;
        RECT 34.230 255.750 35.230 256.200 ;
        RECT 30.880 255.600 38.580 255.750 ;
        RECT 34.230 255.150 35.230 255.600 ;
        RECT 30.880 255.000 38.580 255.150 ;
        RECT 34.230 254.550 35.230 255.000 ;
        RECT 30.880 254.400 38.580 254.550 ;
        RECT 34.230 253.950 35.230 254.400 ;
        RECT 30.880 253.800 38.580 253.950 ;
        RECT 34.230 253.350 35.230 253.800 ;
        RECT 30.880 253.200 38.580 253.350 ;
        RECT 34.230 252.750 35.230 253.200 ;
        RECT 30.880 252.600 38.580 252.750 ;
        RECT 34.230 252.150 35.230 252.600 ;
        RECT 30.880 252.000 38.580 252.150 ;
        RECT 34.230 251.550 35.230 252.000 ;
        RECT 30.880 251.400 38.580 251.550 ;
        RECT 34.230 250.950 35.230 251.400 ;
        RECT 30.880 250.800 38.580 250.950 ;
        RECT 34.230 250.300 35.230 250.800 ;
        RECT 39.480 250.300 39.630 257.850 ;
        RECT 40.080 250.300 40.230 257.850 ;
        RECT 40.680 250.300 40.830 257.850 ;
        RECT 41.280 250.300 41.430 257.850 ;
        RECT 41.880 250.300 42.030 257.850 ;
        RECT 42.480 250.300 42.630 257.850 ;
        RECT 42.780 253.200 43.530 255.000 ;
        RECT 45.930 253.200 46.680 255.000 ;
        RECT 42.780 250.450 46.680 253.200 ;
        RECT 42.780 250.300 43.930 250.450 ;
        RECT 25.530 249.700 43.930 250.300 ;
        RECT 25.530 249.550 26.680 249.700 ;
        RECT 22.780 246.800 26.680 249.550 ;
        RECT 22.780 245.050 23.530 246.800 ;
        RECT 25.930 245.050 26.680 246.800 ;
        RECT 26.830 242.150 26.980 249.700 ;
        RECT 27.430 242.150 27.580 249.700 ;
        RECT 28.030 242.150 28.180 249.700 ;
        RECT 28.630 242.150 28.780 249.700 ;
        RECT 29.230 242.150 29.380 249.700 ;
        RECT 29.830 242.150 29.980 249.700 ;
        RECT 34.230 249.200 35.230 249.700 ;
        RECT 30.880 249.050 38.580 249.200 ;
        RECT 34.230 248.600 35.230 249.050 ;
        RECT 30.880 248.450 38.580 248.600 ;
        RECT 34.230 248.000 35.230 248.450 ;
        RECT 30.880 247.850 38.580 248.000 ;
        RECT 34.230 247.400 35.230 247.850 ;
        RECT 30.880 247.250 38.580 247.400 ;
        RECT 34.230 246.800 35.230 247.250 ;
        RECT 30.880 246.650 38.580 246.800 ;
        RECT 34.230 246.200 35.230 246.650 ;
        RECT 30.880 246.050 38.580 246.200 ;
        RECT 34.230 245.600 35.230 246.050 ;
        RECT 30.880 245.450 38.580 245.600 ;
        RECT 34.230 245.000 35.230 245.450 ;
        RECT 30.880 244.850 38.580 245.000 ;
        RECT 34.230 244.400 35.230 244.850 ;
        RECT 30.880 244.250 38.580 244.400 ;
        RECT 34.230 243.800 35.230 244.250 ;
        RECT 30.880 243.650 38.580 243.800 ;
        RECT 34.230 243.200 35.230 243.650 ;
        RECT 30.880 243.050 38.580 243.200 ;
        RECT 34.230 242.600 35.230 243.050 ;
        RECT 30.880 242.450 38.580 242.600 ;
        RECT 34.230 242.000 35.230 242.450 ;
        RECT 39.480 242.150 39.630 249.700 ;
        RECT 40.080 242.150 40.230 249.700 ;
        RECT 40.680 242.150 40.830 249.700 ;
        RECT 41.280 242.150 41.430 249.700 ;
        RECT 41.880 242.150 42.030 249.700 ;
        RECT 42.480 242.150 42.630 249.700 ;
        RECT 42.780 249.550 43.930 249.700 ;
        RECT 44.580 249.550 44.880 250.450 ;
        RECT 45.530 250.300 46.680 250.450 ;
        RECT 46.830 250.300 46.980 257.850 ;
        RECT 47.430 250.300 47.580 257.850 ;
        RECT 48.030 250.300 48.180 257.850 ;
        RECT 48.630 250.300 48.780 257.850 ;
        RECT 49.230 250.300 49.380 257.850 ;
        RECT 49.830 250.300 49.980 257.850 ;
        RECT 54.230 257.550 55.230 258.000 ;
        RECT 50.880 257.400 58.580 257.550 ;
        RECT 54.230 256.950 55.230 257.400 ;
        RECT 50.880 256.800 58.580 256.950 ;
        RECT 54.230 256.350 55.230 256.800 ;
        RECT 50.880 256.200 58.580 256.350 ;
        RECT 54.230 255.750 55.230 256.200 ;
        RECT 50.880 255.600 58.580 255.750 ;
        RECT 54.230 255.150 55.230 255.600 ;
        RECT 50.880 255.000 58.580 255.150 ;
        RECT 54.230 254.550 55.230 255.000 ;
        RECT 50.880 254.400 58.580 254.550 ;
        RECT 54.230 253.950 55.230 254.400 ;
        RECT 50.880 253.800 58.580 253.950 ;
        RECT 54.230 253.350 55.230 253.800 ;
        RECT 50.880 253.200 58.580 253.350 ;
        RECT 54.230 252.750 55.230 253.200 ;
        RECT 50.880 252.600 58.580 252.750 ;
        RECT 54.230 252.150 55.230 252.600 ;
        RECT 50.880 252.000 58.580 252.150 ;
        RECT 54.230 251.550 55.230 252.000 ;
        RECT 50.880 251.400 58.580 251.550 ;
        RECT 54.230 250.950 55.230 251.400 ;
        RECT 50.880 250.800 58.580 250.950 ;
        RECT 54.230 250.300 55.230 250.800 ;
        RECT 59.480 250.300 59.630 257.850 ;
        RECT 60.080 250.300 60.230 257.850 ;
        RECT 60.680 250.300 60.830 257.850 ;
        RECT 61.280 250.300 61.430 257.850 ;
        RECT 61.880 250.300 62.030 257.850 ;
        RECT 62.480 250.300 62.630 257.850 ;
        RECT 62.780 253.200 63.530 255.000 ;
        RECT 65.930 253.200 66.680 255.000 ;
        RECT 62.780 250.450 66.680 253.200 ;
        RECT 62.780 250.300 63.930 250.450 ;
        RECT 45.530 249.700 63.930 250.300 ;
        RECT 45.530 249.550 46.680 249.700 ;
        RECT 42.780 246.800 46.680 249.550 ;
        RECT 42.780 245.050 43.530 246.800 ;
        RECT 45.930 245.050 46.680 246.800 ;
        RECT 46.830 242.150 46.980 249.700 ;
        RECT 47.430 242.150 47.580 249.700 ;
        RECT 48.030 242.150 48.180 249.700 ;
        RECT 48.630 242.150 48.780 249.700 ;
        RECT 49.230 242.150 49.380 249.700 ;
        RECT 49.830 242.150 49.980 249.700 ;
        RECT 54.230 249.200 55.230 249.700 ;
        RECT 50.880 249.050 58.580 249.200 ;
        RECT 54.230 248.600 55.230 249.050 ;
        RECT 50.880 248.450 58.580 248.600 ;
        RECT 54.230 248.000 55.230 248.450 ;
        RECT 50.880 247.850 58.580 248.000 ;
        RECT 54.230 247.400 55.230 247.850 ;
        RECT 50.880 247.250 58.580 247.400 ;
        RECT 54.230 246.800 55.230 247.250 ;
        RECT 50.880 246.650 58.580 246.800 ;
        RECT 54.230 246.200 55.230 246.650 ;
        RECT 50.880 246.050 58.580 246.200 ;
        RECT 54.230 245.600 55.230 246.050 ;
        RECT 50.880 245.450 58.580 245.600 ;
        RECT 54.230 245.000 55.230 245.450 ;
        RECT 50.880 244.850 58.580 245.000 ;
        RECT 54.230 244.400 55.230 244.850 ;
        RECT 50.880 244.250 58.580 244.400 ;
        RECT 54.230 243.800 55.230 244.250 ;
        RECT 50.880 243.650 58.580 243.800 ;
        RECT 54.230 243.200 55.230 243.650 ;
        RECT 50.880 243.050 58.580 243.200 ;
        RECT 54.230 242.600 55.230 243.050 ;
        RECT 50.880 242.450 58.580 242.600 ;
        RECT 54.230 242.000 55.230 242.450 ;
        RECT 59.480 242.150 59.630 249.700 ;
        RECT 60.080 242.150 60.230 249.700 ;
        RECT 60.680 242.150 60.830 249.700 ;
        RECT 61.280 242.150 61.430 249.700 ;
        RECT 61.880 242.150 62.030 249.700 ;
        RECT 62.480 242.150 62.630 249.700 ;
        RECT 62.780 249.550 63.930 249.700 ;
        RECT 64.580 249.550 64.880 250.450 ;
        RECT 65.530 250.300 66.680 250.450 ;
        RECT 66.830 250.300 66.980 257.850 ;
        RECT 67.430 250.300 67.580 257.850 ;
        RECT 68.030 250.300 68.180 257.850 ;
        RECT 68.630 250.300 68.780 257.850 ;
        RECT 69.230 250.300 69.380 257.850 ;
        RECT 69.830 250.300 69.980 257.850 ;
        RECT 74.230 257.550 75.230 258.000 ;
        RECT 70.880 257.400 78.580 257.550 ;
        RECT 74.230 256.950 75.230 257.400 ;
        RECT 70.880 256.800 78.580 256.950 ;
        RECT 74.230 256.350 75.230 256.800 ;
        RECT 70.880 256.200 78.580 256.350 ;
        RECT 74.230 255.750 75.230 256.200 ;
        RECT 70.880 255.600 78.580 255.750 ;
        RECT 74.230 255.150 75.230 255.600 ;
        RECT 70.880 255.000 78.580 255.150 ;
        RECT 74.230 254.550 75.230 255.000 ;
        RECT 70.880 254.400 78.580 254.550 ;
        RECT 74.230 253.950 75.230 254.400 ;
        RECT 70.880 253.800 78.580 253.950 ;
        RECT 74.230 253.350 75.230 253.800 ;
        RECT 70.880 253.200 78.580 253.350 ;
        RECT 74.230 252.750 75.230 253.200 ;
        RECT 70.880 252.600 78.580 252.750 ;
        RECT 74.230 252.150 75.230 252.600 ;
        RECT 70.880 252.000 78.580 252.150 ;
        RECT 74.230 251.550 75.230 252.000 ;
        RECT 70.880 251.400 78.580 251.550 ;
        RECT 74.230 250.950 75.230 251.400 ;
        RECT 70.880 250.800 78.580 250.950 ;
        RECT 74.230 250.300 75.230 250.800 ;
        RECT 79.480 250.300 79.630 257.850 ;
        RECT 80.080 250.300 80.230 257.850 ;
        RECT 80.680 250.300 80.830 257.850 ;
        RECT 81.280 250.300 81.430 257.850 ;
        RECT 81.880 250.300 82.030 257.850 ;
        RECT 82.480 250.300 82.630 257.850 ;
        RECT 82.780 253.200 83.530 255.000 ;
        RECT 85.930 253.200 86.680 255.000 ;
        RECT 82.780 250.450 86.680 253.200 ;
        RECT 82.780 250.300 83.930 250.450 ;
        RECT 65.530 249.700 83.930 250.300 ;
        RECT 65.530 249.550 66.680 249.700 ;
        RECT 62.780 246.800 66.680 249.550 ;
        RECT 62.780 245.050 63.530 246.800 ;
        RECT 65.930 245.050 66.680 246.800 ;
        RECT 66.830 242.150 66.980 249.700 ;
        RECT 67.430 242.150 67.580 249.700 ;
        RECT 68.030 242.150 68.180 249.700 ;
        RECT 68.630 242.150 68.780 249.700 ;
        RECT 69.230 242.150 69.380 249.700 ;
        RECT 69.830 242.150 69.980 249.700 ;
        RECT 74.230 249.200 75.230 249.700 ;
        RECT 70.880 249.050 78.580 249.200 ;
        RECT 74.230 248.600 75.230 249.050 ;
        RECT 70.880 248.450 78.580 248.600 ;
        RECT 74.230 248.000 75.230 248.450 ;
        RECT 70.880 247.850 78.580 248.000 ;
        RECT 74.230 247.400 75.230 247.850 ;
        RECT 70.880 247.250 78.580 247.400 ;
        RECT 74.230 246.800 75.230 247.250 ;
        RECT 70.880 246.650 78.580 246.800 ;
        RECT 74.230 246.200 75.230 246.650 ;
        RECT 70.880 246.050 78.580 246.200 ;
        RECT 74.230 245.600 75.230 246.050 ;
        RECT 70.880 245.450 78.580 245.600 ;
        RECT 74.230 245.000 75.230 245.450 ;
        RECT 70.880 244.850 78.580 245.000 ;
        RECT 74.230 244.400 75.230 244.850 ;
        RECT 70.880 244.250 78.580 244.400 ;
        RECT 74.230 243.800 75.230 244.250 ;
        RECT 70.880 243.650 78.580 243.800 ;
        RECT 74.230 243.200 75.230 243.650 ;
        RECT 70.880 243.050 78.580 243.200 ;
        RECT 74.230 242.600 75.230 243.050 ;
        RECT 70.880 242.450 78.580 242.600 ;
        RECT 74.230 242.000 75.230 242.450 ;
        RECT 79.480 242.150 79.630 249.700 ;
        RECT 80.080 242.150 80.230 249.700 ;
        RECT 80.680 242.150 80.830 249.700 ;
        RECT 81.280 242.150 81.430 249.700 ;
        RECT 81.880 242.150 82.030 249.700 ;
        RECT 82.480 242.150 82.630 249.700 ;
        RECT 82.780 249.550 83.930 249.700 ;
        RECT 84.580 249.550 84.880 250.450 ;
        RECT 85.530 250.300 86.680 250.450 ;
        RECT 86.830 250.300 86.980 257.850 ;
        RECT 87.430 250.300 87.580 257.850 ;
        RECT 88.030 250.300 88.180 257.850 ;
        RECT 88.630 250.300 88.780 257.850 ;
        RECT 89.230 250.300 89.380 257.850 ;
        RECT 89.830 250.300 89.980 257.850 ;
        RECT 94.230 257.550 95.230 258.000 ;
        RECT 90.880 257.400 98.580 257.550 ;
        RECT 94.230 256.950 95.230 257.400 ;
        RECT 90.880 256.800 98.580 256.950 ;
        RECT 94.230 256.350 95.230 256.800 ;
        RECT 90.880 256.200 98.580 256.350 ;
        RECT 94.230 255.750 95.230 256.200 ;
        RECT 90.880 255.600 98.580 255.750 ;
        RECT 94.230 255.150 95.230 255.600 ;
        RECT 90.880 255.000 98.580 255.150 ;
        RECT 94.230 254.550 95.230 255.000 ;
        RECT 90.880 254.400 98.580 254.550 ;
        RECT 94.230 253.950 95.230 254.400 ;
        RECT 90.880 253.800 98.580 253.950 ;
        RECT 94.230 253.350 95.230 253.800 ;
        RECT 90.880 253.200 98.580 253.350 ;
        RECT 94.230 252.750 95.230 253.200 ;
        RECT 90.880 252.600 98.580 252.750 ;
        RECT 94.230 252.150 95.230 252.600 ;
        RECT 90.880 252.000 98.580 252.150 ;
        RECT 94.230 251.550 95.230 252.000 ;
        RECT 90.880 251.400 98.580 251.550 ;
        RECT 94.230 250.950 95.230 251.400 ;
        RECT 90.880 250.800 98.580 250.950 ;
        RECT 94.230 250.300 95.230 250.800 ;
        RECT 99.480 250.300 99.630 257.850 ;
        RECT 100.080 250.300 100.230 257.850 ;
        RECT 100.680 250.300 100.830 257.850 ;
        RECT 101.280 250.300 101.430 257.850 ;
        RECT 101.880 250.300 102.030 257.850 ;
        RECT 102.480 250.300 102.630 257.850 ;
        RECT 102.780 253.200 103.530 255.000 ;
        RECT 105.930 253.200 106.680 255.000 ;
        RECT 102.780 250.450 106.680 253.200 ;
        RECT 102.780 250.300 103.930 250.450 ;
        RECT 85.530 249.700 103.930 250.300 ;
        RECT 85.530 249.550 86.680 249.700 ;
        RECT 82.780 246.800 86.680 249.550 ;
        RECT 82.780 245.050 83.530 246.800 ;
        RECT 85.930 245.050 86.680 246.800 ;
        RECT 86.830 242.150 86.980 249.700 ;
        RECT 87.430 242.150 87.580 249.700 ;
        RECT 88.030 242.150 88.180 249.700 ;
        RECT 88.630 242.150 88.780 249.700 ;
        RECT 89.230 242.150 89.380 249.700 ;
        RECT 89.830 242.150 89.980 249.700 ;
        RECT 94.230 249.200 95.230 249.700 ;
        RECT 90.880 249.050 98.580 249.200 ;
        RECT 94.230 248.600 95.230 249.050 ;
        RECT 90.880 248.450 98.580 248.600 ;
        RECT 94.230 248.000 95.230 248.450 ;
        RECT 90.880 247.850 98.580 248.000 ;
        RECT 94.230 247.400 95.230 247.850 ;
        RECT 90.880 247.250 98.580 247.400 ;
        RECT 94.230 246.800 95.230 247.250 ;
        RECT 90.880 246.650 98.580 246.800 ;
        RECT 94.230 246.200 95.230 246.650 ;
        RECT 90.880 246.050 98.580 246.200 ;
        RECT 94.230 245.600 95.230 246.050 ;
        RECT 90.880 245.450 98.580 245.600 ;
        RECT 94.230 245.000 95.230 245.450 ;
        RECT 90.880 244.850 98.580 245.000 ;
        RECT 94.230 244.400 95.230 244.850 ;
        RECT 90.880 244.250 98.580 244.400 ;
        RECT 94.230 243.800 95.230 244.250 ;
        RECT 90.880 243.650 98.580 243.800 ;
        RECT 94.230 243.200 95.230 243.650 ;
        RECT 90.880 243.050 98.580 243.200 ;
        RECT 94.230 242.600 95.230 243.050 ;
        RECT 90.880 242.450 98.580 242.600 ;
        RECT 94.230 242.000 95.230 242.450 ;
        RECT 99.480 242.150 99.630 249.700 ;
        RECT 100.080 242.150 100.230 249.700 ;
        RECT 100.680 242.150 100.830 249.700 ;
        RECT 101.280 242.150 101.430 249.700 ;
        RECT 101.880 242.150 102.030 249.700 ;
        RECT 102.480 242.150 102.630 249.700 ;
        RECT 102.780 249.550 103.930 249.700 ;
        RECT 104.580 249.550 104.880 250.450 ;
        RECT 105.530 250.300 106.680 250.450 ;
        RECT 106.830 250.300 106.980 257.850 ;
        RECT 107.430 250.300 107.580 257.850 ;
        RECT 108.030 250.300 108.180 257.850 ;
        RECT 108.630 250.300 108.780 257.850 ;
        RECT 109.230 250.300 109.380 257.850 ;
        RECT 109.830 250.300 109.980 257.850 ;
        RECT 114.230 257.550 115.230 258.000 ;
        RECT 110.880 257.400 118.580 257.550 ;
        RECT 114.230 256.950 115.230 257.400 ;
        RECT 110.880 256.800 118.580 256.950 ;
        RECT 114.230 256.350 115.230 256.800 ;
        RECT 110.880 256.200 118.580 256.350 ;
        RECT 114.230 255.750 115.230 256.200 ;
        RECT 110.880 255.600 118.580 255.750 ;
        RECT 114.230 255.150 115.230 255.600 ;
        RECT 110.880 255.000 118.580 255.150 ;
        RECT 114.230 254.550 115.230 255.000 ;
        RECT 110.880 254.400 118.580 254.550 ;
        RECT 114.230 253.950 115.230 254.400 ;
        RECT 110.880 253.800 118.580 253.950 ;
        RECT 114.230 253.350 115.230 253.800 ;
        RECT 110.880 253.200 118.580 253.350 ;
        RECT 114.230 252.750 115.230 253.200 ;
        RECT 110.880 252.600 118.580 252.750 ;
        RECT 114.230 252.150 115.230 252.600 ;
        RECT 110.880 252.000 118.580 252.150 ;
        RECT 114.230 251.550 115.230 252.000 ;
        RECT 110.880 251.400 118.580 251.550 ;
        RECT 114.230 250.950 115.230 251.400 ;
        RECT 110.880 250.800 118.580 250.950 ;
        RECT 114.230 250.300 115.230 250.800 ;
        RECT 119.480 250.300 119.630 257.850 ;
        RECT 120.080 250.300 120.230 257.850 ;
        RECT 120.680 250.300 120.830 257.850 ;
        RECT 121.280 250.300 121.430 257.850 ;
        RECT 121.880 250.300 122.030 257.850 ;
        RECT 122.480 250.300 122.630 257.850 ;
        RECT 122.780 253.200 123.530 255.000 ;
        RECT 122.780 250.520 124.730 253.200 ;
        RECT 122.780 250.450 131.850 250.520 ;
        RECT 122.780 250.300 123.930 250.450 ;
        RECT 105.530 249.700 123.930 250.300 ;
        RECT 105.530 249.550 106.680 249.700 ;
        RECT 102.780 246.800 106.680 249.550 ;
        RECT 102.780 245.050 103.530 246.800 ;
        RECT 105.930 245.050 106.680 246.800 ;
        RECT 106.830 242.150 106.980 249.700 ;
        RECT 107.430 242.150 107.580 249.700 ;
        RECT 108.030 242.150 108.180 249.700 ;
        RECT 108.630 242.150 108.780 249.700 ;
        RECT 109.230 242.150 109.380 249.700 ;
        RECT 109.830 242.150 109.980 249.700 ;
        RECT 114.230 249.200 115.230 249.700 ;
        RECT 110.880 249.050 118.580 249.200 ;
        RECT 114.230 248.600 115.230 249.050 ;
        RECT 110.880 248.450 118.580 248.600 ;
        RECT 114.230 248.000 115.230 248.450 ;
        RECT 110.880 247.850 118.580 248.000 ;
        RECT 114.230 247.400 115.230 247.850 ;
        RECT 110.880 247.250 118.580 247.400 ;
        RECT 114.230 246.800 115.230 247.250 ;
        RECT 110.880 246.650 118.580 246.800 ;
        RECT 114.230 246.200 115.230 246.650 ;
        RECT 110.880 246.050 118.580 246.200 ;
        RECT 114.230 245.600 115.230 246.050 ;
        RECT 110.880 245.450 118.580 245.600 ;
        RECT 114.230 245.000 115.230 245.450 ;
        RECT 110.880 244.850 118.580 245.000 ;
        RECT 114.230 244.400 115.230 244.850 ;
        RECT 110.880 244.250 118.580 244.400 ;
        RECT 114.230 243.800 115.230 244.250 ;
        RECT 110.880 243.650 118.580 243.800 ;
        RECT 114.230 243.200 115.230 243.650 ;
        RECT 110.880 243.050 118.580 243.200 ;
        RECT 114.230 242.600 115.230 243.050 ;
        RECT 110.880 242.450 118.580 242.600 ;
        RECT 114.230 242.000 115.230 242.450 ;
        RECT 119.480 242.150 119.630 249.700 ;
        RECT 120.080 242.150 120.230 249.700 ;
        RECT 120.680 242.150 120.830 249.700 ;
        RECT 121.280 242.150 121.430 249.700 ;
        RECT 121.880 242.150 122.030 249.700 ;
        RECT 122.480 242.150 122.630 249.700 ;
        RECT 122.780 249.550 123.930 249.700 ;
        RECT 124.580 249.550 131.850 250.450 ;
        RECT 122.780 249.245 131.850 249.550 ;
        RECT 122.780 246.800 124.730 249.245 ;
        RECT 122.780 245.050 123.530 246.800 ;
        RECT 10.880 241.850 18.580 242.000 ;
        RECT 30.880 241.850 38.580 242.000 ;
        RECT 50.880 241.850 58.580 242.000 ;
        RECT 70.880 241.850 78.580 242.000 ;
        RECT 90.880 241.850 98.580 242.000 ;
        RECT 110.880 241.850 118.580 242.000 ;
        RECT 14.230 241.200 15.230 241.850 ;
        RECT 34.230 241.200 35.230 241.850 ;
        RECT 54.230 241.200 55.230 241.850 ;
        RECT 74.230 241.200 75.230 241.850 ;
        RECT 94.230 241.200 95.230 241.850 ;
        RECT 114.230 241.200 115.230 241.850 ;
        RECT 11.530 238.800 17.930 241.200 ;
        RECT 31.530 238.800 37.930 241.200 ;
        RECT 51.530 238.800 57.930 241.200 ;
        RECT 71.530 238.800 77.930 241.200 ;
        RECT 91.530 238.800 97.930 241.200 ;
        RECT 111.530 238.800 117.930 241.200 ;
        RECT 14.230 238.150 15.230 238.800 ;
        RECT 34.230 238.150 35.230 238.800 ;
        RECT 54.230 238.150 55.230 238.800 ;
        RECT 74.230 238.150 75.230 238.800 ;
        RECT 94.230 238.150 95.230 238.800 ;
        RECT 114.230 238.150 115.230 238.800 ;
        RECT 10.880 238.000 18.580 238.150 ;
        RECT 30.880 238.000 38.580 238.150 ;
        RECT 50.880 238.000 58.580 238.150 ;
        RECT 70.880 238.000 78.580 238.150 ;
        RECT 90.880 238.000 98.580 238.150 ;
        RECT 110.880 238.000 118.580 238.150 ;
        RECT 5.930 233.200 6.680 235.000 ;
        RECT 4.730 230.450 6.680 233.200 ;
        RECT 4.730 229.550 4.880 230.450 ;
        RECT 5.530 230.300 6.680 230.450 ;
        RECT 6.830 230.300 6.980 237.850 ;
        RECT 7.430 230.300 7.580 237.850 ;
        RECT 8.030 230.300 8.180 237.850 ;
        RECT 8.630 230.300 8.780 237.850 ;
        RECT 9.230 230.300 9.380 237.850 ;
        RECT 9.830 230.300 9.980 237.850 ;
        RECT 14.230 237.550 15.230 238.000 ;
        RECT 10.880 237.400 18.580 237.550 ;
        RECT 14.230 236.950 15.230 237.400 ;
        RECT 10.880 236.800 18.580 236.950 ;
        RECT 14.230 236.350 15.230 236.800 ;
        RECT 10.880 236.200 18.580 236.350 ;
        RECT 14.230 235.750 15.230 236.200 ;
        RECT 10.880 235.600 18.580 235.750 ;
        RECT 14.230 235.150 15.230 235.600 ;
        RECT 10.880 235.000 18.580 235.150 ;
        RECT 14.230 234.550 15.230 235.000 ;
        RECT 10.880 234.400 18.580 234.550 ;
        RECT 14.230 233.950 15.230 234.400 ;
        RECT 10.880 233.800 18.580 233.950 ;
        RECT 14.230 233.350 15.230 233.800 ;
        RECT 10.880 233.200 18.580 233.350 ;
        RECT 14.230 232.750 15.230 233.200 ;
        RECT 10.880 232.600 18.580 232.750 ;
        RECT 14.230 232.150 15.230 232.600 ;
        RECT 10.880 232.000 18.580 232.150 ;
        RECT 14.230 231.550 15.230 232.000 ;
        RECT 10.880 231.400 18.580 231.550 ;
        RECT 14.230 230.950 15.230 231.400 ;
        RECT 10.880 230.800 18.580 230.950 ;
        RECT 14.230 230.300 15.230 230.800 ;
        RECT 19.480 230.300 19.630 237.850 ;
        RECT 20.080 230.300 20.230 237.850 ;
        RECT 20.680 230.300 20.830 237.850 ;
        RECT 21.280 230.300 21.430 237.850 ;
        RECT 21.880 230.300 22.030 237.850 ;
        RECT 22.480 230.300 22.630 237.850 ;
        RECT 22.780 233.200 23.530 235.000 ;
        RECT 25.930 233.200 26.680 235.000 ;
        RECT 22.780 230.450 26.680 233.200 ;
        RECT 22.780 230.300 23.930 230.450 ;
        RECT 5.530 229.700 23.930 230.300 ;
        RECT 5.530 229.550 6.680 229.700 ;
        RECT 4.730 226.800 6.680 229.550 ;
        RECT 5.930 225.050 6.680 226.800 ;
        RECT 6.830 222.150 6.980 229.700 ;
        RECT 7.430 222.150 7.580 229.700 ;
        RECT 8.030 222.150 8.180 229.700 ;
        RECT 8.630 222.150 8.780 229.700 ;
        RECT 9.230 222.150 9.380 229.700 ;
        RECT 9.830 222.150 9.980 229.700 ;
        RECT 14.230 229.200 15.230 229.700 ;
        RECT 10.880 229.050 18.580 229.200 ;
        RECT 14.230 228.600 15.230 229.050 ;
        RECT 10.880 228.450 18.580 228.600 ;
        RECT 14.230 228.000 15.230 228.450 ;
        RECT 10.880 227.850 18.580 228.000 ;
        RECT 14.230 227.400 15.230 227.850 ;
        RECT 10.880 227.250 18.580 227.400 ;
        RECT 14.230 226.800 15.230 227.250 ;
        RECT 10.880 226.650 18.580 226.800 ;
        RECT 14.230 226.200 15.230 226.650 ;
        RECT 10.880 226.050 18.580 226.200 ;
        RECT 14.230 225.600 15.230 226.050 ;
        RECT 10.880 225.450 18.580 225.600 ;
        RECT 14.230 225.000 15.230 225.450 ;
        RECT 10.880 224.850 18.580 225.000 ;
        RECT 14.230 224.400 15.230 224.850 ;
        RECT 10.880 224.250 18.580 224.400 ;
        RECT 14.230 223.800 15.230 224.250 ;
        RECT 10.880 223.650 18.580 223.800 ;
        RECT 14.230 223.200 15.230 223.650 ;
        RECT 10.880 223.050 18.580 223.200 ;
        RECT 14.230 222.600 15.230 223.050 ;
        RECT 10.880 222.450 18.580 222.600 ;
        RECT 14.230 222.000 15.230 222.450 ;
        RECT 19.480 222.150 19.630 229.700 ;
        RECT 20.080 222.150 20.230 229.700 ;
        RECT 20.680 222.150 20.830 229.700 ;
        RECT 21.280 222.150 21.430 229.700 ;
        RECT 21.880 222.150 22.030 229.700 ;
        RECT 22.480 222.150 22.630 229.700 ;
        RECT 22.780 229.550 23.930 229.700 ;
        RECT 24.580 229.550 24.880 230.450 ;
        RECT 25.530 230.300 26.680 230.450 ;
        RECT 26.830 230.300 26.980 237.850 ;
        RECT 27.430 230.300 27.580 237.850 ;
        RECT 28.030 230.300 28.180 237.850 ;
        RECT 28.630 230.300 28.780 237.850 ;
        RECT 29.230 230.300 29.380 237.850 ;
        RECT 29.830 230.300 29.980 237.850 ;
        RECT 34.230 237.550 35.230 238.000 ;
        RECT 30.880 237.400 38.580 237.550 ;
        RECT 34.230 236.950 35.230 237.400 ;
        RECT 30.880 236.800 38.580 236.950 ;
        RECT 34.230 236.350 35.230 236.800 ;
        RECT 30.880 236.200 38.580 236.350 ;
        RECT 34.230 235.750 35.230 236.200 ;
        RECT 30.880 235.600 38.580 235.750 ;
        RECT 34.230 235.150 35.230 235.600 ;
        RECT 30.880 235.000 38.580 235.150 ;
        RECT 34.230 234.550 35.230 235.000 ;
        RECT 30.880 234.400 38.580 234.550 ;
        RECT 34.230 233.950 35.230 234.400 ;
        RECT 30.880 233.800 38.580 233.950 ;
        RECT 34.230 233.350 35.230 233.800 ;
        RECT 30.880 233.200 38.580 233.350 ;
        RECT 34.230 232.750 35.230 233.200 ;
        RECT 30.880 232.600 38.580 232.750 ;
        RECT 34.230 232.150 35.230 232.600 ;
        RECT 30.880 232.000 38.580 232.150 ;
        RECT 34.230 231.550 35.230 232.000 ;
        RECT 30.880 231.400 38.580 231.550 ;
        RECT 34.230 230.950 35.230 231.400 ;
        RECT 30.880 230.800 38.580 230.950 ;
        RECT 34.230 230.300 35.230 230.800 ;
        RECT 39.480 230.300 39.630 237.850 ;
        RECT 40.080 230.300 40.230 237.850 ;
        RECT 40.680 230.300 40.830 237.850 ;
        RECT 41.280 230.300 41.430 237.850 ;
        RECT 41.880 230.300 42.030 237.850 ;
        RECT 42.480 230.300 42.630 237.850 ;
        RECT 42.780 233.200 43.530 235.000 ;
        RECT 45.930 233.200 46.680 235.000 ;
        RECT 42.780 230.450 46.680 233.200 ;
        RECT 42.780 230.300 43.930 230.450 ;
        RECT 25.530 229.700 43.930 230.300 ;
        RECT 25.530 229.550 26.680 229.700 ;
        RECT 22.780 226.800 26.680 229.550 ;
        RECT 22.780 225.050 23.530 226.800 ;
        RECT 25.930 225.050 26.680 226.800 ;
        RECT 26.830 222.150 26.980 229.700 ;
        RECT 27.430 222.150 27.580 229.700 ;
        RECT 28.030 222.150 28.180 229.700 ;
        RECT 28.630 222.150 28.780 229.700 ;
        RECT 29.230 222.150 29.380 229.700 ;
        RECT 29.830 222.150 29.980 229.700 ;
        RECT 34.230 229.200 35.230 229.700 ;
        RECT 30.880 229.050 38.580 229.200 ;
        RECT 34.230 228.600 35.230 229.050 ;
        RECT 30.880 228.450 38.580 228.600 ;
        RECT 34.230 228.000 35.230 228.450 ;
        RECT 30.880 227.850 38.580 228.000 ;
        RECT 34.230 227.400 35.230 227.850 ;
        RECT 30.880 227.250 38.580 227.400 ;
        RECT 34.230 226.800 35.230 227.250 ;
        RECT 30.880 226.650 38.580 226.800 ;
        RECT 34.230 226.200 35.230 226.650 ;
        RECT 30.880 226.050 38.580 226.200 ;
        RECT 34.230 225.600 35.230 226.050 ;
        RECT 30.880 225.450 38.580 225.600 ;
        RECT 34.230 225.000 35.230 225.450 ;
        RECT 30.880 224.850 38.580 225.000 ;
        RECT 34.230 224.400 35.230 224.850 ;
        RECT 30.880 224.250 38.580 224.400 ;
        RECT 34.230 223.800 35.230 224.250 ;
        RECT 30.880 223.650 38.580 223.800 ;
        RECT 34.230 223.200 35.230 223.650 ;
        RECT 30.880 223.050 38.580 223.200 ;
        RECT 34.230 222.600 35.230 223.050 ;
        RECT 30.880 222.450 38.580 222.600 ;
        RECT 34.230 222.000 35.230 222.450 ;
        RECT 39.480 222.150 39.630 229.700 ;
        RECT 40.080 222.150 40.230 229.700 ;
        RECT 40.680 222.150 40.830 229.700 ;
        RECT 41.280 222.150 41.430 229.700 ;
        RECT 41.880 222.150 42.030 229.700 ;
        RECT 42.480 222.150 42.630 229.700 ;
        RECT 42.780 229.550 43.930 229.700 ;
        RECT 44.580 229.550 44.880 230.450 ;
        RECT 45.530 230.300 46.680 230.450 ;
        RECT 46.830 230.300 46.980 237.850 ;
        RECT 47.430 230.300 47.580 237.850 ;
        RECT 48.030 230.300 48.180 237.850 ;
        RECT 48.630 230.300 48.780 237.850 ;
        RECT 49.230 230.300 49.380 237.850 ;
        RECT 49.830 230.300 49.980 237.850 ;
        RECT 54.230 237.550 55.230 238.000 ;
        RECT 50.880 237.400 58.580 237.550 ;
        RECT 54.230 236.950 55.230 237.400 ;
        RECT 50.880 236.800 58.580 236.950 ;
        RECT 54.230 236.350 55.230 236.800 ;
        RECT 50.880 236.200 58.580 236.350 ;
        RECT 54.230 235.750 55.230 236.200 ;
        RECT 50.880 235.600 58.580 235.750 ;
        RECT 54.230 235.150 55.230 235.600 ;
        RECT 50.880 235.000 58.580 235.150 ;
        RECT 54.230 234.550 55.230 235.000 ;
        RECT 50.880 234.400 58.580 234.550 ;
        RECT 54.230 233.950 55.230 234.400 ;
        RECT 50.880 233.800 58.580 233.950 ;
        RECT 54.230 233.350 55.230 233.800 ;
        RECT 50.880 233.200 58.580 233.350 ;
        RECT 54.230 232.750 55.230 233.200 ;
        RECT 50.880 232.600 58.580 232.750 ;
        RECT 54.230 232.150 55.230 232.600 ;
        RECT 50.880 232.000 58.580 232.150 ;
        RECT 54.230 231.550 55.230 232.000 ;
        RECT 50.880 231.400 58.580 231.550 ;
        RECT 54.230 230.950 55.230 231.400 ;
        RECT 50.880 230.800 58.580 230.950 ;
        RECT 54.230 230.300 55.230 230.800 ;
        RECT 59.480 230.300 59.630 237.850 ;
        RECT 60.080 230.300 60.230 237.850 ;
        RECT 60.680 230.300 60.830 237.850 ;
        RECT 61.280 230.300 61.430 237.850 ;
        RECT 61.880 230.300 62.030 237.850 ;
        RECT 62.480 230.300 62.630 237.850 ;
        RECT 62.780 233.200 63.530 235.000 ;
        RECT 65.930 233.200 66.680 235.000 ;
        RECT 62.780 230.450 66.680 233.200 ;
        RECT 62.780 230.300 63.930 230.450 ;
        RECT 45.530 229.700 63.930 230.300 ;
        RECT 45.530 229.550 46.680 229.700 ;
        RECT 42.780 226.800 46.680 229.550 ;
        RECT 42.780 225.050 43.530 226.800 ;
        RECT 45.930 225.050 46.680 226.800 ;
        RECT 46.830 222.150 46.980 229.700 ;
        RECT 47.430 222.150 47.580 229.700 ;
        RECT 48.030 222.150 48.180 229.700 ;
        RECT 48.630 222.150 48.780 229.700 ;
        RECT 49.230 222.150 49.380 229.700 ;
        RECT 49.830 222.150 49.980 229.700 ;
        RECT 54.230 229.200 55.230 229.700 ;
        RECT 50.880 229.050 58.580 229.200 ;
        RECT 54.230 228.600 55.230 229.050 ;
        RECT 50.880 228.450 58.580 228.600 ;
        RECT 54.230 228.000 55.230 228.450 ;
        RECT 50.880 227.850 58.580 228.000 ;
        RECT 54.230 227.400 55.230 227.850 ;
        RECT 50.880 227.250 58.580 227.400 ;
        RECT 54.230 226.800 55.230 227.250 ;
        RECT 50.880 226.650 58.580 226.800 ;
        RECT 54.230 226.200 55.230 226.650 ;
        RECT 50.880 226.050 58.580 226.200 ;
        RECT 54.230 225.600 55.230 226.050 ;
        RECT 50.880 225.450 58.580 225.600 ;
        RECT 54.230 225.000 55.230 225.450 ;
        RECT 50.880 224.850 58.580 225.000 ;
        RECT 54.230 224.400 55.230 224.850 ;
        RECT 50.880 224.250 58.580 224.400 ;
        RECT 54.230 223.800 55.230 224.250 ;
        RECT 50.880 223.650 58.580 223.800 ;
        RECT 54.230 223.200 55.230 223.650 ;
        RECT 50.880 223.050 58.580 223.200 ;
        RECT 54.230 222.600 55.230 223.050 ;
        RECT 50.880 222.450 58.580 222.600 ;
        RECT 54.230 222.000 55.230 222.450 ;
        RECT 59.480 222.150 59.630 229.700 ;
        RECT 60.080 222.150 60.230 229.700 ;
        RECT 60.680 222.150 60.830 229.700 ;
        RECT 61.280 222.150 61.430 229.700 ;
        RECT 61.880 222.150 62.030 229.700 ;
        RECT 62.480 222.150 62.630 229.700 ;
        RECT 62.780 229.550 63.930 229.700 ;
        RECT 64.580 229.550 64.880 230.450 ;
        RECT 65.530 230.300 66.680 230.450 ;
        RECT 66.830 230.300 66.980 237.850 ;
        RECT 67.430 230.300 67.580 237.850 ;
        RECT 68.030 230.300 68.180 237.850 ;
        RECT 68.630 230.300 68.780 237.850 ;
        RECT 69.230 230.300 69.380 237.850 ;
        RECT 69.830 230.300 69.980 237.850 ;
        RECT 74.230 237.550 75.230 238.000 ;
        RECT 70.880 237.400 78.580 237.550 ;
        RECT 74.230 236.950 75.230 237.400 ;
        RECT 70.880 236.800 78.580 236.950 ;
        RECT 74.230 236.350 75.230 236.800 ;
        RECT 70.880 236.200 78.580 236.350 ;
        RECT 74.230 235.750 75.230 236.200 ;
        RECT 70.880 235.600 78.580 235.750 ;
        RECT 74.230 235.150 75.230 235.600 ;
        RECT 70.880 235.000 78.580 235.150 ;
        RECT 74.230 234.550 75.230 235.000 ;
        RECT 70.880 234.400 78.580 234.550 ;
        RECT 74.230 233.950 75.230 234.400 ;
        RECT 70.880 233.800 78.580 233.950 ;
        RECT 74.230 233.350 75.230 233.800 ;
        RECT 70.880 233.200 78.580 233.350 ;
        RECT 74.230 232.750 75.230 233.200 ;
        RECT 70.880 232.600 78.580 232.750 ;
        RECT 74.230 232.150 75.230 232.600 ;
        RECT 70.880 232.000 78.580 232.150 ;
        RECT 74.230 231.550 75.230 232.000 ;
        RECT 70.880 231.400 78.580 231.550 ;
        RECT 74.230 230.950 75.230 231.400 ;
        RECT 70.880 230.800 78.580 230.950 ;
        RECT 74.230 230.300 75.230 230.800 ;
        RECT 79.480 230.300 79.630 237.850 ;
        RECT 80.080 230.300 80.230 237.850 ;
        RECT 80.680 230.300 80.830 237.850 ;
        RECT 81.280 230.300 81.430 237.850 ;
        RECT 81.880 230.300 82.030 237.850 ;
        RECT 82.480 230.300 82.630 237.850 ;
        RECT 82.780 233.200 83.530 235.000 ;
        RECT 85.930 233.200 86.680 235.000 ;
        RECT 82.780 230.450 86.680 233.200 ;
        RECT 82.780 230.300 83.930 230.450 ;
        RECT 65.530 229.700 83.930 230.300 ;
        RECT 65.530 229.550 66.680 229.700 ;
        RECT 62.780 226.800 66.680 229.550 ;
        RECT 62.780 225.050 63.530 226.800 ;
        RECT 65.930 225.050 66.680 226.800 ;
        RECT 66.830 222.150 66.980 229.700 ;
        RECT 67.430 222.150 67.580 229.700 ;
        RECT 68.030 222.150 68.180 229.700 ;
        RECT 68.630 222.150 68.780 229.700 ;
        RECT 69.230 222.150 69.380 229.700 ;
        RECT 69.830 222.150 69.980 229.700 ;
        RECT 74.230 229.200 75.230 229.700 ;
        RECT 70.880 229.050 78.580 229.200 ;
        RECT 74.230 228.600 75.230 229.050 ;
        RECT 70.880 228.450 78.580 228.600 ;
        RECT 74.230 228.000 75.230 228.450 ;
        RECT 70.880 227.850 78.580 228.000 ;
        RECT 74.230 227.400 75.230 227.850 ;
        RECT 70.880 227.250 78.580 227.400 ;
        RECT 74.230 226.800 75.230 227.250 ;
        RECT 70.880 226.650 78.580 226.800 ;
        RECT 74.230 226.200 75.230 226.650 ;
        RECT 70.880 226.050 78.580 226.200 ;
        RECT 74.230 225.600 75.230 226.050 ;
        RECT 70.880 225.450 78.580 225.600 ;
        RECT 74.230 225.000 75.230 225.450 ;
        RECT 70.880 224.850 78.580 225.000 ;
        RECT 74.230 224.400 75.230 224.850 ;
        RECT 70.880 224.250 78.580 224.400 ;
        RECT 74.230 223.800 75.230 224.250 ;
        RECT 70.880 223.650 78.580 223.800 ;
        RECT 74.230 223.200 75.230 223.650 ;
        RECT 70.880 223.050 78.580 223.200 ;
        RECT 74.230 222.600 75.230 223.050 ;
        RECT 70.880 222.450 78.580 222.600 ;
        RECT 74.230 222.000 75.230 222.450 ;
        RECT 79.480 222.150 79.630 229.700 ;
        RECT 80.080 222.150 80.230 229.700 ;
        RECT 80.680 222.150 80.830 229.700 ;
        RECT 81.280 222.150 81.430 229.700 ;
        RECT 81.880 222.150 82.030 229.700 ;
        RECT 82.480 222.150 82.630 229.700 ;
        RECT 82.780 229.550 83.930 229.700 ;
        RECT 84.580 229.550 84.880 230.450 ;
        RECT 85.530 230.300 86.680 230.450 ;
        RECT 86.830 230.300 86.980 237.850 ;
        RECT 87.430 230.300 87.580 237.850 ;
        RECT 88.030 230.300 88.180 237.850 ;
        RECT 88.630 230.300 88.780 237.850 ;
        RECT 89.230 230.300 89.380 237.850 ;
        RECT 89.830 230.300 89.980 237.850 ;
        RECT 94.230 237.550 95.230 238.000 ;
        RECT 90.880 237.400 98.580 237.550 ;
        RECT 94.230 236.950 95.230 237.400 ;
        RECT 90.880 236.800 98.580 236.950 ;
        RECT 94.230 236.350 95.230 236.800 ;
        RECT 90.880 236.200 98.580 236.350 ;
        RECT 94.230 235.750 95.230 236.200 ;
        RECT 90.880 235.600 98.580 235.750 ;
        RECT 94.230 235.150 95.230 235.600 ;
        RECT 90.880 235.000 98.580 235.150 ;
        RECT 94.230 234.550 95.230 235.000 ;
        RECT 90.880 234.400 98.580 234.550 ;
        RECT 94.230 233.950 95.230 234.400 ;
        RECT 90.880 233.800 98.580 233.950 ;
        RECT 94.230 233.350 95.230 233.800 ;
        RECT 90.880 233.200 98.580 233.350 ;
        RECT 94.230 232.750 95.230 233.200 ;
        RECT 90.880 232.600 98.580 232.750 ;
        RECT 94.230 232.150 95.230 232.600 ;
        RECT 90.880 232.000 98.580 232.150 ;
        RECT 94.230 231.550 95.230 232.000 ;
        RECT 90.880 231.400 98.580 231.550 ;
        RECT 94.230 230.950 95.230 231.400 ;
        RECT 90.880 230.800 98.580 230.950 ;
        RECT 94.230 230.300 95.230 230.800 ;
        RECT 99.480 230.300 99.630 237.850 ;
        RECT 100.080 230.300 100.230 237.850 ;
        RECT 100.680 230.300 100.830 237.850 ;
        RECT 101.280 230.300 101.430 237.850 ;
        RECT 101.880 230.300 102.030 237.850 ;
        RECT 102.480 230.300 102.630 237.850 ;
        RECT 102.780 233.200 103.530 235.000 ;
        RECT 105.930 233.200 106.680 235.000 ;
        RECT 102.780 230.450 106.680 233.200 ;
        RECT 102.780 230.300 103.930 230.450 ;
        RECT 85.530 229.700 103.930 230.300 ;
        RECT 85.530 229.550 86.680 229.700 ;
        RECT 82.780 226.800 86.680 229.550 ;
        RECT 82.780 225.050 83.530 226.800 ;
        RECT 85.930 225.050 86.680 226.800 ;
        RECT 86.830 222.150 86.980 229.700 ;
        RECT 87.430 222.150 87.580 229.700 ;
        RECT 88.030 222.150 88.180 229.700 ;
        RECT 88.630 222.150 88.780 229.700 ;
        RECT 89.230 222.150 89.380 229.700 ;
        RECT 89.830 222.150 89.980 229.700 ;
        RECT 94.230 229.200 95.230 229.700 ;
        RECT 90.880 229.050 98.580 229.200 ;
        RECT 94.230 228.600 95.230 229.050 ;
        RECT 90.880 228.450 98.580 228.600 ;
        RECT 94.230 228.000 95.230 228.450 ;
        RECT 90.880 227.850 98.580 228.000 ;
        RECT 94.230 227.400 95.230 227.850 ;
        RECT 90.880 227.250 98.580 227.400 ;
        RECT 94.230 226.800 95.230 227.250 ;
        RECT 90.880 226.650 98.580 226.800 ;
        RECT 94.230 226.200 95.230 226.650 ;
        RECT 90.880 226.050 98.580 226.200 ;
        RECT 94.230 225.600 95.230 226.050 ;
        RECT 90.880 225.450 98.580 225.600 ;
        RECT 94.230 225.000 95.230 225.450 ;
        RECT 90.880 224.850 98.580 225.000 ;
        RECT 94.230 224.400 95.230 224.850 ;
        RECT 90.880 224.250 98.580 224.400 ;
        RECT 94.230 223.800 95.230 224.250 ;
        RECT 90.880 223.650 98.580 223.800 ;
        RECT 94.230 223.200 95.230 223.650 ;
        RECT 90.880 223.050 98.580 223.200 ;
        RECT 94.230 222.600 95.230 223.050 ;
        RECT 90.880 222.450 98.580 222.600 ;
        RECT 94.230 222.000 95.230 222.450 ;
        RECT 99.480 222.150 99.630 229.700 ;
        RECT 100.080 222.150 100.230 229.700 ;
        RECT 100.680 222.150 100.830 229.700 ;
        RECT 101.280 222.150 101.430 229.700 ;
        RECT 101.880 222.150 102.030 229.700 ;
        RECT 102.480 222.150 102.630 229.700 ;
        RECT 102.780 229.550 103.930 229.700 ;
        RECT 104.580 229.550 104.880 230.450 ;
        RECT 105.530 230.300 106.680 230.450 ;
        RECT 106.830 230.300 106.980 237.850 ;
        RECT 107.430 230.300 107.580 237.850 ;
        RECT 108.030 230.300 108.180 237.850 ;
        RECT 108.630 230.300 108.780 237.850 ;
        RECT 109.230 230.300 109.380 237.850 ;
        RECT 109.830 230.300 109.980 237.850 ;
        RECT 114.230 237.550 115.230 238.000 ;
        RECT 110.880 237.400 118.580 237.550 ;
        RECT 114.230 236.950 115.230 237.400 ;
        RECT 110.880 236.800 118.580 236.950 ;
        RECT 114.230 236.350 115.230 236.800 ;
        RECT 110.880 236.200 118.580 236.350 ;
        RECT 114.230 235.750 115.230 236.200 ;
        RECT 110.880 235.600 118.580 235.750 ;
        RECT 114.230 235.150 115.230 235.600 ;
        RECT 110.880 235.000 118.580 235.150 ;
        RECT 114.230 234.550 115.230 235.000 ;
        RECT 110.880 234.400 118.580 234.550 ;
        RECT 114.230 233.950 115.230 234.400 ;
        RECT 110.880 233.800 118.580 233.950 ;
        RECT 114.230 233.350 115.230 233.800 ;
        RECT 110.880 233.200 118.580 233.350 ;
        RECT 114.230 232.750 115.230 233.200 ;
        RECT 110.880 232.600 118.580 232.750 ;
        RECT 114.230 232.150 115.230 232.600 ;
        RECT 110.880 232.000 118.580 232.150 ;
        RECT 114.230 231.550 115.230 232.000 ;
        RECT 110.880 231.400 118.580 231.550 ;
        RECT 114.230 230.950 115.230 231.400 ;
        RECT 110.880 230.800 118.580 230.950 ;
        RECT 114.230 230.300 115.230 230.800 ;
        RECT 119.480 230.300 119.630 237.850 ;
        RECT 120.080 230.300 120.230 237.850 ;
        RECT 120.680 230.300 120.830 237.850 ;
        RECT 121.280 230.300 121.430 237.850 ;
        RECT 121.880 230.300 122.030 237.850 ;
        RECT 122.480 230.300 122.630 237.850 ;
        RECT 122.780 233.200 123.530 235.000 ;
        RECT 122.780 230.915 124.730 233.200 ;
        RECT 122.780 230.450 131.850 230.915 ;
        RECT 122.780 230.300 123.930 230.450 ;
        RECT 105.530 229.700 123.930 230.300 ;
        RECT 105.530 229.550 106.680 229.700 ;
        RECT 102.780 226.800 106.680 229.550 ;
        RECT 102.780 225.050 103.530 226.800 ;
        RECT 105.930 225.050 106.680 226.800 ;
        RECT 106.830 222.150 106.980 229.700 ;
        RECT 107.430 222.150 107.580 229.700 ;
        RECT 108.030 222.150 108.180 229.700 ;
        RECT 108.630 222.150 108.780 229.700 ;
        RECT 109.230 222.150 109.380 229.700 ;
        RECT 109.830 222.150 109.980 229.700 ;
        RECT 114.230 229.200 115.230 229.700 ;
        RECT 110.880 229.050 118.580 229.200 ;
        RECT 114.230 228.600 115.230 229.050 ;
        RECT 110.880 228.450 118.580 228.600 ;
        RECT 114.230 228.000 115.230 228.450 ;
        RECT 110.880 227.850 118.580 228.000 ;
        RECT 114.230 227.400 115.230 227.850 ;
        RECT 110.880 227.250 118.580 227.400 ;
        RECT 114.230 226.800 115.230 227.250 ;
        RECT 110.880 226.650 118.580 226.800 ;
        RECT 114.230 226.200 115.230 226.650 ;
        RECT 110.880 226.050 118.580 226.200 ;
        RECT 114.230 225.600 115.230 226.050 ;
        RECT 110.880 225.450 118.580 225.600 ;
        RECT 114.230 225.000 115.230 225.450 ;
        RECT 110.880 224.850 118.580 225.000 ;
        RECT 114.230 224.400 115.230 224.850 ;
        RECT 110.880 224.250 118.580 224.400 ;
        RECT 114.230 223.800 115.230 224.250 ;
        RECT 110.880 223.650 118.580 223.800 ;
        RECT 114.230 223.200 115.230 223.650 ;
        RECT 110.880 223.050 118.580 223.200 ;
        RECT 114.230 222.600 115.230 223.050 ;
        RECT 110.880 222.450 118.580 222.600 ;
        RECT 114.230 222.000 115.230 222.450 ;
        RECT 119.480 222.150 119.630 229.700 ;
        RECT 120.080 222.150 120.230 229.700 ;
        RECT 120.680 222.150 120.830 229.700 ;
        RECT 121.280 222.150 121.430 229.700 ;
        RECT 121.880 222.150 122.030 229.700 ;
        RECT 122.480 222.150 122.630 229.700 ;
        RECT 122.780 229.550 123.930 229.700 ;
        RECT 124.580 229.640 131.850 230.450 ;
        RECT 124.580 229.550 124.730 229.640 ;
        RECT 122.780 226.800 124.730 229.550 ;
        RECT 122.780 225.050 123.530 226.800 ;
        RECT 10.880 221.850 18.580 222.000 ;
        RECT 30.880 221.850 38.580 222.000 ;
        RECT 50.880 221.850 58.580 222.000 ;
        RECT 70.880 221.850 78.580 222.000 ;
        RECT 90.880 221.850 98.580 222.000 ;
        RECT 110.880 221.850 118.580 222.000 ;
        RECT 14.230 221.200 15.230 221.850 ;
        RECT 34.230 221.200 35.230 221.850 ;
        RECT 54.230 221.200 55.230 221.850 ;
        RECT 74.230 221.200 75.230 221.850 ;
        RECT 94.230 221.200 95.230 221.850 ;
        RECT 114.230 221.200 115.230 221.850 ;
        RECT 11.530 218.800 17.930 221.200 ;
        RECT 31.530 218.800 37.930 221.200 ;
        RECT 51.530 218.800 57.930 221.200 ;
        RECT 71.530 218.800 77.930 221.200 ;
        RECT 91.530 218.800 97.930 221.200 ;
        RECT 111.530 218.800 117.930 221.200 ;
        RECT 14.230 218.150 15.230 218.800 ;
        RECT 34.230 218.150 35.230 218.800 ;
        RECT 54.230 218.150 55.230 218.800 ;
        RECT 74.230 218.150 75.230 218.800 ;
        RECT 94.230 218.150 95.230 218.800 ;
        RECT 114.230 218.150 115.230 218.800 ;
        RECT 10.880 218.000 18.580 218.150 ;
        RECT 30.880 218.000 38.580 218.150 ;
        RECT 50.880 218.000 58.580 218.150 ;
        RECT 70.880 218.000 78.580 218.150 ;
        RECT 90.880 218.000 98.580 218.150 ;
        RECT 110.880 218.000 118.580 218.150 ;
        RECT 5.930 213.200 6.680 215.000 ;
        RECT 4.730 210.450 6.680 213.200 ;
        RECT 4.730 209.550 4.880 210.450 ;
        RECT 5.530 210.300 6.680 210.450 ;
        RECT 6.830 210.300 6.980 217.850 ;
        RECT 7.430 210.300 7.580 217.850 ;
        RECT 8.030 210.300 8.180 217.850 ;
        RECT 8.630 210.300 8.780 217.850 ;
        RECT 9.230 210.300 9.380 217.850 ;
        RECT 9.830 210.300 9.980 217.850 ;
        RECT 14.230 217.550 15.230 218.000 ;
        RECT 10.880 217.400 18.580 217.550 ;
        RECT 14.230 216.950 15.230 217.400 ;
        RECT 10.880 216.800 18.580 216.950 ;
        RECT 14.230 216.350 15.230 216.800 ;
        RECT 10.880 216.200 18.580 216.350 ;
        RECT 14.230 215.750 15.230 216.200 ;
        RECT 10.880 215.600 18.580 215.750 ;
        RECT 14.230 215.150 15.230 215.600 ;
        RECT 10.880 215.000 18.580 215.150 ;
        RECT 14.230 214.550 15.230 215.000 ;
        RECT 10.880 214.400 18.580 214.550 ;
        RECT 14.230 213.950 15.230 214.400 ;
        RECT 10.880 213.800 18.580 213.950 ;
        RECT 14.230 213.350 15.230 213.800 ;
        RECT 10.880 213.200 18.580 213.350 ;
        RECT 14.230 212.750 15.230 213.200 ;
        RECT 10.880 212.600 18.580 212.750 ;
        RECT 14.230 212.150 15.230 212.600 ;
        RECT 10.880 212.000 18.580 212.150 ;
        RECT 14.230 211.550 15.230 212.000 ;
        RECT 10.880 211.400 18.580 211.550 ;
        RECT 14.230 210.950 15.230 211.400 ;
        RECT 10.880 210.800 18.580 210.950 ;
        RECT 14.230 210.300 15.230 210.800 ;
        RECT 19.480 210.300 19.630 217.850 ;
        RECT 20.080 210.300 20.230 217.850 ;
        RECT 20.680 210.300 20.830 217.850 ;
        RECT 21.280 210.300 21.430 217.850 ;
        RECT 21.880 210.300 22.030 217.850 ;
        RECT 22.480 210.300 22.630 217.850 ;
        RECT 22.780 213.200 23.530 215.000 ;
        RECT 25.930 213.200 26.680 215.000 ;
        RECT 22.780 210.450 26.680 213.200 ;
        RECT 22.780 210.300 23.930 210.450 ;
        RECT 5.530 209.700 23.930 210.300 ;
        RECT 5.530 209.550 6.680 209.700 ;
        RECT 4.730 206.800 6.680 209.550 ;
        RECT 5.930 205.050 6.680 206.800 ;
        RECT 6.830 202.150 6.980 209.700 ;
        RECT 7.430 202.150 7.580 209.700 ;
        RECT 8.030 202.150 8.180 209.700 ;
        RECT 8.630 202.150 8.780 209.700 ;
        RECT 9.230 202.150 9.380 209.700 ;
        RECT 9.830 202.150 9.980 209.700 ;
        RECT 14.230 209.200 15.230 209.700 ;
        RECT 10.880 209.050 18.580 209.200 ;
        RECT 14.230 208.600 15.230 209.050 ;
        RECT 10.880 208.450 18.580 208.600 ;
        RECT 14.230 208.000 15.230 208.450 ;
        RECT 10.880 207.850 18.580 208.000 ;
        RECT 14.230 207.400 15.230 207.850 ;
        RECT 10.880 207.250 18.580 207.400 ;
        RECT 14.230 206.800 15.230 207.250 ;
        RECT 10.880 206.650 18.580 206.800 ;
        RECT 14.230 206.200 15.230 206.650 ;
        RECT 10.880 206.050 18.580 206.200 ;
        RECT 14.230 205.600 15.230 206.050 ;
        RECT 10.880 205.450 18.580 205.600 ;
        RECT 14.230 205.000 15.230 205.450 ;
        RECT 10.880 204.850 18.580 205.000 ;
        RECT 14.230 204.400 15.230 204.850 ;
        RECT 10.880 204.250 18.580 204.400 ;
        RECT 14.230 203.800 15.230 204.250 ;
        RECT 10.880 203.650 18.580 203.800 ;
        RECT 14.230 203.200 15.230 203.650 ;
        RECT 10.880 203.050 18.580 203.200 ;
        RECT 14.230 202.600 15.230 203.050 ;
        RECT 10.880 202.450 18.580 202.600 ;
        RECT 14.230 202.000 15.230 202.450 ;
        RECT 19.480 202.150 19.630 209.700 ;
        RECT 20.080 202.150 20.230 209.700 ;
        RECT 20.680 202.150 20.830 209.700 ;
        RECT 21.280 202.150 21.430 209.700 ;
        RECT 21.880 202.150 22.030 209.700 ;
        RECT 22.480 202.150 22.630 209.700 ;
        RECT 22.780 209.550 23.930 209.700 ;
        RECT 24.580 209.550 24.880 210.450 ;
        RECT 25.530 210.300 26.680 210.450 ;
        RECT 26.830 210.300 26.980 217.850 ;
        RECT 27.430 210.300 27.580 217.850 ;
        RECT 28.030 210.300 28.180 217.850 ;
        RECT 28.630 210.300 28.780 217.850 ;
        RECT 29.230 210.300 29.380 217.850 ;
        RECT 29.830 210.300 29.980 217.850 ;
        RECT 34.230 217.550 35.230 218.000 ;
        RECT 30.880 217.400 38.580 217.550 ;
        RECT 34.230 216.950 35.230 217.400 ;
        RECT 30.880 216.800 38.580 216.950 ;
        RECT 34.230 216.350 35.230 216.800 ;
        RECT 30.880 216.200 38.580 216.350 ;
        RECT 34.230 215.750 35.230 216.200 ;
        RECT 30.880 215.600 38.580 215.750 ;
        RECT 34.230 215.150 35.230 215.600 ;
        RECT 30.880 215.000 38.580 215.150 ;
        RECT 34.230 214.550 35.230 215.000 ;
        RECT 30.880 214.400 38.580 214.550 ;
        RECT 34.230 213.950 35.230 214.400 ;
        RECT 30.880 213.800 38.580 213.950 ;
        RECT 34.230 213.350 35.230 213.800 ;
        RECT 30.880 213.200 38.580 213.350 ;
        RECT 34.230 212.750 35.230 213.200 ;
        RECT 30.880 212.600 38.580 212.750 ;
        RECT 34.230 212.150 35.230 212.600 ;
        RECT 30.880 212.000 38.580 212.150 ;
        RECT 34.230 211.550 35.230 212.000 ;
        RECT 30.880 211.400 38.580 211.550 ;
        RECT 34.230 210.950 35.230 211.400 ;
        RECT 30.880 210.800 38.580 210.950 ;
        RECT 34.230 210.300 35.230 210.800 ;
        RECT 39.480 210.300 39.630 217.850 ;
        RECT 40.080 210.300 40.230 217.850 ;
        RECT 40.680 210.300 40.830 217.850 ;
        RECT 41.280 210.300 41.430 217.850 ;
        RECT 41.880 210.300 42.030 217.850 ;
        RECT 42.480 210.300 42.630 217.850 ;
        RECT 42.780 213.200 43.530 215.000 ;
        RECT 45.930 213.200 46.680 215.000 ;
        RECT 42.780 210.450 46.680 213.200 ;
        RECT 42.780 210.300 43.930 210.450 ;
        RECT 25.530 209.700 43.930 210.300 ;
        RECT 25.530 209.550 26.680 209.700 ;
        RECT 22.780 206.800 26.680 209.550 ;
        RECT 22.780 205.050 23.530 206.800 ;
        RECT 25.930 205.050 26.680 206.800 ;
        RECT 26.830 202.150 26.980 209.700 ;
        RECT 27.430 202.150 27.580 209.700 ;
        RECT 28.030 202.150 28.180 209.700 ;
        RECT 28.630 202.150 28.780 209.700 ;
        RECT 29.230 202.150 29.380 209.700 ;
        RECT 29.830 202.150 29.980 209.700 ;
        RECT 34.230 209.200 35.230 209.700 ;
        RECT 30.880 209.050 38.580 209.200 ;
        RECT 34.230 208.600 35.230 209.050 ;
        RECT 30.880 208.450 38.580 208.600 ;
        RECT 34.230 208.000 35.230 208.450 ;
        RECT 30.880 207.850 38.580 208.000 ;
        RECT 34.230 207.400 35.230 207.850 ;
        RECT 30.880 207.250 38.580 207.400 ;
        RECT 34.230 206.800 35.230 207.250 ;
        RECT 30.880 206.650 38.580 206.800 ;
        RECT 34.230 206.200 35.230 206.650 ;
        RECT 30.880 206.050 38.580 206.200 ;
        RECT 34.230 205.600 35.230 206.050 ;
        RECT 30.880 205.450 38.580 205.600 ;
        RECT 34.230 205.000 35.230 205.450 ;
        RECT 30.880 204.850 38.580 205.000 ;
        RECT 34.230 204.400 35.230 204.850 ;
        RECT 30.880 204.250 38.580 204.400 ;
        RECT 34.230 203.800 35.230 204.250 ;
        RECT 30.880 203.650 38.580 203.800 ;
        RECT 34.230 203.200 35.230 203.650 ;
        RECT 30.880 203.050 38.580 203.200 ;
        RECT 34.230 202.600 35.230 203.050 ;
        RECT 30.880 202.450 38.580 202.600 ;
        RECT 34.230 202.000 35.230 202.450 ;
        RECT 39.480 202.150 39.630 209.700 ;
        RECT 40.080 202.150 40.230 209.700 ;
        RECT 40.680 202.150 40.830 209.700 ;
        RECT 41.280 202.150 41.430 209.700 ;
        RECT 41.880 202.150 42.030 209.700 ;
        RECT 42.480 202.150 42.630 209.700 ;
        RECT 42.780 209.550 43.930 209.700 ;
        RECT 44.580 209.550 44.880 210.450 ;
        RECT 45.530 210.300 46.680 210.450 ;
        RECT 46.830 210.300 46.980 217.850 ;
        RECT 47.430 210.300 47.580 217.850 ;
        RECT 48.030 210.300 48.180 217.850 ;
        RECT 48.630 210.300 48.780 217.850 ;
        RECT 49.230 210.300 49.380 217.850 ;
        RECT 49.830 210.300 49.980 217.850 ;
        RECT 54.230 217.550 55.230 218.000 ;
        RECT 50.880 217.400 58.580 217.550 ;
        RECT 54.230 216.950 55.230 217.400 ;
        RECT 50.880 216.800 58.580 216.950 ;
        RECT 54.230 216.350 55.230 216.800 ;
        RECT 50.880 216.200 58.580 216.350 ;
        RECT 54.230 215.750 55.230 216.200 ;
        RECT 50.880 215.600 58.580 215.750 ;
        RECT 54.230 215.150 55.230 215.600 ;
        RECT 50.880 215.000 58.580 215.150 ;
        RECT 54.230 214.550 55.230 215.000 ;
        RECT 50.880 214.400 58.580 214.550 ;
        RECT 54.230 213.950 55.230 214.400 ;
        RECT 50.880 213.800 58.580 213.950 ;
        RECT 54.230 213.350 55.230 213.800 ;
        RECT 50.880 213.200 58.580 213.350 ;
        RECT 54.230 212.750 55.230 213.200 ;
        RECT 50.880 212.600 58.580 212.750 ;
        RECT 54.230 212.150 55.230 212.600 ;
        RECT 50.880 212.000 58.580 212.150 ;
        RECT 54.230 211.550 55.230 212.000 ;
        RECT 50.880 211.400 58.580 211.550 ;
        RECT 54.230 210.950 55.230 211.400 ;
        RECT 50.880 210.800 58.580 210.950 ;
        RECT 54.230 210.300 55.230 210.800 ;
        RECT 59.480 210.300 59.630 217.850 ;
        RECT 60.080 210.300 60.230 217.850 ;
        RECT 60.680 210.300 60.830 217.850 ;
        RECT 61.280 210.300 61.430 217.850 ;
        RECT 61.880 210.300 62.030 217.850 ;
        RECT 62.480 210.300 62.630 217.850 ;
        RECT 62.780 213.200 63.530 215.000 ;
        RECT 65.930 213.200 66.680 215.000 ;
        RECT 62.780 210.450 66.680 213.200 ;
        RECT 62.780 210.300 63.930 210.450 ;
        RECT 45.530 209.700 63.930 210.300 ;
        RECT 45.530 209.550 46.680 209.700 ;
        RECT 42.780 206.800 46.680 209.550 ;
        RECT 42.780 205.050 43.530 206.800 ;
        RECT 45.930 205.050 46.680 206.800 ;
        RECT 46.830 202.150 46.980 209.700 ;
        RECT 47.430 202.150 47.580 209.700 ;
        RECT 48.030 202.150 48.180 209.700 ;
        RECT 48.630 202.150 48.780 209.700 ;
        RECT 49.230 202.150 49.380 209.700 ;
        RECT 49.830 202.150 49.980 209.700 ;
        RECT 54.230 209.200 55.230 209.700 ;
        RECT 50.880 209.050 58.580 209.200 ;
        RECT 54.230 208.600 55.230 209.050 ;
        RECT 50.880 208.450 58.580 208.600 ;
        RECT 54.230 208.000 55.230 208.450 ;
        RECT 50.880 207.850 58.580 208.000 ;
        RECT 54.230 207.400 55.230 207.850 ;
        RECT 50.880 207.250 58.580 207.400 ;
        RECT 54.230 206.800 55.230 207.250 ;
        RECT 50.880 206.650 58.580 206.800 ;
        RECT 54.230 206.200 55.230 206.650 ;
        RECT 50.880 206.050 58.580 206.200 ;
        RECT 54.230 205.600 55.230 206.050 ;
        RECT 50.880 205.450 58.580 205.600 ;
        RECT 54.230 205.000 55.230 205.450 ;
        RECT 50.880 204.850 58.580 205.000 ;
        RECT 54.230 204.400 55.230 204.850 ;
        RECT 50.880 204.250 58.580 204.400 ;
        RECT 54.230 203.800 55.230 204.250 ;
        RECT 50.880 203.650 58.580 203.800 ;
        RECT 54.230 203.200 55.230 203.650 ;
        RECT 50.880 203.050 58.580 203.200 ;
        RECT 54.230 202.600 55.230 203.050 ;
        RECT 50.880 202.450 58.580 202.600 ;
        RECT 54.230 202.000 55.230 202.450 ;
        RECT 59.480 202.150 59.630 209.700 ;
        RECT 60.080 202.150 60.230 209.700 ;
        RECT 60.680 202.150 60.830 209.700 ;
        RECT 61.280 202.150 61.430 209.700 ;
        RECT 61.880 202.150 62.030 209.700 ;
        RECT 62.480 202.150 62.630 209.700 ;
        RECT 62.780 209.550 63.930 209.700 ;
        RECT 64.580 209.550 64.880 210.450 ;
        RECT 65.530 210.300 66.680 210.450 ;
        RECT 66.830 210.300 66.980 217.850 ;
        RECT 67.430 210.300 67.580 217.850 ;
        RECT 68.030 210.300 68.180 217.850 ;
        RECT 68.630 210.300 68.780 217.850 ;
        RECT 69.230 210.300 69.380 217.850 ;
        RECT 69.830 210.300 69.980 217.850 ;
        RECT 74.230 217.550 75.230 218.000 ;
        RECT 70.880 217.400 78.580 217.550 ;
        RECT 74.230 216.950 75.230 217.400 ;
        RECT 70.880 216.800 78.580 216.950 ;
        RECT 74.230 216.350 75.230 216.800 ;
        RECT 70.880 216.200 78.580 216.350 ;
        RECT 74.230 215.750 75.230 216.200 ;
        RECT 70.880 215.600 78.580 215.750 ;
        RECT 74.230 215.150 75.230 215.600 ;
        RECT 70.880 215.000 78.580 215.150 ;
        RECT 74.230 214.550 75.230 215.000 ;
        RECT 70.880 214.400 78.580 214.550 ;
        RECT 74.230 213.950 75.230 214.400 ;
        RECT 70.880 213.800 78.580 213.950 ;
        RECT 74.230 213.350 75.230 213.800 ;
        RECT 70.880 213.200 78.580 213.350 ;
        RECT 74.230 212.750 75.230 213.200 ;
        RECT 70.880 212.600 78.580 212.750 ;
        RECT 74.230 212.150 75.230 212.600 ;
        RECT 70.880 212.000 78.580 212.150 ;
        RECT 74.230 211.550 75.230 212.000 ;
        RECT 70.880 211.400 78.580 211.550 ;
        RECT 74.230 210.950 75.230 211.400 ;
        RECT 70.880 210.800 78.580 210.950 ;
        RECT 74.230 210.300 75.230 210.800 ;
        RECT 79.480 210.300 79.630 217.850 ;
        RECT 80.080 210.300 80.230 217.850 ;
        RECT 80.680 210.300 80.830 217.850 ;
        RECT 81.280 210.300 81.430 217.850 ;
        RECT 81.880 210.300 82.030 217.850 ;
        RECT 82.480 210.300 82.630 217.850 ;
        RECT 82.780 213.200 83.530 215.000 ;
        RECT 85.930 213.200 86.680 215.000 ;
        RECT 82.780 210.450 86.680 213.200 ;
        RECT 82.780 210.300 83.930 210.450 ;
        RECT 65.530 209.700 83.930 210.300 ;
        RECT 65.530 209.550 66.680 209.700 ;
        RECT 62.780 206.800 66.680 209.550 ;
        RECT 62.780 205.050 63.530 206.800 ;
        RECT 65.930 205.050 66.680 206.800 ;
        RECT 66.830 202.150 66.980 209.700 ;
        RECT 67.430 202.150 67.580 209.700 ;
        RECT 68.030 202.150 68.180 209.700 ;
        RECT 68.630 202.150 68.780 209.700 ;
        RECT 69.230 202.150 69.380 209.700 ;
        RECT 69.830 202.150 69.980 209.700 ;
        RECT 74.230 209.200 75.230 209.700 ;
        RECT 70.880 209.050 78.580 209.200 ;
        RECT 74.230 208.600 75.230 209.050 ;
        RECT 70.880 208.450 78.580 208.600 ;
        RECT 74.230 208.000 75.230 208.450 ;
        RECT 70.880 207.850 78.580 208.000 ;
        RECT 74.230 207.400 75.230 207.850 ;
        RECT 70.880 207.250 78.580 207.400 ;
        RECT 74.230 206.800 75.230 207.250 ;
        RECT 70.880 206.650 78.580 206.800 ;
        RECT 74.230 206.200 75.230 206.650 ;
        RECT 70.880 206.050 78.580 206.200 ;
        RECT 74.230 205.600 75.230 206.050 ;
        RECT 70.880 205.450 78.580 205.600 ;
        RECT 74.230 205.000 75.230 205.450 ;
        RECT 70.880 204.850 78.580 205.000 ;
        RECT 74.230 204.400 75.230 204.850 ;
        RECT 70.880 204.250 78.580 204.400 ;
        RECT 74.230 203.800 75.230 204.250 ;
        RECT 70.880 203.650 78.580 203.800 ;
        RECT 74.230 203.200 75.230 203.650 ;
        RECT 70.880 203.050 78.580 203.200 ;
        RECT 74.230 202.600 75.230 203.050 ;
        RECT 70.880 202.450 78.580 202.600 ;
        RECT 74.230 202.000 75.230 202.450 ;
        RECT 79.480 202.150 79.630 209.700 ;
        RECT 80.080 202.150 80.230 209.700 ;
        RECT 80.680 202.150 80.830 209.700 ;
        RECT 81.280 202.150 81.430 209.700 ;
        RECT 81.880 202.150 82.030 209.700 ;
        RECT 82.480 202.150 82.630 209.700 ;
        RECT 82.780 209.550 83.930 209.700 ;
        RECT 84.580 209.550 84.880 210.450 ;
        RECT 85.530 210.300 86.680 210.450 ;
        RECT 86.830 210.300 86.980 217.850 ;
        RECT 87.430 210.300 87.580 217.850 ;
        RECT 88.030 210.300 88.180 217.850 ;
        RECT 88.630 210.300 88.780 217.850 ;
        RECT 89.230 210.300 89.380 217.850 ;
        RECT 89.830 210.300 89.980 217.850 ;
        RECT 94.230 217.550 95.230 218.000 ;
        RECT 90.880 217.400 98.580 217.550 ;
        RECT 94.230 216.950 95.230 217.400 ;
        RECT 90.880 216.800 98.580 216.950 ;
        RECT 94.230 216.350 95.230 216.800 ;
        RECT 90.880 216.200 98.580 216.350 ;
        RECT 94.230 215.750 95.230 216.200 ;
        RECT 90.880 215.600 98.580 215.750 ;
        RECT 94.230 215.150 95.230 215.600 ;
        RECT 90.880 215.000 98.580 215.150 ;
        RECT 94.230 214.550 95.230 215.000 ;
        RECT 90.880 214.400 98.580 214.550 ;
        RECT 94.230 213.950 95.230 214.400 ;
        RECT 90.880 213.800 98.580 213.950 ;
        RECT 94.230 213.350 95.230 213.800 ;
        RECT 90.880 213.200 98.580 213.350 ;
        RECT 94.230 212.750 95.230 213.200 ;
        RECT 90.880 212.600 98.580 212.750 ;
        RECT 94.230 212.150 95.230 212.600 ;
        RECT 90.880 212.000 98.580 212.150 ;
        RECT 94.230 211.550 95.230 212.000 ;
        RECT 90.880 211.400 98.580 211.550 ;
        RECT 94.230 210.950 95.230 211.400 ;
        RECT 90.880 210.800 98.580 210.950 ;
        RECT 94.230 210.300 95.230 210.800 ;
        RECT 99.480 210.300 99.630 217.850 ;
        RECT 100.080 210.300 100.230 217.850 ;
        RECT 100.680 210.300 100.830 217.850 ;
        RECT 101.280 210.300 101.430 217.850 ;
        RECT 101.880 210.300 102.030 217.850 ;
        RECT 102.480 210.300 102.630 217.850 ;
        RECT 102.780 213.200 103.530 215.000 ;
        RECT 105.930 213.200 106.680 215.000 ;
        RECT 102.780 210.450 106.680 213.200 ;
        RECT 102.780 210.300 103.930 210.450 ;
        RECT 85.530 209.700 103.930 210.300 ;
        RECT 85.530 209.550 86.680 209.700 ;
        RECT 82.780 206.800 86.680 209.550 ;
        RECT 82.780 205.050 83.530 206.800 ;
        RECT 85.930 205.050 86.680 206.800 ;
        RECT 86.830 202.150 86.980 209.700 ;
        RECT 87.430 202.150 87.580 209.700 ;
        RECT 88.030 202.150 88.180 209.700 ;
        RECT 88.630 202.150 88.780 209.700 ;
        RECT 89.230 202.150 89.380 209.700 ;
        RECT 89.830 202.150 89.980 209.700 ;
        RECT 94.230 209.200 95.230 209.700 ;
        RECT 90.880 209.050 98.580 209.200 ;
        RECT 94.230 208.600 95.230 209.050 ;
        RECT 90.880 208.450 98.580 208.600 ;
        RECT 94.230 208.000 95.230 208.450 ;
        RECT 90.880 207.850 98.580 208.000 ;
        RECT 94.230 207.400 95.230 207.850 ;
        RECT 90.880 207.250 98.580 207.400 ;
        RECT 94.230 206.800 95.230 207.250 ;
        RECT 90.880 206.650 98.580 206.800 ;
        RECT 94.230 206.200 95.230 206.650 ;
        RECT 90.880 206.050 98.580 206.200 ;
        RECT 94.230 205.600 95.230 206.050 ;
        RECT 90.880 205.450 98.580 205.600 ;
        RECT 94.230 205.000 95.230 205.450 ;
        RECT 90.880 204.850 98.580 205.000 ;
        RECT 94.230 204.400 95.230 204.850 ;
        RECT 90.880 204.250 98.580 204.400 ;
        RECT 94.230 203.800 95.230 204.250 ;
        RECT 90.880 203.650 98.580 203.800 ;
        RECT 94.230 203.200 95.230 203.650 ;
        RECT 90.880 203.050 98.580 203.200 ;
        RECT 94.230 202.600 95.230 203.050 ;
        RECT 90.880 202.450 98.580 202.600 ;
        RECT 94.230 202.000 95.230 202.450 ;
        RECT 99.480 202.150 99.630 209.700 ;
        RECT 100.080 202.150 100.230 209.700 ;
        RECT 100.680 202.150 100.830 209.700 ;
        RECT 101.280 202.150 101.430 209.700 ;
        RECT 101.880 202.150 102.030 209.700 ;
        RECT 102.480 202.150 102.630 209.700 ;
        RECT 102.780 209.550 103.930 209.700 ;
        RECT 104.580 209.550 104.880 210.450 ;
        RECT 105.530 210.300 106.680 210.450 ;
        RECT 106.830 210.300 106.980 217.850 ;
        RECT 107.430 210.300 107.580 217.850 ;
        RECT 108.030 210.300 108.180 217.850 ;
        RECT 108.630 210.300 108.780 217.850 ;
        RECT 109.230 210.300 109.380 217.850 ;
        RECT 109.830 210.300 109.980 217.850 ;
        RECT 114.230 217.550 115.230 218.000 ;
        RECT 110.880 217.400 118.580 217.550 ;
        RECT 114.230 216.950 115.230 217.400 ;
        RECT 110.880 216.800 118.580 216.950 ;
        RECT 114.230 216.350 115.230 216.800 ;
        RECT 110.880 216.200 118.580 216.350 ;
        RECT 114.230 215.750 115.230 216.200 ;
        RECT 110.880 215.600 118.580 215.750 ;
        RECT 114.230 215.150 115.230 215.600 ;
        RECT 110.880 215.000 118.580 215.150 ;
        RECT 114.230 214.550 115.230 215.000 ;
        RECT 110.880 214.400 118.580 214.550 ;
        RECT 114.230 213.950 115.230 214.400 ;
        RECT 110.880 213.800 118.580 213.950 ;
        RECT 114.230 213.350 115.230 213.800 ;
        RECT 110.880 213.200 118.580 213.350 ;
        RECT 114.230 212.750 115.230 213.200 ;
        RECT 110.880 212.600 118.580 212.750 ;
        RECT 114.230 212.150 115.230 212.600 ;
        RECT 110.880 212.000 118.580 212.150 ;
        RECT 114.230 211.550 115.230 212.000 ;
        RECT 110.880 211.400 118.580 211.550 ;
        RECT 114.230 210.950 115.230 211.400 ;
        RECT 110.880 210.800 118.580 210.950 ;
        RECT 114.230 210.300 115.230 210.800 ;
        RECT 119.480 210.300 119.630 217.850 ;
        RECT 120.080 210.300 120.230 217.850 ;
        RECT 120.680 210.300 120.830 217.850 ;
        RECT 121.280 210.300 121.430 217.850 ;
        RECT 121.880 210.300 122.030 217.850 ;
        RECT 122.480 210.300 122.630 217.850 ;
        RECT 122.780 213.200 123.530 215.000 ;
        RECT 122.780 210.450 124.730 213.200 ;
        RECT 122.780 210.300 123.930 210.450 ;
        RECT 105.530 209.700 123.930 210.300 ;
        RECT 105.530 209.550 106.680 209.700 ;
        RECT 102.780 206.800 106.680 209.550 ;
        RECT 102.780 205.050 103.530 206.800 ;
        RECT 105.930 205.050 106.680 206.800 ;
        RECT 106.830 202.150 106.980 209.700 ;
        RECT 107.430 202.150 107.580 209.700 ;
        RECT 108.030 202.150 108.180 209.700 ;
        RECT 108.630 202.150 108.780 209.700 ;
        RECT 109.230 202.150 109.380 209.700 ;
        RECT 109.830 202.150 109.980 209.700 ;
        RECT 114.230 209.200 115.230 209.700 ;
        RECT 110.880 209.050 118.580 209.200 ;
        RECT 114.230 208.600 115.230 209.050 ;
        RECT 110.880 208.450 118.580 208.600 ;
        RECT 114.230 208.000 115.230 208.450 ;
        RECT 110.880 207.850 118.580 208.000 ;
        RECT 114.230 207.400 115.230 207.850 ;
        RECT 110.880 207.250 118.580 207.400 ;
        RECT 114.230 206.800 115.230 207.250 ;
        RECT 110.880 206.650 118.580 206.800 ;
        RECT 114.230 206.200 115.230 206.650 ;
        RECT 110.880 206.050 118.580 206.200 ;
        RECT 114.230 205.600 115.230 206.050 ;
        RECT 110.880 205.450 118.580 205.600 ;
        RECT 114.230 205.000 115.230 205.450 ;
        RECT 110.880 204.850 118.580 205.000 ;
        RECT 114.230 204.400 115.230 204.850 ;
        RECT 110.880 204.250 118.580 204.400 ;
        RECT 114.230 203.800 115.230 204.250 ;
        RECT 110.880 203.650 118.580 203.800 ;
        RECT 114.230 203.200 115.230 203.650 ;
        RECT 110.880 203.050 118.580 203.200 ;
        RECT 114.230 202.600 115.230 203.050 ;
        RECT 110.880 202.450 118.580 202.600 ;
        RECT 114.230 202.000 115.230 202.450 ;
        RECT 119.480 202.150 119.630 209.700 ;
        RECT 120.080 202.150 120.230 209.700 ;
        RECT 120.680 202.150 120.830 209.700 ;
        RECT 121.280 202.150 121.430 209.700 ;
        RECT 121.880 202.150 122.030 209.700 ;
        RECT 122.480 202.150 122.630 209.700 ;
        RECT 122.780 209.550 123.930 209.700 ;
        RECT 124.580 209.625 124.730 210.450 ;
        RECT 124.580 209.550 131.850 209.625 ;
        RECT 122.780 208.350 131.850 209.550 ;
        RECT 122.780 206.800 124.730 208.350 ;
        RECT 122.780 205.050 123.530 206.800 ;
        RECT 10.880 201.850 18.580 202.000 ;
        RECT 30.880 201.850 38.580 202.000 ;
        RECT 50.880 201.850 58.580 202.000 ;
        RECT 70.880 201.850 78.580 202.000 ;
        RECT 90.880 201.850 98.580 202.000 ;
        RECT 110.880 201.850 118.580 202.000 ;
        RECT 14.230 201.200 15.230 201.850 ;
        RECT 34.230 201.200 35.230 201.850 ;
        RECT 54.230 201.200 55.230 201.850 ;
        RECT 74.230 201.200 75.230 201.850 ;
        RECT 94.230 201.200 95.230 201.850 ;
        RECT 114.230 201.200 115.230 201.850 ;
        RECT 11.530 200.000 17.930 201.200 ;
        RECT 31.530 200.000 37.930 201.200 ;
        RECT 51.530 200.000 57.930 201.200 ;
        RECT 71.530 200.000 77.930 201.200 ;
        RECT 91.530 200.000 97.930 201.200 ;
        RECT 111.530 200.000 117.930 201.200 ;
        RECT 9.340 176.350 11.675 177.050 ;
        RECT 10.110 174.410 11.985 174.770 ;
        RECT 12.335 174.415 14.215 174.775 ;
        RECT 11.530 138.800 17.930 140.000 ;
        RECT 31.530 138.800 37.930 140.000 ;
        RECT 51.530 138.800 57.930 140.000 ;
        RECT 71.530 138.800 77.930 140.000 ;
        RECT 91.530 138.800 97.930 140.000 ;
        RECT 111.530 138.800 117.930 140.000 ;
        RECT 14.230 138.150 15.230 138.800 ;
        RECT 34.230 138.150 35.230 138.800 ;
        RECT 54.230 138.150 55.230 138.800 ;
        RECT 74.230 138.150 75.230 138.800 ;
        RECT 94.230 138.150 95.230 138.800 ;
        RECT 114.230 138.150 115.230 138.800 ;
        RECT 10.880 138.000 18.580 138.150 ;
        RECT 30.880 138.000 38.580 138.150 ;
        RECT 50.880 138.000 58.580 138.150 ;
        RECT 70.880 138.000 78.580 138.150 ;
        RECT 90.880 138.000 98.580 138.150 ;
        RECT 110.880 138.000 118.580 138.150 ;
        RECT 5.930 133.200 6.680 135.000 ;
        RECT 4.730 130.450 6.680 133.200 ;
        RECT 4.730 129.550 4.880 130.450 ;
        RECT 5.530 130.300 6.680 130.450 ;
        RECT 6.830 130.300 6.980 137.850 ;
        RECT 7.430 130.300 7.580 137.850 ;
        RECT 8.030 130.300 8.180 137.850 ;
        RECT 8.630 130.300 8.780 137.850 ;
        RECT 9.230 130.300 9.380 137.850 ;
        RECT 9.830 130.300 9.980 137.850 ;
        RECT 14.230 137.550 15.230 138.000 ;
        RECT 10.880 137.400 18.580 137.550 ;
        RECT 14.230 136.950 15.230 137.400 ;
        RECT 10.880 136.800 18.580 136.950 ;
        RECT 14.230 136.350 15.230 136.800 ;
        RECT 10.880 136.200 18.580 136.350 ;
        RECT 14.230 135.750 15.230 136.200 ;
        RECT 10.880 135.600 18.580 135.750 ;
        RECT 14.230 135.150 15.230 135.600 ;
        RECT 10.880 135.000 18.580 135.150 ;
        RECT 14.230 134.550 15.230 135.000 ;
        RECT 10.880 134.400 18.580 134.550 ;
        RECT 14.230 133.950 15.230 134.400 ;
        RECT 10.880 133.800 18.580 133.950 ;
        RECT 14.230 133.350 15.230 133.800 ;
        RECT 10.880 133.200 18.580 133.350 ;
        RECT 14.230 132.750 15.230 133.200 ;
        RECT 10.880 132.600 18.580 132.750 ;
        RECT 14.230 132.150 15.230 132.600 ;
        RECT 10.880 132.000 18.580 132.150 ;
        RECT 14.230 131.550 15.230 132.000 ;
        RECT 10.880 131.400 18.580 131.550 ;
        RECT 14.230 130.950 15.230 131.400 ;
        RECT 10.880 130.800 18.580 130.950 ;
        RECT 14.230 130.300 15.230 130.800 ;
        RECT 19.480 130.300 19.630 137.850 ;
        RECT 20.080 130.300 20.230 137.850 ;
        RECT 20.680 130.300 20.830 137.850 ;
        RECT 21.280 130.300 21.430 137.850 ;
        RECT 21.880 130.300 22.030 137.850 ;
        RECT 22.480 130.300 22.630 137.850 ;
        RECT 22.780 133.200 23.530 135.000 ;
        RECT 25.930 133.200 26.680 135.000 ;
        RECT 22.780 130.450 26.680 133.200 ;
        RECT 22.780 130.300 23.930 130.450 ;
        RECT 5.530 129.700 23.930 130.300 ;
        RECT 5.530 129.550 6.680 129.700 ;
        RECT 4.730 126.800 6.680 129.550 ;
        RECT 5.930 125.050 6.680 126.800 ;
        RECT 6.830 122.150 6.980 129.700 ;
        RECT 7.430 122.150 7.580 129.700 ;
        RECT 8.030 122.150 8.180 129.700 ;
        RECT 8.630 122.150 8.780 129.700 ;
        RECT 9.230 122.150 9.380 129.700 ;
        RECT 9.830 122.150 9.980 129.700 ;
        RECT 14.230 129.200 15.230 129.700 ;
        RECT 10.880 129.050 18.580 129.200 ;
        RECT 14.230 128.600 15.230 129.050 ;
        RECT 10.880 128.450 18.580 128.600 ;
        RECT 14.230 128.000 15.230 128.450 ;
        RECT 10.880 127.850 18.580 128.000 ;
        RECT 14.230 127.400 15.230 127.850 ;
        RECT 10.880 127.250 18.580 127.400 ;
        RECT 14.230 126.800 15.230 127.250 ;
        RECT 10.880 126.650 18.580 126.800 ;
        RECT 14.230 126.200 15.230 126.650 ;
        RECT 10.880 126.050 18.580 126.200 ;
        RECT 14.230 125.600 15.230 126.050 ;
        RECT 10.880 125.450 18.580 125.600 ;
        RECT 14.230 125.000 15.230 125.450 ;
        RECT 10.880 124.850 18.580 125.000 ;
        RECT 14.230 124.400 15.230 124.850 ;
        RECT 10.880 124.250 18.580 124.400 ;
        RECT 14.230 123.800 15.230 124.250 ;
        RECT 10.880 123.650 18.580 123.800 ;
        RECT 14.230 123.200 15.230 123.650 ;
        RECT 10.880 123.050 18.580 123.200 ;
        RECT 14.230 122.600 15.230 123.050 ;
        RECT 10.880 122.450 18.580 122.600 ;
        RECT 14.230 122.000 15.230 122.450 ;
        RECT 19.480 122.150 19.630 129.700 ;
        RECT 20.080 122.150 20.230 129.700 ;
        RECT 20.680 122.150 20.830 129.700 ;
        RECT 21.280 122.150 21.430 129.700 ;
        RECT 21.880 122.150 22.030 129.700 ;
        RECT 22.480 122.150 22.630 129.700 ;
        RECT 22.780 129.550 23.930 129.700 ;
        RECT 24.580 129.550 24.880 130.450 ;
        RECT 25.530 130.300 26.680 130.450 ;
        RECT 26.830 130.300 26.980 137.850 ;
        RECT 27.430 130.300 27.580 137.850 ;
        RECT 28.030 130.300 28.180 137.850 ;
        RECT 28.630 130.300 28.780 137.850 ;
        RECT 29.230 130.300 29.380 137.850 ;
        RECT 29.830 130.300 29.980 137.850 ;
        RECT 34.230 137.550 35.230 138.000 ;
        RECT 30.880 137.400 38.580 137.550 ;
        RECT 34.230 136.950 35.230 137.400 ;
        RECT 30.880 136.800 38.580 136.950 ;
        RECT 34.230 136.350 35.230 136.800 ;
        RECT 30.880 136.200 38.580 136.350 ;
        RECT 34.230 135.750 35.230 136.200 ;
        RECT 30.880 135.600 38.580 135.750 ;
        RECT 34.230 135.150 35.230 135.600 ;
        RECT 30.880 135.000 38.580 135.150 ;
        RECT 34.230 134.550 35.230 135.000 ;
        RECT 30.880 134.400 38.580 134.550 ;
        RECT 34.230 133.950 35.230 134.400 ;
        RECT 30.880 133.800 38.580 133.950 ;
        RECT 34.230 133.350 35.230 133.800 ;
        RECT 30.880 133.200 38.580 133.350 ;
        RECT 34.230 132.750 35.230 133.200 ;
        RECT 30.880 132.600 38.580 132.750 ;
        RECT 34.230 132.150 35.230 132.600 ;
        RECT 30.880 132.000 38.580 132.150 ;
        RECT 34.230 131.550 35.230 132.000 ;
        RECT 30.880 131.400 38.580 131.550 ;
        RECT 34.230 130.950 35.230 131.400 ;
        RECT 30.880 130.800 38.580 130.950 ;
        RECT 34.230 130.300 35.230 130.800 ;
        RECT 39.480 130.300 39.630 137.850 ;
        RECT 40.080 130.300 40.230 137.850 ;
        RECT 40.680 130.300 40.830 137.850 ;
        RECT 41.280 130.300 41.430 137.850 ;
        RECT 41.880 130.300 42.030 137.850 ;
        RECT 42.480 130.300 42.630 137.850 ;
        RECT 42.780 133.200 43.530 135.000 ;
        RECT 45.930 133.200 46.680 135.000 ;
        RECT 42.780 130.450 46.680 133.200 ;
        RECT 42.780 130.300 43.930 130.450 ;
        RECT 25.530 129.700 43.930 130.300 ;
        RECT 25.530 129.550 26.680 129.700 ;
        RECT 22.780 126.800 26.680 129.550 ;
        RECT 22.780 125.050 23.530 126.800 ;
        RECT 25.930 125.050 26.680 126.800 ;
        RECT 26.830 122.150 26.980 129.700 ;
        RECT 27.430 122.150 27.580 129.700 ;
        RECT 28.030 122.150 28.180 129.700 ;
        RECT 28.630 122.150 28.780 129.700 ;
        RECT 29.230 122.150 29.380 129.700 ;
        RECT 29.830 122.150 29.980 129.700 ;
        RECT 34.230 129.200 35.230 129.700 ;
        RECT 30.880 129.050 38.580 129.200 ;
        RECT 34.230 128.600 35.230 129.050 ;
        RECT 30.880 128.450 38.580 128.600 ;
        RECT 34.230 128.000 35.230 128.450 ;
        RECT 30.880 127.850 38.580 128.000 ;
        RECT 34.230 127.400 35.230 127.850 ;
        RECT 30.880 127.250 38.580 127.400 ;
        RECT 34.230 126.800 35.230 127.250 ;
        RECT 30.880 126.650 38.580 126.800 ;
        RECT 34.230 126.200 35.230 126.650 ;
        RECT 30.880 126.050 38.580 126.200 ;
        RECT 34.230 125.600 35.230 126.050 ;
        RECT 30.880 125.450 38.580 125.600 ;
        RECT 34.230 125.000 35.230 125.450 ;
        RECT 30.880 124.850 38.580 125.000 ;
        RECT 34.230 124.400 35.230 124.850 ;
        RECT 30.880 124.250 38.580 124.400 ;
        RECT 34.230 123.800 35.230 124.250 ;
        RECT 30.880 123.650 38.580 123.800 ;
        RECT 34.230 123.200 35.230 123.650 ;
        RECT 30.880 123.050 38.580 123.200 ;
        RECT 34.230 122.600 35.230 123.050 ;
        RECT 30.880 122.450 38.580 122.600 ;
        RECT 34.230 122.000 35.230 122.450 ;
        RECT 39.480 122.150 39.630 129.700 ;
        RECT 40.080 122.150 40.230 129.700 ;
        RECT 40.680 122.150 40.830 129.700 ;
        RECT 41.280 122.150 41.430 129.700 ;
        RECT 41.880 122.150 42.030 129.700 ;
        RECT 42.480 122.150 42.630 129.700 ;
        RECT 42.780 129.550 43.930 129.700 ;
        RECT 44.580 129.550 44.880 130.450 ;
        RECT 45.530 130.300 46.680 130.450 ;
        RECT 46.830 130.300 46.980 137.850 ;
        RECT 47.430 130.300 47.580 137.850 ;
        RECT 48.030 130.300 48.180 137.850 ;
        RECT 48.630 130.300 48.780 137.850 ;
        RECT 49.230 130.300 49.380 137.850 ;
        RECT 49.830 130.300 49.980 137.850 ;
        RECT 54.230 137.550 55.230 138.000 ;
        RECT 50.880 137.400 58.580 137.550 ;
        RECT 54.230 136.950 55.230 137.400 ;
        RECT 50.880 136.800 58.580 136.950 ;
        RECT 54.230 136.350 55.230 136.800 ;
        RECT 50.880 136.200 58.580 136.350 ;
        RECT 54.230 135.750 55.230 136.200 ;
        RECT 50.880 135.600 58.580 135.750 ;
        RECT 54.230 135.150 55.230 135.600 ;
        RECT 50.880 135.000 58.580 135.150 ;
        RECT 54.230 134.550 55.230 135.000 ;
        RECT 50.880 134.400 58.580 134.550 ;
        RECT 54.230 133.950 55.230 134.400 ;
        RECT 50.880 133.800 58.580 133.950 ;
        RECT 54.230 133.350 55.230 133.800 ;
        RECT 50.880 133.200 58.580 133.350 ;
        RECT 54.230 132.750 55.230 133.200 ;
        RECT 50.880 132.600 58.580 132.750 ;
        RECT 54.230 132.150 55.230 132.600 ;
        RECT 50.880 132.000 58.580 132.150 ;
        RECT 54.230 131.550 55.230 132.000 ;
        RECT 50.880 131.400 58.580 131.550 ;
        RECT 54.230 130.950 55.230 131.400 ;
        RECT 50.880 130.800 58.580 130.950 ;
        RECT 54.230 130.300 55.230 130.800 ;
        RECT 59.480 130.300 59.630 137.850 ;
        RECT 60.080 130.300 60.230 137.850 ;
        RECT 60.680 130.300 60.830 137.850 ;
        RECT 61.280 130.300 61.430 137.850 ;
        RECT 61.880 130.300 62.030 137.850 ;
        RECT 62.480 130.300 62.630 137.850 ;
        RECT 62.780 133.200 63.530 135.000 ;
        RECT 65.930 133.200 66.680 135.000 ;
        RECT 62.780 130.450 66.680 133.200 ;
        RECT 62.780 130.300 63.930 130.450 ;
        RECT 45.530 129.700 63.930 130.300 ;
        RECT 45.530 129.550 46.680 129.700 ;
        RECT 42.780 126.800 46.680 129.550 ;
        RECT 42.780 125.050 43.530 126.800 ;
        RECT 45.930 125.050 46.680 126.800 ;
        RECT 46.830 122.150 46.980 129.700 ;
        RECT 47.430 122.150 47.580 129.700 ;
        RECT 48.030 122.150 48.180 129.700 ;
        RECT 48.630 122.150 48.780 129.700 ;
        RECT 49.230 122.150 49.380 129.700 ;
        RECT 49.830 122.150 49.980 129.700 ;
        RECT 54.230 129.200 55.230 129.700 ;
        RECT 50.880 129.050 58.580 129.200 ;
        RECT 54.230 128.600 55.230 129.050 ;
        RECT 50.880 128.450 58.580 128.600 ;
        RECT 54.230 128.000 55.230 128.450 ;
        RECT 50.880 127.850 58.580 128.000 ;
        RECT 54.230 127.400 55.230 127.850 ;
        RECT 50.880 127.250 58.580 127.400 ;
        RECT 54.230 126.800 55.230 127.250 ;
        RECT 50.880 126.650 58.580 126.800 ;
        RECT 54.230 126.200 55.230 126.650 ;
        RECT 50.880 126.050 58.580 126.200 ;
        RECT 54.230 125.600 55.230 126.050 ;
        RECT 50.880 125.450 58.580 125.600 ;
        RECT 54.230 125.000 55.230 125.450 ;
        RECT 50.880 124.850 58.580 125.000 ;
        RECT 54.230 124.400 55.230 124.850 ;
        RECT 50.880 124.250 58.580 124.400 ;
        RECT 54.230 123.800 55.230 124.250 ;
        RECT 50.880 123.650 58.580 123.800 ;
        RECT 54.230 123.200 55.230 123.650 ;
        RECT 50.880 123.050 58.580 123.200 ;
        RECT 54.230 122.600 55.230 123.050 ;
        RECT 50.880 122.450 58.580 122.600 ;
        RECT 54.230 122.000 55.230 122.450 ;
        RECT 59.480 122.150 59.630 129.700 ;
        RECT 60.080 122.150 60.230 129.700 ;
        RECT 60.680 122.150 60.830 129.700 ;
        RECT 61.280 122.150 61.430 129.700 ;
        RECT 61.880 122.150 62.030 129.700 ;
        RECT 62.480 122.150 62.630 129.700 ;
        RECT 62.780 129.550 63.930 129.700 ;
        RECT 64.580 129.550 64.880 130.450 ;
        RECT 65.530 130.300 66.680 130.450 ;
        RECT 66.830 130.300 66.980 137.850 ;
        RECT 67.430 130.300 67.580 137.850 ;
        RECT 68.030 130.300 68.180 137.850 ;
        RECT 68.630 130.300 68.780 137.850 ;
        RECT 69.230 130.300 69.380 137.850 ;
        RECT 69.830 130.300 69.980 137.850 ;
        RECT 74.230 137.550 75.230 138.000 ;
        RECT 70.880 137.400 78.580 137.550 ;
        RECT 74.230 136.950 75.230 137.400 ;
        RECT 70.880 136.800 78.580 136.950 ;
        RECT 74.230 136.350 75.230 136.800 ;
        RECT 70.880 136.200 78.580 136.350 ;
        RECT 74.230 135.750 75.230 136.200 ;
        RECT 70.880 135.600 78.580 135.750 ;
        RECT 74.230 135.150 75.230 135.600 ;
        RECT 70.880 135.000 78.580 135.150 ;
        RECT 74.230 134.550 75.230 135.000 ;
        RECT 70.880 134.400 78.580 134.550 ;
        RECT 74.230 133.950 75.230 134.400 ;
        RECT 70.880 133.800 78.580 133.950 ;
        RECT 74.230 133.350 75.230 133.800 ;
        RECT 70.880 133.200 78.580 133.350 ;
        RECT 74.230 132.750 75.230 133.200 ;
        RECT 70.880 132.600 78.580 132.750 ;
        RECT 74.230 132.150 75.230 132.600 ;
        RECT 70.880 132.000 78.580 132.150 ;
        RECT 74.230 131.550 75.230 132.000 ;
        RECT 70.880 131.400 78.580 131.550 ;
        RECT 74.230 130.950 75.230 131.400 ;
        RECT 70.880 130.800 78.580 130.950 ;
        RECT 74.230 130.300 75.230 130.800 ;
        RECT 79.480 130.300 79.630 137.850 ;
        RECT 80.080 130.300 80.230 137.850 ;
        RECT 80.680 130.300 80.830 137.850 ;
        RECT 81.280 130.300 81.430 137.850 ;
        RECT 81.880 130.300 82.030 137.850 ;
        RECT 82.480 130.300 82.630 137.850 ;
        RECT 82.780 133.200 83.530 135.000 ;
        RECT 85.930 133.200 86.680 135.000 ;
        RECT 82.780 130.450 86.680 133.200 ;
        RECT 82.780 130.300 83.930 130.450 ;
        RECT 65.530 129.700 83.930 130.300 ;
        RECT 65.530 129.550 66.680 129.700 ;
        RECT 62.780 126.800 66.680 129.550 ;
        RECT 62.780 125.050 63.530 126.800 ;
        RECT 65.930 125.050 66.680 126.800 ;
        RECT 66.830 122.150 66.980 129.700 ;
        RECT 67.430 122.150 67.580 129.700 ;
        RECT 68.030 122.150 68.180 129.700 ;
        RECT 68.630 122.150 68.780 129.700 ;
        RECT 69.230 122.150 69.380 129.700 ;
        RECT 69.830 122.150 69.980 129.700 ;
        RECT 74.230 129.200 75.230 129.700 ;
        RECT 70.880 129.050 78.580 129.200 ;
        RECT 74.230 128.600 75.230 129.050 ;
        RECT 70.880 128.450 78.580 128.600 ;
        RECT 74.230 128.000 75.230 128.450 ;
        RECT 70.880 127.850 78.580 128.000 ;
        RECT 74.230 127.400 75.230 127.850 ;
        RECT 70.880 127.250 78.580 127.400 ;
        RECT 74.230 126.800 75.230 127.250 ;
        RECT 70.880 126.650 78.580 126.800 ;
        RECT 74.230 126.200 75.230 126.650 ;
        RECT 70.880 126.050 78.580 126.200 ;
        RECT 74.230 125.600 75.230 126.050 ;
        RECT 70.880 125.450 78.580 125.600 ;
        RECT 74.230 125.000 75.230 125.450 ;
        RECT 70.880 124.850 78.580 125.000 ;
        RECT 74.230 124.400 75.230 124.850 ;
        RECT 70.880 124.250 78.580 124.400 ;
        RECT 74.230 123.800 75.230 124.250 ;
        RECT 70.880 123.650 78.580 123.800 ;
        RECT 74.230 123.200 75.230 123.650 ;
        RECT 70.880 123.050 78.580 123.200 ;
        RECT 74.230 122.600 75.230 123.050 ;
        RECT 70.880 122.450 78.580 122.600 ;
        RECT 74.230 122.000 75.230 122.450 ;
        RECT 79.480 122.150 79.630 129.700 ;
        RECT 80.080 122.150 80.230 129.700 ;
        RECT 80.680 122.150 80.830 129.700 ;
        RECT 81.280 122.150 81.430 129.700 ;
        RECT 81.880 122.150 82.030 129.700 ;
        RECT 82.480 122.150 82.630 129.700 ;
        RECT 82.780 129.550 83.930 129.700 ;
        RECT 84.580 129.550 84.880 130.450 ;
        RECT 85.530 130.300 86.680 130.450 ;
        RECT 86.830 130.300 86.980 137.850 ;
        RECT 87.430 130.300 87.580 137.850 ;
        RECT 88.030 130.300 88.180 137.850 ;
        RECT 88.630 130.300 88.780 137.850 ;
        RECT 89.230 130.300 89.380 137.850 ;
        RECT 89.830 130.300 89.980 137.850 ;
        RECT 94.230 137.550 95.230 138.000 ;
        RECT 90.880 137.400 98.580 137.550 ;
        RECT 94.230 136.950 95.230 137.400 ;
        RECT 90.880 136.800 98.580 136.950 ;
        RECT 94.230 136.350 95.230 136.800 ;
        RECT 90.880 136.200 98.580 136.350 ;
        RECT 94.230 135.750 95.230 136.200 ;
        RECT 90.880 135.600 98.580 135.750 ;
        RECT 94.230 135.150 95.230 135.600 ;
        RECT 90.880 135.000 98.580 135.150 ;
        RECT 94.230 134.550 95.230 135.000 ;
        RECT 90.880 134.400 98.580 134.550 ;
        RECT 94.230 133.950 95.230 134.400 ;
        RECT 90.880 133.800 98.580 133.950 ;
        RECT 94.230 133.350 95.230 133.800 ;
        RECT 90.880 133.200 98.580 133.350 ;
        RECT 94.230 132.750 95.230 133.200 ;
        RECT 90.880 132.600 98.580 132.750 ;
        RECT 94.230 132.150 95.230 132.600 ;
        RECT 90.880 132.000 98.580 132.150 ;
        RECT 94.230 131.550 95.230 132.000 ;
        RECT 90.880 131.400 98.580 131.550 ;
        RECT 94.230 130.950 95.230 131.400 ;
        RECT 90.880 130.800 98.580 130.950 ;
        RECT 94.230 130.300 95.230 130.800 ;
        RECT 99.480 130.300 99.630 137.850 ;
        RECT 100.080 130.300 100.230 137.850 ;
        RECT 100.680 130.300 100.830 137.850 ;
        RECT 101.280 130.300 101.430 137.850 ;
        RECT 101.880 130.300 102.030 137.850 ;
        RECT 102.480 130.300 102.630 137.850 ;
        RECT 102.780 133.200 103.530 135.000 ;
        RECT 105.930 133.200 106.680 135.000 ;
        RECT 102.780 130.450 106.680 133.200 ;
        RECT 102.780 130.300 103.930 130.450 ;
        RECT 85.530 129.700 103.930 130.300 ;
        RECT 85.530 129.550 86.680 129.700 ;
        RECT 82.780 126.800 86.680 129.550 ;
        RECT 82.780 125.050 83.530 126.800 ;
        RECT 85.930 125.050 86.680 126.800 ;
        RECT 86.830 122.150 86.980 129.700 ;
        RECT 87.430 122.150 87.580 129.700 ;
        RECT 88.030 122.150 88.180 129.700 ;
        RECT 88.630 122.150 88.780 129.700 ;
        RECT 89.230 122.150 89.380 129.700 ;
        RECT 89.830 122.150 89.980 129.700 ;
        RECT 94.230 129.200 95.230 129.700 ;
        RECT 90.880 129.050 98.580 129.200 ;
        RECT 94.230 128.600 95.230 129.050 ;
        RECT 90.880 128.450 98.580 128.600 ;
        RECT 94.230 128.000 95.230 128.450 ;
        RECT 90.880 127.850 98.580 128.000 ;
        RECT 94.230 127.400 95.230 127.850 ;
        RECT 90.880 127.250 98.580 127.400 ;
        RECT 94.230 126.800 95.230 127.250 ;
        RECT 90.880 126.650 98.580 126.800 ;
        RECT 94.230 126.200 95.230 126.650 ;
        RECT 90.880 126.050 98.580 126.200 ;
        RECT 94.230 125.600 95.230 126.050 ;
        RECT 90.880 125.450 98.580 125.600 ;
        RECT 94.230 125.000 95.230 125.450 ;
        RECT 90.880 124.850 98.580 125.000 ;
        RECT 94.230 124.400 95.230 124.850 ;
        RECT 90.880 124.250 98.580 124.400 ;
        RECT 94.230 123.800 95.230 124.250 ;
        RECT 90.880 123.650 98.580 123.800 ;
        RECT 94.230 123.200 95.230 123.650 ;
        RECT 90.880 123.050 98.580 123.200 ;
        RECT 94.230 122.600 95.230 123.050 ;
        RECT 90.880 122.450 98.580 122.600 ;
        RECT 94.230 122.000 95.230 122.450 ;
        RECT 99.480 122.150 99.630 129.700 ;
        RECT 100.080 122.150 100.230 129.700 ;
        RECT 100.680 122.150 100.830 129.700 ;
        RECT 101.280 122.150 101.430 129.700 ;
        RECT 101.880 122.150 102.030 129.700 ;
        RECT 102.480 122.150 102.630 129.700 ;
        RECT 102.780 129.550 103.930 129.700 ;
        RECT 104.580 129.550 104.880 130.450 ;
        RECT 105.530 130.300 106.680 130.450 ;
        RECT 106.830 130.300 106.980 137.850 ;
        RECT 107.430 130.300 107.580 137.850 ;
        RECT 108.030 130.300 108.180 137.850 ;
        RECT 108.630 130.300 108.780 137.850 ;
        RECT 109.230 130.300 109.380 137.850 ;
        RECT 109.830 130.300 109.980 137.850 ;
        RECT 114.230 137.550 115.230 138.000 ;
        RECT 110.880 137.400 118.580 137.550 ;
        RECT 114.230 136.950 115.230 137.400 ;
        RECT 110.880 136.800 118.580 136.950 ;
        RECT 114.230 136.350 115.230 136.800 ;
        RECT 110.880 136.200 118.580 136.350 ;
        RECT 114.230 135.750 115.230 136.200 ;
        RECT 110.880 135.600 118.580 135.750 ;
        RECT 114.230 135.150 115.230 135.600 ;
        RECT 110.880 135.000 118.580 135.150 ;
        RECT 114.230 134.550 115.230 135.000 ;
        RECT 110.880 134.400 118.580 134.550 ;
        RECT 114.230 133.950 115.230 134.400 ;
        RECT 110.880 133.800 118.580 133.950 ;
        RECT 114.230 133.350 115.230 133.800 ;
        RECT 110.880 133.200 118.580 133.350 ;
        RECT 114.230 132.750 115.230 133.200 ;
        RECT 110.880 132.600 118.580 132.750 ;
        RECT 114.230 132.150 115.230 132.600 ;
        RECT 110.880 132.000 118.580 132.150 ;
        RECT 114.230 131.550 115.230 132.000 ;
        RECT 110.880 131.400 118.580 131.550 ;
        RECT 114.230 130.950 115.230 131.400 ;
        RECT 110.880 130.800 118.580 130.950 ;
        RECT 114.230 130.300 115.230 130.800 ;
        RECT 119.480 130.300 119.630 137.850 ;
        RECT 120.080 130.300 120.230 137.850 ;
        RECT 120.680 130.300 120.830 137.850 ;
        RECT 121.280 130.300 121.430 137.850 ;
        RECT 121.880 130.300 122.030 137.850 ;
        RECT 122.480 130.300 122.630 137.850 ;
        RECT 122.780 133.200 123.530 135.000 ;
        RECT 122.780 130.775 124.730 133.200 ;
        RECT 122.780 130.450 131.850 130.775 ;
        RECT 122.780 130.300 123.930 130.450 ;
        RECT 105.530 129.700 123.930 130.300 ;
        RECT 105.530 129.550 106.680 129.700 ;
        RECT 102.780 126.800 106.680 129.550 ;
        RECT 102.780 125.050 103.530 126.800 ;
        RECT 105.930 125.050 106.680 126.800 ;
        RECT 106.830 122.150 106.980 129.700 ;
        RECT 107.430 122.150 107.580 129.700 ;
        RECT 108.030 122.150 108.180 129.700 ;
        RECT 108.630 122.150 108.780 129.700 ;
        RECT 109.230 122.150 109.380 129.700 ;
        RECT 109.830 122.150 109.980 129.700 ;
        RECT 114.230 129.200 115.230 129.700 ;
        RECT 110.880 129.050 118.580 129.200 ;
        RECT 114.230 128.600 115.230 129.050 ;
        RECT 110.880 128.450 118.580 128.600 ;
        RECT 114.230 128.000 115.230 128.450 ;
        RECT 110.880 127.850 118.580 128.000 ;
        RECT 114.230 127.400 115.230 127.850 ;
        RECT 110.880 127.250 118.580 127.400 ;
        RECT 114.230 126.800 115.230 127.250 ;
        RECT 110.880 126.650 118.580 126.800 ;
        RECT 114.230 126.200 115.230 126.650 ;
        RECT 110.880 126.050 118.580 126.200 ;
        RECT 114.230 125.600 115.230 126.050 ;
        RECT 110.880 125.450 118.580 125.600 ;
        RECT 114.230 125.000 115.230 125.450 ;
        RECT 110.880 124.850 118.580 125.000 ;
        RECT 114.230 124.400 115.230 124.850 ;
        RECT 110.880 124.250 118.580 124.400 ;
        RECT 114.230 123.800 115.230 124.250 ;
        RECT 110.880 123.650 118.580 123.800 ;
        RECT 114.230 123.200 115.230 123.650 ;
        RECT 110.880 123.050 118.580 123.200 ;
        RECT 114.230 122.600 115.230 123.050 ;
        RECT 110.880 122.450 118.580 122.600 ;
        RECT 114.230 122.000 115.230 122.450 ;
        RECT 119.480 122.150 119.630 129.700 ;
        RECT 120.080 122.150 120.230 129.700 ;
        RECT 120.680 122.150 120.830 129.700 ;
        RECT 121.280 122.150 121.430 129.700 ;
        RECT 121.880 122.150 122.030 129.700 ;
        RECT 122.480 122.150 122.630 129.700 ;
        RECT 122.780 129.550 123.930 129.700 ;
        RECT 124.580 129.550 131.850 130.450 ;
        RECT 122.780 129.500 131.850 129.550 ;
        RECT 122.780 126.800 124.730 129.500 ;
        RECT 122.780 125.050 123.530 126.800 ;
        RECT 10.880 121.850 18.580 122.000 ;
        RECT 30.880 121.850 38.580 122.000 ;
        RECT 50.880 121.850 58.580 122.000 ;
        RECT 70.880 121.850 78.580 122.000 ;
        RECT 90.880 121.850 98.580 122.000 ;
        RECT 110.880 121.850 118.580 122.000 ;
        RECT 14.230 121.200 15.230 121.850 ;
        RECT 34.230 121.200 35.230 121.850 ;
        RECT 54.230 121.200 55.230 121.850 ;
        RECT 74.230 121.200 75.230 121.850 ;
        RECT 94.230 121.200 95.230 121.850 ;
        RECT 114.230 121.200 115.230 121.850 ;
        RECT 11.530 118.800 17.930 121.200 ;
        RECT 31.530 118.800 37.930 121.200 ;
        RECT 51.530 118.800 57.930 121.200 ;
        RECT 71.530 118.800 77.930 121.200 ;
        RECT 91.530 118.800 97.930 121.200 ;
        RECT 111.530 118.800 117.930 121.200 ;
        RECT 14.230 118.150 15.230 118.800 ;
        RECT 34.230 118.150 35.230 118.800 ;
        RECT 54.230 118.150 55.230 118.800 ;
        RECT 74.230 118.150 75.230 118.800 ;
        RECT 94.230 118.150 95.230 118.800 ;
        RECT 114.230 118.150 115.230 118.800 ;
        RECT 10.880 118.000 18.580 118.150 ;
        RECT 30.880 118.000 38.580 118.150 ;
        RECT 50.880 118.000 58.580 118.150 ;
        RECT 70.880 118.000 78.580 118.150 ;
        RECT 90.880 118.000 98.580 118.150 ;
        RECT 110.880 118.000 118.580 118.150 ;
        RECT 5.930 113.200 6.680 115.000 ;
        RECT 4.730 110.450 6.680 113.200 ;
        RECT 4.730 109.550 4.880 110.450 ;
        RECT 5.530 110.300 6.680 110.450 ;
        RECT 6.830 110.300 6.980 117.850 ;
        RECT 7.430 110.300 7.580 117.850 ;
        RECT 8.030 110.300 8.180 117.850 ;
        RECT 8.630 110.300 8.780 117.850 ;
        RECT 9.230 110.300 9.380 117.850 ;
        RECT 9.830 110.300 9.980 117.850 ;
        RECT 14.230 117.550 15.230 118.000 ;
        RECT 10.880 117.400 18.580 117.550 ;
        RECT 14.230 116.950 15.230 117.400 ;
        RECT 10.880 116.800 18.580 116.950 ;
        RECT 14.230 116.350 15.230 116.800 ;
        RECT 10.880 116.200 18.580 116.350 ;
        RECT 14.230 115.750 15.230 116.200 ;
        RECT 10.880 115.600 18.580 115.750 ;
        RECT 14.230 115.150 15.230 115.600 ;
        RECT 10.880 115.000 18.580 115.150 ;
        RECT 14.230 114.550 15.230 115.000 ;
        RECT 10.880 114.400 18.580 114.550 ;
        RECT 14.230 113.950 15.230 114.400 ;
        RECT 10.880 113.800 18.580 113.950 ;
        RECT 14.230 113.350 15.230 113.800 ;
        RECT 10.880 113.200 18.580 113.350 ;
        RECT 14.230 112.750 15.230 113.200 ;
        RECT 10.880 112.600 18.580 112.750 ;
        RECT 14.230 112.150 15.230 112.600 ;
        RECT 10.880 112.000 18.580 112.150 ;
        RECT 14.230 111.550 15.230 112.000 ;
        RECT 10.880 111.400 18.580 111.550 ;
        RECT 14.230 110.950 15.230 111.400 ;
        RECT 10.880 110.800 18.580 110.950 ;
        RECT 14.230 110.300 15.230 110.800 ;
        RECT 19.480 110.300 19.630 117.850 ;
        RECT 20.080 110.300 20.230 117.850 ;
        RECT 20.680 110.300 20.830 117.850 ;
        RECT 21.280 110.300 21.430 117.850 ;
        RECT 21.880 110.300 22.030 117.850 ;
        RECT 22.480 110.300 22.630 117.850 ;
        RECT 22.780 113.200 23.530 115.000 ;
        RECT 25.930 113.200 26.680 115.000 ;
        RECT 22.780 110.450 26.680 113.200 ;
        RECT 22.780 110.300 23.930 110.450 ;
        RECT 5.530 109.700 23.930 110.300 ;
        RECT 5.530 109.550 6.680 109.700 ;
        RECT 4.730 106.800 6.680 109.550 ;
        RECT 5.930 105.050 6.680 106.800 ;
        RECT 6.830 102.150 6.980 109.700 ;
        RECT 7.430 102.150 7.580 109.700 ;
        RECT 8.030 102.150 8.180 109.700 ;
        RECT 8.630 102.150 8.780 109.700 ;
        RECT 9.230 102.150 9.380 109.700 ;
        RECT 9.830 102.150 9.980 109.700 ;
        RECT 14.230 109.200 15.230 109.700 ;
        RECT 10.880 109.050 18.580 109.200 ;
        RECT 14.230 108.600 15.230 109.050 ;
        RECT 10.880 108.450 18.580 108.600 ;
        RECT 14.230 108.000 15.230 108.450 ;
        RECT 10.880 107.850 18.580 108.000 ;
        RECT 14.230 107.400 15.230 107.850 ;
        RECT 10.880 107.250 18.580 107.400 ;
        RECT 14.230 106.800 15.230 107.250 ;
        RECT 10.880 106.650 18.580 106.800 ;
        RECT 14.230 106.200 15.230 106.650 ;
        RECT 10.880 106.050 18.580 106.200 ;
        RECT 14.230 105.600 15.230 106.050 ;
        RECT 10.880 105.450 18.580 105.600 ;
        RECT 14.230 105.000 15.230 105.450 ;
        RECT 10.880 104.850 18.580 105.000 ;
        RECT 14.230 104.400 15.230 104.850 ;
        RECT 10.880 104.250 18.580 104.400 ;
        RECT 14.230 103.800 15.230 104.250 ;
        RECT 10.880 103.650 18.580 103.800 ;
        RECT 14.230 103.200 15.230 103.650 ;
        RECT 10.880 103.050 18.580 103.200 ;
        RECT 14.230 102.600 15.230 103.050 ;
        RECT 10.880 102.450 18.580 102.600 ;
        RECT 14.230 102.000 15.230 102.450 ;
        RECT 19.480 102.150 19.630 109.700 ;
        RECT 20.080 102.150 20.230 109.700 ;
        RECT 20.680 102.150 20.830 109.700 ;
        RECT 21.280 102.150 21.430 109.700 ;
        RECT 21.880 102.150 22.030 109.700 ;
        RECT 22.480 102.150 22.630 109.700 ;
        RECT 22.780 109.550 23.930 109.700 ;
        RECT 24.580 109.550 24.880 110.450 ;
        RECT 25.530 110.300 26.680 110.450 ;
        RECT 26.830 110.300 26.980 117.850 ;
        RECT 27.430 110.300 27.580 117.850 ;
        RECT 28.030 110.300 28.180 117.850 ;
        RECT 28.630 110.300 28.780 117.850 ;
        RECT 29.230 110.300 29.380 117.850 ;
        RECT 29.830 110.300 29.980 117.850 ;
        RECT 34.230 117.550 35.230 118.000 ;
        RECT 30.880 117.400 38.580 117.550 ;
        RECT 34.230 116.950 35.230 117.400 ;
        RECT 30.880 116.800 38.580 116.950 ;
        RECT 34.230 116.350 35.230 116.800 ;
        RECT 30.880 116.200 38.580 116.350 ;
        RECT 34.230 115.750 35.230 116.200 ;
        RECT 30.880 115.600 38.580 115.750 ;
        RECT 34.230 115.150 35.230 115.600 ;
        RECT 30.880 115.000 38.580 115.150 ;
        RECT 34.230 114.550 35.230 115.000 ;
        RECT 30.880 114.400 38.580 114.550 ;
        RECT 34.230 113.950 35.230 114.400 ;
        RECT 30.880 113.800 38.580 113.950 ;
        RECT 34.230 113.350 35.230 113.800 ;
        RECT 30.880 113.200 38.580 113.350 ;
        RECT 34.230 112.750 35.230 113.200 ;
        RECT 30.880 112.600 38.580 112.750 ;
        RECT 34.230 112.150 35.230 112.600 ;
        RECT 30.880 112.000 38.580 112.150 ;
        RECT 34.230 111.550 35.230 112.000 ;
        RECT 30.880 111.400 38.580 111.550 ;
        RECT 34.230 110.950 35.230 111.400 ;
        RECT 30.880 110.800 38.580 110.950 ;
        RECT 34.230 110.300 35.230 110.800 ;
        RECT 39.480 110.300 39.630 117.850 ;
        RECT 40.080 110.300 40.230 117.850 ;
        RECT 40.680 110.300 40.830 117.850 ;
        RECT 41.280 110.300 41.430 117.850 ;
        RECT 41.880 110.300 42.030 117.850 ;
        RECT 42.480 110.300 42.630 117.850 ;
        RECT 42.780 113.200 43.530 115.000 ;
        RECT 45.930 113.200 46.680 115.000 ;
        RECT 42.780 110.450 46.680 113.200 ;
        RECT 42.780 110.300 43.930 110.450 ;
        RECT 25.530 109.700 43.930 110.300 ;
        RECT 25.530 109.550 26.680 109.700 ;
        RECT 22.780 106.800 26.680 109.550 ;
        RECT 22.780 105.050 23.530 106.800 ;
        RECT 25.930 105.050 26.680 106.800 ;
        RECT 26.830 102.150 26.980 109.700 ;
        RECT 27.430 102.150 27.580 109.700 ;
        RECT 28.030 102.150 28.180 109.700 ;
        RECT 28.630 102.150 28.780 109.700 ;
        RECT 29.230 102.150 29.380 109.700 ;
        RECT 29.830 102.150 29.980 109.700 ;
        RECT 34.230 109.200 35.230 109.700 ;
        RECT 30.880 109.050 38.580 109.200 ;
        RECT 34.230 108.600 35.230 109.050 ;
        RECT 30.880 108.450 38.580 108.600 ;
        RECT 34.230 108.000 35.230 108.450 ;
        RECT 30.880 107.850 38.580 108.000 ;
        RECT 34.230 107.400 35.230 107.850 ;
        RECT 30.880 107.250 38.580 107.400 ;
        RECT 34.230 106.800 35.230 107.250 ;
        RECT 30.880 106.650 38.580 106.800 ;
        RECT 34.230 106.200 35.230 106.650 ;
        RECT 30.880 106.050 38.580 106.200 ;
        RECT 34.230 105.600 35.230 106.050 ;
        RECT 30.880 105.450 38.580 105.600 ;
        RECT 34.230 105.000 35.230 105.450 ;
        RECT 30.880 104.850 38.580 105.000 ;
        RECT 34.230 104.400 35.230 104.850 ;
        RECT 30.880 104.250 38.580 104.400 ;
        RECT 34.230 103.800 35.230 104.250 ;
        RECT 30.880 103.650 38.580 103.800 ;
        RECT 34.230 103.200 35.230 103.650 ;
        RECT 30.880 103.050 38.580 103.200 ;
        RECT 34.230 102.600 35.230 103.050 ;
        RECT 30.880 102.450 38.580 102.600 ;
        RECT 34.230 102.000 35.230 102.450 ;
        RECT 39.480 102.150 39.630 109.700 ;
        RECT 40.080 102.150 40.230 109.700 ;
        RECT 40.680 102.150 40.830 109.700 ;
        RECT 41.280 102.150 41.430 109.700 ;
        RECT 41.880 102.150 42.030 109.700 ;
        RECT 42.480 102.150 42.630 109.700 ;
        RECT 42.780 109.550 43.930 109.700 ;
        RECT 44.580 109.550 44.880 110.450 ;
        RECT 45.530 110.300 46.680 110.450 ;
        RECT 46.830 110.300 46.980 117.850 ;
        RECT 47.430 110.300 47.580 117.850 ;
        RECT 48.030 110.300 48.180 117.850 ;
        RECT 48.630 110.300 48.780 117.850 ;
        RECT 49.230 110.300 49.380 117.850 ;
        RECT 49.830 110.300 49.980 117.850 ;
        RECT 54.230 117.550 55.230 118.000 ;
        RECT 50.880 117.400 58.580 117.550 ;
        RECT 54.230 116.950 55.230 117.400 ;
        RECT 50.880 116.800 58.580 116.950 ;
        RECT 54.230 116.350 55.230 116.800 ;
        RECT 50.880 116.200 58.580 116.350 ;
        RECT 54.230 115.750 55.230 116.200 ;
        RECT 50.880 115.600 58.580 115.750 ;
        RECT 54.230 115.150 55.230 115.600 ;
        RECT 50.880 115.000 58.580 115.150 ;
        RECT 54.230 114.550 55.230 115.000 ;
        RECT 50.880 114.400 58.580 114.550 ;
        RECT 54.230 113.950 55.230 114.400 ;
        RECT 50.880 113.800 58.580 113.950 ;
        RECT 54.230 113.350 55.230 113.800 ;
        RECT 50.880 113.200 58.580 113.350 ;
        RECT 54.230 112.750 55.230 113.200 ;
        RECT 50.880 112.600 58.580 112.750 ;
        RECT 54.230 112.150 55.230 112.600 ;
        RECT 50.880 112.000 58.580 112.150 ;
        RECT 54.230 111.550 55.230 112.000 ;
        RECT 50.880 111.400 58.580 111.550 ;
        RECT 54.230 110.950 55.230 111.400 ;
        RECT 50.880 110.800 58.580 110.950 ;
        RECT 54.230 110.300 55.230 110.800 ;
        RECT 59.480 110.300 59.630 117.850 ;
        RECT 60.080 110.300 60.230 117.850 ;
        RECT 60.680 110.300 60.830 117.850 ;
        RECT 61.280 110.300 61.430 117.850 ;
        RECT 61.880 110.300 62.030 117.850 ;
        RECT 62.480 110.300 62.630 117.850 ;
        RECT 62.780 113.200 63.530 115.000 ;
        RECT 65.930 113.200 66.680 115.000 ;
        RECT 62.780 110.450 66.680 113.200 ;
        RECT 62.780 110.300 63.930 110.450 ;
        RECT 45.530 109.700 63.930 110.300 ;
        RECT 45.530 109.550 46.680 109.700 ;
        RECT 42.780 106.800 46.680 109.550 ;
        RECT 42.780 105.050 43.530 106.800 ;
        RECT 45.930 105.050 46.680 106.800 ;
        RECT 46.830 102.150 46.980 109.700 ;
        RECT 47.430 102.150 47.580 109.700 ;
        RECT 48.030 102.150 48.180 109.700 ;
        RECT 48.630 102.150 48.780 109.700 ;
        RECT 49.230 102.150 49.380 109.700 ;
        RECT 49.830 102.150 49.980 109.700 ;
        RECT 54.230 109.200 55.230 109.700 ;
        RECT 50.880 109.050 58.580 109.200 ;
        RECT 54.230 108.600 55.230 109.050 ;
        RECT 50.880 108.450 58.580 108.600 ;
        RECT 54.230 108.000 55.230 108.450 ;
        RECT 50.880 107.850 58.580 108.000 ;
        RECT 54.230 107.400 55.230 107.850 ;
        RECT 50.880 107.250 58.580 107.400 ;
        RECT 54.230 106.800 55.230 107.250 ;
        RECT 50.880 106.650 58.580 106.800 ;
        RECT 54.230 106.200 55.230 106.650 ;
        RECT 50.880 106.050 58.580 106.200 ;
        RECT 54.230 105.600 55.230 106.050 ;
        RECT 50.880 105.450 58.580 105.600 ;
        RECT 54.230 105.000 55.230 105.450 ;
        RECT 50.880 104.850 58.580 105.000 ;
        RECT 54.230 104.400 55.230 104.850 ;
        RECT 50.880 104.250 58.580 104.400 ;
        RECT 54.230 103.800 55.230 104.250 ;
        RECT 50.880 103.650 58.580 103.800 ;
        RECT 54.230 103.200 55.230 103.650 ;
        RECT 50.880 103.050 58.580 103.200 ;
        RECT 54.230 102.600 55.230 103.050 ;
        RECT 50.880 102.450 58.580 102.600 ;
        RECT 54.230 102.000 55.230 102.450 ;
        RECT 59.480 102.150 59.630 109.700 ;
        RECT 60.080 102.150 60.230 109.700 ;
        RECT 60.680 102.150 60.830 109.700 ;
        RECT 61.280 102.150 61.430 109.700 ;
        RECT 61.880 102.150 62.030 109.700 ;
        RECT 62.480 102.150 62.630 109.700 ;
        RECT 62.780 109.550 63.930 109.700 ;
        RECT 64.580 109.550 64.880 110.450 ;
        RECT 65.530 110.300 66.680 110.450 ;
        RECT 66.830 110.300 66.980 117.850 ;
        RECT 67.430 110.300 67.580 117.850 ;
        RECT 68.030 110.300 68.180 117.850 ;
        RECT 68.630 110.300 68.780 117.850 ;
        RECT 69.230 110.300 69.380 117.850 ;
        RECT 69.830 110.300 69.980 117.850 ;
        RECT 74.230 117.550 75.230 118.000 ;
        RECT 70.880 117.400 78.580 117.550 ;
        RECT 74.230 116.950 75.230 117.400 ;
        RECT 70.880 116.800 78.580 116.950 ;
        RECT 74.230 116.350 75.230 116.800 ;
        RECT 70.880 116.200 78.580 116.350 ;
        RECT 74.230 115.750 75.230 116.200 ;
        RECT 70.880 115.600 78.580 115.750 ;
        RECT 74.230 115.150 75.230 115.600 ;
        RECT 70.880 115.000 78.580 115.150 ;
        RECT 74.230 114.550 75.230 115.000 ;
        RECT 70.880 114.400 78.580 114.550 ;
        RECT 74.230 113.950 75.230 114.400 ;
        RECT 70.880 113.800 78.580 113.950 ;
        RECT 74.230 113.350 75.230 113.800 ;
        RECT 70.880 113.200 78.580 113.350 ;
        RECT 74.230 112.750 75.230 113.200 ;
        RECT 70.880 112.600 78.580 112.750 ;
        RECT 74.230 112.150 75.230 112.600 ;
        RECT 70.880 112.000 78.580 112.150 ;
        RECT 74.230 111.550 75.230 112.000 ;
        RECT 70.880 111.400 78.580 111.550 ;
        RECT 74.230 110.950 75.230 111.400 ;
        RECT 70.880 110.800 78.580 110.950 ;
        RECT 74.230 110.300 75.230 110.800 ;
        RECT 79.480 110.300 79.630 117.850 ;
        RECT 80.080 110.300 80.230 117.850 ;
        RECT 80.680 110.300 80.830 117.850 ;
        RECT 81.280 110.300 81.430 117.850 ;
        RECT 81.880 110.300 82.030 117.850 ;
        RECT 82.480 110.300 82.630 117.850 ;
        RECT 82.780 113.200 83.530 115.000 ;
        RECT 85.930 113.200 86.680 115.000 ;
        RECT 82.780 110.450 86.680 113.200 ;
        RECT 82.780 110.300 83.930 110.450 ;
        RECT 65.530 109.700 83.930 110.300 ;
        RECT 65.530 109.550 66.680 109.700 ;
        RECT 62.780 106.800 66.680 109.550 ;
        RECT 62.780 105.050 63.530 106.800 ;
        RECT 65.930 105.050 66.680 106.800 ;
        RECT 66.830 102.150 66.980 109.700 ;
        RECT 67.430 102.150 67.580 109.700 ;
        RECT 68.030 102.150 68.180 109.700 ;
        RECT 68.630 102.150 68.780 109.700 ;
        RECT 69.230 102.150 69.380 109.700 ;
        RECT 69.830 102.150 69.980 109.700 ;
        RECT 74.230 109.200 75.230 109.700 ;
        RECT 70.880 109.050 78.580 109.200 ;
        RECT 74.230 108.600 75.230 109.050 ;
        RECT 70.880 108.450 78.580 108.600 ;
        RECT 74.230 108.000 75.230 108.450 ;
        RECT 70.880 107.850 78.580 108.000 ;
        RECT 74.230 107.400 75.230 107.850 ;
        RECT 70.880 107.250 78.580 107.400 ;
        RECT 74.230 106.800 75.230 107.250 ;
        RECT 70.880 106.650 78.580 106.800 ;
        RECT 74.230 106.200 75.230 106.650 ;
        RECT 70.880 106.050 78.580 106.200 ;
        RECT 74.230 105.600 75.230 106.050 ;
        RECT 70.880 105.450 78.580 105.600 ;
        RECT 74.230 105.000 75.230 105.450 ;
        RECT 70.880 104.850 78.580 105.000 ;
        RECT 74.230 104.400 75.230 104.850 ;
        RECT 70.880 104.250 78.580 104.400 ;
        RECT 74.230 103.800 75.230 104.250 ;
        RECT 70.880 103.650 78.580 103.800 ;
        RECT 74.230 103.200 75.230 103.650 ;
        RECT 70.880 103.050 78.580 103.200 ;
        RECT 74.230 102.600 75.230 103.050 ;
        RECT 70.880 102.450 78.580 102.600 ;
        RECT 74.230 102.000 75.230 102.450 ;
        RECT 79.480 102.150 79.630 109.700 ;
        RECT 80.080 102.150 80.230 109.700 ;
        RECT 80.680 102.150 80.830 109.700 ;
        RECT 81.280 102.150 81.430 109.700 ;
        RECT 81.880 102.150 82.030 109.700 ;
        RECT 82.480 102.150 82.630 109.700 ;
        RECT 82.780 109.550 83.930 109.700 ;
        RECT 84.580 109.550 84.880 110.450 ;
        RECT 85.530 110.300 86.680 110.450 ;
        RECT 86.830 110.300 86.980 117.850 ;
        RECT 87.430 110.300 87.580 117.850 ;
        RECT 88.030 110.300 88.180 117.850 ;
        RECT 88.630 110.300 88.780 117.850 ;
        RECT 89.230 110.300 89.380 117.850 ;
        RECT 89.830 110.300 89.980 117.850 ;
        RECT 94.230 117.550 95.230 118.000 ;
        RECT 90.880 117.400 98.580 117.550 ;
        RECT 94.230 116.950 95.230 117.400 ;
        RECT 90.880 116.800 98.580 116.950 ;
        RECT 94.230 116.350 95.230 116.800 ;
        RECT 90.880 116.200 98.580 116.350 ;
        RECT 94.230 115.750 95.230 116.200 ;
        RECT 90.880 115.600 98.580 115.750 ;
        RECT 94.230 115.150 95.230 115.600 ;
        RECT 90.880 115.000 98.580 115.150 ;
        RECT 94.230 114.550 95.230 115.000 ;
        RECT 90.880 114.400 98.580 114.550 ;
        RECT 94.230 113.950 95.230 114.400 ;
        RECT 90.880 113.800 98.580 113.950 ;
        RECT 94.230 113.350 95.230 113.800 ;
        RECT 90.880 113.200 98.580 113.350 ;
        RECT 94.230 112.750 95.230 113.200 ;
        RECT 90.880 112.600 98.580 112.750 ;
        RECT 94.230 112.150 95.230 112.600 ;
        RECT 90.880 112.000 98.580 112.150 ;
        RECT 94.230 111.550 95.230 112.000 ;
        RECT 90.880 111.400 98.580 111.550 ;
        RECT 94.230 110.950 95.230 111.400 ;
        RECT 90.880 110.800 98.580 110.950 ;
        RECT 94.230 110.300 95.230 110.800 ;
        RECT 99.480 110.300 99.630 117.850 ;
        RECT 100.080 110.300 100.230 117.850 ;
        RECT 100.680 110.300 100.830 117.850 ;
        RECT 101.280 110.300 101.430 117.850 ;
        RECT 101.880 110.300 102.030 117.850 ;
        RECT 102.480 110.300 102.630 117.850 ;
        RECT 102.780 113.200 103.530 115.000 ;
        RECT 105.930 113.200 106.680 115.000 ;
        RECT 102.780 110.450 106.680 113.200 ;
        RECT 102.780 110.300 103.930 110.450 ;
        RECT 85.530 109.700 103.930 110.300 ;
        RECT 85.530 109.550 86.680 109.700 ;
        RECT 82.780 106.800 86.680 109.550 ;
        RECT 82.780 105.050 83.530 106.800 ;
        RECT 85.930 105.050 86.680 106.800 ;
        RECT 86.830 102.150 86.980 109.700 ;
        RECT 87.430 102.150 87.580 109.700 ;
        RECT 88.030 102.150 88.180 109.700 ;
        RECT 88.630 102.150 88.780 109.700 ;
        RECT 89.230 102.150 89.380 109.700 ;
        RECT 89.830 102.150 89.980 109.700 ;
        RECT 94.230 109.200 95.230 109.700 ;
        RECT 90.880 109.050 98.580 109.200 ;
        RECT 94.230 108.600 95.230 109.050 ;
        RECT 90.880 108.450 98.580 108.600 ;
        RECT 94.230 108.000 95.230 108.450 ;
        RECT 90.880 107.850 98.580 108.000 ;
        RECT 94.230 107.400 95.230 107.850 ;
        RECT 90.880 107.250 98.580 107.400 ;
        RECT 94.230 106.800 95.230 107.250 ;
        RECT 90.880 106.650 98.580 106.800 ;
        RECT 94.230 106.200 95.230 106.650 ;
        RECT 90.880 106.050 98.580 106.200 ;
        RECT 94.230 105.600 95.230 106.050 ;
        RECT 90.880 105.450 98.580 105.600 ;
        RECT 94.230 105.000 95.230 105.450 ;
        RECT 90.880 104.850 98.580 105.000 ;
        RECT 94.230 104.400 95.230 104.850 ;
        RECT 90.880 104.250 98.580 104.400 ;
        RECT 94.230 103.800 95.230 104.250 ;
        RECT 90.880 103.650 98.580 103.800 ;
        RECT 94.230 103.200 95.230 103.650 ;
        RECT 90.880 103.050 98.580 103.200 ;
        RECT 94.230 102.600 95.230 103.050 ;
        RECT 90.880 102.450 98.580 102.600 ;
        RECT 94.230 102.000 95.230 102.450 ;
        RECT 99.480 102.150 99.630 109.700 ;
        RECT 100.080 102.150 100.230 109.700 ;
        RECT 100.680 102.150 100.830 109.700 ;
        RECT 101.280 102.150 101.430 109.700 ;
        RECT 101.880 102.150 102.030 109.700 ;
        RECT 102.480 102.150 102.630 109.700 ;
        RECT 102.780 109.550 103.930 109.700 ;
        RECT 104.580 109.550 104.880 110.450 ;
        RECT 105.530 110.300 106.680 110.450 ;
        RECT 106.830 110.300 106.980 117.850 ;
        RECT 107.430 110.300 107.580 117.850 ;
        RECT 108.030 110.300 108.180 117.850 ;
        RECT 108.630 110.300 108.780 117.850 ;
        RECT 109.230 110.300 109.380 117.850 ;
        RECT 109.830 110.300 109.980 117.850 ;
        RECT 114.230 117.550 115.230 118.000 ;
        RECT 110.880 117.400 118.580 117.550 ;
        RECT 114.230 116.950 115.230 117.400 ;
        RECT 110.880 116.800 118.580 116.950 ;
        RECT 114.230 116.350 115.230 116.800 ;
        RECT 110.880 116.200 118.580 116.350 ;
        RECT 114.230 115.750 115.230 116.200 ;
        RECT 110.880 115.600 118.580 115.750 ;
        RECT 114.230 115.150 115.230 115.600 ;
        RECT 110.880 115.000 118.580 115.150 ;
        RECT 114.230 114.550 115.230 115.000 ;
        RECT 110.880 114.400 118.580 114.550 ;
        RECT 114.230 113.950 115.230 114.400 ;
        RECT 110.880 113.800 118.580 113.950 ;
        RECT 114.230 113.350 115.230 113.800 ;
        RECT 110.880 113.200 118.580 113.350 ;
        RECT 114.230 112.750 115.230 113.200 ;
        RECT 110.880 112.600 118.580 112.750 ;
        RECT 114.230 112.150 115.230 112.600 ;
        RECT 110.880 112.000 118.580 112.150 ;
        RECT 114.230 111.550 115.230 112.000 ;
        RECT 110.880 111.400 118.580 111.550 ;
        RECT 114.230 110.950 115.230 111.400 ;
        RECT 110.880 110.800 118.580 110.950 ;
        RECT 114.230 110.300 115.230 110.800 ;
        RECT 119.480 110.300 119.630 117.850 ;
        RECT 120.080 110.300 120.230 117.850 ;
        RECT 120.680 110.300 120.830 117.850 ;
        RECT 121.280 110.300 121.430 117.850 ;
        RECT 121.880 110.300 122.030 117.850 ;
        RECT 122.480 110.300 122.630 117.850 ;
        RECT 122.780 113.200 123.530 115.000 ;
        RECT 122.780 110.450 124.730 113.200 ;
        RECT 122.780 110.300 123.930 110.450 ;
        RECT 105.530 109.700 123.930 110.300 ;
        RECT 105.530 109.550 106.680 109.700 ;
        RECT 102.780 106.800 106.680 109.550 ;
        RECT 102.780 105.050 103.530 106.800 ;
        RECT 105.930 105.050 106.680 106.800 ;
        RECT 106.830 102.150 106.980 109.700 ;
        RECT 107.430 102.150 107.580 109.700 ;
        RECT 108.030 102.150 108.180 109.700 ;
        RECT 108.630 102.150 108.780 109.700 ;
        RECT 109.230 102.150 109.380 109.700 ;
        RECT 109.830 102.150 109.980 109.700 ;
        RECT 114.230 109.200 115.230 109.700 ;
        RECT 110.880 109.050 118.580 109.200 ;
        RECT 114.230 108.600 115.230 109.050 ;
        RECT 110.880 108.450 118.580 108.600 ;
        RECT 114.230 108.000 115.230 108.450 ;
        RECT 110.880 107.850 118.580 108.000 ;
        RECT 114.230 107.400 115.230 107.850 ;
        RECT 110.880 107.250 118.580 107.400 ;
        RECT 114.230 106.800 115.230 107.250 ;
        RECT 110.880 106.650 118.580 106.800 ;
        RECT 114.230 106.200 115.230 106.650 ;
        RECT 110.880 106.050 118.580 106.200 ;
        RECT 114.230 105.600 115.230 106.050 ;
        RECT 110.880 105.450 118.580 105.600 ;
        RECT 114.230 105.000 115.230 105.450 ;
        RECT 110.880 104.850 118.580 105.000 ;
        RECT 114.230 104.400 115.230 104.850 ;
        RECT 110.880 104.250 118.580 104.400 ;
        RECT 114.230 103.800 115.230 104.250 ;
        RECT 110.880 103.650 118.580 103.800 ;
        RECT 114.230 103.200 115.230 103.650 ;
        RECT 110.880 103.050 118.580 103.200 ;
        RECT 114.230 102.600 115.230 103.050 ;
        RECT 110.880 102.450 118.580 102.600 ;
        RECT 114.230 102.000 115.230 102.450 ;
        RECT 119.480 102.150 119.630 109.700 ;
        RECT 120.080 102.150 120.230 109.700 ;
        RECT 120.680 102.150 120.830 109.700 ;
        RECT 121.280 102.150 121.430 109.700 ;
        RECT 121.880 102.150 122.030 109.700 ;
        RECT 122.480 102.150 122.630 109.700 ;
        RECT 122.780 109.550 123.930 109.700 ;
        RECT 124.580 109.980 124.730 110.450 ;
        RECT 124.580 109.550 131.850 109.980 ;
        RECT 122.780 108.705 131.850 109.550 ;
        RECT 122.780 106.800 124.730 108.705 ;
        RECT 122.780 105.050 123.530 106.800 ;
        RECT 10.880 101.850 18.580 102.000 ;
        RECT 30.880 101.850 38.580 102.000 ;
        RECT 50.880 101.850 58.580 102.000 ;
        RECT 70.880 101.850 78.580 102.000 ;
        RECT 90.880 101.850 98.580 102.000 ;
        RECT 110.880 101.850 118.580 102.000 ;
        RECT 14.230 101.200 15.230 101.850 ;
        RECT 34.230 101.200 35.230 101.850 ;
        RECT 54.230 101.200 55.230 101.850 ;
        RECT 74.230 101.200 75.230 101.850 ;
        RECT 94.230 101.200 95.230 101.850 ;
        RECT 114.230 101.200 115.230 101.850 ;
        RECT 11.530 98.800 17.930 101.200 ;
        RECT 31.530 98.800 37.930 101.200 ;
        RECT 51.530 98.800 57.930 101.200 ;
        RECT 71.530 98.800 77.930 101.200 ;
        RECT 91.530 98.800 97.930 101.200 ;
        RECT 111.530 98.800 117.930 101.200 ;
        RECT 14.230 98.150 15.230 98.800 ;
        RECT 34.230 98.150 35.230 98.800 ;
        RECT 54.230 98.150 55.230 98.800 ;
        RECT 74.230 98.150 75.230 98.800 ;
        RECT 94.230 98.150 95.230 98.800 ;
        RECT 114.230 98.150 115.230 98.800 ;
        RECT 10.880 98.000 18.580 98.150 ;
        RECT 30.880 98.000 38.580 98.150 ;
        RECT 50.880 98.000 58.580 98.150 ;
        RECT 70.880 98.000 78.580 98.150 ;
        RECT 90.880 98.000 98.580 98.150 ;
        RECT 110.880 98.000 118.580 98.150 ;
        RECT 5.930 93.200 6.680 95.000 ;
        RECT 4.730 90.450 6.680 93.200 ;
        RECT 4.730 89.550 4.880 90.450 ;
        RECT 5.530 90.300 6.680 90.450 ;
        RECT 6.830 90.300 6.980 97.850 ;
        RECT 7.430 90.300 7.580 97.850 ;
        RECT 8.030 90.300 8.180 97.850 ;
        RECT 8.630 90.300 8.780 97.850 ;
        RECT 9.230 90.300 9.380 97.850 ;
        RECT 9.830 90.300 9.980 97.850 ;
        RECT 14.230 97.550 15.230 98.000 ;
        RECT 10.880 97.400 18.580 97.550 ;
        RECT 14.230 96.950 15.230 97.400 ;
        RECT 10.880 96.800 18.580 96.950 ;
        RECT 14.230 96.350 15.230 96.800 ;
        RECT 10.880 96.200 18.580 96.350 ;
        RECT 14.230 95.750 15.230 96.200 ;
        RECT 10.880 95.600 18.580 95.750 ;
        RECT 14.230 95.150 15.230 95.600 ;
        RECT 10.880 95.000 18.580 95.150 ;
        RECT 14.230 94.550 15.230 95.000 ;
        RECT 10.880 94.400 18.580 94.550 ;
        RECT 14.230 93.950 15.230 94.400 ;
        RECT 10.880 93.800 18.580 93.950 ;
        RECT 14.230 93.350 15.230 93.800 ;
        RECT 10.880 93.200 18.580 93.350 ;
        RECT 14.230 92.750 15.230 93.200 ;
        RECT 10.880 92.600 18.580 92.750 ;
        RECT 14.230 92.150 15.230 92.600 ;
        RECT 10.880 92.000 18.580 92.150 ;
        RECT 14.230 91.550 15.230 92.000 ;
        RECT 10.880 91.400 18.580 91.550 ;
        RECT 14.230 90.950 15.230 91.400 ;
        RECT 10.880 90.800 18.580 90.950 ;
        RECT 14.230 90.300 15.230 90.800 ;
        RECT 19.480 90.300 19.630 97.850 ;
        RECT 20.080 90.300 20.230 97.850 ;
        RECT 20.680 90.300 20.830 97.850 ;
        RECT 21.280 90.300 21.430 97.850 ;
        RECT 21.880 90.300 22.030 97.850 ;
        RECT 22.480 90.300 22.630 97.850 ;
        RECT 22.780 93.200 23.530 95.000 ;
        RECT 25.930 93.200 26.680 95.000 ;
        RECT 22.780 90.450 26.680 93.200 ;
        RECT 22.780 90.300 23.930 90.450 ;
        RECT 5.530 89.700 23.930 90.300 ;
        RECT 5.530 89.550 6.680 89.700 ;
        RECT 4.730 86.800 6.680 89.550 ;
        RECT 5.930 85.050 6.680 86.800 ;
        RECT 6.830 82.150 6.980 89.700 ;
        RECT 7.430 82.150 7.580 89.700 ;
        RECT 8.030 82.150 8.180 89.700 ;
        RECT 8.630 82.150 8.780 89.700 ;
        RECT 9.230 82.150 9.380 89.700 ;
        RECT 9.830 82.150 9.980 89.700 ;
        RECT 14.230 89.200 15.230 89.700 ;
        RECT 10.880 89.050 18.580 89.200 ;
        RECT 14.230 88.600 15.230 89.050 ;
        RECT 10.880 88.450 18.580 88.600 ;
        RECT 14.230 88.000 15.230 88.450 ;
        RECT 10.880 87.850 18.580 88.000 ;
        RECT 14.230 87.400 15.230 87.850 ;
        RECT 10.880 87.250 18.580 87.400 ;
        RECT 14.230 86.800 15.230 87.250 ;
        RECT 10.880 86.650 18.580 86.800 ;
        RECT 14.230 86.200 15.230 86.650 ;
        RECT 10.880 86.050 18.580 86.200 ;
        RECT 14.230 85.600 15.230 86.050 ;
        RECT 10.880 85.450 18.580 85.600 ;
        RECT 14.230 85.000 15.230 85.450 ;
        RECT 10.880 84.850 18.580 85.000 ;
        RECT 14.230 84.400 15.230 84.850 ;
        RECT 10.880 84.250 18.580 84.400 ;
        RECT 14.230 83.800 15.230 84.250 ;
        RECT 10.880 83.650 18.580 83.800 ;
        RECT 14.230 83.200 15.230 83.650 ;
        RECT 10.880 83.050 18.580 83.200 ;
        RECT 14.230 82.600 15.230 83.050 ;
        RECT 10.880 82.450 18.580 82.600 ;
        RECT 14.230 82.000 15.230 82.450 ;
        RECT 19.480 82.150 19.630 89.700 ;
        RECT 20.080 82.150 20.230 89.700 ;
        RECT 20.680 82.150 20.830 89.700 ;
        RECT 21.280 82.150 21.430 89.700 ;
        RECT 21.880 82.150 22.030 89.700 ;
        RECT 22.480 82.150 22.630 89.700 ;
        RECT 22.780 89.550 23.930 89.700 ;
        RECT 24.580 89.550 24.880 90.450 ;
        RECT 25.530 90.300 26.680 90.450 ;
        RECT 26.830 90.300 26.980 97.850 ;
        RECT 27.430 90.300 27.580 97.850 ;
        RECT 28.030 90.300 28.180 97.850 ;
        RECT 28.630 90.300 28.780 97.850 ;
        RECT 29.230 90.300 29.380 97.850 ;
        RECT 29.830 90.300 29.980 97.850 ;
        RECT 34.230 97.550 35.230 98.000 ;
        RECT 30.880 97.400 38.580 97.550 ;
        RECT 34.230 96.950 35.230 97.400 ;
        RECT 30.880 96.800 38.580 96.950 ;
        RECT 34.230 96.350 35.230 96.800 ;
        RECT 30.880 96.200 38.580 96.350 ;
        RECT 34.230 95.750 35.230 96.200 ;
        RECT 30.880 95.600 38.580 95.750 ;
        RECT 34.230 95.150 35.230 95.600 ;
        RECT 30.880 95.000 38.580 95.150 ;
        RECT 34.230 94.550 35.230 95.000 ;
        RECT 30.880 94.400 38.580 94.550 ;
        RECT 34.230 93.950 35.230 94.400 ;
        RECT 30.880 93.800 38.580 93.950 ;
        RECT 34.230 93.350 35.230 93.800 ;
        RECT 30.880 93.200 38.580 93.350 ;
        RECT 34.230 92.750 35.230 93.200 ;
        RECT 30.880 92.600 38.580 92.750 ;
        RECT 34.230 92.150 35.230 92.600 ;
        RECT 30.880 92.000 38.580 92.150 ;
        RECT 34.230 91.550 35.230 92.000 ;
        RECT 30.880 91.400 38.580 91.550 ;
        RECT 34.230 90.950 35.230 91.400 ;
        RECT 30.880 90.800 38.580 90.950 ;
        RECT 34.230 90.300 35.230 90.800 ;
        RECT 39.480 90.300 39.630 97.850 ;
        RECT 40.080 90.300 40.230 97.850 ;
        RECT 40.680 90.300 40.830 97.850 ;
        RECT 41.280 90.300 41.430 97.850 ;
        RECT 41.880 90.300 42.030 97.850 ;
        RECT 42.480 90.300 42.630 97.850 ;
        RECT 42.780 93.200 43.530 95.000 ;
        RECT 45.930 93.200 46.680 95.000 ;
        RECT 42.780 90.450 46.680 93.200 ;
        RECT 42.780 90.300 43.930 90.450 ;
        RECT 25.530 89.700 43.930 90.300 ;
        RECT 25.530 89.550 26.680 89.700 ;
        RECT 22.780 86.800 26.680 89.550 ;
        RECT 22.780 85.050 23.530 86.800 ;
        RECT 25.930 85.050 26.680 86.800 ;
        RECT 26.830 82.150 26.980 89.700 ;
        RECT 27.430 82.150 27.580 89.700 ;
        RECT 28.030 82.150 28.180 89.700 ;
        RECT 28.630 82.150 28.780 89.700 ;
        RECT 29.230 82.150 29.380 89.700 ;
        RECT 29.830 82.150 29.980 89.700 ;
        RECT 34.230 89.200 35.230 89.700 ;
        RECT 30.880 89.050 38.580 89.200 ;
        RECT 34.230 88.600 35.230 89.050 ;
        RECT 30.880 88.450 38.580 88.600 ;
        RECT 34.230 88.000 35.230 88.450 ;
        RECT 30.880 87.850 38.580 88.000 ;
        RECT 34.230 87.400 35.230 87.850 ;
        RECT 30.880 87.250 38.580 87.400 ;
        RECT 34.230 86.800 35.230 87.250 ;
        RECT 30.880 86.650 38.580 86.800 ;
        RECT 34.230 86.200 35.230 86.650 ;
        RECT 30.880 86.050 38.580 86.200 ;
        RECT 34.230 85.600 35.230 86.050 ;
        RECT 30.880 85.450 38.580 85.600 ;
        RECT 34.230 85.000 35.230 85.450 ;
        RECT 30.880 84.850 38.580 85.000 ;
        RECT 34.230 84.400 35.230 84.850 ;
        RECT 30.880 84.250 38.580 84.400 ;
        RECT 34.230 83.800 35.230 84.250 ;
        RECT 30.880 83.650 38.580 83.800 ;
        RECT 34.230 83.200 35.230 83.650 ;
        RECT 30.880 83.050 38.580 83.200 ;
        RECT 34.230 82.600 35.230 83.050 ;
        RECT 30.880 82.450 38.580 82.600 ;
        RECT 34.230 82.000 35.230 82.450 ;
        RECT 39.480 82.150 39.630 89.700 ;
        RECT 40.080 82.150 40.230 89.700 ;
        RECT 40.680 82.150 40.830 89.700 ;
        RECT 41.280 82.150 41.430 89.700 ;
        RECT 41.880 82.150 42.030 89.700 ;
        RECT 42.480 82.150 42.630 89.700 ;
        RECT 42.780 89.550 43.930 89.700 ;
        RECT 44.580 89.550 44.880 90.450 ;
        RECT 45.530 90.300 46.680 90.450 ;
        RECT 46.830 90.300 46.980 97.850 ;
        RECT 47.430 90.300 47.580 97.850 ;
        RECT 48.030 90.300 48.180 97.850 ;
        RECT 48.630 90.300 48.780 97.850 ;
        RECT 49.230 90.300 49.380 97.850 ;
        RECT 49.830 90.300 49.980 97.850 ;
        RECT 54.230 97.550 55.230 98.000 ;
        RECT 50.880 97.400 58.580 97.550 ;
        RECT 54.230 96.950 55.230 97.400 ;
        RECT 50.880 96.800 58.580 96.950 ;
        RECT 54.230 96.350 55.230 96.800 ;
        RECT 50.880 96.200 58.580 96.350 ;
        RECT 54.230 95.750 55.230 96.200 ;
        RECT 50.880 95.600 58.580 95.750 ;
        RECT 54.230 95.150 55.230 95.600 ;
        RECT 50.880 95.000 58.580 95.150 ;
        RECT 54.230 94.550 55.230 95.000 ;
        RECT 50.880 94.400 58.580 94.550 ;
        RECT 54.230 93.950 55.230 94.400 ;
        RECT 50.880 93.800 58.580 93.950 ;
        RECT 54.230 93.350 55.230 93.800 ;
        RECT 50.880 93.200 58.580 93.350 ;
        RECT 54.230 92.750 55.230 93.200 ;
        RECT 50.880 92.600 58.580 92.750 ;
        RECT 54.230 92.150 55.230 92.600 ;
        RECT 50.880 92.000 58.580 92.150 ;
        RECT 54.230 91.550 55.230 92.000 ;
        RECT 50.880 91.400 58.580 91.550 ;
        RECT 54.230 90.950 55.230 91.400 ;
        RECT 50.880 90.800 58.580 90.950 ;
        RECT 54.230 90.300 55.230 90.800 ;
        RECT 59.480 90.300 59.630 97.850 ;
        RECT 60.080 90.300 60.230 97.850 ;
        RECT 60.680 90.300 60.830 97.850 ;
        RECT 61.280 90.300 61.430 97.850 ;
        RECT 61.880 90.300 62.030 97.850 ;
        RECT 62.480 90.300 62.630 97.850 ;
        RECT 62.780 93.200 63.530 95.000 ;
        RECT 65.930 93.200 66.680 95.000 ;
        RECT 62.780 90.450 66.680 93.200 ;
        RECT 62.780 90.300 63.930 90.450 ;
        RECT 45.530 89.700 63.930 90.300 ;
        RECT 45.530 89.550 46.680 89.700 ;
        RECT 42.780 86.800 46.680 89.550 ;
        RECT 42.780 85.050 43.530 86.800 ;
        RECT 45.930 85.050 46.680 86.800 ;
        RECT 46.830 82.150 46.980 89.700 ;
        RECT 47.430 82.150 47.580 89.700 ;
        RECT 48.030 82.150 48.180 89.700 ;
        RECT 48.630 82.150 48.780 89.700 ;
        RECT 49.230 82.150 49.380 89.700 ;
        RECT 49.830 82.150 49.980 89.700 ;
        RECT 54.230 89.200 55.230 89.700 ;
        RECT 50.880 89.050 58.580 89.200 ;
        RECT 54.230 88.600 55.230 89.050 ;
        RECT 50.880 88.450 58.580 88.600 ;
        RECT 54.230 88.000 55.230 88.450 ;
        RECT 50.880 87.850 58.580 88.000 ;
        RECT 54.230 87.400 55.230 87.850 ;
        RECT 50.880 87.250 58.580 87.400 ;
        RECT 54.230 86.800 55.230 87.250 ;
        RECT 50.880 86.650 58.580 86.800 ;
        RECT 54.230 86.200 55.230 86.650 ;
        RECT 50.880 86.050 58.580 86.200 ;
        RECT 54.230 85.600 55.230 86.050 ;
        RECT 50.880 85.450 58.580 85.600 ;
        RECT 54.230 85.000 55.230 85.450 ;
        RECT 50.880 84.850 58.580 85.000 ;
        RECT 54.230 84.400 55.230 84.850 ;
        RECT 50.880 84.250 58.580 84.400 ;
        RECT 54.230 83.800 55.230 84.250 ;
        RECT 50.880 83.650 58.580 83.800 ;
        RECT 54.230 83.200 55.230 83.650 ;
        RECT 50.880 83.050 58.580 83.200 ;
        RECT 54.230 82.600 55.230 83.050 ;
        RECT 50.880 82.450 58.580 82.600 ;
        RECT 54.230 82.000 55.230 82.450 ;
        RECT 59.480 82.150 59.630 89.700 ;
        RECT 60.080 82.150 60.230 89.700 ;
        RECT 60.680 82.150 60.830 89.700 ;
        RECT 61.280 82.150 61.430 89.700 ;
        RECT 61.880 82.150 62.030 89.700 ;
        RECT 62.480 82.150 62.630 89.700 ;
        RECT 62.780 89.550 63.930 89.700 ;
        RECT 64.580 89.550 64.880 90.450 ;
        RECT 65.530 90.300 66.680 90.450 ;
        RECT 66.830 90.300 66.980 97.850 ;
        RECT 67.430 90.300 67.580 97.850 ;
        RECT 68.030 90.300 68.180 97.850 ;
        RECT 68.630 90.300 68.780 97.850 ;
        RECT 69.230 90.300 69.380 97.850 ;
        RECT 69.830 90.300 69.980 97.850 ;
        RECT 74.230 97.550 75.230 98.000 ;
        RECT 70.880 97.400 78.580 97.550 ;
        RECT 74.230 96.950 75.230 97.400 ;
        RECT 70.880 96.800 78.580 96.950 ;
        RECT 74.230 96.350 75.230 96.800 ;
        RECT 70.880 96.200 78.580 96.350 ;
        RECT 74.230 95.750 75.230 96.200 ;
        RECT 70.880 95.600 78.580 95.750 ;
        RECT 74.230 95.150 75.230 95.600 ;
        RECT 70.880 95.000 78.580 95.150 ;
        RECT 74.230 94.550 75.230 95.000 ;
        RECT 70.880 94.400 78.580 94.550 ;
        RECT 74.230 93.950 75.230 94.400 ;
        RECT 70.880 93.800 78.580 93.950 ;
        RECT 74.230 93.350 75.230 93.800 ;
        RECT 70.880 93.200 78.580 93.350 ;
        RECT 74.230 92.750 75.230 93.200 ;
        RECT 70.880 92.600 78.580 92.750 ;
        RECT 74.230 92.150 75.230 92.600 ;
        RECT 70.880 92.000 78.580 92.150 ;
        RECT 74.230 91.550 75.230 92.000 ;
        RECT 70.880 91.400 78.580 91.550 ;
        RECT 74.230 90.950 75.230 91.400 ;
        RECT 70.880 90.800 78.580 90.950 ;
        RECT 74.230 90.300 75.230 90.800 ;
        RECT 79.480 90.300 79.630 97.850 ;
        RECT 80.080 90.300 80.230 97.850 ;
        RECT 80.680 90.300 80.830 97.850 ;
        RECT 81.280 90.300 81.430 97.850 ;
        RECT 81.880 90.300 82.030 97.850 ;
        RECT 82.480 90.300 82.630 97.850 ;
        RECT 82.780 93.200 83.530 95.000 ;
        RECT 85.930 93.200 86.680 95.000 ;
        RECT 82.780 90.450 86.680 93.200 ;
        RECT 82.780 90.300 83.930 90.450 ;
        RECT 65.530 89.700 83.930 90.300 ;
        RECT 65.530 89.550 66.680 89.700 ;
        RECT 62.780 86.800 66.680 89.550 ;
        RECT 62.780 85.050 63.530 86.800 ;
        RECT 65.930 85.050 66.680 86.800 ;
        RECT 66.830 82.150 66.980 89.700 ;
        RECT 67.430 82.150 67.580 89.700 ;
        RECT 68.030 82.150 68.180 89.700 ;
        RECT 68.630 82.150 68.780 89.700 ;
        RECT 69.230 82.150 69.380 89.700 ;
        RECT 69.830 82.150 69.980 89.700 ;
        RECT 74.230 89.200 75.230 89.700 ;
        RECT 70.880 89.050 78.580 89.200 ;
        RECT 74.230 88.600 75.230 89.050 ;
        RECT 70.880 88.450 78.580 88.600 ;
        RECT 74.230 88.000 75.230 88.450 ;
        RECT 70.880 87.850 78.580 88.000 ;
        RECT 74.230 87.400 75.230 87.850 ;
        RECT 70.880 87.250 78.580 87.400 ;
        RECT 74.230 86.800 75.230 87.250 ;
        RECT 70.880 86.650 78.580 86.800 ;
        RECT 74.230 86.200 75.230 86.650 ;
        RECT 70.880 86.050 78.580 86.200 ;
        RECT 74.230 85.600 75.230 86.050 ;
        RECT 70.880 85.450 78.580 85.600 ;
        RECT 74.230 85.000 75.230 85.450 ;
        RECT 70.880 84.850 78.580 85.000 ;
        RECT 74.230 84.400 75.230 84.850 ;
        RECT 70.880 84.250 78.580 84.400 ;
        RECT 74.230 83.800 75.230 84.250 ;
        RECT 70.880 83.650 78.580 83.800 ;
        RECT 74.230 83.200 75.230 83.650 ;
        RECT 70.880 83.050 78.580 83.200 ;
        RECT 74.230 82.600 75.230 83.050 ;
        RECT 70.880 82.450 78.580 82.600 ;
        RECT 74.230 82.000 75.230 82.450 ;
        RECT 79.480 82.150 79.630 89.700 ;
        RECT 80.080 82.150 80.230 89.700 ;
        RECT 80.680 82.150 80.830 89.700 ;
        RECT 81.280 82.150 81.430 89.700 ;
        RECT 81.880 82.150 82.030 89.700 ;
        RECT 82.480 82.150 82.630 89.700 ;
        RECT 82.780 89.550 83.930 89.700 ;
        RECT 84.580 89.550 84.880 90.450 ;
        RECT 85.530 90.300 86.680 90.450 ;
        RECT 86.830 90.300 86.980 97.850 ;
        RECT 87.430 90.300 87.580 97.850 ;
        RECT 88.030 90.300 88.180 97.850 ;
        RECT 88.630 90.300 88.780 97.850 ;
        RECT 89.230 90.300 89.380 97.850 ;
        RECT 89.830 90.300 89.980 97.850 ;
        RECT 94.230 97.550 95.230 98.000 ;
        RECT 90.880 97.400 98.580 97.550 ;
        RECT 94.230 96.950 95.230 97.400 ;
        RECT 90.880 96.800 98.580 96.950 ;
        RECT 94.230 96.350 95.230 96.800 ;
        RECT 90.880 96.200 98.580 96.350 ;
        RECT 94.230 95.750 95.230 96.200 ;
        RECT 90.880 95.600 98.580 95.750 ;
        RECT 94.230 95.150 95.230 95.600 ;
        RECT 90.880 95.000 98.580 95.150 ;
        RECT 94.230 94.550 95.230 95.000 ;
        RECT 90.880 94.400 98.580 94.550 ;
        RECT 94.230 93.950 95.230 94.400 ;
        RECT 90.880 93.800 98.580 93.950 ;
        RECT 94.230 93.350 95.230 93.800 ;
        RECT 90.880 93.200 98.580 93.350 ;
        RECT 94.230 92.750 95.230 93.200 ;
        RECT 90.880 92.600 98.580 92.750 ;
        RECT 94.230 92.150 95.230 92.600 ;
        RECT 90.880 92.000 98.580 92.150 ;
        RECT 94.230 91.550 95.230 92.000 ;
        RECT 90.880 91.400 98.580 91.550 ;
        RECT 94.230 90.950 95.230 91.400 ;
        RECT 90.880 90.800 98.580 90.950 ;
        RECT 94.230 90.300 95.230 90.800 ;
        RECT 99.480 90.300 99.630 97.850 ;
        RECT 100.080 90.300 100.230 97.850 ;
        RECT 100.680 90.300 100.830 97.850 ;
        RECT 101.280 90.300 101.430 97.850 ;
        RECT 101.880 90.300 102.030 97.850 ;
        RECT 102.480 90.300 102.630 97.850 ;
        RECT 102.780 93.200 103.530 95.000 ;
        RECT 105.930 93.200 106.680 95.000 ;
        RECT 102.780 90.450 106.680 93.200 ;
        RECT 102.780 90.300 103.930 90.450 ;
        RECT 85.530 89.700 103.930 90.300 ;
        RECT 85.530 89.550 86.680 89.700 ;
        RECT 82.780 86.800 86.680 89.550 ;
        RECT 82.780 85.050 83.530 86.800 ;
        RECT 85.930 85.050 86.680 86.800 ;
        RECT 86.830 82.150 86.980 89.700 ;
        RECT 87.430 82.150 87.580 89.700 ;
        RECT 88.030 82.150 88.180 89.700 ;
        RECT 88.630 82.150 88.780 89.700 ;
        RECT 89.230 82.150 89.380 89.700 ;
        RECT 89.830 82.150 89.980 89.700 ;
        RECT 94.230 89.200 95.230 89.700 ;
        RECT 90.880 89.050 98.580 89.200 ;
        RECT 94.230 88.600 95.230 89.050 ;
        RECT 90.880 88.450 98.580 88.600 ;
        RECT 94.230 88.000 95.230 88.450 ;
        RECT 90.880 87.850 98.580 88.000 ;
        RECT 94.230 87.400 95.230 87.850 ;
        RECT 90.880 87.250 98.580 87.400 ;
        RECT 94.230 86.800 95.230 87.250 ;
        RECT 90.880 86.650 98.580 86.800 ;
        RECT 94.230 86.200 95.230 86.650 ;
        RECT 90.880 86.050 98.580 86.200 ;
        RECT 94.230 85.600 95.230 86.050 ;
        RECT 90.880 85.450 98.580 85.600 ;
        RECT 94.230 85.000 95.230 85.450 ;
        RECT 90.880 84.850 98.580 85.000 ;
        RECT 94.230 84.400 95.230 84.850 ;
        RECT 90.880 84.250 98.580 84.400 ;
        RECT 94.230 83.800 95.230 84.250 ;
        RECT 90.880 83.650 98.580 83.800 ;
        RECT 94.230 83.200 95.230 83.650 ;
        RECT 90.880 83.050 98.580 83.200 ;
        RECT 94.230 82.600 95.230 83.050 ;
        RECT 90.880 82.450 98.580 82.600 ;
        RECT 94.230 82.000 95.230 82.450 ;
        RECT 99.480 82.150 99.630 89.700 ;
        RECT 100.080 82.150 100.230 89.700 ;
        RECT 100.680 82.150 100.830 89.700 ;
        RECT 101.280 82.150 101.430 89.700 ;
        RECT 101.880 82.150 102.030 89.700 ;
        RECT 102.480 82.150 102.630 89.700 ;
        RECT 102.780 89.550 103.930 89.700 ;
        RECT 104.580 89.550 104.880 90.450 ;
        RECT 105.530 90.300 106.680 90.450 ;
        RECT 106.830 90.300 106.980 97.850 ;
        RECT 107.430 90.300 107.580 97.850 ;
        RECT 108.030 90.300 108.180 97.850 ;
        RECT 108.630 90.300 108.780 97.850 ;
        RECT 109.230 90.300 109.380 97.850 ;
        RECT 109.830 90.300 109.980 97.850 ;
        RECT 114.230 97.550 115.230 98.000 ;
        RECT 110.880 97.400 118.580 97.550 ;
        RECT 114.230 96.950 115.230 97.400 ;
        RECT 110.880 96.800 118.580 96.950 ;
        RECT 114.230 96.350 115.230 96.800 ;
        RECT 110.880 96.200 118.580 96.350 ;
        RECT 114.230 95.750 115.230 96.200 ;
        RECT 110.880 95.600 118.580 95.750 ;
        RECT 114.230 95.150 115.230 95.600 ;
        RECT 110.880 95.000 118.580 95.150 ;
        RECT 114.230 94.550 115.230 95.000 ;
        RECT 110.880 94.400 118.580 94.550 ;
        RECT 114.230 93.950 115.230 94.400 ;
        RECT 110.880 93.800 118.580 93.950 ;
        RECT 114.230 93.350 115.230 93.800 ;
        RECT 110.880 93.200 118.580 93.350 ;
        RECT 114.230 92.750 115.230 93.200 ;
        RECT 110.880 92.600 118.580 92.750 ;
        RECT 114.230 92.150 115.230 92.600 ;
        RECT 110.880 92.000 118.580 92.150 ;
        RECT 114.230 91.550 115.230 92.000 ;
        RECT 110.880 91.400 118.580 91.550 ;
        RECT 114.230 90.950 115.230 91.400 ;
        RECT 110.880 90.800 118.580 90.950 ;
        RECT 114.230 90.300 115.230 90.800 ;
        RECT 119.480 90.300 119.630 97.850 ;
        RECT 120.080 90.300 120.230 97.850 ;
        RECT 120.680 90.300 120.830 97.850 ;
        RECT 121.280 90.300 121.430 97.850 ;
        RECT 121.880 90.300 122.030 97.850 ;
        RECT 122.480 90.300 122.630 97.850 ;
        RECT 122.780 93.200 123.530 95.000 ;
        RECT 122.780 91.030 124.730 93.200 ;
        RECT 122.780 90.450 131.850 91.030 ;
        RECT 122.780 90.300 123.930 90.450 ;
        RECT 105.530 89.700 123.930 90.300 ;
        RECT 105.530 89.550 106.680 89.700 ;
        RECT 102.780 86.800 106.680 89.550 ;
        RECT 102.780 85.050 103.530 86.800 ;
        RECT 105.930 85.050 106.680 86.800 ;
        RECT 106.830 82.150 106.980 89.700 ;
        RECT 107.430 82.150 107.580 89.700 ;
        RECT 108.030 82.150 108.180 89.700 ;
        RECT 108.630 82.150 108.780 89.700 ;
        RECT 109.230 82.150 109.380 89.700 ;
        RECT 109.830 82.150 109.980 89.700 ;
        RECT 114.230 89.200 115.230 89.700 ;
        RECT 110.880 89.050 118.580 89.200 ;
        RECT 114.230 88.600 115.230 89.050 ;
        RECT 110.880 88.450 118.580 88.600 ;
        RECT 114.230 88.000 115.230 88.450 ;
        RECT 110.880 87.850 118.580 88.000 ;
        RECT 114.230 87.400 115.230 87.850 ;
        RECT 110.880 87.250 118.580 87.400 ;
        RECT 114.230 86.800 115.230 87.250 ;
        RECT 110.880 86.650 118.580 86.800 ;
        RECT 114.230 86.200 115.230 86.650 ;
        RECT 110.880 86.050 118.580 86.200 ;
        RECT 114.230 85.600 115.230 86.050 ;
        RECT 110.880 85.450 118.580 85.600 ;
        RECT 114.230 85.000 115.230 85.450 ;
        RECT 110.880 84.850 118.580 85.000 ;
        RECT 114.230 84.400 115.230 84.850 ;
        RECT 110.880 84.250 118.580 84.400 ;
        RECT 114.230 83.800 115.230 84.250 ;
        RECT 110.880 83.650 118.580 83.800 ;
        RECT 114.230 83.200 115.230 83.650 ;
        RECT 110.880 83.050 118.580 83.200 ;
        RECT 114.230 82.600 115.230 83.050 ;
        RECT 110.880 82.450 118.580 82.600 ;
        RECT 114.230 82.000 115.230 82.450 ;
        RECT 119.480 82.150 119.630 89.700 ;
        RECT 120.080 82.150 120.230 89.700 ;
        RECT 120.680 82.150 120.830 89.700 ;
        RECT 121.280 82.150 121.430 89.700 ;
        RECT 121.880 82.150 122.030 89.700 ;
        RECT 122.480 82.150 122.630 89.700 ;
        RECT 122.780 89.550 123.930 89.700 ;
        RECT 124.580 89.755 131.850 90.450 ;
        RECT 124.580 89.550 124.730 89.755 ;
        RECT 122.780 86.800 124.730 89.550 ;
        RECT 122.780 85.050 123.530 86.800 ;
        RECT 10.880 81.850 18.580 82.000 ;
        RECT 30.880 81.850 38.580 82.000 ;
        RECT 50.880 81.850 58.580 82.000 ;
        RECT 70.880 81.850 78.580 82.000 ;
        RECT 90.880 81.850 98.580 82.000 ;
        RECT 110.880 81.850 118.580 82.000 ;
        RECT 14.230 81.200 15.230 81.850 ;
        RECT 34.230 81.200 35.230 81.850 ;
        RECT 54.230 81.200 55.230 81.850 ;
        RECT 74.230 81.200 75.230 81.850 ;
        RECT 94.230 81.200 95.230 81.850 ;
        RECT 114.230 81.200 115.230 81.850 ;
        RECT 11.530 78.800 17.930 81.200 ;
        RECT 31.530 78.800 37.930 81.200 ;
        RECT 51.530 78.800 57.930 81.200 ;
        RECT 71.530 78.800 77.930 81.200 ;
        RECT 91.530 78.800 97.930 81.200 ;
        RECT 111.530 78.800 117.930 81.200 ;
        RECT 14.230 78.150 15.230 78.800 ;
        RECT 34.230 78.150 35.230 78.800 ;
        RECT 54.230 78.150 55.230 78.800 ;
        RECT 74.230 78.150 75.230 78.800 ;
        RECT 94.230 78.150 95.230 78.800 ;
        RECT 114.230 78.150 115.230 78.800 ;
        RECT 10.880 78.000 18.580 78.150 ;
        RECT 30.880 78.000 38.580 78.150 ;
        RECT 50.880 78.000 58.580 78.150 ;
        RECT 70.880 78.000 78.580 78.150 ;
        RECT 90.880 78.000 98.580 78.150 ;
        RECT 110.880 78.000 118.580 78.150 ;
        RECT 5.930 73.200 6.680 75.000 ;
        RECT 4.730 70.450 6.680 73.200 ;
        RECT 4.730 69.550 4.880 70.450 ;
        RECT 5.530 70.300 6.680 70.450 ;
        RECT 6.830 70.300 6.980 77.850 ;
        RECT 7.430 70.300 7.580 77.850 ;
        RECT 8.030 70.300 8.180 77.850 ;
        RECT 8.630 70.300 8.780 77.850 ;
        RECT 9.230 70.300 9.380 77.850 ;
        RECT 9.830 70.300 9.980 77.850 ;
        RECT 14.230 77.550 15.230 78.000 ;
        RECT 10.880 77.400 18.580 77.550 ;
        RECT 14.230 76.950 15.230 77.400 ;
        RECT 10.880 76.800 18.580 76.950 ;
        RECT 14.230 76.350 15.230 76.800 ;
        RECT 10.880 76.200 18.580 76.350 ;
        RECT 14.230 75.750 15.230 76.200 ;
        RECT 10.880 75.600 18.580 75.750 ;
        RECT 14.230 75.150 15.230 75.600 ;
        RECT 10.880 75.000 18.580 75.150 ;
        RECT 14.230 74.550 15.230 75.000 ;
        RECT 10.880 74.400 18.580 74.550 ;
        RECT 14.230 73.950 15.230 74.400 ;
        RECT 10.880 73.800 18.580 73.950 ;
        RECT 14.230 73.350 15.230 73.800 ;
        RECT 10.880 73.200 18.580 73.350 ;
        RECT 14.230 72.750 15.230 73.200 ;
        RECT 10.880 72.600 18.580 72.750 ;
        RECT 14.230 72.150 15.230 72.600 ;
        RECT 10.880 72.000 18.580 72.150 ;
        RECT 14.230 71.550 15.230 72.000 ;
        RECT 10.880 71.400 18.580 71.550 ;
        RECT 14.230 70.950 15.230 71.400 ;
        RECT 10.880 70.800 18.580 70.950 ;
        RECT 14.230 70.300 15.230 70.800 ;
        RECT 19.480 70.300 19.630 77.850 ;
        RECT 20.080 70.300 20.230 77.850 ;
        RECT 20.680 70.300 20.830 77.850 ;
        RECT 21.280 70.300 21.430 77.850 ;
        RECT 21.880 70.300 22.030 77.850 ;
        RECT 22.480 70.300 22.630 77.850 ;
        RECT 22.780 73.200 23.530 75.000 ;
        RECT 25.930 73.200 26.680 75.000 ;
        RECT 22.780 70.450 26.680 73.200 ;
        RECT 22.780 70.300 23.930 70.450 ;
        RECT 5.530 69.700 23.930 70.300 ;
        RECT 5.530 69.550 6.680 69.700 ;
        RECT 4.730 66.800 6.680 69.550 ;
        RECT 5.930 65.050 6.680 66.800 ;
        RECT 6.830 62.150 6.980 69.700 ;
        RECT 7.430 62.150 7.580 69.700 ;
        RECT 8.030 62.150 8.180 69.700 ;
        RECT 8.630 62.150 8.780 69.700 ;
        RECT 9.230 62.150 9.380 69.700 ;
        RECT 9.830 62.150 9.980 69.700 ;
        RECT 14.230 69.200 15.230 69.700 ;
        RECT 10.880 69.050 18.580 69.200 ;
        RECT 14.230 68.600 15.230 69.050 ;
        RECT 10.880 68.450 18.580 68.600 ;
        RECT 14.230 68.000 15.230 68.450 ;
        RECT 10.880 67.850 18.580 68.000 ;
        RECT 14.230 67.400 15.230 67.850 ;
        RECT 10.880 67.250 18.580 67.400 ;
        RECT 14.230 66.800 15.230 67.250 ;
        RECT 10.880 66.650 18.580 66.800 ;
        RECT 14.230 66.200 15.230 66.650 ;
        RECT 10.880 66.050 18.580 66.200 ;
        RECT 14.230 65.600 15.230 66.050 ;
        RECT 10.880 65.450 18.580 65.600 ;
        RECT 14.230 65.000 15.230 65.450 ;
        RECT 10.880 64.850 18.580 65.000 ;
        RECT 14.230 64.400 15.230 64.850 ;
        RECT 10.880 64.250 18.580 64.400 ;
        RECT 14.230 63.800 15.230 64.250 ;
        RECT 10.880 63.650 18.580 63.800 ;
        RECT 14.230 63.200 15.230 63.650 ;
        RECT 10.880 63.050 18.580 63.200 ;
        RECT 14.230 62.600 15.230 63.050 ;
        RECT 10.880 62.450 18.580 62.600 ;
        RECT 14.230 62.000 15.230 62.450 ;
        RECT 19.480 62.150 19.630 69.700 ;
        RECT 20.080 62.150 20.230 69.700 ;
        RECT 20.680 62.150 20.830 69.700 ;
        RECT 21.280 62.150 21.430 69.700 ;
        RECT 21.880 62.150 22.030 69.700 ;
        RECT 22.480 62.150 22.630 69.700 ;
        RECT 22.780 69.550 23.930 69.700 ;
        RECT 24.580 69.550 24.880 70.450 ;
        RECT 25.530 70.300 26.680 70.450 ;
        RECT 26.830 70.300 26.980 77.850 ;
        RECT 27.430 70.300 27.580 77.850 ;
        RECT 28.030 70.300 28.180 77.850 ;
        RECT 28.630 70.300 28.780 77.850 ;
        RECT 29.230 70.300 29.380 77.850 ;
        RECT 29.830 70.300 29.980 77.850 ;
        RECT 34.230 77.550 35.230 78.000 ;
        RECT 30.880 77.400 38.580 77.550 ;
        RECT 34.230 76.950 35.230 77.400 ;
        RECT 30.880 76.800 38.580 76.950 ;
        RECT 34.230 76.350 35.230 76.800 ;
        RECT 30.880 76.200 38.580 76.350 ;
        RECT 34.230 75.750 35.230 76.200 ;
        RECT 30.880 75.600 38.580 75.750 ;
        RECT 34.230 75.150 35.230 75.600 ;
        RECT 30.880 75.000 38.580 75.150 ;
        RECT 34.230 74.550 35.230 75.000 ;
        RECT 30.880 74.400 38.580 74.550 ;
        RECT 34.230 73.950 35.230 74.400 ;
        RECT 30.880 73.800 38.580 73.950 ;
        RECT 34.230 73.350 35.230 73.800 ;
        RECT 30.880 73.200 38.580 73.350 ;
        RECT 34.230 72.750 35.230 73.200 ;
        RECT 30.880 72.600 38.580 72.750 ;
        RECT 34.230 72.150 35.230 72.600 ;
        RECT 30.880 72.000 38.580 72.150 ;
        RECT 34.230 71.550 35.230 72.000 ;
        RECT 30.880 71.400 38.580 71.550 ;
        RECT 34.230 70.950 35.230 71.400 ;
        RECT 30.880 70.800 38.580 70.950 ;
        RECT 34.230 70.300 35.230 70.800 ;
        RECT 39.480 70.300 39.630 77.850 ;
        RECT 40.080 70.300 40.230 77.850 ;
        RECT 40.680 70.300 40.830 77.850 ;
        RECT 41.280 70.300 41.430 77.850 ;
        RECT 41.880 70.300 42.030 77.850 ;
        RECT 42.480 70.300 42.630 77.850 ;
        RECT 42.780 73.200 43.530 75.000 ;
        RECT 45.930 73.200 46.680 75.000 ;
        RECT 42.780 70.450 46.680 73.200 ;
        RECT 42.780 70.300 43.930 70.450 ;
        RECT 25.530 69.700 43.930 70.300 ;
        RECT 25.530 69.550 26.680 69.700 ;
        RECT 22.780 66.800 26.680 69.550 ;
        RECT 22.780 65.050 23.530 66.800 ;
        RECT 25.930 65.050 26.680 66.800 ;
        RECT 26.830 62.150 26.980 69.700 ;
        RECT 27.430 62.150 27.580 69.700 ;
        RECT 28.030 62.150 28.180 69.700 ;
        RECT 28.630 62.150 28.780 69.700 ;
        RECT 29.230 62.150 29.380 69.700 ;
        RECT 29.830 62.150 29.980 69.700 ;
        RECT 34.230 69.200 35.230 69.700 ;
        RECT 30.880 69.050 38.580 69.200 ;
        RECT 34.230 68.600 35.230 69.050 ;
        RECT 30.880 68.450 38.580 68.600 ;
        RECT 34.230 68.000 35.230 68.450 ;
        RECT 30.880 67.850 38.580 68.000 ;
        RECT 34.230 67.400 35.230 67.850 ;
        RECT 30.880 67.250 38.580 67.400 ;
        RECT 34.230 66.800 35.230 67.250 ;
        RECT 30.880 66.650 38.580 66.800 ;
        RECT 34.230 66.200 35.230 66.650 ;
        RECT 30.880 66.050 38.580 66.200 ;
        RECT 34.230 65.600 35.230 66.050 ;
        RECT 30.880 65.450 38.580 65.600 ;
        RECT 34.230 65.000 35.230 65.450 ;
        RECT 30.880 64.850 38.580 65.000 ;
        RECT 34.230 64.400 35.230 64.850 ;
        RECT 30.880 64.250 38.580 64.400 ;
        RECT 34.230 63.800 35.230 64.250 ;
        RECT 30.880 63.650 38.580 63.800 ;
        RECT 34.230 63.200 35.230 63.650 ;
        RECT 30.880 63.050 38.580 63.200 ;
        RECT 34.230 62.600 35.230 63.050 ;
        RECT 30.880 62.450 38.580 62.600 ;
        RECT 34.230 62.000 35.230 62.450 ;
        RECT 39.480 62.150 39.630 69.700 ;
        RECT 40.080 62.150 40.230 69.700 ;
        RECT 40.680 62.150 40.830 69.700 ;
        RECT 41.280 62.150 41.430 69.700 ;
        RECT 41.880 62.150 42.030 69.700 ;
        RECT 42.480 62.150 42.630 69.700 ;
        RECT 42.780 69.550 43.930 69.700 ;
        RECT 44.580 69.550 44.880 70.450 ;
        RECT 45.530 70.300 46.680 70.450 ;
        RECT 46.830 70.300 46.980 77.850 ;
        RECT 47.430 70.300 47.580 77.850 ;
        RECT 48.030 70.300 48.180 77.850 ;
        RECT 48.630 70.300 48.780 77.850 ;
        RECT 49.230 70.300 49.380 77.850 ;
        RECT 49.830 70.300 49.980 77.850 ;
        RECT 54.230 77.550 55.230 78.000 ;
        RECT 50.880 77.400 58.580 77.550 ;
        RECT 54.230 76.950 55.230 77.400 ;
        RECT 50.880 76.800 58.580 76.950 ;
        RECT 54.230 76.350 55.230 76.800 ;
        RECT 50.880 76.200 58.580 76.350 ;
        RECT 54.230 75.750 55.230 76.200 ;
        RECT 50.880 75.600 58.580 75.750 ;
        RECT 54.230 75.150 55.230 75.600 ;
        RECT 50.880 75.000 58.580 75.150 ;
        RECT 54.230 74.550 55.230 75.000 ;
        RECT 50.880 74.400 58.580 74.550 ;
        RECT 54.230 73.950 55.230 74.400 ;
        RECT 50.880 73.800 58.580 73.950 ;
        RECT 54.230 73.350 55.230 73.800 ;
        RECT 50.880 73.200 58.580 73.350 ;
        RECT 54.230 72.750 55.230 73.200 ;
        RECT 50.880 72.600 58.580 72.750 ;
        RECT 54.230 72.150 55.230 72.600 ;
        RECT 50.880 72.000 58.580 72.150 ;
        RECT 54.230 71.550 55.230 72.000 ;
        RECT 50.880 71.400 58.580 71.550 ;
        RECT 54.230 70.950 55.230 71.400 ;
        RECT 50.880 70.800 58.580 70.950 ;
        RECT 54.230 70.300 55.230 70.800 ;
        RECT 59.480 70.300 59.630 77.850 ;
        RECT 60.080 70.300 60.230 77.850 ;
        RECT 60.680 70.300 60.830 77.850 ;
        RECT 61.280 70.300 61.430 77.850 ;
        RECT 61.880 70.300 62.030 77.850 ;
        RECT 62.480 70.300 62.630 77.850 ;
        RECT 62.780 73.200 63.530 75.000 ;
        RECT 65.930 73.200 66.680 75.000 ;
        RECT 62.780 70.450 66.680 73.200 ;
        RECT 62.780 70.300 63.930 70.450 ;
        RECT 45.530 69.700 63.930 70.300 ;
        RECT 45.530 69.550 46.680 69.700 ;
        RECT 42.780 66.800 46.680 69.550 ;
        RECT 42.780 65.050 43.530 66.800 ;
        RECT 45.930 65.050 46.680 66.800 ;
        RECT 46.830 62.150 46.980 69.700 ;
        RECT 47.430 62.150 47.580 69.700 ;
        RECT 48.030 62.150 48.180 69.700 ;
        RECT 48.630 62.150 48.780 69.700 ;
        RECT 49.230 62.150 49.380 69.700 ;
        RECT 49.830 62.150 49.980 69.700 ;
        RECT 54.230 69.200 55.230 69.700 ;
        RECT 50.880 69.050 58.580 69.200 ;
        RECT 54.230 68.600 55.230 69.050 ;
        RECT 50.880 68.450 58.580 68.600 ;
        RECT 54.230 68.000 55.230 68.450 ;
        RECT 50.880 67.850 58.580 68.000 ;
        RECT 54.230 67.400 55.230 67.850 ;
        RECT 50.880 67.250 58.580 67.400 ;
        RECT 54.230 66.800 55.230 67.250 ;
        RECT 50.880 66.650 58.580 66.800 ;
        RECT 54.230 66.200 55.230 66.650 ;
        RECT 50.880 66.050 58.580 66.200 ;
        RECT 54.230 65.600 55.230 66.050 ;
        RECT 50.880 65.450 58.580 65.600 ;
        RECT 54.230 65.000 55.230 65.450 ;
        RECT 50.880 64.850 58.580 65.000 ;
        RECT 54.230 64.400 55.230 64.850 ;
        RECT 50.880 64.250 58.580 64.400 ;
        RECT 54.230 63.800 55.230 64.250 ;
        RECT 50.880 63.650 58.580 63.800 ;
        RECT 54.230 63.200 55.230 63.650 ;
        RECT 50.880 63.050 58.580 63.200 ;
        RECT 54.230 62.600 55.230 63.050 ;
        RECT 50.880 62.450 58.580 62.600 ;
        RECT 54.230 62.000 55.230 62.450 ;
        RECT 59.480 62.150 59.630 69.700 ;
        RECT 60.080 62.150 60.230 69.700 ;
        RECT 60.680 62.150 60.830 69.700 ;
        RECT 61.280 62.150 61.430 69.700 ;
        RECT 61.880 62.150 62.030 69.700 ;
        RECT 62.480 62.150 62.630 69.700 ;
        RECT 62.780 69.550 63.930 69.700 ;
        RECT 64.580 69.550 64.880 70.450 ;
        RECT 65.530 70.300 66.680 70.450 ;
        RECT 66.830 70.300 66.980 77.850 ;
        RECT 67.430 70.300 67.580 77.850 ;
        RECT 68.030 70.300 68.180 77.850 ;
        RECT 68.630 70.300 68.780 77.850 ;
        RECT 69.230 70.300 69.380 77.850 ;
        RECT 69.830 70.300 69.980 77.850 ;
        RECT 74.230 77.550 75.230 78.000 ;
        RECT 70.880 77.400 78.580 77.550 ;
        RECT 74.230 76.950 75.230 77.400 ;
        RECT 70.880 76.800 78.580 76.950 ;
        RECT 74.230 76.350 75.230 76.800 ;
        RECT 70.880 76.200 78.580 76.350 ;
        RECT 74.230 75.750 75.230 76.200 ;
        RECT 70.880 75.600 78.580 75.750 ;
        RECT 74.230 75.150 75.230 75.600 ;
        RECT 70.880 75.000 78.580 75.150 ;
        RECT 74.230 74.550 75.230 75.000 ;
        RECT 70.880 74.400 78.580 74.550 ;
        RECT 74.230 73.950 75.230 74.400 ;
        RECT 70.880 73.800 78.580 73.950 ;
        RECT 74.230 73.350 75.230 73.800 ;
        RECT 70.880 73.200 78.580 73.350 ;
        RECT 74.230 72.750 75.230 73.200 ;
        RECT 70.880 72.600 78.580 72.750 ;
        RECT 74.230 72.150 75.230 72.600 ;
        RECT 70.880 72.000 78.580 72.150 ;
        RECT 74.230 71.550 75.230 72.000 ;
        RECT 70.880 71.400 78.580 71.550 ;
        RECT 74.230 70.950 75.230 71.400 ;
        RECT 70.880 70.800 78.580 70.950 ;
        RECT 74.230 70.300 75.230 70.800 ;
        RECT 79.480 70.300 79.630 77.850 ;
        RECT 80.080 70.300 80.230 77.850 ;
        RECT 80.680 70.300 80.830 77.850 ;
        RECT 81.280 70.300 81.430 77.850 ;
        RECT 81.880 70.300 82.030 77.850 ;
        RECT 82.480 70.300 82.630 77.850 ;
        RECT 82.780 73.200 83.530 75.000 ;
        RECT 85.930 73.200 86.680 75.000 ;
        RECT 82.780 70.450 86.680 73.200 ;
        RECT 82.780 70.300 83.930 70.450 ;
        RECT 65.530 69.700 83.930 70.300 ;
        RECT 65.530 69.550 66.680 69.700 ;
        RECT 62.780 66.800 66.680 69.550 ;
        RECT 62.780 65.050 63.530 66.800 ;
        RECT 65.930 65.050 66.680 66.800 ;
        RECT 66.830 62.150 66.980 69.700 ;
        RECT 67.430 62.150 67.580 69.700 ;
        RECT 68.030 62.150 68.180 69.700 ;
        RECT 68.630 62.150 68.780 69.700 ;
        RECT 69.230 62.150 69.380 69.700 ;
        RECT 69.830 62.150 69.980 69.700 ;
        RECT 74.230 69.200 75.230 69.700 ;
        RECT 70.880 69.050 78.580 69.200 ;
        RECT 74.230 68.600 75.230 69.050 ;
        RECT 70.880 68.450 78.580 68.600 ;
        RECT 74.230 68.000 75.230 68.450 ;
        RECT 70.880 67.850 78.580 68.000 ;
        RECT 74.230 67.400 75.230 67.850 ;
        RECT 70.880 67.250 78.580 67.400 ;
        RECT 74.230 66.800 75.230 67.250 ;
        RECT 70.880 66.650 78.580 66.800 ;
        RECT 74.230 66.200 75.230 66.650 ;
        RECT 70.880 66.050 78.580 66.200 ;
        RECT 74.230 65.600 75.230 66.050 ;
        RECT 70.880 65.450 78.580 65.600 ;
        RECT 74.230 65.000 75.230 65.450 ;
        RECT 70.880 64.850 78.580 65.000 ;
        RECT 74.230 64.400 75.230 64.850 ;
        RECT 70.880 64.250 78.580 64.400 ;
        RECT 74.230 63.800 75.230 64.250 ;
        RECT 70.880 63.650 78.580 63.800 ;
        RECT 74.230 63.200 75.230 63.650 ;
        RECT 70.880 63.050 78.580 63.200 ;
        RECT 74.230 62.600 75.230 63.050 ;
        RECT 70.880 62.450 78.580 62.600 ;
        RECT 74.230 62.000 75.230 62.450 ;
        RECT 79.480 62.150 79.630 69.700 ;
        RECT 80.080 62.150 80.230 69.700 ;
        RECT 80.680 62.150 80.830 69.700 ;
        RECT 81.280 62.150 81.430 69.700 ;
        RECT 81.880 62.150 82.030 69.700 ;
        RECT 82.480 62.150 82.630 69.700 ;
        RECT 82.780 69.550 83.930 69.700 ;
        RECT 84.580 69.550 84.880 70.450 ;
        RECT 85.530 70.300 86.680 70.450 ;
        RECT 86.830 70.300 86.980 77.850 ;
        RECT 87.430 70.300 87.580 77.850 ;
        RECT 88.030 70.300 88.180 77.850 ;
        RECT 88.630 70.300 88.780 77.850 ;
        RECT 89.230 70.300 89.380 77.850 ;
        RECT 89.830 70.300 89.980 77.850 ;
        RECT 94.230 77.550 95.230 78.000 ;
        RECT 90.880 77.400 98.580 77.550 ;
        RECT 94.230 76.950 95.230 77.400 ;
        RECT 90.880 76.800 98.580 76.950 ;
        RECT 94.230 76.350 95.230 76.800 ;
        RECT 90.880 76.200 98.580 76.350 ;
        RECT 94.230 75.750 95.230 76.200 ;
        RECT 90.880 75.600 98.580 75.750 ;
        RECT 94.230 75.150 95.230 75.600 ;
        RECT 90.880 75.000 98.580 75.150 ;
        RECT 94.230 74.550 95.230 75.000 ;
        RECT 90.880 74.400 98.580 74.550 ;
        RECT 94.230 73.950 95.230 74.400 ;
        RECT 90.880 73.800 98.580 73.950 ;
        RECT 94.230 73.350 95.230 73.800 ;
        RECT 90.880 73.200 98.580 73.350 ;
        RECT 94.230 72.750 95.230 73.200 ;
        RECT 90.880 72.600 98.580 72.750 ;
        RECT 94.230 72.150 95.230 72.600 ;
        RECT 90.880 72.000 98.580 72.150 ;
        RECT 94.230 71.550 95.230 72.000 ;
        RECT 90.880 71.400 98.580 71.550 ;
        RECT 94.230 70.950 95.230 71.400 ;
        RECT 90.880 70.800 98.580 70.950 ;
        RECT 94.230 70.300 95.230 70.800 ;
        RECT 99.480 70.300 99.630 77.850 ;
        RECT 100.080 70.300 100.230 77.850 ;
        RECT 100.680 70.300 100.830 77.850 ;
        RECT 101.280 70.300 101.430 77.850 ;
        RECT 101.880 70.300 102.030 77.850 ;
        RECT 102.480 70.300 102.630 77.850 ;
        RECT 102.780 73.200 103.530 75.000 ;
        RECT 105.930 73.200 106.680 75.000 ;
        RECT 102.780 70.450 106.680 73.200 ;
        RECT 102.780 70.300 103.930 70.450 ;
        RECT 85.530 69.700 103.930 70.300 ;
        RECT 85.530 69.550 86.680 69.700 ;
        RECT 82.780 66.800 86.680 69.550 ;
        RECT 82.780 65.050 83.530 66.800 ;
        RECT 85.930 65.050 86.680 66.800 ;
        RECT 86.830 62.150 86.980 69.700 ;
        RECT 87.430 62.150 87.580 69.700 ;
        RECT 88.030 62.150 88.180 69.700 ;
        RECT 88.630 62.150 88.780 69.700 ;
        RECT 89.230 62.150 89.380 69.700 ;
        RECT 89.830 62.150 89.980 69.700 ;
        RECT 94.230 69.200 95.230 69.700 ;
        RECT 90.880 69.050 98.580 69.200 ;
        RECT 94.230 68.600 95.230 69.050 ;
        RECT 90.880 68.450 98.580 68.600 ;
        RECT 94.230 68.000 95.230 68.450 ;
        RECT 90.880 67.850 98.580 68.000 ;
        RECT 94.230 67.400 95.230 67.850 ;
        RECT 90.880 67.250 98.580 67.400 ;
        RECT 94.230 66.800 95.230 67.250 ;
        RECT 90.880 66.650 98.580 66.800 ;
        RECT 94.230 66.200 95.230 66.650 ;
        RECT 90.880 66.050 98.580 66.200 ;
        RECT 94.230 65.600 95.230 66.050 ;
        RECT 90.880 65.450 98.580 65.600 ;
        RECT 94.230 65.000 95.230 65.450 ;
        RECT 90.880 64.850 98.580 65.000 ;
        RECT 94.230 64.400 95.230 64.850 ;
        RECT 90.880 64.250 98.580 64.400 ;
        RECT 94.230 63.800 95.230 64.250 ;
        RECT 90.880 63.650 98.580 63.800 ;
        RECT 94.230 63.200 95.230 63.650 ;
        RECT 90.880 63.050 98.580 63.200 ;
        RECT 94.230 62.600 95.230 63.050 ;
        RECT 90.880 62.450 98.580 62.600 ;
        RECT 94.230 62.000 95.230 62.450 ;
        RECT 99.480 62.150 99.630 69.700 ;
        RECT 100.080 62.150 100.230 69.700 ;
        RECT 100.680 62.150 100.830 69.700 ;
        RECT 101.280 62.150 101.430 69.700 ;
        RECT 101.880 62.150 102.030 69.700 ;
        RECT 102.480 62.150 102.630 69.700 ;
        RECT 102.780 69.550 103.930 69.700 ;
        RECT 104.580 69.550 104.880 70.450 ;
        RECT 105.530 70.300 106.680 70.450 ;
        RECT 106.830 70.300 106.980 77.850 ;
        RECT 107.430 70.300 107.580 77.850 ;
        RECT 108.030 70.300 108.180 77.850 ;
        RECT 108.630 70.300 108.780 77.850 ;
        RECT 109.230 70.300 109.380 77.850 ;
        RECT 109.830 70.300 109.980 77.850 ;
        RECT 114.230 77.550 115.230 78.000 ;
        RECT 110.880 77.400 118.580 77.550 ;
        RECT 114.230 76.950 115.230 77.400 ;
        RECT 110.880 76.800 118.580 76.950 ;
        RECT 114.230 76.350 115.230 76.800 ;
        RECT 110.880 76.200 118.580 76.350 ;
        RECT 114.230 75.750 115.230 76.200 ;
        RECT 110.880 75.600 118.580 75.750 ;
        RECT 114.230 75.150 115.230 75.600 ;
        RECT 110.880 75.000 118.580 75.150 ;
        RECT 114.230 74.550 115.230 75.000 ;
        RECT 110.880 74.400 118.580 74.550 ;
        RECT 114.230 73.950 115.230 74.400 ;
        RECT 110.880 73.800 118.580 73.950 ;
        RECT 114.230 73.350 115.230 73.800 ;
        RECT 110.880 73.200 118.580 73.350 ;
        RECT 114.230 72.750 115.230 73.200 ;
        RECT 110.880 72.600 118.580 72.750 ;
        RECT 114.230 72.150 115.230 72.600 ;
        RECT 110.880 72.000 118.580 72.150 ;
        RECT 114.230 71.550 115.230 72.000 ;
        RECT 110.880 71.400 118.580 71.550 ;
        RECT 114.230 70.950 115.230 71.400 ;
        RECT 110.880 70.800 118.580 70.950 ;
        RECT 114.230 70.300 115.230 70.800 ;
        RECT 119.480 70.300 119.630 77.850 ;
        RECT 120.080 70.300 120.230 77.850 ;
        RECT 120.680 70.300 120.830 77.850 ;
        RECT 121.280 70.300 121.430 77.850 ;
        RECT 121.880 70.300 122.030 77.850 ;
        RECT 122.480 70.300 122.630 77.850 ;
        RECT 122.780 73.200 123.530 75.000 ;
        RECT 122.780 70.495 124.730 73.200 ;
        RECT 122.780 70.450 131.850 70.495 ;
        RECT 122.780 70.300 123.930 70.450 ;
        RECT 105.530 69.700 123.930 70.300 ;
        RECT 105.530 69.550 106.680 69.700 ;
        RECT 102.780 66.800 106.680 69.550 ;
        RECT 102.780 65.050 103.530 66.800 ;
        RECT 105.930 65.050 106.680 66.800 ;
        RECT 106.830 62.150 106.980 69.700 ;
        RECT 107.430 62.150 107.580 69.700 ;
        RECT 108.030 62.150 108.180 69.700 ;
        RECT 108.630 62.150 108.780 69.700 ;
        RECT 109.230 62.150 109.380 69.700 ;
        RECT 109.830 62.150 109.980 69.700 ;
        RECT 114.230 69.200 115.230 69.700 ;
        RECT 110.880 69.050 118.580 69.200 ;
        RECT 114.230 68.600 115.230 69.050 ;
        RECT 110.880 68.450 118.580 68.600 ;
        RECT 114.230 68.000 115.230 68.450 ;
        RECT 110.880 67.850 118.580 68.000 ;
        RECT 114.230 67.400 115.230 67.850 ;
        RECT 110.880 67.250 118.580 67.400 ;
        RECT 114.230 66.800 115.230 67.250 ;
        RECT 110.880 66.650 118.580 66.800 ;
        RECT 114.230 66.200 115.230 66.650 ;
        RECT 110.880 66.050 118.580 66.200 ;
        RECT 114.230 65.600 115.230 66.050 ;
        RECT 110.880 65.450 118.580 65.600 ;
        RECT 114.230 65.000 115.230 65.450 ;
        RECT 110.880 64.850 118.580 65.000 ;
        RECT 114.230 64.400 115.230 64.850 ;
        RECT 110.880 64.250 118.580 64.400 ;
        RECT 114.230 63.800 115.230 64.250 ;
        RECT 110.880 63.650 118.580 63.800 ;
        RECT 114.230 63.200 115.230 63.650 ;
        RECT 110.880 63.050 118.580 63.200 ;
        RECT 114.230 62.600 115.230 63.050 ;
        RECT 110.880 62.450 118.580 62.600 ;
        RECT 114.230 62.000 115.230 62.450 ;
        RECT 119.480 62.150 119.630 69.700 ;
        RECT 120.080 62.150 120.230 69.700 ;
        RECT 120.680 62.150 120.830 69.700 ;
        RECT 121.280 62.150 121.430 69.700 ;
        RECT 121.880 62.150 122.030 69.700 ;
        RECT 122.480 62.150 122.630 69.700 ;
        RECT 122.780 69.550 123.930 69.700 ;
        RECT 124.580 69.550 131.850 70.450 ;
        RECT 122.780 69.220 131.850 69.550 ;
        RECT 122.780 66.800 124.730 69.220 ;
        RECT 122.780 65.050 123.530 66.800 ;
        RECT 10.880 61.850 18.580 62.000 ;
        RECT 30.880 61.850 38.580 62.000 ;
        RECT 50.880 61.850 58.580 62.000 ;
        RECT 70.880 61.850 78.580 62.000 ;
        RECT 90.880 61.850 98.580 62.000 ;
        RECT 110.880 61.850 118.580 62.000 ;
        RECT 14.230 61.200 15.230 61.850 ;
        RECT 34.230 61.200 35.230 61.850 ;
        RECT 54.230 61.200 55.230 61.850 ;
        RECT 74.230 61.200 75.230 61.850 ;
        RECT 94.230 61.200 95.230 61.850 ;
        RECT 114.230 61.200 115.230 61.850 ;
        RECT 11.530 58.800 17.930 61.200 ;
        RECT 31.530 58.800 37.930 61.200 ;
        RECT 51.530 58.800 57.930 61.200 ;
        RECT 71.530 58.800 77.930 61.200 ;
        RECT 91.530 58.800 97.930 61.200 ;
        RECT 111.530 58.800 117.930 61.200 ;
        RECT 14.230 58.150 15.230 58.800 ;
        RECT 34.230 58.150 35.230 58.800 ;
        RECT 54.230 58.150 55.230 58.800 ;
        RECT 74.230 58.150 75.230 58.800 ;
        RECT 94.230 58.150 95.230 58.800 ;
        RECT 114.230 58.150 115.230 58.800 ;
        RECT 10.880 58.000 18.580 58.150 ;
        RECT 30.880 58.000 38.580 58.150 ;
        RECT 50.880 58.000 58.580 58.150 ;
        RECT 70.880 58.000 78.580 58.150 ;
        RECT 90.880 58.000 98.580 58.150 ;
        RECT 110.880 58.000 118.580 58.150 ;
        RECT 5.930 53.200 6.680 55.000 ;
        RECT 4.730 50.450 6.680 53.200 ;
        RECT 4.730 49.550 4.880 50.450 ;
        RECT 5.530 50.300 6.680 50.450 ;
        RECT 6.830 50.300 6.980 57.850 ;
        RECT 7.430 50.300 7.580 57.850 ;
        RECT 8.030 50.300 8.180 57.850 ;
        RECT 8.630 50.300 8.780 57.850 ;
        RECT 9.230 50.300 9.380 57.850 ;
        RECT 9.830 50.300 9.980 57.850 ;
        RECT 14.230 57.550 15.230 58.000 ;
        RECT 10.880 57.400 18.580 57.550 ;
        RECT 14.230 56.950 15.230 57.400 ;
        RECT 10.880 56.800 18.580 56.950 ;
        RECT 14.230 56.350 15.230 56.800 ;
        RECT 10.880 56.200 18.580 56.350 ;
        RECT 14.230 55.750 15.230 56.200 ;
        RECT 10.880 55.600 18.580 55.750 ;
        RECT 14.230 55.150 15.230 55.600 ;
        RECT 10.880 55.000 18.580 55.150 ;
        RECT 14.230 54.550 15.230 55.000 ;
        RECT 10.880 54.400 18.580 54.550 ;
        RECT 14.230 53.950 15.230 54.400 ;
        RECT 10.880 53.800 18.580 53.950 ;
        RECT 14.230 53.350 15.230 53.800 ;
        RECT 10.880 53.200 18.580 53.350 ;
        RECT 14.230 52.750 15.230 53.200 ;
        RECT 10.880 52.600 18.580 52.750 ;
        RECT 14.230 52.150 15.230 52.600 ;
        RECT 10.880 52.000 18.580 52.150 ;
        RECT 14.230 51.550 15.230 52.000 ;
        RECT 10.880 51.400 18.580 51.550 ;
        RECT 14.230 50.950 15.230 51.400 ;
        RECT 10.880 50.800 18.580 50.950 ;
        RECT 14.230 50.300 15.230 50.800 ;
        RECT 19.480 50.300 19.630 57.850 ;
        RECT 20.080 50.300 20.230 57.850 ;
        RECT 20.680 50.300 20.830 57.850 ;
        RECT 21.280 50.300 21.430 57.850 ;
        RECT 21.880 50.300 22.030 57.850 ;
        RECT 22.480 50.300 22.630 57.850 ;
        RECT 22.780 53.200 23.530 55.000 ;
        RECT 25.930 53.200 26.680 55.000 ;
        RECT 22.780 50.450 26.680 53.200 ;
        RECT 22.780 50.300 23.930 50.450 ;
        RECT 5.530 49.700 23.930 50.300 ;
        RECT 5.530 49.550 6.680 49.700 ;
        RECT 4.730 46.800 6.680 49.550 ;
        RECT 5.930 45.050 6.680 46.800 ;
        RECT 6.830 42.150 6.980 49.700 ;
        RECT 7.430 42.150 7.580 49.700 ;
        RECT 8.030 42.150 8.180 49.700 ;
        RECT 8.630 42.150 8.780 49.700 ;
        RECT 9.230 42.150 9.380 49.700 ;
        RECT 9.830 42.150 9.980 49.700 ;
        RECT 14.230 49.200 15.230 49.700 ;
        RECT 10.880 49.050 18.580 49.200 ;
        RECT 14.230 48.600 15.230 49.050 ;
        RECT 10.880 48.450 18.580 48.600 ;
        RECT 14.230 48.000 15.230 48.450 ;
        RECT 10.880 47.850 18.580 48.000 ;
        RECT 14.230 47.400 15.230 47.850 ;
        RECT 10.880 47.250 18.580 47.400 ;
        RECT 14.230 46.800 15.230 47.250 ;
        RECT 10.880 46.650 18.580 46.800 ;
        RECT 14.230 46.200 15.230 46.650 ;
        RECT 10.880 46.050 18.580 46.200 ;
        RECT 14.230 45.600 15.230 46.050 ;
        RECT 10.880 45.450 18.580 45.600 ;
        RECT 14.230 45.000 15.230 45.450 ;
        RECT 10.880 44.850 18.580 45.000 ;
        RECT 14.230 44.400 15.230 44.850 ;
        RECT 10.880 44.250 18.580 44.400 ;
        RECT 14.230 43.800 15.230 44.250 ;
        RECT 10.880 43.650 18.580 43.800 ;
        RECT 14.230 43.200 15.230 43.650 ;
        RECT 10.880 43.050 18.580 43.200 ;
        RECT 14.230 42.600 15.230 43.050 ;
        RECT 10.880 42.450 18.580 42.600 ;
        RECT 14.230 42.000 15.230 42.450 ;
        RECT 19.480 42.150 19.630 49.700 ;
        RECT 20.080 42.150 20.230 49.700 ;
        RECT 20.680 42.150 20.830 49.700 ;
        RECT 21.280 42.150 21.430 49.700 ;
        RECT 21.880 42.150 22.030 49.700 ;
        RECT 22.480 42.150 22.630 49.700 ;
        RECT 22.780 49.550 23.930 49.700 ;
        RECT 24.580 49.550 24.880 50.450 ;
        RECT 25.530 50.300 26.680 50.450 ;
        RECT 26.830 50.300 26.980 57.850 ;
        RECT 27.430 50.300 27.580 57.850 ;
        RECT 28.030 50.300 28.180 57.850 ;
        RECT 28.630 50.300 28.780 57.850 ;
        RECT 29.230 50.300 29.380 57.850 ;
        RECT 29.830 50.300 29.980 57.850 ;
        RECT 34.230 57.550 35.230 58.000 ;
        RECT 30.880 57.400 38.580 57.550 ;
        RECT 34.230 56.950 35.230 57.400 ;
        RECT 30.880 56.800 38.580 56.950 ;
        RECT 34.230 56.350 35.230 56.800 ;
        RECT 30.880 56.200 38.580 56.350 ;
        RECT 34.230 55.750 35.230 56.200 ;
        RECT 30.880 55.600 38.580 55.750 ;
        RECT 34.230 55.150 35.230 55.600 ;
        RECT 30.880 55.000 38.580 55.150 ;
        RECT 34.230 54.550 35.230 55.000 ;
        RECT 30.880 54.400 38.580 54.550 ;
        RECT 34.230 53.950 35.230 54.400 ;
        RECT 30.880 53.800 38.580 53.950 ;
        RECT 34.230 53.350 35.230 53.800 ;
        RECT 30.880 53.200 38.580 53.350 ;
        RECT 34.230 52.750 35.230 53.200 ;
        RECT 30.880 52.600 38.580 52.750 ;
        RECT 34.230 52.150 35.230 52.600 ;
        RECT 30.880 52.000 38.580 52.150 ;
        RECT 34.230 51.550 35.230 52.000 ;
        RECT 30.880 51.400 38.580 51.550 ;
        RECT 34.230 50.950 35.230 51.400 ;
        RECT 30.880 50.800 38.580 50.950 ;
        RECT 34.230 50.300 35.230 50.800 ;
        RECT 39.480 50.300 39.630 57.850 ;
        RECT 40.080 50.300 40.230 57.850 ;
        RECT 40.680 50.300 40.830 57.850 ;
        RECT 41.280 50.300 41.430 57.850 ;
        RECT 41.880 50.300 42.030 57.850 ;
        RECT 42.480 50.300 42.630 57.850 ;
        RECT 42.780 53.200 43.530 55.000 ;
        RECT 45.930 53.200 46.680 55.000 ;
        RECT 42.780 50.450 46.680 53.200 ;
        RECT 42.780 50.300 43.930 50.450 ;
        RECT 25.530 49.700 43.930 50.300 ;
        RECT 25.530 49.550 26.680 49.700 ;
        RECT 22.780 46.800 26.680 49.550 ;
        RECT 22.780 45.050 23.530 46.800 ;
        RECT 25.930 45.050 26.680 46.800 ;
        RECT 26.830 42.150 26.980 49.700 ;
        RECT 27.430 42.150 27.580 49.700 ;
        RECT 28.030 42.150 28.180 49.700 ;
        RECT 28.630 42.150 28.780 49.700 ;
        RECT 29.230 42.150 29.380 49.700 ;
        RECT 29.830 42.150 29.980 49.700 ;
        RECT 34.230 49.200 35.230 49.700 ;
        RECT 30.880 49.050 38.580 49.200 ;
        RECT 34.230 48.600 35.230 49.050 ;
        RECT 30.880 48.450 38.580 48.600 ;
        RECT 34.230 48.000 35.230 48.450 ;
        RECT 30.880 47.850 38.580 48.000 ;
        RECT 34.230 47.400 35.230 47.850 ;
        RECT 30.880 47.250 38.580 47.400 ;
        RECT 34.230 46.800 35.230 47.250 ;
        RECT 30.880 46.650 38.580 46.800 ;
        RECT 34.230 46.200 35.230 46.650 ;
        RECT 30.880 46.050 38.580 46.200 ;
        RECT 34.230 45.600 35.230 46.050 ;
        RECT 30.880 45.450 38.580 45.600 ;
        RECT 34.230 45.000 35.230 45.450 ;
        RECT 30.880 44.850 38.580 45.000 ;
        RECT 34.230 44.400 35.230 44.850 ;
        RECT 30.880 44.250 38.580 44.400 ;
        RECT 34.230 43.800 35.230 44.250 ;
        RECT 30.880 43.650 38.580 43.800 ;
        RECT 34.230 43.200 35.230 43.650 ;
        RECT 30.880 43.050 38.580 43.200 ;
        RECT 34.230 42.600 35.230 43.050 ;
        RECT 30.880 42.450 38.580 42.600 ;
        RECT 34.230 42.000 35.230 42.450 ;
        RECT 39.480 42.150 39.630 49.700 ;
        RECT 40.080 42.150 40.230 49.700 ;
        RECT 40.680 42.150 40.830 49.700 ;
        RECT 41.280 42.150 41.430 49.700 ;
        RECT 41.880 42.150 42.030 49.700 ;
        RECT 42.480 42.150 42.630 49.700 ;
        RECT 42.780 49.550 43.930 49.700 ;
        RECT 44.580 49.550 44.880 50.450 ;
        RECT 45.530 50.300 46.680 50.450 ;
        RECT 46.830 50.300 46.980 57.850 ;
        RECT 47.430 50.300 47.580 57.850 ;
        RECT 48.030 50.300 48.180 57.850 ;
        RECT 48.630 50.300 48.780 57.850 ;
        RECT 49.230 50.300 49.380 57.850 ;
        RECT 49.830 50.300 49.980 57.850 ;
        RECT 54.230 57.550 55.230 58.000 ;
        RECT 50.880 57.400 58.580 57.550 ;
        RECT 54.230 56.950 55.230 57.400 ;
        RECT 50.880 56.800 58.580 56.950 ;
        RECT 54.230 56.350 55.230 56.800 ;
        RECT 50.880 56.200 58.580 56.350 ;
        RECT 54.230 55.750 55.230 56.200 ;
        RECT 50.880 55.600 58.580 55.750 ;
        RECT 54.230 55.150 55.230 55.600 ;
        RECT 50.880 55.000 58.580 55.150 ;
        RECT 54.230 54.550 55.230 55.000 ;
        RECT 50.880 54.400 58.580 54.550 ;
        RECT 54.230 53.950 55.230 54.400 ;
        RECT 50.880 53.800 58.580 53.950 ;
        RECT 54.230 53.350 55.230 53.800 ;
        RECT 50.880 53.200 58.580 53.350 ;
        RECT 54.230 52.750 55.230 53.200 ;
        RECT 50.880 52.600 58.580 52.750 ;
        RECT 54.230 52.150 55.230 52.600 ;
        RECT 50.880 52.000 58.580 52.150 ;
        RECT 54.230 51.550 55.230 52.000 ;
        RECT 50.880 51.400 58.580 51.550 ;
        RECT 54.230 50.950 55.230 51.400 ;
        RECT 50.880 50.800 58.580 50.950 ;
        RECT 54.230 50.300 55.230 50.800 ;
        RECT 59.480 50.300 59.630 57.850 ;
        RECT 60.080 50.300 60.230 57.850 ;
        RECT 60.680 50.300 60.830 57.850 ;
        RECT 61.280 50.300 61.430 57.850 ;
        RECT 61.880 50.300 62.030 57.850 ;
        RECT 62.480 50.300 62.630 57.850 ;
        RECT 62.780 53.200 63.530 55.000 ;
        RECT 65.930 53.200 66.680 55.000 ;
        RECT 62.780 50.450 66.680 53.200 ;
        RECT 62.780 50.300 63.930 50.450 ;
        RECT 45.530 49.700 63.930 50.300 ;
        RECT 45.530 49.550 46.680 49.700 ;
        RECT 42.780 46.800 46.680 49.550 ;
        RECT 42.780 45.050 43.530 46.800 ;
        RECT 45.930 45.050 46.680 46.800 ;
        RECT 46.830 42.150 46.980 49.700 ;
        RECT 47.430 42.150 47.580 49.700 ;
        RECT 48.030 42.150 48.180 49.700 ;
        RECT 48.630 42.150 48.780 49.700 ;
        RECT 49.230 42.150 49.380 49.700 ;
        RECT 49.830 42.150 49.980 49.700 ;
        RECT 54.230 49.200 55.230 49.700 ;
        RECT 50.880 49.050 58.580 49.200 ;
        RECT 54.230 48.600 55.230 49.050 ;
        RECT 50.880 48.450 58.580 48.600 ;
        RECT 54.230 48.000 55.230 48.450 ;
        RECT 50.880 47.850 58.580 48.000 ;
        RECT 54.230 47.400 55.230 47.850 ;
        RECT 50.880 47.250 58.580 47.400 ;
        RECT 54.230 46.800 55.230 47.250 ;
        RECT 50.880 46.650 58.580 46.800 ;
        RECT 54.230 46.200 55.230 46.650 ;
        RECT 50.880 46.050 58.580 46.200 ;
        RECT 54.230 45.600 55.230 46.050 ;
        RECT 50.880 45.450 58.580 45.600 ;
        RECT 54.230 45.000 55.230 45.450 ;
        RECT 50.880 44.850 58.580 45.000 ;
        RECT 54.230 44.400 55.230 44.850 ;
        RECT 50.880 44.250 58.580 44.400 ;
        RECT 54.230 43.800 55.230 44.250 ;
        RECT 50.880 43.650 58.580 43.800 ;
        RECT 54.230 43.200 55.230 43.650 ;
        RECT 50.880 43.050 58.580 43.200 ;
        RECT 54.230 42.600 55.230 43.050 ;
        RECT 50.880 42.450 58.580 42.600 ;
        RECT 54.230 42.000 55.230 42.450 ;
        RECT 59.480 42.150 59.630 49.700 ;
        RECT 60.080 42.150 60.230 49.700 ;
        RECT 60.680 42.150 60.830 49.700 ;
        RECT 61.280 42.150 61.430 49.700 ;
        RECT 61.880 42.150 62.030 49.700 ;
        RECT 62.480 42.150 62.630 49.700 ;
        RECT 62.780 49.550 63.930 49.700 ;
        RECT 64.580 49.550 64.880 50.450 ;
        RECT 65.530 50.300 66.680 50.450 ;
        RECT 66.830 50.300 66.980 57.850 ;
        RECT 67.430 50.300 67.580 57.850 ;
        RECT 68.030 50.300 68.180 57.850 ;
        RECT 68.630 50.300 68.780 57.850 ;
        RECT 69.230 50.300 69.380 57.850 ;
        RECT 69.830 50.300 69.980 57.850 ;
        RECT 74.230 57.550 75.230 58.000 ;
        RECT 70.880 57.400 78.580 57.550 ;
        RECT 74.230 56.950 75.230 57.400 ;
        RECT 70.880 56.800 78.580 56.950 ;
        RECT 74.230 56.350 75.230 56.800 ;
        RECT 70.880 56.200 78.580 56.350 ;
        RECT 74.230 55.750 75.230 56.200 ;
        RECT 70.880 55.600 78.580 55.750 ;
        RECT 74.230 55.150 75.230 55.600 ;
        RECT 70.880 55.000 78.580 55.150 ;
        RECT 74.230 54.550 75.230 55.000 ;
        RECT 70.880 54.400 78.580 54.550 ;
        RECT 74.230 53.950 75.230 54.400 ;
        RECT 70.880 53.800 78.580 53.950 ;
        RECT 74.230 53.350 75.230 53.800 ;
        RECT 70.880 53.200 78.580 53.350 ;
        RECT 74.230 52.750 75.230 53.200 ;
        RECT 70.880 52.600 78.580 52.750 ;
        RECT 74.230 52.150 75.230 52.600 ;
        RECT 70.880 52.000 78.580 52.150 ;
        RECT 74.230 51.550 75.230 52.000 ;
        RECT 70.880 51.400 78.580 51.550 ;
        RECT 74.230 50.950 75.230 51.400 ;
        RECT 70.880 50.800 78.580 50.950 ;
        RECT 74.230 50.300 75.230 50.800 ;
        RECT 79.480 50.300 79.630 57.850 ;
        RECT 80.080 50.300 80.230 57.850 ;
        RECT 80.680 50.300 80.830 57.850 ;
        RECT 81.280 50.300 81.430 57.850 ;
        RECT 81.880 50.300 82.030 57.850 ;
        RECT 82.480 50.300 82.630 57.850 ;
        RECT 82.780 53.200 83.530 55.000 ;
        RECT 85.930 53.200 86.680 55.000 ;
        RECT 82.780 50.450 86.680 53.200 ;
        RECT 82.780 50.300 83.930 50.450 ;
        RECT 65.530 49.700 83.930 50.300 ;
        RECT 65.530 49.550 66.680 49.700 ;
        RECT 62.780 46.800 66.680 49.550 ;
        RECT 62.780 45.050 63.530 46.800 ;
        RECT 65.930 45.050 66.680 46.800 ;
        RECT 66.830 42.150 66.980 49.700 ;
        RECT 67.430 42.150 67.580 49.700 ;
        RECT 68.030 42.150 68.180 49.700 ;
        RECT 68.630 42.150 68.780 49.700 ;
        RECT 69.230 42.150 69.380 49.700 ;
        RECT 69.830 42.150 69.980 49.700 ;
        RECT 74.230 49.200 75.230 49.700 ;
        RECT 70.880 49.050 78.580 49.200 ;
        RECT 74.230 48.600 75.230 49.050 ;
        RECT 70.880 48.450 78.580 48.600 ;
        RECT 74.230 48.000 75.230 48.450 ;
        RECT 70.880 47.850 78.580 48.000 ;
        RECT 74.230 47.400 75.230 47.850 ;
        RECT 70.880 47.250 78.580 47.400 ;
        RECT 74.230 46.800 75.230 47.250 ;
        RECT 70.880 46.650 78.580 46.800 ;
        RECT 74.230 46.200 75.230 46.650 ;
        RECT 70.880 46.050 78.580 46.200 ;
        RECT 74.230 45.600 75.230 46.050 ;
        RECT 70.880 45.450 78.580 45.600 ;
        RECT 74.230 45.000 75.230 45.450 ;
        RECT 70.880 44.850 78.580 45.000 ;
        RECT 74.230 44.400 75.230 44.850 ;
        RECT 70.880 44.250 78.580 44.400 ;
        RECT 74.230 43.800 75.230 44.250 ;
        RECT 70.880 43.650 78.580 43.800 ;
        RECT 74.230 43.200 75.230 43.650 ;
        RECT 70.880 43.050 78.580 43.200 ;
        RECT 74.230 42.600 75.230 43.050 ;
        RECT 70.880 42.450 78.580 42.600 ;
        RECT 74.230 42.000 75.230 42.450 ;
        RECT 79.480 42.150 79.630 49.700 ;
        RECT 80.080 42.150 80.230 49.700 ;
        RECT 80.680 42.150 80.830 49.700 ;
        RECT 81.280 42.150 81.430 49.700 ;
        RECT 81.880 42.150 82.030 49.700 ;
        RECT 82.480 42.150 82.630 49.700 ;
        RECT 82.780 49.550 83.930 49.700 ;
        RECT 84.580 49.550 84.880 50.450 ;
        RECT 85.530 50.300 86.680 50.450 ;
        RECT 86.830 50.300 86.980 57.850 ;
        RECT 87.430 50.300 87.580 57.850 ;
        RECT 88.030 50.300 88.180 57.850 ;
        RECT 88.630 50.300 88.780 57.850 ;
        RECT 89.230 50.300 89.380 57.850 ;
        RECT 89.830 50.300 89.980 57.850 ;
        RECT 94.230 57.550 95.230 58.000 ;
        RECT 90.880 57.400 98.580 57.550 ;
        RECT 94.230 56.950 95.230 57.400 ;
        RECT 90.880 56.800 98.580 56.950 ;
        RECT 94.230 56.350 95.230 56.800 ;
        RECT 90.880 56.200 98.580 56.350 ;
        RECT 94.230 55.750 95.230 56.200 ;
        RECT 90.880 55.600 98.580 55.750 ;
        RECT 94.230 55.150 95.230 55.600 ;
        RECT 90.880 55.000 98.580 55.150 ;
        RECT 94.230 54.550 95.230 55.000 ;
        RECT 90.880 54.400 98.580 54.550 ;
        RECT 94.230 53.950 95.230 54.400 ;
        RECT 90.880 53.800 98.580 53.950 ;
        RECT 94.230 53.350 95.230 53.800 ;
        RECT 90.880 53.200 98.580 53.350 ;
        RECT 94.230 52.750 95.230 53.200 ;
        RECT 90.880 52.600 98.580 52.750 ;
        RECT 94.230 52.150 95.230 52.600 ;
        RECT 90.880 52.000 98.580 52.150 ;
        RECT 94.230 51.550 95.230 52.000 ;
        RECT 90.880 51.400 98.580 51.550 ;
        RECT 94.230 50.950 95.230 51.400 ;
        RECT 90.880 50.800 98.580 50.950 ;
        RECT 94.230 50.300 95.230 50.800 ;
        RECT 99.480 50.300 99.630 57.850 ;
        RECT 100.080 50.300 100.230 57.850 ;
        RECT 100.680 50.300 100.830 57.850 ;
        RECT 101.280 50.300 101.430 57.850 ;
        RECT 101.880 50.300 102.030 57.850 ;
        RECT 102.480 50.300 102.630 57.850 ;
        RECT 102.780 53.200 103.530 55.000 ;
        RECT 105.930 53.200 106.680 55.000 ;
        RECT 102.780 50.450 106.680 53.200 ;
        RECT 102.780 50.300 103.930 50.450 ;
        RECT 85.530 49.700 103.930 50.300 ;
        RECT 85.530 49.550 86.680 49.700 ;
        RECT 82.780 46.800 86.680 49.550 ;
        RECT 82.780 45.050 83.530 46.800 ;
        RECT 85.930 45.050 86.680 46.800 ;
        RECT 86.830 42.150 86.980 49.700 ;
        RECT 87.430 42.150 87.580 49.700 ;
        RECT 88.030 42.150 88.180 49.700 ;
        RECT 88.630 42.150 88.780 49.700 ;
        RECT 89.230 42.150 89.380 49.700 ;
        RECT 89.830 42.150 89.980 49.700 ;
        RECT 94.230 49.200 95.230 49.700 ;
        RECT 90.880 49.050 98.580 49.200 ;
        RECT 94.230 48.600 95.230 49.050 ;
        RECT 90.880 48.450 98.580 48.600 ;
        RECT 94.230 48.000 95.230 48.450 ;
        RECT 90.880 47.850 98.580 48.000 ;
        RECT 94.230 47.400 95.230 47.850 ;
        RECT 90.880 47.250 98.580 47.400 ;
        RECT 94.230 46.800 95.230 47.250 ;
        RECT 90.880 46.650 98.580 46.800 ;
        RECT 94.230 46.200 95.230 46.650 ;
        RECT 90.880 46.050 98.580 46.200 ;
        RECT 94.230 45.600 95.230 46.050 ;
        RECT 90.880 45.450 98.580 45.600 ;
        RECT 94.230 45.000 95.230 45.450 ;
        RECT 90.880 44.850 98.580 45.000 ;
        RECT 94.230 44.400 95.230 44.850 ;
        RECT 90.880 44.250 98.580 44.400 ;
        RECT 94.230 43.800 95.230 44.250 ;
        RECT 90.880 43.650 98.580 43.800 ;
        RECT 94.230 43.200 95.230 43.650 ;
        RECT 90.880 43.050 98.580 43.200 ;
        RECT 94.230 42.600 95.230 43.050 ;
        RECT 90.880 42.450 98.580 42.600 ;
        RECT 94.230 42.000 95.230 42.450 ;
        RECT 99.480 42.150 99.630 49.700 ;
        RECT 100.080 42.150 100.230 49.700 ;
        RECT 100.680 42.150 100.830 49.700 ;
        RECT 101.280 42.150 101.430 49.700 ;
        RECT 101.880 42.150 102.030 49.700 ;
        RECT 102.480 42.150 102.630 49.700 ;
        RECT 102.780 49.550 103.930 49.700 ;
        RECT 104.580 49.550 104.880 50.450 ;
        RECT 105.530 50.300 106.680 50.450 ;
        RECT 106.830 50.300 106.980 57.850 ;
        RECT 107.430 50.300 107.580 57.850 ;
        RECT 108.030 50.300 108.180 57.850 ;
        RECT 108.630 50.300 108.780 57.850 ;
        RECT 109.230 50.300 109.380 57.850 ;
        RECT 109.830 50.300 109.980 57.850 ;
        RECT 114.230 57.550 115.230 58.000 ;
        RECT 110.880 57.400 118.580 57.550 ;
        RECT 114.230 56.950 115.230 57.400 ;
        RECT 110.880 56.800 118.580 56.950 ;
        RECT 114.230 56.350 115.230 56.800 ;
        RECT 110.880 56.200 118.580 56.350 ;
        RECT 114.230 55.750 115.230 56.200 ;
        RECT 110.880 55.600 118.580 55.750 ;
        RECT 114.230 55.150 115.230 55.600 ;
        RECT 110.880 55.000 118.580 55.150 ;
        RECT 114.230 54.550 115.230 55.000 ;
        RECT 110.880 54.400 118.580 54.550 ;
        RECT 114.230 53.950 115.230 54.400 ;
        RECT 110.880 53.800 118.580 53.950 ;
        RECT 114.230 53.350 115.230 53.800 ;
        RECT 110.880 53.200 118.580 53.350 ;
        RECT 114.230 52.750 115.230 53.200 ;
        RECT 110.880 52.600 118.580 52.750 ;
        RECT 114.230 52.150 115.230 52.600 ;
        RECT 110.880 52.000 118.580 52.150 ;
        RECT 114.230 51.550 115.230 52.000 ;
        RECT 110.880 51.400 118.580 51.550 ;
        RECT 114.230 50.950 115.230 51.400 ;
        RECT 110.880 50.800 118.580 50.950 ;
        RECT 114.230 50.300 115.230 50.800 ;
        RECT 119.480 50.300 119.630 57.850 ;
        RECT 120.080 50.300 120.230 57.850 ;
        RECT 120.680 50.300 120.830 57.850 ;
        RECT 121.280 50.300 121.430 57.850 ;
        RECT 121.880 50.300 122.030 57.850 ;
        RECT 122.480 50.300 122.630 57.850 ;
        RECT 122.780 53.200 123.530 55.000 ;
        RECT 122.780 51.405 124.730 53.200 ;
        RECT 122.780 50.450 131.850 51.405 ;
        RECT 122.780 50.300 123.930 50.450 ;
        RECT 105.530 49.700 123.930 50.300 ;
        RECT 105.530 49.550 106.680 49.700 ;
        RECT 102.780 46.800 106.680 49.550 ;
        RECT 102.780 45.050 103.530 46.800 ;
        RECT 105.930 45.050 106.680 46.800 ;
        RECT 106.830 42.150 106.980 49.700 ;
        RECT 107.430 42.150 107.580 49.700 ;
        RECT 108.030 42.150 108.180 49.700 ;
        RECT 108.630 42.150 108.780 49.700 ;
        RECT 109.230 42.150 109.380 49.700 ;
        RECT 109.830 42.150 109.980 49.700 ;
        RECT 114.230 49.200 115.230 49.700 ;
        RECT 110.880 49.050 118.580 49.200 ;
        RECT 114.230 48.600 115.230 49.050 ;
        RECT 110.880 48.450 118.580 48.600 ;
        RECT 114.230 48.000 115.230 48.450 ;
        RECT 110.880 47.850 118.580 48.000 ;
        RECT 114.230 47.400 115.230 47.850 ;
        RECT 110.880 47.250 118.580 47.400 ;
        RECT 114.230 46.800 115.230 47.250 ;
        RECT 110.880 46.650 118.580 46.800 ;
        RECT 114.230 46.200 115.230 46.650 ;
        RECT 110.880 46.050 118.580 46.200 ;
        RECT 114.230 45.600 115.230 46.050 ;
        RECT 110.880 45.450 118.580 45.600 ;
        RECT 114.230 45.000 115.230 45.450 ;
        RECT 110.880 44.850 118.580 45.000 ;
        RECT 114.230 44.400 115.230 44.850 ;
        RECT 110.880 44.250 118.580 44.400 ;
        RECT 114.230 43.800 115.230 44.250 ;
        RECT 110.880 43.650 118.580 43.800 ;
        RECT 114.230 43.200 115.230 43.650 ;
        RECT 110.880 43.050 118.580 43.200 ;
        RECT 114.230 42.600 115.230 43.050 ;
        RECT 110.880 42.450 118.580 42.600 ;
        RECT 114.230 42.000 115.230 42.450 ;
        RECT 119.480 42.150 119.630 49.700 ;
        RECT 120.080 42.150 120.230 49.700 ;
        RECT 120.680 42.150 120.830 49.700 ;
        RECT 121.280 42.150 121.430 49.700 ;
        RECT 121.880 42.150 122.030 49.700 ;
        RECT 122.480 42.150 122.630 49.700 ;
        RECT 122.780 49.550 123.930 49.700 ;
        RECT 124.580 50.130 131.850 50.450 ;
        RECT 124.580 49.550 124.730 50.130 ;
        RECT 122.780 46.800 124.730 49.550 ;
        RECT 122.780 45.050 123.530 46.800 ;
        RECT 10.880 41.850 18.580 42.000 ;
        RECT 30.880 41.850 38.580 42.000 ;
        RECT 50.880 41.850 58.580 42.000 ;
        RECT 70.880 41.850 78.580 42.000 ;
        RECT 90.880 41.850 98.580 42.000 ;
        RECT 110.880 41.850 118.580 42.000 ;
        RECT 14.230 41.200 15.230 41.850 ;
        RECT 34.230 41.200 35.230 41.850 ;
        RECT 54.230 41.200 55.230 41.850 ;
        RECT 74.230 41.200 75.230 41.850 ;
        RECT 94.230 41.200 95.230 41.850 ;
        RECT 114.230 41.200 115.230 41.850 ;
        RECT 11.530 38.800 17.930 41.200 ;
        RECT 31.530 38.800 37.930 41.200 ;
        RECT 51.530 38.800 57.930 41.200 ;
        RECT 71.530 38.800 77.930 41.200 ;
        RECT 91.530 38.800 97.930 41.200 ;
        RECT 111.530 38.800 117.930 41.200 ;
        RECT 14.230 38.150 15.230 38.800 ;
        RECT 34.230 38.150 35.230 38.800 ;
        RECT 54.230 38.150 55.230 38.800 ;
        RECT 74.230 38.150 75.230 38.800 ;
        RECT 94.230 38.150 95.230 38.800 ;
        RECT 114.230 38.150 115.230 38.800 ;
        RECT 10.880 38.000 18.580 38.150 ;
        RECT 30.880 38.000 38.580 38.150 ;
        RECT 50.880 38.000 58.580 38.150 ;
        RECT 70.880 38.000 78.580 38.150 ;
        RECT 90.880 38.000 98.580 38.150 ;
        RECT 110.880 38.000 118.580 38.150 ;
        RECT 5.930 33.200 6.680 35.000 ;
        RECT 4.730 30.450 6.680 33.200 ;
        RECT 4.730 29.550 4.880 30.450 ;
        RECT 5.530 30.300 6.680 30.450 ;
        RECT 6.830 30.300 6.980 37.850 ;
        RECT 7.430 30.300 7.580 37.850 ;
        RECT 8.030 30.300 8.180 37.850 ;
        RECT 8.630 30.300 8.780 37.850 ;
        RECT 9.230 30.300 9.380 37.850 ;
        RECT 9.830 30.300 9.980 37.850 ;
        RECT 14.230 37.550 15.230 38.000 ;
        RECT 10.880 37.400 18.580 37.550 ;
        RECT 14.230 36.950 15.230 37.400 ;
        RECT 10.880 36.800 18.580 36.950 ;
        RECT 14.230 36.350 15.230 36.800 ;
        RECT 10.880 36.200 18.580 36.350 ;
        RECT 14.230 35.750 15.230 36.200 ;
        RECT 10.880 35.600 18.580 35.750 ;
        RECT 14.230 35.150 15.230 35.600 ;
        RECT 10.880 35.000 18.580 35.150 ;
        RECT 14.230 34.550 15.230 35.000 ;
        RECT 10.880 34.400 18.580 34.550 ;
        RECT 14.230 33.950 15.230 34.400 ;
        RECT 10.880 33.800 18.580 33.950 ;
        RECT 14.230 33.350 15.230 33.800 ;
        RECT 10.880 33.200 18.580 33.350 ;
        RECT 14.230 32.750 15.230 33.200 ;
        RECT 10.880 32.600 18.580 32.750 ;
        RECT 14.230 32.150 15.230 32.600 ;
        RECT 10.880 32.000 18.580 32.150 ;
        RECT 14.230 31.550 15.230 32.000 ;
        RECT 10.880 31.400 18.580 31.550 ;
        RECT 14.230 30.950 15.230 31.400 ;
        RECT 10.880 30.800 18.580 30.950 ;
        RECT 14.230 30.300 15.230 30.800 ;
        RECT 19.480 30.300 19.630 37.850 ;
        RECT 20.080 30.300 20.230 37.850 ;
        RECT 20.680 30.300 20.830 37.850 ;
        RECT 21.280 30.300 21.430 37.850 ;
        RECT 21.880 30.300 22.030 37.850 ;
        RECT 22.480 30.300 22.630 37.850 ;
        RECT 22.780 33.200 23.530 35.000 ;
        RECT 25.930 33.200 26.680 35.000 ;
        RECT 22.780 30.450 26.680 33.200 ;
        RECT 22.780 30.300 23.930 30.450 ;
        RECT 5.530 29.700 23.930 30.300 ;
        RECT 5.530 29.550 6.680 29.700 ;
        RECT 4.730 26.800 6.680 29.550 ;
        RECT 5.930 25.050 6.680 26.800 ;
        RECT 6.830 22.150 6.980 29.700 ;
        RECT 7.430 22.150 7.580 29.700 ;
        RECT 8.030 22.150 8.180 29.700 ;
        RECT 8.630 22.150 8.780 29.700 ;
        RECT 9.230 22.150 9.380 29.700 ;
        RECT 9.830 22.150 9.980 29.700 ;
        RECT 14.230 29.200 15.230 29.700 ;
        RECT 10.880 29.050 18.580 29.200 ;
        RECT 14.230 28.600 15.230 29.050 ;
        RECT 10.880 28.450 18.580 28.600 ;
        RECT 14.230 28.000 15.230 28.450 ;
        RECT 10.880 27.850 18.580 28.000 ;
        RECT 14.230 27.400 15.230 27.850 ;
        RECT 10.880 27.250 18.580 27.400 ;
        RECT 14.230 26.800 15.230 27.250 ;
        RECT 10.880 26.650 18.580 26.800 ;
        RECT 14.230 26.200 15.230 26.650 ;
        RECT 10.880 26.050 18.580 26.200 ;
        RECT 14.230 25.600 15.230 26.050 ;
        RECT 10.880 25.450 18.580 25.600 ;
        RECT 14.230 25.000 15.230 25.450 ;
        RECT 10.880 24.850 18.580 25.000 ;
        RECT 14.230 24.400 15.230 24.850 ;
        RECT 10.880 24.250 18.580 24.400 ;
        RECT 14.230 23.800 15.230 24.250 ;
        RECT 10.880 23.650 18.580 23.800 ;
        RECT 14.230 23.200 15.230 23.650 ;
        RECT 10.880 23.050 18.580 23.200 ;
        RECT 14.230 22.600 15.230 23.050 ;
        RECT 10.880 22.450 18.580 22.600 ;
        RECT 14.230 22.000 15.230 22.450 ;
        RECT 19.480 22.150 19.630 29.700 ;
        RECT 20.080 22.150 20.230 29.700 ;
        RECT 20.680 22.150 20.830 29.700 ;
        RECT 21.280 22.150 21.430 29.700 ;
        RECT 21.880 22.150 22.030 29.700 ;
        RECT 22.480 22.150 22.630 29.700 ;
        RECT 22.780 29.550 23.930 29.700 ;
        RECT 24.580 29.550 24.880 30.450 ;
        RECT 25.530 30.300 26.680 30.450 ;
        RECT 26.830 30.300 26.980 37.850 ;
        RECT 27.430 30.300 27.580 37.850 ;
        RECT 28.030 30.300 28.180 37.850 ;
        RECT 28.630 30.300 28.780 37.850 ;
        RECT 29.230 30.300 29.380 37.850 ;
        RECT 29.830 30.300 29.980 37.850 ;
        RECT 34.230 37.550 35.230 38.000 ;
        RECT 30.880 37.400 38.580 37.550 ;
        RECT 34.230 36.950 35.230 37.400 ;
        RECT 30.880 36.800 38.580 36.950 ;
        RECT 34.230 36.350 35.230 36.800 ;
        RECT 30.880 36.200 38.580 36.350 ;
        RECT 34.230 35.750 35.230 36.200 ;
        RECT 30.880 35.600 38.580 35.750 ;
        RECT 34.230 35.150 35.230 35.600 ;
        RECT 30.880 35.000 38.580 35.150 ;
        RECT 34.230 34.550 35.230 35.000 ;
        RECT 30.880 34.400 38.580 34.550 ;
        RECT 34.230 33.950 35.230 34.400 ;
        RECT 30.880 33.800 38.580 33.950 ;
        RECT 34.230 33.350 35.230 33.800 ;
        RECT 30.880 33.200 38.580 33.350 ;
        RECT 34.230 32.750 35.230 33.200 ;
        RECT 30.880 32.600 38.580 32.750 ;
        RECT 34.230 32.150 35.230 32.600 ;
        RECT 30.880 32.000 38.580 32.150 ;
        RECT 34.230 31.550 35.230 32.000 ;
        RECT 30.880 31.400 38.580 31.550 ;
        RECT 34.230 30.950 35.230 31.400 ;
        RECT 30.880 30.800 38.580 30.950 ;
        RECT 34.230 30.300 35.230 30.800 ;
        RECT 39.480 30.300 39.630 37.850 ;
        RECT 40.080 30.300 40.230 37.850 ;
        RECT 40.680 30.300 40.830 37.850 ;
        RECT 41.280 30.300 41.430 37.850 ;
        RECT 41.880 30.300 42.030 37.850 ;
        RECT 42.480 30.300 42.630 37.850 ;
        RECT 42.780 33.200 43.530 35.000 ;
        RECT 45.930 33.200 46.680 35.000 ;
        RECT 42.780 30.450 46.680 33.200 ;
        RECT 42.780 30.300 43.930 30.450 ;
        RECT 25.530 29.700 43.930 30.300 ;
        RECT 25.530 29.550 26.680 29.700 ;
        RECT 22.780 26.800 26.680 29.550 ;
        RECT 22.780 25.050 23.530 26.800 ;
        RECT 25.930 25.050 26.680 26.800 ;
        RECT 26.830 22.150 26.980 29.700 ;
        RECT 27.430 22.150 27.580 29.700 ;
        RECT 28.030 22.150 28.180 29.700 ;
        RECT 28.630 22.150 28.780 29.700 ;
        RECT 29.230 22.150 29.380 29.700 ;
        RECT 29.830 22.150 29.980 29.700 ;
        RECT 34.230 29.200 35.230 29.700 ;
        RECT 30.880 29.050 38.580 29.200 ;
        RECT 34.230 28.600 35.230 29.050 ;
        RECT 30.880 28.450 38.580 28.600 ;
        RECT 34.230 28.000 35.230 28.450 ;
        RECT 30.880 27.850 38.580 28.000 ;
        RECT 34.230 27.400 35.230 27.850 ;
        RECT 30.880 27.250 38.580 27.400 ;
        RECT 34.230 26.800 35.230 27.250 ;
        RECT 30.880 26.650 38.580 26.800 ;
        RECT 34.230 26.200 35.230 26.650 ;
        RECT 30.880 26.050 38.580 26.200 ;
        RECT 34.230 25.600 35.230 26.050 ;
        RECT 30.880 25.450 38.580 25.600 ;
        RECT 34.230 25.000 35.230 25.450 ;
        RECT 30.880 24.850 38.580 25.000 ;
        RECT 34.230 24.400 35.230 24.850 ;
        RECT 30.880 24.250 38.580 24.400 ;
        RECT 34.230 23.800 35.230 24.250 ;
        RECT 30.880 23.650 38.580 23.800 ;
        RECT 34.230 23.200 35.230 23.650 ;
        RECT 30.880 23.050 38.580 23.200 ;
        RECT 34.230 22.600 35.230 23.050 ;
        RECT 30.880 22.450 38.580 22.600 ;
        RECT 34.230 22.000 35.230 22.450 ;
        RECT 39.480 22.150 39.630 29.700 ;
        RECT 40.080 22.150 40.230 29.700 ;
        RECT 40.680 22.150 40.830 29.700 ;
        RECT 41.280 22.150 41.430 29.700 ;
        RECT 41.880 22.150 42.030 29.700 ;
        RECT 42.480 22.150 42.630 29.700 ;
        RECT 42.780 29.550 43.930 29.700 ;
        RECT 44.580 29.550 44.880 30.450 ;
        RECT 45.530 30.300 46.680 30.450 ;
        RECT 46.830 30.300 46.980 37.850 ;
        RECT 47.430 30.300 47.580 37.850 ;
        RECT 48.030 30.300 48.180 37.850 ;
        RECT 48.630 30.300 48.780 37.850 ;
        RECT 49.230 30.300 49.380 37.850 ;
        RECT 49.830 30.300 49.980 37.850 ;
        RECT 54.230 37.550 55.230 38.000 ;
        RECT 50.880 37.400 58.580 37.550 ;
        RECT 54.230 36.950 55.230 37.400 ;
        RECT 50.880 36.800 58.580 36.950 ;
        RECT 54.230 36.350 55.230 36.800 ;
        RECT 50.880 36.200 58.580 36.350 ;
        RECT 54.230 35.750 55.230 36.200 ;
        RECT 50.880 35.600 58.580 35.750 ;
        RECT 54.230 35.150 55.230 35.600 ;
        RECT 50.880 35.000 58.580 35.150 ;
        RECT 54.230 34.550 55.230 35.000 ;
        RECT 50.880 34.400 58.580 34.550 ;
        RECT 54.230 33.950 55.230 34.400 ;
        RECT 50.880 33.800 58.580 33.950 ;
        RECT 54.230 33.350 55.230 33.800 ;
        RECT 50.880 33.200 58.580 33.350 ;
        RECT 54.230 32.750 55.230 33.200 ;
        RECT 50.880 32.600 58.580 32.750 ;
        RECT 54.230 32.150 55.230 32.600 ;
        RECT 50.880 32.000 58.580 32.150 ;
        RECT 54.230 31.550 55.230 32.000 ;
        RECT 50.880 31.400 58.580 31.550 ;
        RECT 54.230 30.950 55.230 31.400 ;
        RECT 50.880 30.800 58.580 30.950 ;
        RECT 54.230 30.300 55.230 30.800 ;
        RECT 59.480 30.300 59.630 37.850 ;
        RECT 60.080 30.300 60.230 37.850 ;
        RECT 60.680 30.300 60.830 37.850 ;
        RECT 61.280 30.300 61.430 37.850 ;
        RECT 61.880 30.300 62.030 37.850 ;
        RECT 62.480 30.300 62.630 37.850 ;
        RECT 62.780 33.200 63.530 35.000 ;
        RECT 65.930 33.200 66.680 35.000 ;
        RECT 62.780 30.450 66.680 33.200 ;
        RECT 62.780 30.300 63.930 30.450 ;
        RECT 45.530 29.700 63.930 30.300 ;
        RECT 45.530 29.550 46.680 29.700 ;
        RECT 42.780 26.800 46.680 29.550 ;
        RECT 42.780 25.050 43.530 26.800 ;
        RECT 45.930 25.050 46.680 26.800 ;
        RECT 46.830 22.150 46.980 29.700 ;
        RECT 47.430 22.150 47.580 29.700 ;
        RECT 48.030 22.150 48.180 29.700 ;
        RECT 48.630 22.150 48.780 29.700 ;
        RECT 49.230 22.150 49.380 29.700 ;
        RECT 49.830 22.150 49.980 29.700 ;
        RECT 54.230 29.200 55.230 29.700 ;
        RECT 50.880 29.050 58.580 29.200 ;
        RECT 54.230 28.600 55.230 29.050 ;
        RECT 50.880 28.450 58.580 28.600 ;
        RECT 54.230 28.000 55.230 28.450 ;
        RECT 50.880 27.850 58.580 28.000 ;
        RECT 54.230 27.400 55.230 27.850 ;
        RECT 50.880 27.250 58.580 27.400 ;
        RECT 54.230 26.800 55.230 27.250 ;
        RECT 50.880 26.650 58.580 26.800 ;
        RECT 54.230 26.200 55.230 26.650 ;
        RECT 50.880 26.050 58.580 26.200 ;
        RECT 54.230 25.600 55.230 26.050 ;
        RECT 50.880 25.450 58.580 25.600 ;
        RECT 54.230 25.000 55.230 25.450 ;
        RECT 50.880 24.850 58.580 25.000 ;
        RECT 54.230 24.400 55.230 24.850 ;
        RECT 50.880 24.250 58.580 24.400 ;
        RECT 54.230 23.800 55.230 24.250 ;
        RECT 50.880 23.650 58.580 23.800 ;
        RECT 54.230 23.200 55.230 23.650 ;
        RECT 50.880 23.050 58.580 23.200 ;
        RECT 54.230 22.600 55.230 23.050 ;
        RECT 50.880 22.450 58.580 22.600 ;
        RECT 54.230 22.000 55.230 22.450 ;
        RECT 59.480 22.150 59.630 29.700 ;
        RECT 60.080 22.150 60.230 29.700 ;
        RECT 60.680 22.150 60.830 29.700 ;
        RECT 61.280 22.150 61.430 29.700 ;
        RECT 61.880 22.150 62.030 29.700 ;
        RECT 62.480 22.150 62.630 29.700 ;
        RECT 62.780 29.550 63.930 29.700 ;
        RECT 64.580 29.550 64.880 30.450 ;
        RECT 65.530 30.300 66.680 30.450 ;
        RECT 66.830 30.300 66.980 37.850 ;
        RECT 67.430 30.300 67.580 37.850 ;
        RECT 68.030 30.300 68.180 37.850 ;
        RECT 68.630 30.300 68.780 37.850 ;
        RECT 69.230 30.300 69.380 37.850 ;
        RECT 69.830 30.300 69.980 37.850 ;
        RECT 74.230 37.550 75.230 38.000 ;
        RECT 70.880 37.400 78.580 37.550 ;
        RECT 74.230 36.950 75.230 37.400 ;
        RECT 70.880 36.800 78.580 36.950 ;
        RECT 74.230 36.350 75.230 36.800 ;
        RECT 70.880 36.200 78.580 36.350 ;
        RECT 74.230 35.750 75.230 36.200 ;
        RECT 70.880 35.600 78.580 35.750 ;
        RECT 74.230 35.150 75.230 35.600 ;
        RECT 70.880 35.000 78.580 35.150 ;
        RECT 74.230 34.550 75.230 35.000 ;
        RECT 70.880 34.400 78.580 34.550 ;
        RECT 74.230 33.950 75.230 34.400 ;
        RECT 70.880 33.800 78.580 33.950 ;
        RECT 74.230 33.350 75.230 33.800 ;
        RECT 70.880 33.200 78.580 33.350 ;
        RECT 74.230 32.750 75.230 33.200 ;
        RECT 70.880 32.600 78.580 32.750 ;
        RECT 74.230 32.150 75.230 32.600 ;
        RECT 70.880 32.000 78.580 32.150 ;
        RECT 74.230 31.550 75.230 32.000 ;
        RECT 70.880 31.400 78.580 31.550 ;
        RECT 74.230 30.950 75.230 31.400 ;
        RECT 70.880 30.800 78.580 30.950 ;
        RECT 74.230 30.300 75.230 30.800 ;
        RECT 79.480 30.300 79.630 37.850 ;
        RECT 80.080 30.300 80.230 37.850 ;
        RECT 80.680 30.300 80.830 37.850 ;
        RECT 81.280 30.300 81.430 37.850 ;
        RECT 81.880 30.300 82.030 37.850 ;
        RECT 82.480 30.300 82.630 37.850 ;
        RECT 82.780 33.200 83.530 35.000 ;
        RECT 85.930 33.200 86.680 35.000 ;
        RECT 82.780 30.450 86.680 33.200 ;
        RECT 82.780 30.300 83.930 30.450 ;
        RECT 65.530 29.700 83.930 30.300 ;
        RECT 65.530 29.550 66.680 29.700 ;
        RECT 62.780 26.800 66.680 29.550 ;
        RECT 62.780 25.050 63.530 26.800 ;
        RECT 65.930 25.050 66.680 26.800 ;
        RECT 66.830 22.150 66.980 29.700 ;
        RECT 67.430 22.150 67.580 29.700 ;
        RECT 68.030 22.150 68.180 29.700 ;
        RECT 68.630 22.150 68.780 29.700 ;
        RECT 69.230 22.150 69.380 29.700 ;
        RECT 69.830 22.150 69.980 29.700 ;
        RECT 74.230 29.200 75.230 29.700 ;
        RECT 70.880 29.050 78.580 29.200 ;
        RECT 74.230 28.600 75.230 29.050 ;
        RECT 70.880 28.450 78.580 28.600 ;
        RECT 74.230 28.000 75.230 28.450 ;
        RECT 70.880 27.850 78.580 28.000 ;
        RECT 74.230 27.400 75.230 27.850 ;
        RECT 70.880 27.250 78.580 27.400 ;
        RECT 74.230 26.800 75.230 27.250 ;
        RECT 70.880 26.650 78.580 26.800 ;
        RECT 74.230 26.200 75.230 26.650 ;
        RECT 70.880 26.050 78.580 26.200 ;
        RECT 74.230 25.600 75.230 26.050 ;
        RECT 70.880 25.450 78.580 25.600 ;
        RECT 74.230 25.000 75.230 25.450 ;
        RECT 70.880 24.850 78.580 25.000 ;
        RECT 74.230 24.400 75.230 24.850 ;
        RECT 70.880 24.250 78.580 24.400 ;
        RECT 74.230 23.800 75.230 24.250 ;
        RECT 70.880 23.650 78.580 23.800 ;
        RECT 74.230 23.200 75.230 23.650 ;
        RECT 70.880 23.050 78.580 23.200 ;
        RECT 74.230 22.600 75.230 23.050 ;
        RECT 70.880 22.450 78.580 22.600 ;
        RECT 74.230 22.000 75.230 22.450 ;
        RECT 79.480 22.150 79.630 29.700 ;
        RECT 80.080 22.150 80.230 29.700 ;
        RECT 80.680 22.150 80.830 29.700 ;
        RECT 81.280 22.150 81.430 29.700 ;
        RECT 81.880 22.150 82.030 29.700 ;
        RECT 82.480 22.150 82.630 29.700 ;
        RECT 82.780 29.550 83.930 29.700 ;
        RECT 84.580 29.550 84.880 30.450 ;
        RECT 85.530 30.300 86.680 30.450 ;
        RECT 86.830 30.300 86.980 37.850 ;
        RECT 87.430 30.300 87.580 37.850 ;
        RECT 88.030 30.300 88.180 37.850 ;
        RECT 88.630 30.300 88.780 37.850 ;
        RECT 89.230 30.300 89.380 37.850 ;
        RECT 89.830 30.300 89.980 37.850 ;
        RECT 94.230 37.550 95.230 38.000 ;
        RECT 90.880 37.400 98.580 37.550 ;
        RECT 94.230 36.950 95.230 37.400 ;
        RECT 90.880 36.800 98.580 36.950 ;
        RECT 94.230 36.350 95.230 36.800 ;
        RECT 90.880 36.200 98.580 36.350 ;
        RECT 94.230 35.750 95.230 36.200 ;
        RECT 90.880 35.600 98.580 35.750 ;
        RECT 94.230 35.150 95.230 35.600 ;
        RECT 90.880 35.000 98.580 35.150 ;
        RECT 94.230 34.550 95.230 35.000 ;
        RECT 90.880 34.400 98.580 34.550 ;
        RECT 94.230 33.950 95.230 34.400 ;
        RECT 90.880 33.800 98.580 33.950 ;
        RECT 94.230 33.350 95.230 33.800 ;
        RECT 90.880 33.200 98.580 33.350 ;
        RECT 94.230 32.750 95.230 33.200 ;
        RECT 90.880 32.600 98.580 32.750 ;
        RECT 94.230 32.150 95.230 32.600 ;
        RECT 90.880 32.000 98.580 32.150 ;
        RECT 94.230 31.550 95.230 32.000 ;
        RECT 90.880 31.400 98.580 31.550 ;
        RECT 94.230 30.950 95.230 31.400 ;
        RECT 90.880 30.800 98.580 30.950 ;
        RECT 94.230 30.300 95.230 30.800 ;
        RECT 99.480 30.300 99.630 37.850 ;
        RECT 100.080 30.300 100.230 37.850 ;
        RECT 100.680 30.300 100.830 37.850 ;
        RECT 101.280 30.300 101.430 37.850 ;
        RECT 101.880 30.300 102.030 37.850 ;
        RECT 102.480 30.300 102.630 37.850 ;
        RECT 102.780 33.200 103.530 35.000 ;
        RECT 105.930 33.200 106.680 35.000 ;
        RECT 102.780 30.450 106.680 33.200 ;
        RECT 102.780 30.300 103.930 30.450 ;
        RECT 85.530 29.700 103.930 30.300 ;
        RECT 85.530 29.550 86.680 29.700 ;
        RECT 82.780 26.800 86.680 29.550 ;
        RECT 82.780 25.050 83.530 26.800 ;
        RECT 85.930 25.050 86.680 26.800 ;
        RECT 86.830 22.150 86.980 29.700 ;
        RECT 87.430 22.150 87.580 29.700 ;
        RECT 88.030 22.150 88.180 29.700 ;
        RECT 88.630 22.150 88.780 29.700 ;
        RECT 89.230 22.150 89.380 29.700 ;
        RECT 89.830 22.150 89.980 29.700 ;
        RECT 94.230 29.200 95.230 29.700 ;
        RECT 90.880 29.050 98.580 29.200 ;
        RECT 94.230 28.600 95.230 29.050 ;
        RECT 90.880 28.450 98.580 28.600 ;
        RECT 94.230 28.000 95.230 28.450 ;
        RECT 90.880 27.850 98.580 28.000 ;
        RECT 94.230 27.400 95.230 27.850 ;
        RECT 90.880 27.250 98.580 27.400 ;
        RECT 94.230 26.800 95.230 27.250 ;
        RECT 90.880 26.650 98.580 26.800 ;
        RECT 94.230 26.200 95.230 26.650 ;
        RECT 90.880 26.050 98.580 26.200 ;
        RECT 94.230 25.600 95.230 26.050 ;
        RECT 90.880 25.450 98.580 25.600 ;
        RECT 94.230 25.000 95.230 25.450 ;
        RECT 90.880 24.850 98.580 25.000 ;
        RECT 94.230 24.400 95.230 24.850 ;
        RECT 90.880 24.250 98.580 24.400 ;
        RECT 94.230 23.800 95.230 24.250 ;
        RECT 90.880 23.650 98.580 23.800 ;
        RECT 94.230 23.200 95.230 23.650 ;
        RECT 90.880 23.050 98.580 23.200 ;
        RECT 94.230 22.600 95.230 23.050 ;
        RECT 90.880 22.450 98.580 22.600 ;
        RECT 94.230 22.000 95.230 22.450 ;
        RECT 99.480 22.150 99.630 29.700 ;
        RECT 100.080 22.150 100.230 29.700 ;
        RECT 100.680 22.150 100.830 29.700 ;
        RECT 101.280 22.150 101.430 29.700 ;
        RECT 101.880 22.150 102.030 29.700 ;
        RECT 102.480 22.150 102.630 29.700 ;
        RECT 102.780 29.550 103.930 29.700 ;
        RECT 104.580 29.550 104.880 30.450 ;
        RECT 105.530 30.300 106.680 30.450 ;
        RECT 106.830 30.300 106.980 37.850 ;
        RECT 107.430 30.300 107.580 37.850 ;
        RECT 108.030 30.300 108.180 37.850 ;
        RECT 108.630 30.300 108.780 37.850 ;
        RECT 109.230 30.300 109.380 37.850 ;
        RECT 109.830 30.300 109.980 37.850 ;
        RECT 114.230 37.550 115.230 38.000 ;
        RECT 110.880 37.400 118.580 37.550 ;
        RECT 114.230 36.950 115.230 37.400 ;
        RECT 110.880 36.800 118.580 36.950 ;
        RECT 114.230 36.350 115.230 36.800 ;
        RECT 110.880 36.200 118.580 36.350 ;
        RECT 114.230 35.750 115.230 36.200 ;
        RECT 110.880 35.600 118.580 35.750 ;
        RECT 114.230 35.150 115.230 35.600 ;
        RECT 110.880 35.000 118.580 35.150 ;
        RECT 114.230 34.550 115.230 35.000 ;
        RECT 110.880 34.400 118.580 34.550 ;
        RECT 114.230 33.950 115.230 34.400 ;
        RECT 110.880 33.800 118.580 33.950 ;
        RECT 114.230 33.350 115.230 33.800 ;
        RECT 110.880 33.200 118.580 33.350 ;
        RECT 114.230 32.750 115.230 33.200 ;
        RECT 110.880 32.600 118.580 32.750 ;
        RECT 114.230 32.150 115.230 32.600 ;
        RECT 110.880 32.000 118.580 32.150 ;
        RECT 114.230 31.550 115.230 32.000 ;
        RECT 110.880 31.400 118.580 31.550 ;
        RECT 114.230 30.950 115.230 31.400 ;
        RECT 110.880 30.800 118.580 30.950 ;
        RECT 114.230 30.300 115.230 30.800 ;
        RECT 119.480 30.300 119.630 37.850 ;
        RECT 120.080 30.300 120.230 37.850 ;
        RECT 120.680 30.300 120.830 37.850 ;
        RECT 121.280 30.300 121.430 37.850 ;
        RECT 121.880 30.300 122.030 37.850 ;
        RECT 122.480 30.300 122.630 37.850 ;
        RECT 122.780 33.200 123.530 35.000 ;
        RECT 122.780 31.585 124.730 33.200 ;
        RECT 122.780 30.450 131.850 31.585 ;
        RECT 122.780 30.300 123.930 30.450 ;
        RECT 105.530 29.700 123.930 30.300 ;
        RECT 105.530 29.550 106.680 29.700 ;
        RECT 102.780 26.800 106.680 29.550 ;
        RECT 102.780 25.050 103.530 26.800 ;
        RECT 105.930 25.050 106.680 26.800 ;
        RECT 106.830 22.150 106.980 29.700 ;
        RECT 107.430 22.150 107.580 29.700 ;
        RECT 108.030 22.150 108.180 29.700 ;
        RECT 108.630 22.150 108.780 29.700 ;
        RECT 109.230 22.150 109.380 29.700 ;
        RECT 109.830 22.150 109.980 29.700 ;
        RECT 114.230 29.200 115.230 29.700 ;
        RECT 110.880 29.050 118.580 29.200 ;
        RECT 114.230 28.600 115.230 29.050 ;
        RECT 110.880 28.450 118.580 28.600 ;
        RECT 114.230 28.000 115.230 28.450 ;
        RECT 110.880 27.850 118.580 28.000 ;
        RECT 114.230 27.400 115.230 27.850 ;
        RECT 110.880 27.250 118.580 27.400 ;
        RECT 114.230 26.800 115.230 27.250 ;
        RECT 110.880 26.650 118.580 26.800 ;
        RECT 114.230 26.200 115.230 26.650 ;
        RECT 110.880 26.050 118.580 26.200 ;
        RECT 114.230 25.600 115.230 26.050 ;
        RECT 110.880 25.450 118.580 25.600 ;
        RECT 114.230 25.000 115.230 25.450 ;
        RECT 110.880 24.850 118.580 25.000 ;
        RECT 114.230 24.400 115.230 24.850 ;
        RECT 110.880 24.250 118.580 24.400 ;
        RECT 114.230 23.800 115.230 24.250 ;
        RECT 110.880 23.650 118.580 23.800 ;
        RECT 114.230 23.200 115.230 23.650 ;
        RECT 110.880 23.050 118.580 23.200 ;
        RECT 114.230 22.600 115.230 23.050 ;
        RECT 110.880 22.450 118.580 22.600 ;
        RECT 114.230 22.000 115.230 22.450 ;
        RECT 119.480 22.150 119.630 29.700 ;
        RECT 120.080 22.150 120.230 29.700 ;
        RECT 120.680 22.150 120.830 29.700 ;
        RECT 121.280 22.150 121.430 29.700 ;
        RECT 121.880 22.150 122.030 29.700 ;
        RECT 122.480 22.150 122.630 29.700 ;
        RECT 122.780 29.550 123.930 29.700 ;
        RECT 124.580 30.310 131.850 30.450 ;
        RECT 124.580 29.550 124.730 30.310 ;
        RECT 122.780 26.800 124.730 29.550 ;
        RECT 122.780 25.050 123.530 26.800 ;
        RECT 10.880 21.850 18.580 22.000 ;
        RECT 30.880 21.850 38.580 22.000 ;
        RECT 50.880 21.850 58.580 22.000 ;
        RECT 70.880 21.850 78.580 22.000 ;
        RECT 90.880 21.850 98.580 22.000 ;
        RECT 110.880 21.850 118.580 22.000 ;
        RECT 14.230 21.200 15.230 21.850 ;
        RECT 34.230 21.200 35.230 21.850 ;
        RECT 54.230 21.200 55.230 21.850 ;
        RECT 74.230 21.200 75.230 21.850 ;
        RECT 94.230 21.200 95.230 21.850 ;
        RECT 114.230 21.200 115.230 21.850 ;
        RECT 11.530 18.800 17.930 21.200 ;
        RECT 31.530 18.800 37.930 21.200 ;
        RECT 51.530 18.800 57.930 21.200 ;
        RECT 71.530 18.800 77.930 21.200 ;
        RECT 91.530 18.800 97.930 21.200 ;
        RECT 111.530 18.800 117.930 21.200 ;
        RECT 14.230 18.150 15.230 18.800 ;
        RECT 34.230 18.150 35.230 18.800 ;
        RECT 54.230 18.150 55.230 18.800 ;
        RECT 74.230 18.150 75.230 18.800 ;
        RECT 94.230 18.150 95.230 18.800 ;
        RECT 114.230 18.150 115.230 18.800 ;
        RECT 10.880 18.000 18.580 18.150 ;
        RECT 30.880 18.000 38.580 18.150 ;
        RECT 50.880 18.000 58.580 18.150 ;
        RECT 70.880 18.000 78.580 18.150 ;
        RECT 90.880 18.000 98.580 18.150 ;
        RECT 110.880 18.000 118.580 18.150 ;
        RECT 5.930 13.200 6.680 15.000 ;
        RECT 4.730 10.450 6.680 13.200 ;
        RECT 4.730 9.550 4.880 10.450 ;
        RECT 5.530 10.300 6.680 10.450 ;
        RECT 6.830 10.300 6.980 17.850 ;
        RECT 7.430 10.300 7.580 17.850 ;
        RECT 8.030 10.300 8.180 17.850 ;
        RECT 8.630 10.300 8.780 17.850 ;
        RECT 9.230 10.300 9.380 17.850 ;
        RECT 9.830 10.300 9.980 17.850 ;
        RECT 14.230 17.550 15.230 18.000 ;
        RECT 10.880 17.400 18.580 17.550 ;
        RECT 14.230 16.950 15.230 17.400 ;
        RECT 10.880 16.800 18.580 16.950 ;
        RECT 14.230 16.350 15.230 16.800 ;
        RECT 10.880 16.200 18.580 16.350 ;
        RECT 14.230 15.750 15.230 16.200 ;
        RECT 10.880 15.600 18.580 15.750 ;
        RECT 14.230 15.150 15.230 15.600 ;
        RECT 10.880 15.000 18.580 15.150 ;
        RECT 14.230 14.550 15.230 15.000 ;
        RECT 10.880 14.400 18.580 14.550 ;
        RECT 14.230 13.950 15.230 14.400 ;
        RECT 10.880 13.800 18.580 13.950 ;
        RECT 14.230 13.350 15.230 13.800 ;
        RECT 10.880 13.200 18.580 13.350 ;
        RECT 14.230 12.750 15.230 13.200 ;
        RECT 10.880 12.600 18.580 12.750 ;
        RECT 14.230 12.150 15.230 12.600 ;
        RECT 10.880 12.000 18.580 12.150 ;
        RECT 14.230 11.550 15.230 12.000 ;
        RECT 10.880 11.400 18.580 11.550 ;
        RECT 14.230 10.950 15.230 11.400 ;
        RECT 10.880 10.800 18.580 10.950 ;
        RECT 14.230 10.300 15.230 10.800 ;
        RECT 19.480 10.300 19.630 17.850 ;
        RECT 20.080 10.300 20.230 17.850 ;
        RECT 20.680 10.300 20.830 17.850 ;
        RECT 21.280 10.300 21.430 17.850 ;
        RECT 21.880 10.300 22.030 17.850 ;
        RECT 22.480 10.300 22.630 17.850 ;
        RECT 22.780 13.200 23.530 15.000 ;
        RECT 25.930 13.200 26.680 15.000 ;
        RECT 22.780 10.450 26.680 13.200 ;
        RECT 22.780 10.300 23.930 10.450 ;
        RECT 5.530 9.700 23.930 10.300 ;
        RECT 5.530 9.550 6.680 9.700 ;
        RECT 4.730 6.800 6.680 9.550 ;
        RECT 5.930 5.050 6.680 6.800 ;
        RECT 6.830 2.150 6.980 9.700 ;
        RECT 7.430 2.150 7.580 9.700 ;
        RECT 8.030 2.150 8.180 9.700 ;
        RECT 8.630 2.150 8.780 9.700 ;
        RECT 9.230 2.150 9.380 9.700 ;
        RECT 9.830 2.150 9.980 9.700 ;
        RECT 14.230 9.200 15.230 9.700 ;
        RECT 10.880 9.050 18.580 9.200 ;
        RECT 14.230 8.600 15.230 9.050 ;
        RECT 10.880 8.450 18.580 8.600 ;
        RECT 14.230 8.000 15.230 8.450 ;
        RECT 10.880 7.850 18.580 8.000 ;
        RECT 14.230 7.400 15.230 7.850 ;
        RECT 10.880 7.250 18.580 7.400 ;
        RECT 14.230 6.800 15.230 7.250 ;
        RECT 10.880 6.650 18.580 6.800 ;
        RECT 14.230 6.200 15.230 6.650 ;
        RECT 10.880 6.050 18.580 6.200 ;
        RECT 14.230 5.600 15.230 6.050 ;
        RECT 10.880 5.450 18.580 5.600 ;
        RECT 14.230 5.000 15.230 5.450 ;
        RECT 10.880 4.850 18.580 5.000 ;
        RECT 14.230 4.400 15.230 4.850 ;
        RECT 10.880 4.250 18.580 4.400 ;
        RECT 14.230 3.800 15.230 4.250 ;
        RECT 10.880 3.650 18.580 3.800 ;
        RECT 14.230 3.200 15.230 3.650 ;
        RECT 10.880 3.050 18.580 3.200 ;
        RECT 14.230 2.600 15.230 3.050 ;
        RECT 10.880 2.450 18.580 2.600 ;
        RECT 14.230 2.000 15.230 2.450 ;
        RECT 19.480 2.150 19.630 9.700 ;
        RECT 20.080 2.150 20.230 9.700 ;
        RECT 20.680 2.150 20.830 9.700 ;
        RECT 21.280 2.150 21.430 9.700 ;
        RECT 21.880 2.150 22.030 9.700 ;
        RECT 22.480 2.150 22.630 9.700 ;
        RECT 22.780 9.550 23.930 9.700 ;
        RECT 24.580 9.550 24.880 10.450 ;
        RECT 25.530 10.300 26.680 10.450 ;
        RECT 26.830 10.300 26.980 17.850 ;
        RECT 27.430 10.300 27.580 17.850 ;
        RECT 28.030 10.300 28.180 17.850 ;
        RECT 28.630 10.300 28.780 17.850 ;
        RECT 29.230 10.300 29.380 17.850 ;
        RECT 29.830 10.300 29.980 17.850 ;
        RECT 34.230 17.550 35.230 18.000 ;
        RECT 30.880 17.400 38.580 17.550 ;
        RECT 34.230 16.950 35.230 17.400 ;
        RECT 30.880 16.800 38.580 16.950 ;
        RECT 34.230 16.350 35.230 16.800 ;
        RECT 30.880 16.200 38.580 16.350 ;
        RECT 34.230 15.750 35.230 16.200 ;
        RECT 30.880 15.600 38.580 15.750 ;
        RECT 34.230 15.150 35.230 15.600 ;
        RECT 30.880 15.000 38.580 15.150 ;
        RECT 34.230 14.550 35.230 15.000 ;
        RECT 30.880 14.400 38.580 14.550 ;
        RECT 34.230 13.950 35.230 14.400 ;
        RECT 30.880 13.800 38.580 13.950 ;
        RECT 34.230 13.350 35.230 13.800 ;
        RECT 30.880 13.200 38.580 13.350 ;
        RECT 34.230 12.750 35.230 13.200 ;
        RECT 30.880 12.600 38.580 12.750 ;
        RECT 34.230 12.150 35.230 12.600 ;
        RECT 30.880 12.000 38.580 12.150 ;
        RECT 34.230 11.550 35.230 12.000 ;
        RECT 30.880 11.400 38.580 11.550 ;
        RECT 34.230 10.950 35.230 11.400 ;
        RECT 30.880 10.800 38.580 10.950 ;
        RECT 34.230 10.300 35.230 10.800 ;
        RECT 39.480 10.300 39.630 17.850 ;
        RECT 40.080 10.300 40.230 17.850 ;
        RECT 40.680 10.300 40.830 17.850 ;
        RECT 41.280 10.300 41.430 17.850 ;
        RECT 41.880 10.300 42.030 17.850 ;
        RECT 42.480 10.300 42.630 17.850 ;
        RECT 42.780 13.200 43.530 15.000 ;
        RECT 45.930 13.200 46.680 15.000 ;
        RECT 42.780 10.450 46.680 13.200 ;
        RECT 42.780 10.300 43.930 10.450 ;
        RECT 25.530 9.700 43.930 10.300 ;
        RECT 25.530 9.550 26.680 9.700 ;
        RECT 22.780 6.800 26.680 9.550 ;
        RECT 22.780 5.050 23.530 6.800 ;
        RECT 25.930 5.050 26.680 6.800 ;
        RECT 26.830 2.150 26.980 9.700 ;
        RECT 27.430 2.150 27.580 9.700 ;
        RECT 28.030 2.150 28.180 9.700 ;
        RECT 28.630 2.150 28.780 9.700 ;
        RECT 29.230 2.150 29.380 9.700 ;
        RECT 29.830 2.150 29.980 9.700 ;
        RECT 34.230 9.200 35.230 9.700 ;
        RECT 30.880 9.050 38.580 9.200 ;
        RECT 34.230 8.600 35.230 9.050 ;
        RECT 30.880 8.450 38.580 8.600 ;
        RECT 34.230 8.000 35.230 8.450 ;
        RECT 30.880 7.850 38.580 8.000 ;
        RECT 34.230 7.400 35.230 7.850 ;
        RECT 30.880 7.250 38.580 7.400 ;
        RECT 34.230 6.800 35.230 7.250 ;
        RECT 30.880 6.650 38.580 6.800 ;
        RECT 34.230 6.200 35.230 6.650 ;
        RECT 30.880 6.050 38.580 6.200 ;
        RECT 34.230 5.600 35.230 6.050 ;
        RECT 30.880 5.450 38.580 5.600 ;
        RECT 34.230 5.000 35.230 5.450 ;
        RECT 30.880 4.850 38.580 5.000 ;
        RECT 34.230 4.400 35.230 4.850 ;
        RECT 30.880 4.250 38.580 4.400 ;
        RECT 34.230 3.800 35.230 4.250 ;
        RECT 30.880 3.650 38.580 3.800 ;
        RECT 34.230 3.200 35.230 3.650 ;
        RECT 30.880 3.050 38.580 3.200 ;
        RECT 34.230 2.600 35.230 3.050 ;
        RECT 30.880 2.450 38.580 2.600 ;
        RECT 34.230 2.000 35.230 2.450 ;
        RECT 39.480 2.150 39.630 9.700 ;
        RECT 40.080 2.150 40.230 9.700 ;
        RECT 40.680 2.150 40.830 9.700 ;
        RECT 41.280 2.150 41.430 9.700 ;
        RECT 41.880 2.150 42.030 9.700 ;
        RECT 42.480 2.150 42.630 9.700 ;
        RECT 42.780 9.550 43.930 9.700 ;
        RECT 44.580 9.550 44.880 10.450 ;
        RECT 45.530 10.300 46.680 10.450 ;
        RECT 46.830 10.300 46.980 17.850 ;
        RECT 47.430 10.300 47.580 17.850 ;
        RECT 48.030 10.300 48.180 17.850 ;
        RECT 48.630 10.300 48.780 17.850 ;
        RECT 49.230 10.300 49.380 17.850 ;
        RECT 49.830 10.300 49.980 17.850 ;
        RECT 54.230 17.550 55.230 18.000 ;
        RECT 50.880 17.400 58.580 17.550 ;
        RECT 54.230 16.950 55.230 17.400 ;
        RECT 50.880 16.800 58.580 16.950 ;
        RECT 54.230 16.350 55.230 16.800 ;
        RECT 50.880 16.200 58.580 16.350 ;
        RECT 54.230 15.750 55.230 16.200 ;
        RECT 50.880 15.600 58.580 15.750 ;
        RECT 54.230 15.150 55.230 15.600 ;
        RECT 50.880 15.000 58.580 15.150 ;
        RECT 54.230 14.550 55.230 15.000 ;
        RECT 50.880 14.400 58.580 14.550 ;
        RECT 54.230 13.950 55.230 14.400 ;
        RECT 50.880 13.800 58.580 13.950 ;
        RECT 54.230 13.350 55.230 13.800 ;
        RECT 50.880 13.200 58.580 13.350 ;
        RECT 54.230 12.750 55.230 13.200 ;
        RECT 50.880 12.600 58.580 12.750 ;
        RECT 54.230 12.150 55.230 12.600 ;
        RECT 50.880 12.000 58.580 12.150 ;
        RECT 54.230 11.550 55.230 12.000 ;
        RECT 50.880 11.400 58.580 11.550 ;
        RECT 54.230 10.950 55.230 11.400 ;
        RECT 50.880 10.800 58.580 10.950 ;
        RECT 54.230 10.300 55.230 10.800 ;
        RECT 59.480 10.300 59.630 17.850 ;
        RECT 60.080 10.300 60.230 17.850 ;
        RECT 60.680 10.300 60.830 17.850 ;
        RECT 61.280 10.300 61.430 17.850 ;
        RECT 61.880 10.300 62.030 17.850 ;
        RECT 62.480 10.300 62.630 17.850 ;
        RECT 62.780 13.200 63.530 15.000 ;
        RECT 65.930 13.200 66.680 15.000 ;
        RECT 62.780 10.450 66.680 13.200 ;
        RECT 62.780 10.300 63.930 10.450 ;
        RECT 45.530 9.700 63.930 10.300 ;
        RECT 45.530 9.550 46.680 9.700 ;
        RECT 42.780 6.800 46.680 9.550 ;
        RECT 42.780 5.050 43.530 6.800 ;
        RECT 45.930 5.050 46.680 6.800 ;
        RECT 46.830 2.150 46.980 9.700 ;
        RECT 47.430 2.150 47.580 9.700 ;
        RECT 48.030 2.150 48.180 9.700 ;
        RECT 48.630 2.150 48.780 9.700 ;
        RECT 49.230 2.150 49.380 9.700 ;
        RECT 49.830 2.150 49.980 9.700 ;
        RECT 54.230 9.200 55.230 9.700 ;
        RECT 50.880 9.050 58.580 9.200 ;
        RECT 54.230 8.600 55.230 9.050 ;
        RECT 50.880 8.450 58.580 8.600 ;
        RECT 54.230 8.000 55.230 8.450 ;
        RECT 50.880 7.850 58.580 8.000 ;
        RECT 54.230 7.400 55.230 7.850 ;
        RECT 50.880 7.250 58.580 7.400 ;
        RECT 54.230 6.800 55.230 7.250 ;
        RECT 50.880 6.650 58.580 6.800 ;
        RECT 54.230 6.200 55.230 6.650 ;
        RECT 50.880 6.050 58.580 6.200 ;
        RECT 54.230 5.600 55.230 6.050 ;
        RECT 50.880 5.450 58.580 5.600 ;
        RECT 54.230 5.000 55.230 5.450 ;
        RECT 50.880 4.850 58.580 5.000 ;
        RECT 54.230 4.400 55.230 4.850 ;
        RECT 50.880 4.250 58.580 4.400 ;
        RECT 54.230 3.800 55.230 4.250 ;
        RECT 50.880 3.650 58.580 3.800 ;
        RECT 54.230 3.200 55.230 3.650 ;
        RECT 50.880 3.050 58.580 3.200 ;
        RECT 54.230 2.600 55.230 3.050 ;
        RECT 50.880 2.450 58.580 2.600 ;
        RECT 54.230 2.000 55.230 2.450 ;
        RECT 59.480 2.150 59.630 9.700 ;
        RECT 60.080 2.150 60.230 9.700 ;
        RECT 60.680 2.150 60.830 9.700 ;
        RECT 61.280 2.150 61.430 9.700 ;
        RECT 61.880 2.150 62.030 9.700 ;
        RECT 62.480 2.150 62.630 9.700 ;
        RECT 62.780 9.550 63.930 9.700 ;
        RECT 64.580 9.550 64.880 10.450 ;
        RECT 65.530 10.300 66.680 10.450 ;
        RECT 66.830 10.300 66.980 17.850 ;
        RECT 67.430 10.300 67.580 17.850 ;
        RECT 68.030 10.300 68.180 17.850 ;
        RECT 68.630 10.300 68.780 17.850 ;
        RECT 69.230 10.300 69.380 17.850 ;
        RECT 69.830 10.300 69.980 17.850 ;
        RECT 74.230 17.550 75.230 18.000 ;
        RECT 70.880 17.400 78.580 17.550 ;
        RECT 74.230 16.950 75.230 17.400 ;
        RECT 70.880 16.800 78.580 16.950 ;
        RECT 74.230 16.350 75.230 16.800 ;
        RECT 70.880 16.200 78.580 16.350 ;
        RECT 74.230 15.750 75.230 16.200 ;
        RECT 70.880 15.600 78.580 15.750 ;
        RECT 74.230 15.150 75.230 15.600 ;
        RECT 70.880 15.000 78.580 15.150 ;
        RECT 74.230 14.550 75.230 15.000 ;
        RECT 70.880 14.400 78.580 14.550 ;
        RECT 74.230 13.950 75.230 14.400 ;
        RECT 70.880 13.800 78.580 13.950 ;
        RECT 74.230 13.350 75.230 13.800 ;
        RECT 70.880 13.200 78.580 13.350 ;
        RECT 74.230 12.750 75.230 13.200 ;
        RECT 70.880 12.600 78.580 12.750 ;
        RECT 74.230 12.150 75.230 12.600 ;
        RECT 70.880 12.000 78.580 12.150 ;
        RECT 74.230 11.550 75.230 12.000 ;
        RECT 70.880 11.400 78.580 11.550 ;
        RECT 74.230 10.950 75.230 11.400 ;
        RECT 70.880 10.800 78.580 10.950 ;
        RECT 74.230 10.300 75.230 10.800 ;
        RECT 79.480 10.300 79.630 17.850 ;
        RECT 80.080 10.300 80.230 17.850 ;
        RECT 80.680 10.300 80.830 17.850 ;
        RECT 81.280 10.300 81.430 17.850 ;
        RECT 81.880 10.300 82.030 17.850 ;
        RECT 82.480 10.300 82.630 17.850 ;
        RECT 82.780 13.200 83.530 15.000 ;
        RECT 85.930 13.200 86.680 15.000 ;
        RECT 82.780 10.450 86.680 13.200 ;
        RECT 82.780 10.300 83.930 10.450 ;
        RECT 65.530 9.700 83.930 10.300 ;
        RECT 65.530 9.550 66.680 9.700 ;
        RECT 62.780 6.800 66.680 9.550 ;
        RECT 62.780 5.050 63.530 6.800 ;
        RECT 65.930 5.050 66.680 6.800 ;
        RECT 66.830 2.150 66.980 9.700 ;
        RECT 67.430 2.150 67.580 9.700 ;
        RECT 68.030 2.150 68.180 9.700 ;
        RECT 68.630 2.150 68.780 9.700 ;
        RECT 69.230 2.150 69.380 9.700 ;
        RECT 69.830 2.150 69.980 9.700 ;
        RECT 74.230 9.200 75.230 9.700 ;
        RECT 70.880 9.050 78.580 9.200 ;
        RECT 74.230 8.600 75.230 9.050 ;
        RECT 70.880 8.450 78.580 8.600 ;
        RECT 74.230 8.000 75.230 8.450 ;
        RECT 70.880 7.850 78.580 8.000 ;
        RECT 74.230 7.400 75.230 7.850 ;
        RECT 70.880 7.250 78.580 7.400 ;
        RECT 74.230 6.800 75.230 7.250 ;
        RECT 70.880 6.650 78.580 6.800 ;
        RECT 74.230 6.200 75.230 6.650 ;
        RECT 70.880 6.050 78.580 6.200 ;
        RECT 74.230 5.600 75.230 6.050 ;
        RECT 70.880 5.450 78.580 5.600 ;
        RECT 74.230 5.000 75.230 5.450 ;
        RECT 70.880 4.850 78.580 5.000 ;
        RECT 74.230 4.400 75.230 4.850 ;
        RECT 70.880 4.250 78.580 4.400 ;
        RECT 74.230 3.800 75.230 4.250 ;
        RECT 70.880 3.650 78.580 3.800 ;
        RECT 74.230 3.200 75.230 3.650 ;
        RECT 70.880 3.050 78.580 3.200 ;
        RECT 74.230 2.600 75.230 3.050 ;
        RECT 70.880 2.450 78.580 2.600 ;
        RECT 74.230 2.000 75.230 2.450 ;
        RECT 79.480 2.150 79.630 9.700 ;
        RECT 80.080 2.150 80.230 9.700 ;
        RECT 80.680 2.150 80.830 9.700 ;
        RECT 81.280 2.150 81.430 9.700 ;
        RECT 81.880 2.150 82.030 9.700 ;
        RECT 82.480 2.150 82.630 9.700 ;
        RECT 82.780 9.550 83.930 9.700 ;
        RECT 84.580 9.550 84.880 10.450 ;
        RECT 85.530 10.300 86.680 10.450 ;
        RECT 86.830 10.300 86.980 17.850 ;
        RECT 87.430 10.300 87.580 17.850 ;
        RECT 88.030 10.300 88.180 17.850 ;
        RECT 88.630 10.300 88.780 17.850 ;
        RECT 89.230 10.300 89.380 17.850 ;
        RECT 89.830 10.300 89.980 17.850 ;
        RECT 94.230 17.550 95.230 18.000 ;
        RECT 90.880 17.400 98.580 17.550 ;
        RECT 94.230 16.950 95.230 17.400 ;
        RECT 90.880 16.800 98.580 16.950 ;
        RECT 94.230 16.350 95.230 16.800 ;
        RECT 90.880 16.200 98.580 16.350 ;
        RECT 94.230 15.750 95.230 16.200 ;
        RECT 90.880 15.600 98.580 15.750 ;
        RECT 94.230 15.150 95.230 15.600 ;
        RECT 90.880 15.000 98.580 15.150 ;
        RECT 94.230 14.550 95.230 15.000 ;
        RECT 90.880 14.400 98.580 14.550 ;
        RECT 94.230 13.950 95.230 14.400 ;
        RECT 90.880 13.800 98.580 13.950 ;
        RECT 94.230 13.350 95.230 13.800 ;
        RECT 90.880 13.200 98.580 13.350 ;
        RECT 94.230 12.750 95.230 13.200 ;
        RECT 90.880 12.600 98.580 12.750 ;
        RECT 94.230 12.150 95.230 12.600 ;
        RECT 90.880 12.000 98.580 12.150 ;
        RECT 94.230 11.550 95.230 12.000 ;
        RECT 90.880 11.400 98.580 11.550 ;
        RECT 94.230 10.950 95.230 11.400 ;
        RECT 90.880 10.800 98.580 10.950 ;
        RECT 94.230 10.300 95.230 10.800 ;
        RECT 99.480 10.300 99.630 17.850 ;
        RECT 100.080 10.300 100.230 17.850 ;
        RECT 100.680 10.300 100.830 17.850 ;
        RECT 101.280 10.300 101.430 17.850 ;
        RECT 101.880 10.300 102.030 17.850 ;
        RECT 102.480 10.300 102.630 17.850 ;
        RECT 102.780 13.200 103.530 15.000 ;
        RECT 105.930 13.200 106.680 15.000 ;
        RECT 102.780 10.450 106.680 13.200 ;
        RECT 102.780 10.300 103.930 10.450 ;
        RECT 85.530 9.700 103.930 10.300 ;
        RECT 85.530 9.550 86.680 9.700 ;
        RECT 82.780 6.800 86.680 9.550 ;
        RECT 82.780 5.050 83.530 6.800 ;
        RECT 85.930 5.050 86.680 6.800 ;
        RECT 86.830 2.150 86.980 9.700 ;
        RECT 87.430 2.150 87.580 9.700 ;
        RECT 88.030 2.150 88.180 9.700 ;
        RECT 88.630 2.150 88.780 9.700 ;
        RECT 89.230 2.150 89.380 9.700 ;
        RECT 89.830 2.150 89.980 9.700 ;
        RECT 94.230 9.200 95.230 9.700 ;
        RECT 90.880 9.050 98.580 9.200 ;
        RECT 94.230 8.600 95.230 9.050 ;
        RECT 90.880 8.450 98.580 8.600 ;
        RECT 94.230 8.000 95.230 8.450 ;
        RECT 90.880 7.850 98.580 8.000 ;
        RECT 94.230 7.400 95.230 7.850 ;
        RECT 90.880 7.250 98.580 7.400 ;
        RECT 94.230 6.800 95.230 7.250 ;
        RECT 90.880 6.650 98.580 6.800 ;
        RECT 94.230 6.200 95.230 6.650 ;
        RECT 90.880 6.050 98.580 6.200 ;
        RECT 94.230 5.600 95.230 6.050 ;
        RECT 90.880 5.450 98.580 5.600 ;
        RECT 94.230 5.000 95.230 5.450 ;
        RECT 90.880 4.850 98.580 5.000 ;
        RECT 94.230 4.400 95.230 4.850 ;
        RECT 90.880 4.250 98.580 4.400 ;
        RECT 94.230 3.800 95.230 4.250 ;
        RECT 90.880 3.650 98.580 3.800 ;
        RECT 94.230 3.200 95.230 3.650 ;
        RECT 90.880 3.050 98.580 3.200 ;
        RECT 94.230 2.600 95.230 3.050 ;
        RECT 90.880 2.450 98.580 2.600 ;
        RECT 94.230 2.000 95.230 2.450 ;
        RECT 99.480 2.150 99.630 9.700 ;
        RECT 100.080 2.150 100.230 9.700 ;
        RECT 100.680 2.150 100.830 9.700 ;
        RECT 101.280 2.150 101.430 9.700 ;
        RECT 101.880 2.150 102.030 9.700 ;
        RECT 102.480 2.150 102.630 9.700 ;
        RECT 102.780 9.550 103.930 9.700 ;
        RECT 104.580 9.550 104.880 10.450 ;
        RECT 105.530 10.300 106.680 10.450 ;
        RECT 106.830 10.300 106.980 17.850 ;
        RECT 107.430 10.300 107.580 17.850 ;
        RECT 108.030 10.300 108.180 17.850 ;
        RECT 108.630 10.300 108.780 17.850 ;
        RECT 109.230 10.300 109.380 17.850 ;
        RECT 109.830 10.300 109.980 17.850 ;
        RECT 114.230 17.550 115.230 18.000 ;
        RECT 110.880 17.400 118.580 17.550 ;
        RECT 114.230 16.950 115.230 17.400 ;
        RECT 110.880 16.800 118.580 16.950 ;
        RECT 114.230 16.350 115.230 16.800 ;
        RECT 110.880 16.200 118.580 16.350 ;
        RECT 114.230 15.750 115.230 16.200 ;
        RECT 110.880 15.600 118.580 15.750 ;
        RECT 114.230 15.150 115.230 15.600 ;
        RECT 110.880 15.000 118.580 15.150 ;
        RECT 114.230 14.550 115.230 15.000 ;
        RECT 110.880 14.400 118.580 14.550 ;
        RECT 114.230 13.950 115.230 14.400 ;
        RECT 110.880 13.800 118.580 13.950 ;
        RECT 114.230 13.350 115.230 13.800 ;
        RECT 110.880 13.200 118.580 13.350 ;
        RECT 114.230 12.750 115.230 13.200 ;
        RECT 110.880 12.600 118.580 12.750 ;
        RECT 114.230 12.150 115.230 12.600 ;
        RECT 110.880 12.000 118.580 12.150 ;
        RECT 114.230 11.550 115.230 12.000 ;
        RECT 110.880 11.400 118.580 11.550 ;
        RECT 114.230 10.950 115.230 11.400 ;
        RECT 110.880 10.800 118.580 10.950 ;
        RECT 114.230 10.300 115.230 10.800 ;
        RECT 119.480 10.300 119.630 17.850 ;
        RECT 120.080 10.300 120.230 17.850 ;
        RECT 120.680 10.300 120.830 17.850 ;
        RECT 121.280 10.300 121.430 17.850 ;
        RECT 121.880 10.300 122.030 17.850 ;
        RECT 122.480 10.300 122.630 17.850 ;
        RECT 122.780 13.200 123.530 15.000 ;
        RECT 122.780 11.525 124.730 13.200 ;
        RECT 122.780 10.450 131.850 11.525 ;
        RECT 122.780 10.300 123.930 10.450 ;
        RECT 105.530 9.700 123.930 10.300 ;
        RECT 105.530 9.550 106.680 9.700 ;
        RECT 102.780 6.800 106.680 9.550 ;
        RECT 102.780 5.050 103.530 6.800 ;
        RECT 105.930 5.050 106.680 6.800 ;
        RECT 106.830 2.150 106.980 9.700 ;
        RECT 107.430 2.150 107.580 9.700 ;
        RECT 108.030 2.150 108.180 9.700 ;
        RECT 108.630 2.150 108.780 9.700 ;
        RECT 109.230 2.150 109.380 9.700 ;
        RECT 109.830 2.150 109.980 9.700 ;
        RECT 114.230 9.200 115.230 9.700 ;
        RECT 110.880 9.050 118.580 9.200 ;
        RECT 114.230 8.600 115.230 9.050 ;
        RECT 110.880 8.450 118.580 8.600 ;
        RECT 114.230 8.000 115.230 8.450 ;
        RECT 110.880 7.850 118.580 8.000 ;
        RECT 114.230 7.400 115.230 7.850 ;
        RECT 110.880 7.250 118.580 7.400 ;
        RECT 114.230 6.800 115.230 7.250 ;
        RECT 110.880 6.650 118.580 6.800 ;
        RECT 114.230 6.200 115.230 6.650 ;
        RECT 110.880 6.050 118.580 6.200 ;
        RECT 114.230 5.600 115.230 6.050 ;
        RECT 110.880 5.450 118.580 5.600 ;
        RECT 114.230 5.000 115.230 5.450 ;
        RECT 110.880 4.850 118.580 5.000 ;
        RECT 114.230 4.400 115.230 4.850 ;
        RECT 110.880 4.250 118.580 4.400 ;
        RECT 114.230 3.800 115.230 4.250 ;
        RECT 110.880 3.650 118.580 3.800 ;
        RECT 114.230 3.200 115.230 3.650 ;
        RECT 110.880 3.050 118.580 3.200 ;
        RECT 114.230 2.600 115.230 3.050 ;
        RECT 110.880 2.450 118.580 2.600 ;
        RECT 114.230 2.000 115.230 2.450 ;
        RECT 119.480 2.150 119.630 9.700 ;
        RECT 120.080 2.150 120.230 9.700 ;
        RECT 120.680 2.150 120.830 9.700 ;
        RECT 121.280 2.150 121.430 9.700 ;
        RECT 121.880 2.150 122.030 9.700 ;
        RECT 122.480 2.150 122.630 9.700 ;
        RECT 122.780 9.550 123.930 9.700 ;
        RECT 124.580 10.250 131.850 10.450 ;
        RECT 124.580 9.550 124.730 10.250 ;
        RECT 122.780 6.800 124.730 9.550 ;
        RECT 122.780 5.050 123.530 6.800 ;
        RECT 10.880 1.850 18.580 2.000 ;
        RECT 30.880 1.850 38.580 2.000 ;
        RECT 50.880 1.850 58.580 2.000 ;
        RECT 70.880 1.850 78.580 2.000 ;
        RECT 90.880 1.850 98.580 2.000 ;
        RECT 110.880 1.850 118.580 2.000 ;
        RECT 14.230 1.200 15.230 1.850 ;
        RECT 34.230 1.200 35.230 1.850 ;
        RECT 54.230 1.200 55.230 1.850 ;
        RECT 74.230 1.200 75.230 1.850 ;
        RECT 94.230 1.200 95.230 1.850 ;
        RECT 114.230 1.200 115.230 1.850 ;
        RECT 11.530 0.000 17.930 1.200 ;
        RECT 31.530 0.000 37.930 1.200 ;
        RECT 51.530 0.000 57.930 1.200 ;
        RECT 71.530 0.000 77.930 1.200 ;
        RECT 91.530 0.000 97.930 1.200 ;
        RECT 111.530 0.000 117.930 1.200 ;
      LAYER via ;
        RECT 11.630 338.900 12.630 339.900 ;
        RECT 12.780 338.900 13.780 339.900 ;
        RECT 13.930 338.900 15.530 339.900 ;
        RECT 15.680 338.900 16.680 339.900 ;
        RECT 16.830 338.900 17.830 339.900 ;
        RECT 31.630 338.900 32.630 339.900 ;
        RECT 32.780 338.900 33.780 339.900 ;
        RECT 33.930 338.900 35.530 339.900 ;
        RECT 35.680 338.900 36.680 339.900 ;
        RECT 36.830 338.900 37.830 339.900 ;
        RECT 51.630 338.900 52.630 339.900 ;
        RECT 52.780 338.900 53.780 339.900 ;
        RECT 53.930 338.900 55.530 339.900 ;
        RECT 55.680 338.900 56.680 339.900 ;
        RECT 56.830 338.900 57.830 339.900 ;
        RECT 71.630 338.900 72.630 339.900 ;
        RECT 72.780 338.900 73.780 339.900 ;
        RECT 73.930 338.900 75.530 339.900 ;
        RECT 75.680 338.900 76.680 339.900 ;
        RECT 76.830 338.900 77.830 339.900 ;
        RECT 91.630 338.900 92.630 339.900 ;
        RECT 92.780 338.900 93.780 339.900 ;
        RECT 93.930 338.900 95.530 339.900 ;
        RECT 95.680 338.900 96.680 339.900 ;
        RECT 96.830 338.900 97.830 339.900 ;
        RECT 111.630 338.900 112.630 339.900 ;
        RECT 112.780 338.900 113.780 339.900 ;
        RECT 113.930 338.900 115.530 339.900 ;
        RECT 115.680 338.900 116.680 339.900 ;
        RECT 116.830 338.900 117.830 339.900 ;
        RECT 4.830 332.400 5.530 333.100 ;
        RECT 4.830 331.550 5.530 332.250 ;
        RECT 4.830 330.700 5.530 331.400 ;
        RECT 23.930 332.400 24.630 333.100 ;
        RECT 24.830 332.400 25.530 333.100 ;
        RECT 23.930 331.550 24.630 332.250 ;
        RECT 24.830 331.550 25.530 332.250 ;
        RECT 23.930 330.700 24.630 331.400 ;
        RECT 24.830 330.700 25.530 331.400 ;
        RECT 4.830 328.600 5.530 329.300 ;
        RECT 4.830 327.750 5.530 328.450 ;
        RECT 4.830 326.900 5.530 327.600 ;
        RECT 43.930 332.400 44.630 333.100 ;
        RECT 44.830 332.400 45.530 333.100 ;
        RECT 43.930 331.550 44.630 332.250 ;
        RECT 44.830 331.550 45.530 332.250 ;
        RECT 43.930 330.700 44.630 331.400 ;
        RECT 44.830 330.700 45.530 331.400 ;
        RECT 23.930 328.600 24.630 329.300 ;
        RECT 24.830 328.600 25.530 329.300 ;
        RECT 23.930 327.750 24.630 328.450 ;
        RECT 24.830 327.750 25.530 328.450 ;
        RECT 23.930 326.900 24.630 327.600 ;
        RECT 24.830 326.900 25.530 327.600 ;
        RECT 63.930 332.400 64.630 333.100 ;
        RECT 64.830 332.400 65.530 333.100 ;
        RECT 63.930 331.550 64.630 332.250 ;
        RECT 64.830 331.550 65.530 332.250 ;
        RECT 63.930 330.700 64.630 331.400 ;
        RECT 64.830 330.700 65.530 331.400 ;
        RECT 43.930 328.600 44.630 329.300 ;
        RECT 44.830 328.600 45.530 329.300 ;
        RECT 43.930 327.750 44.630 328.450 ;
        RECT 44.830 327.750 45.530 328.450 ;
        RECT 43.930 326.900 44.630 327.600 ;
        RECT 44.830 326.900 45.530 327.600 ;
        RECT 83.930 332.400 84.630 333.100 ;
        RECT 84.830 332.400 85.530 333.100 ;
        RECT 83.930 331.550 84.630 332.250 ;
        RECT 84.830 331.550 85.530 332.250 ;
        RECT 83.930 330.700 84.630 331.400 ;
        RECT 84.830 330.700 85.530 331.400 ;
        RECT 63.930 328.600 64.630 329.300 ;
        RECT 64.830 328.600 65.530 329.300 ;
        RECT 63.930 327.750 64.630 328.450 ;
        RECT 64.830 327.750 65.530 328.450 ;
        RECT 63.930 326.900 64.630 327.600 ;
        RECT 64.830 326.900 65.530 327.600 ;
        RECT 103.930 332.400 104.630 333.100 ;
        RECT 104.830 332.400 105.530 333.100 ;
        RECT 103.930 331.550 104.630 332.250 ;
        RECT 104.830 331.550 105.530 332.250 ;
        RECT 103.930 330.700 104.630 331.400 ;
        RECT 104.830 330.700 105.530 331.400 ;
        RECT 83.930 328.600 84.630 329.300 ;
        RECT 84.830 328.600 85.530 329.300 ;
        RECT 83.930 327.750 84.630 328.450 ;
        RECT 84.830 327.750 85.530 328.450 ;
        RECT 83.930 326.900 84.630 327.600 ;
        RECT 84.830 326.900 85.530 327.600 ;
        RECT 123.930 332.400 124.630 333.100 ;
        RECT 123.930 331.550 124.630 332.250 ;
        RECT 123.930 330.700 124.630 331.400 ;
        RECT 103.930 328.600 104.630 329.300 ;
        RECT 104.830 328.600 105.530 329.300 ;
        RECT 103.930 327.750 104.630 328.450 ;
        RECT 104.830 327.750 105.530 328.450 ;
        RECT 103.930 326.900 104.630 327.600 ;
        RECT 104.830 326.900 105.530 327.600 ;
        RECT 130.050 329.975 130.410 330.355 ;
        RECT 130.680 329.975 131.040 330.355 ;
        RECT 131.280 329.975 131.640 330.355 ;
        RECT 130.050 329.385 130.410 329.765 ;
        RECT 130.680 329.385 131.040 329.765 ;
        RECT 131.280 329.385 131.640 329.765 ;
        RECT 123.930 328.600 124.630 329.300 ;
        RECT 123.930 327.750 124.630 328.450 ;
        RECT 123.930 326.900 124.630 327.600 ;
        RECT 11.630 320.100 12.630 321.100 ;
        RECT 12.730 320.100 13.730 321.100 ;
        RECT 13.880 320.100 15.480 321.100 ;
        RECT 15.680 320.100 16.680 321.100 ;
        RECT 16.830 320.100 17.830 321.100 ;
        RECT 11.630 318.900 12.630 319.900 ;
        RECT 12.780 318.900 13.780 319.900 ;
        RECT 13.930 318.900 15.530 319.900 ;
        RECT 15.680 318.900 16.680 319.900 ;
        RECT 16.830 318.900 17.830 319.900 ;
        RECT 31.630 320.100 32.630 321.100 ;
        RECT 32.730 320.100 33.730 321.100 ;
        RECT 33.880 320.100 35.480 321.100 ;
        RECT 35.680 320.100 36.680 321.100 ;
        RECT 36.830 320.100 37.830 321.100 ;
        RECT 31.630 318.900 32.630 319.900 ;
        RECT 32.780 318.900 33.780 319.900 ;
        RECT 33.930 318.900 35.530 319.900 ;
        RECT 35.680 318.900 36.680 319.900 ;
        RECT 36.830 318.900 37.830 319.900 ;
        RECT 51.630 320.100 52.630 321.100 ;
        RECT 52.730 320.100 53.730 321.100 ;
        RECT 53.880 320.100 55.480 321.100 ;
        RECT 55.680 320.100 56.680 321.100 ;
        RECT 56.830 320.100 57.830 321.100 ;
        RECT 51.630 318.900 52.630 319.900 ;
        RECT 52.780 318.900 53.780 319.900 ;
        RECT 53.930 318.900 55.530 319.900 ;
        RECT 55.680 318.900 56.680 319.900 ;
        RECT 56.830 318.900 57.830 319.900 ;
        RECT 71.630 320.100 72.630 321.100 ;
        RECT 72.730 320.100 73.730 321.100 ;
        RECT 73.880 320.100 75.480 321.100 ;
        RECT 75.680 320.100 76.680 321.100 ;
        RECT 76.830 320.100 77.830 321.100 ;
        RECT 71.630 318.900 72.630 319.900 ;
        RECT 72.780 318.900 73.780 319.900 ;
        RECT 73.930 318.900 75.530 319.900 ;
        RECT 75.680 318.900 76.680 319.900 ;
        RECT 76.830 318.900 77.830 319.900 ;
        RECT 91.630 320.100 92.630 321.100 ;
        RECT 92.730 320.100 93.730 321.100 ;
        RECT 93.880 320.100 95.480 321.100 ;
        RECT 95.680 320.100 96.680 321.100 ;
        RECT 96.830 320.100 97.830 321.100 ;
        RECT 91.630 318.900 92.630 319.900 ;
        RECT 92.780 318.900 93.780 319.900 ;
        RECT 93.930 318.900 95.530 319.900 ;
        RECT 95.680 318.900 96.680 319.900 ;
        RECT 96.830 318.900 97.830 319.900 ;
        RECT 111.630 320.100 112.630 321.100 ;
        RECT 112.730 320.100 113.730 321.100 ;
        RECT 113.880 320.100 115.480 321.100 ;
        RECT 115.680 320.100 116.680 321.100 ;
        RECT 116.830 320.100 117.830 321.100 ;
        RECT 111.630 318.900 112.630 319.900 ;
        RECT 112.780 318.900 113.780 319.900 ;
        RECT 113.930 318.900 115.530 319.900 ;
        RECT 115.680 318.900 116.680 319.900 ;
        RECT 116.830 318.900 117.830 319.900 ;
        RECT 4.830 312.400 5.530 313.100 ;
        RECT 4.830 311.550 5.530 312.250 ;
        RECT 4.830 310.700 5.530 311.400 ;
        RECT 23.930 312.400 24.630 313.100 ;
        RECT 24.830 312.400 25.530 313.100 ;
        RECT 23.930 311.550 24.630 312.250 ;
        RECT 24.830 311.550 25.530 312.250 ;
        RECT 23.930 310.700 24.630 311.400 ;
        RECT 24.830 310.700 25.530 311.400 ;
        RECT 4.830 308.600 5.530 309.300 ;
        RECT 4.830 307.750 5.530 308.450 ;
        RECT 4.830 306.900 5.530 307.600 ;
        RECT 43.930 312.400 44.630 313.100 ;
        RECT 44.830 312.400 45.530 313.100 ;
        RECT 43.930 311.550 44.630 312.250 ;
        RECT 44.830 311.550 45.530 312.250 ;
        RECT 43.930 310.700 44.630 311.400 ;
        RECT 44.830 310.700 45.530 311.400 ;
        RECT 23.930 308.600 24.630 309.300 ;
        RECT 24.830 308.600 25.530 309.300 ;
        RECT 23.930 307.750 24.630 308.450 ;
        RECT 24.830 307.750 25.530 308.450 ;
        RECT 23.930 306.900 24.630 307.600 ;
        RECT 24.830 306.900 25.530 307.600 ;
        RECT 63.930 312.400 64.630 313.100 ;
        RECT 64.830 312.400 65.530 313.100 ;
        RECT 63.930 311.550 64.630 312.250 ;
        RECT 64.830 311.550 65.530 312.250 ;
        RECT 63.930 310.700 64.630 311.400 ;
        RECT 64.830 310.700 65.530 311.400 ;
        RECT 43.930 308.600 44.630 309.300 ;
        RECT 44.830 308.600 45.530 309.300 ;
        RECT 43.930 307.750 44.630 308.450 ;
        RECT 44.830 307.750 45.530 308.450 ;
        RECT 43.930 306.900 44.630 307.600 ;
        RECT 44.830 306.900 45.530 307.600 ;
        RECT 83.930 312.400 84.630 313.100 ;
        RECT 84.830 312.400 85.530 313.100 ;
        RECT 83.930 311.550 84.630 312.250 ;
        RECT 84.830 311.550 85.530 312.250 ;
        RECT 83.930 310.700 84.630 311.400 ;
        RECT 84.830 310.700 85.530 311.400 ;
        RECT 63.930 308.600 64.630 309.300 ;
        RECT 64.830 308.600 65.530 309.300 ;
        RECT 63.930 307.750 64.630 308.450 ;
        RECT 64.830 307.750 65.530 308.450 ;
        RECT 63.930 306.900 64.630 307.600 ;
        RECT 64.830 306.900 65.530 307.600 ;
        RECT 103.930 312.400 104.630 313.100 ;
        RECT 104.830 312.400 105.530 313.100 ;
        RECT 103.930 311.550 104.630 312.250 ;
        RECT 104.830 311.550 105.530 312.250 ;
        RECT 103.930 310.700 104.630 311.400 ;
        RECT 104.830 310.700 105.530 311.400 ;
        RECT 83.930 308.600 84.630 309.300 ;
        RECT 84.830 308.600 85.530 309.300 ;
        RECT 83.930 307.750 84.630 308.450 ;
        RECT 84.830 307.750 85.530 308.450 ;
        RECT 83.930 306.900 84.630 307.600 ;
        RECT 84.830 306.900 85.530 307.600 ;
        RECT 123.930 312.400 124.630 313.100 ;
        RECT 123.930 311.550 124.630 312.250 ;
        RECT 123.930 310.700 124.630 311.400 ;
        RECT 103.930 308.600 104.630 309.300 ;
        RECT 104.830 308.600 105.530 309.300 ;
        RECT 103.930 307.750 104.630 308.450 ;
        RECT 104.830 307.750 105.530 308.450 ;
        RECT 103.930 306.900 104.630 307.600 ;
        RECT 104.830 306.900 105.530 307.600 ;
        RECT 130.050 309.910 130.410 310.290 ;
        RECT 130.680 309.910 131.040 310.290 ;
        RECT 131.280 309.910 131.640 310.290 ;
        RECT 130.050 309.320 130.410 309.700 ;
        RECT 130.680 309.320 131.040 309.700 ;
        RECT 131.280 309.320 131.640 309.700 ;
        RECT 123.930 308.600 124.630 309.300 ;
        RECT 123.930 307.750 124.630 308.450 ;
        RECT 123.930 306.900 124.630 307.600 ;
        RECT 11.630 300.100 12.630 301.100 ;
        RECT 12.730 300.100 13.730 301.100 ;
        RECT 13.880 300.100 15.480 301.100 ;
        RECT 15.680 300.100 16.680 301.100 ;
        RECT 16.830 300.100 17.830 301.100 ;
        RECT 11.630 298.900 12.630 299.900 ;
        RECT 12.780 298.900 13.780 299.900 ;
        RECT 13.930 298.900 15.530 299.900 ;
        RECT 15.680 298.900 16.680 299.900 ;
        RECT 16.830 298.900 17.830 299.900 ;
        RECT 31.630 300.100 32.630 301.100 ;
        RECT 32.730 300.100 33.730 301.100 ;
        RECT 33.880 300.100 35.480 301.100 ;
        RECT 35.680 300.100 36.680 301.100 ;
        RECT 36.830 300.100 37.830 301.100 ;
        RECT 31.630 298.900 32.630 299.900 ;
        RECT 32.780 298.900 33.780 299.900 ;
        RECT 33.930 298.900 35.530 299.900 ;
        RECT 35.680 298.900 36.680 299.900 ;
        RECT 36.830 298.900 37.830 299.900 ;
        RECT 51.630 300.100 52.630 301.100 ;
        RECT 52.730 300.100 53.730 301.100 ;
        RECT 53.880 300.100 55.480 301.100 ;
        RECT 55.680 300.100 56.680 301.100 ;
        RECT 56.830 300.100 57.830 301.100 ;
        RECT 51.630 298.900 52.630 299.900 ;
        RECT 52.780 298.900 53.780 299.900 ;
        RECT 53.930 298.900 55.530 299.900 ;
        RECT 55.680 298.900 56.680 299.900 ;
        RECT 56.830 298.900 57.830 299.900 ;
        RECT 71.630 300.100 72.630 301.100 ;
        RECT 72.730 300.100 73.730 301.100 ;
        RECT 73.880 300.100 75.480 301.100 ;
        RECT 75.680 300.100 76.680 301.100 ;
        RECT 76.830 300.100 77.830 301.100 ;
        RECT 71.630 298.900 72.630 299.900 ;
        RECT 72.780 298.900 73.780 299.900 ;
        RECT 73.930 298.900 75.530 299.900 ;
        RECT 75.680 298.900 76.680 299.900 ;
        RECT 76.830 298.900 77.830 299.900 ;
        RECT 91.630 300.100 92.630 301.100 ;
        RECT 92.730 300.100 93.730 301.100 ;
        RECT 93.880 300.100 95.480 301.100 ;
        RECT 95.680 300.100 96.680 301.100 ;
        RECT 96.830 300.100 97.830 301.100 ;
        RECT 91.630 298.900 92.630 299.900 ;
        RECT 92.780 298.900 93.780 299.900 ;
        RECT 93.930 298.900 95.530 299.900 ;
        RECT 95.680 298.900 96.680 299.900 ;
        RECT 96.830 298.900 97.830 299.900 ;
        RECT 111.630 300.100 112.630 301.100 ;
        RECT 112.730 300.100 113.730 301.100 ;
        RECT 113.880 300.100 115.480 301.100 ;
        RECT 115.680 300.100 116.680 301.100 ;
        RECT 116.830 300.100 117.830 301.100 ;
        RECT 111.630 298.900 112.630 299.900 ;
        RECT 112.780 298.900 113.780 299.900 ;
        RECT 113.930 298.900 115.530 299.900 ;
        RECT 115.680 298.900 116.680 299.900 ;
        RECT 116.830 298.900 117.830 299.900 ;
        RECT 4.830 292.400 5.530 293.100 ;
        RECT 4.830 291.550 5.530 292.250 ;
        RECT 4.830 290.700 5.530 291.400 ;
        RECT 23.930 292.400 24.630 293.100 ;
        RECT 24.830 292.400 25.530 293.100 ;
        RECT 23.930 291.550 24.630 292.250 ;
        RECT 24.830 291.550 25.530 292.250 ;
        RECT 23.930 290.700 24.630 291.400 ;
        RECT 24.830 290.700 25.530 291.400 ;
        RECT 4.830 288.600 5.530 289.300 ;
        RECT 4.830 287.750 5.530 288.450 ;
        RECT 4.830 286.900 5.530 287.600 ;
        RECT 43.930 292.400 44.630 293.100 ;
        RECT 44.830 292.400 45.530 293.100 ;
        RECT 43.930 291.550 44.630 292.250 ;
        RECT 44.830 291.550 45.530 292.250 ;
        RECT 43.930 290.700 44.630 291.400 ;
        RECT 44.830 290.700 45.530 291.400 ;
        RECT 23.930 288.600 24.630 289.300 ;
        RECT 24.830 288.600 25.530 289.300 ;
        RECT 23.930 287.750 24.630 288.450 ;
        RECT 24.830 287.750 25.530 288.450 ;
        RECT 23.930 286.900 24.630 287.600 ;
        RECT 24.830 286.900 25.530 287.600 ;
        RECT 63.930 292.400 64.630 293.100 ;
        RECT 64.830 292.400 65.530 293.100 ;
        RECT 63.930 291.550 64.630 292.250 ;
        RECT 64.830 291.550 65.530 292.250 ;
        RECT 63.930 290.700 64.630 291.400 ;
        RECT 64.830 290.700 65.530 291.400 ;
        RECT 43.930 288.600 44.630 289.300 ;
        RECT 44.830 288.600 45.530 289.300 ;
        RECT 43.930 287.750 44.630 288.450 ;
        RECT 44.830 287.750 45.530 288.450 ;
        RECT 43.930 286.900 44.630 287.600 ;
        RECT 44.830 286.900 45.530 287.600 ;
        RECT 83.930 292.400 84.630 293.100 ;
        RECT 84.830 292.400 85.530 293.100 ;
        RECT 83.930 291.550 84.630 292.250 ;
        RECT 84.830 291.550 85.530 292.250 ;
        RECT 83.930 290.700 84.630 291.400 ;
        RECT 84.830 290.700 85.530 291.400 ;
        RECT 63.930 288.600 64.630 289.300 ;
        RECT 64.830 288.600 65.530 289.300 ;
        RECT 63.930 287.750 64.630 288.450 ;
        RECT 64.830 287.750 65.530 288.450 ;
        RECT 63.930 286.900 64.630 287.600 ;
        RECT 64.830 286.900 65.530 287.600 ;
        RECT 103.930 292.400 104.630 293.100 ;
        RECT 104.830 292.400 105.530 293.100 ;
        RECT 103.930 291.550 104.630 292.250 ;
        RECT 104.830 291.550 105.530 292.250 ;
        RECT 103.930 290.700 104.630 291.400 ;
        RECT 104.830 290.700 105.530 291.400 ;
        RECT 83.930 288.600 84.630 289.300 ;
        RECT 84.830 288.600 85.530 289.300 ;
        RECT 83.930 287.750 84.630 288.450 ;
        RECT 84.830 287.750 85.530 288.450 ;
        RECT 83.930 286.900 84.630 287.600 ;
        RECT 84.830 286.900 85.530 287.600 ;
        RECT 123.930 292.400 124.630 293.100 ;
        RECT 123.930 291.550 124.630 292.250 ;
        RECT 123.930 290.700 124.630 291.400 ;
        RECT 103.930 288.600 104.630 289.300 ;
        RECT 104.830 288.600 105.530 289.300 ;
        RECT 103.930 287.750 104.630 288.450 ;
        RECT 104.830 287.750 105.530 288.450 ;
        RECT 103.930 286.900 104.630 287.600 ;
        RECT 104.830 286.900 105.530 287.600 ;
        RECT 130.050 289.905 130.410 290.285 ;
        RECT 130.680 289.905 131.040 290.285 ;
        RECT 131.280 289.905 131.640 290.285 ;
        RECT 130.050 289.315 130.410 289.695 ;
        RECT 130.680 289.315 131.040 289.695 ;
        RECT 131.280 289.315 131.640 289.695 ;
        RECT 123.930 288.600 124.630 289.300 ;
        RECT 123.930 287.750 124.630 288.450 ;
        RECT 123.930 286.900 124.630 287.600 ;
        RECT 11.630 280.100 12.630 281.100 ;
        RECT 12.730 280.100 13.730 281.100 ;
        RECT 13.880 280.100 15.480 281.100 ;
        RECT 15.680 280.100 16.680 281.100 ;
        RECT 16.830 280.100 17.830 281.100 ;
        RECT 11.630 278.900 12.630 279.900 ;
        RECT 12.780 278.900 13.780 279.900 ;
        RECT 13.930 278.900 15.530 279.900 ;
        RECT 15.680 278.900 16.680 279.900 ;
        RECT 16.830 278.900 17.830 279.900 ;
        RECT 31.630 280.100 32.630 281.100 ;
        RECT 32.730 280.100 33.730 281.100 ;
        RECT 33.880 280.100 35.480 281.100 ;
        RECT 35.680 280.100 36.680 281.100 ;
        RECT 36.830 280.100 37.830 281.100 ;
        RECT 31.630 278.900 32.630 279.900 ;
        RECT 32.780 278.900 33.780 279.900 ;
        RECT 33.930 278.900 35.530 279.900 ;
        RECT 35.680 278.900 36.680 279.900 ;
        RECT 36.830 278.900 37.830 279.900 ;
        RECT 51.630 280.100 52.630 281.100 ;
        RECT 52.730 280.100 53.730 281.100 ;
        RECT 53.880 280.100 55.480 281.100 ;
        RECT 55.680 280.100 56.680 281.100 ;
        RECT 56.830 280.100 57.830 281.100 ;
        RECT 51.630 278.900 52.630 279.900 ;
        RECT 52.780 278.900 53.780 279.900 ;
        RECT 53.930 278.900 55.530 279.900 ;
        RECT 55.680 278.900 56.680 279.900 ;
        RECT 56.830 278.900 57.830 279.900 ;
        RECT 71.630 280.100 72.630 281.100 ;
        RECT 72.730 280.100 73.730 281.100 ;
        RECT 73.880 280.100 75.480 281.100 ;
        RECT 75.680 280.100 76.680 281.100 ;
        RECT 76.830 280.100 77.830 281.100 ;
        RECT 71.630 278.900 72.630 279.900 ;
        RECT 72.780 278.900 73.780 279.900 ;
        RECT 73.930 278.900 75.530 279.900 ;
        RECT 75.680 278.900 76.680 279.900 ;
        RECT 76.830 278.900 77.830 279.900 ;
        RECT 91.630 280.100 92.630 281.100 ;
        RECT 92.730 280.100 93.730 281.100 ;
        RECT 93.880 280.100 95.480 281.100 ;
        RECT 95.680 280.100 96.680 281.100 ;
        RECT 96.830 280.100 97.830 281.100 ;
        RECT 91.630 278.900 92.630 279.900 ;
        RECT 92.780 278.900 93.780 279.900 ;
        RECT 93.930 278.900 95.530 279.900 ;
        RECT 95.680 278.900 96.680 279.900 ;
        RECT 96.830 278.900 97.830 279.900 ;
        RECT 111.630 280.100 112.630 281.100 ;
        RECT 112.730 280.100 113.730 281.100 ;
        RECT 113.880 280.100 115.480 281.100 ;
        RECT 115.680 280.100 116.680 281.100 ;
        RECT 116.830 280.100 117.830 281.100 ;
        RECT 111.630 278.900 112.630 279.900 ;
        RECT 112.780 278.900 113.780 279.900 ;
        RECT 113.930 278.900 115.530 279.900 ;
        RECT 115.680 278.900 116.680 279.900 ;
        RECT 116.830 278.900 117.830 279.900 ;
        RECT 4.830 272.400 5.530 273.100 ;
        RECT 4.830 271.550 5.530 272.250 ;
        RECT 4.830 270.700 5.530 271.400 ;
        RECT 23.930 272.400 24.630 273.100 ;
        RECT 24.830 272.400 25.530 273.100 ;
        RECT 23.930 271.550 24.630 272.250 ;
        RECT 24.830 271.550 25.530 272.250 ;
        RECT 23.930 270.700 24.630 271.400 ;
        RECT 24.830 270.700 25.530 271.400 ;
        RECT 4.830 268.600 5.530 269.300 ;
        RECT 4.830 267.750 5.530 268.450 ;
        RECT 4.830 266.900 5.530 267.600 ;
        RECT 43.930 272.400 44.630 273.100 ;
        RECT 44.830 272.400 45.530 273.100 ;
        RECT 43.930 271.550 44.630 272.250 ;
        RECT 44.830 271.550 45.530 272.250 ;
        RECT 43.930 270.700 44.630 271.400 ;
        RECT 44.830 270.700 45.530 271.400 ;
        RECT 23.930 268.600 24.630 269.300 ;
        RECT 24.830 268.600 25.530 269.300 ;
        RECT 23.930 267.750 24.630 268.450 ;
        RECT 24.830 267.750 25.530 268.450 ;
        RECT 23.930 266.900 24.630 267.600 ;
        RECT 24.830 266.900 25.530 267.600 ;
        RECT 63.930 272.400 64.630 273.100 ;
        RECT 64.830 272.400 65.530 273.100 ;
        RECT 63.930 271.550 64.630 272.250 ;
        RECT 64.830 271.550 65.530 272.250 ;
        RECT 63.930 270.700 64.630 271.400 ;
        RECT 64.830 270.700 65.530 271.400 ;
        RECT 43.930 268.600 44.630 269.300 ;
        RECT 44.830 268.600 45.530 269.300 ;
        RECT 43.930 267.750 44.630 268.450 ;
        RECT 44.830 267.750 45.530 268.450 ;
        RECT 43.930 266.900 44.630 267.600 ;
        RECT 44.830 266.900 45.530 267.600 ;
        RECT 83.930 272.400 84.630 273.100 ;
        RECT 84.830 272.400 85.530 273.100 ;
        RECT 83.930 271.550 84.630 272.250 ;
        RECT 84.830 271.550 85.530 272.250 ;
        RECT 83.930 270.700 84.630 271.400 ;
        RECT 84.830 270.700 85.530 271.400 ;
        RECT 63.930 268.600 64.630 269.300 ;
        RECT 64.830 268.600 65.530 269.300 ;
        RECT 63.930 267.750 64.630 268.450 ;
        RECT 64.830 267.750 65.530 268.450 ;
        RECT 63.930 266.900 64.630 267.600 ;
        RECT 64.830 266.900 65.530 267.600 ;
        RECT 103.930 272.400 104.630 273.100 ;
        RECT 104.830 272.400 105.530 273.100 ;
        RECT 103.930 271.550 104.630 272.250 ;
        RECT 104.830 271.550 105.530 272.250 ;
        RECT 103.930 270.700 104.630 271.400 ;
        RECT 104.830 270.700 105.530 271.400 ;
        RECT 83.930 268.600 84.630 269.300 ;
        RECT 84.830 268.600 85.530 269.300 ;
        RECT 83.930 267.750 84.630 268.450 ;
        RECT 84.830 267.750 85.530 268.450 ;
        RECT 83.930 266.900 84.630 267.600 ;
        RECT 84.830 266.900 85.530 267.600 ;
        RECT 123.930 272.400 124.630 273.100 ;
        RECT 123.930 271.550 124.630 272.250 ;
        RECT 123.930 270.700 124.630 271.400 ;
        RECT 103.930 268.600 104.630 269.300 ;
        RECT 104.830 268.600 105.530 269.300 ;
        RECT 103.930 267.750 104.630 268.450 ;
        RECT 104.830 267.750 105.530 268.450 ;
        RECT 103.930 266.900 104.630 267.600 ;
        RECT 104.830 266.900 105.530 267.600 ;
        RECT 130.050 270.100 130.410 270.480 ;
        RECT 130.680 270.100 131.040 270.480 ;
        RECT 131.280 270.100 131.640 270.480 ;
        RECT 130.050 269.510 130.410 269.890 ;
        RECT 130.680 269.510 131.040 269.890 ;
        RECT 131.280 269.510 131.640 269.890 ;
        RECT 123.930 268.600 124.630 269.300 ;
        RECT 123.930 267.750 124.630 268.450 ;
        RECT 123.930 266.900 124.630 267.600 ;
        RECT 11.630 260.100 12.630 261.100 ;
        RECT 12.730 260.100 13.730 261.100 ;
        RECT 13.880 260.100 15.480 261.100 ;
        RECT 15.680 260.100 16.680 261.100 ;
        RECT 16.830 260.100 17.830 261.100 ;
        RECT 11.630 258.900 12.630 259.900 ;
        RECT 12.780 258.900 13.780 259.900 ;
        RECT 13.930 258.900 15.530 259.900 ;
        RECT 15.680 258.900 16.680 259.900 ;
        RECT 16.830 258.900 17.830 259.900 ;
        RECT 31.630 260.100 32.630 261.100 ;
        RECT 32.730 260.100 33.730 261.100 ;
        RECT 33.880 260.100 35.480 261.100 ;
        RECT 35.680 260.100 36.680 261.100 ;
        RECT 36.830 260.100 37.830 261.100 ;
        RECT 31.630 258.900 32.630 259.900 ;
        RECT 32.780 258.900 33.780 259.900 ;
        RECT 33.930 258.900 35.530 259.900 ;
        RECT 35.680 258.900 36.680 259.900 ;
        RECT 36.830 258.900 37.830 259.900 ;
        RECT 51.630 260.100 52.630 261.100 ;
        RECT 52.730 260.100 53.730 261.100 ;
        RECT 53.880 260.100 55.480 261.100 ;
        RECT 55.680 260.100 56.680 261.100 ;
        RECT 56.830 260.100 57.830 261.100 ;
        RECT 51.630 258.900 52.630 259.900 ;
        RECT 52.780 258.900 53.780 259.900 ;
        RECT 53.930 258.900 55.530 259.900 ;
        RECT 55.680 258.900 56.680 259.900 ;
        RECT 56.830 258.900 57.830 259.900 ;
        RECT 71.630 260.100 72.630 261.100 ;
        RECT 72.730 260.100 73.730 261.100 ;
        RECT 73.880 260.100 75.480 261.100 ;
        RECT 75.680 260.100 76.680 261.100 ;
        RECT 76.830 260.100 77.830 261.100 ;
        RECT 71.630 258.900 72.630 259.900 ;
        RECT 72.780 258.900 73.780 259.900 ;
        RECT 73.930 258.900 75.530 259.900 ;
        RECT 75.680 258.900 76.680 259.900 ;
        RECT 76.830 258.900 77.830 259.900 ;
        RECT 91.630 260.100 92.630 261.100 ;
        RECT 92.730 260.100 93.730 261.100 ;
        RECT 93.880 260.100 95.480 261.100 ;
        RECT 95.680 260.100 96.680 261.100 ;
        RECT 96.830 260.100 97.830 261.100 ;
        RECT 91.630 258.900 92.630 259.900 ;
        RECT 92.780 258.900 93.780 259.900 ;
        RECT 93.930 258.900 95.530 259.900 ;
        RECT 95.680 258.900 96.680 259.900 ;
        RECT 96.830 258.900 97.830 259.900 ;
        RECT 111.630 260.100 112.630 261.100 ;
        RECT 112.730 260.100 113.730 261.100 ;
        RECT 113.880 260.100 115.480 261.100 ;
        RECT 115.680 260.100 116.680 261.100 ;
        RECT 116.830 260.100 117.830 261.100 ;
        RECT 111.630 258.900 112.630 259.900 ;
        RECT 112.780 258.900 113.780 259.900 ;
        RECT 113.930 258.900 115.530 259.900 ;
        RECT 115.680 258.900 116.680 259.900 ;
        RECT 116.830 258.900 117.830 259.900 ;
        RECT 4.830 252.400 5.530 253.100 ;
        RECT 4.830 251.550 5.530 252.250 ;
        RECT 4.830 250.700 5.530 251.400 ;
        RECT 23.930 252.400 24.630 253.100 ;
        RECT 24.830 252.400 25.530 253.100 ;
        RECT 23.930 251.550 24.630 252.250 ;
        RECT 24.830 251.550 25.530 252.250 ;
        RECT 23.930 250.700 24.630 251.400 ;
        RECT 24.830 250.700 25.530 251.400 ;
        RECT 4.830 248.600 5.530 249.300 ;
        RECT 4.830 247.750 5.530 248.450 ;
        RECT 4.830 246.900 5.530 247.600 ;
        RECT 43.930 252.400 44.630 253.100 ;
        RECT 44.830 252.400 45.530 253.100 ;
        RECT 43.930 251.550 44.630 252.250 ;
        RECT 44.830 251.550 45.530 252.250 ;
        RECT 43.930 250.700 44.630 251.400 ;
        RECT 44.830 250.700 45.530 251.400 ;
        RECT 23.930 248.600 24.630 249.300 ;
        RECT 24.830 248.600 25.530 249.300 ;
        RECT 23.930 247.750 24.630 248.450 ;
        RECT 24.830 247.750 25.530 248.450 ;
        RECT 23.930 246.900 24.630 247.600 ;
        RECT 24.830 246.900 25.530 247.600 ;
        RECT 63.930 252.400 64.630 253.100 ;
        RECT 64.830 252.400 65.530 253.100 ;
        RECT 63.930 251.550 64.630 252.250 ;
        RECT 64.830 251.550 65.530 252.250 ;
        RECT 63.930 250.700 64.630 251.400 ;
        RECT 64.830 250.700 65.530 251.400 ;
        RECT 43.930 248.600 44.630 249.300 ;
        RECT 44.830 248.600 45.530 249.300 ;
        RECT 43.930 247.750 44.630 248.450 ;
        RECT 44.830 247.750 45.530 248.450 ;
        RECT 43.930 246.900 44.630 247.600 ;
        RECT 44.830 246.900 45.530 247.600 ;
        RECT 83.930 252.400 84.630 253.100 ;
        RECT 84.830 252.400 85.530 253.100 ;
        RECT 83.930 251.550 84.630 252.250 ;
        RECT 84.830 251.550 85.530 252.250 ;
        RECT 83.930 250.700 84.630 251.400 ;
        RECT 84.830 250.700 85.530 251.400 ;
        RECT 63.930 248.600 64.630 249.300 ;
        RECT 64.830 248.600 65.530 249.300 ;
        RECT 63.930 247.750 64.630 248.450 ;
        RECT 64.830 247.750 65.530 248.450 ;
        RECT 63.930 246.900 64.630 247.600 ;
        RECT 64.830 246.900 65.530 247.600 ;
        RECT 103.930 252.400 104.630 253.100 ;
        RECT 104.830 252.400 105.530 253.100 ;
        RECT 103.930 251.550 104.630 252.250 ;
        RECT 104.830 251.550 105.530 252.250 ;
        RECT 103.930 250.700 104.630 251.400 ;
        RECT 104.830 250.700 105.530 251.400 ;
        RECT 83.930 248.600 84.630 249.300 ;
        RECT 84.830 248.600 85.530 249.300 ;
        RECT 83.930 247.750 84.630 248.450 ;
        RECT 84.830 247.750 85.530 248.450 ;
        RECT 83.930 246.900 84.630 247.600 ;
        RECT 84.830 246.900 85.530 247.600 ;
        RECT 123.930 252.400 124.630 253.100 ;
        RECT 123.930 251.550 124.630 252.250 ;
        RECT 123.930 250.700 124.630 251.400 ;
        RECT 103.930 248.600 104.630 249.300 ;
        RECT 104.830 248.600 105.530 249.300 ;
        RECT 103.930 247.750 104.630 248.450 ;
        RECT 104.830 247.750 105.530 248.450 ;
        RECT 103.930 246.900 104.630 247.600 ;
        RECT 104.830 246.900 105.530 247.600 ;
        RECT 130.050 250.015 130.410 250.395 ;
        RECT 130.680 250.015 131.040 250.395 ;
        RECT 131.280 250.015 131.640 250.395 ;
        RECT 130.050 249.425 130.410 249.805 ;
        RECT 130.680 249.425 131.040 249.805 ;
        RECT 131.280 249.425 131.640 249.805 ;
        RECT 123.930 248.600 124.630 249.300 ;
        RECT 123.930 247.750 124.630 248.450 ;
        RECT 123.930 246.900 124.630 247.600 ;
        RECT 11.630 240.100 12.630 241.100 ;
        RECT 12.730 240.100 13.730 241.100 ;
        RECT 13.880 240.100 15.480 241.100 ;
        RECT 15.680 240.100 16.680 241.100 ;
        RECT 16.830 240.100 17.830 241.100 ;
        RECT 11.630 238.900 12.630 239.900 ;
        RECT 12.780 238.900 13.780 239.900 ;
        RECT 13.930 238.900 15.530 239.900 ;
        RECT 15.680 238.900 16.680 239.900 ;
        RECT 16.830 238.900 17.830 239.900 ;
        RECT 31.630 240.100 32.630 241.100 ;
        RECT 32.730 240.100 33.730 241.100 ;
        RECT 33.880 240.100 35.480 241.100 ;
        RECT 35.680 240.100 36.680 241.100 ;
        RECT 36.830 240.100 37.830 241.100 ;
        RECT 31.630 238.900 32.630 239.900 ;
        RECT 32.780 238.900 33.780 239.900 ;
        RECT 33.930 238.900 35.530 239.900 ;
        RECT 35.680 238.900 36.680 239.900 ;
        RECT 36.830 238.900 37.830 239.900 ;
        RECT 51.630 240.100 52.630 241.100 ;
        RECT 52.730 240.100 53.730 241.100 ;
        RECT 53.880 240.100 55.480 241.100 ;
        RECT 55.680 240.100 56.680 241.100 ;
        RECT 56.830 240.100 57.830 241.100 ;
        RECT 51.630 238.900 52.630 239.900 ;
        RECT 52.780 238.900 53.780 239.900 ;
        RECT 53.930 238.900 55.530 239.900 ;
        RECT 55.680 238.900 56.680 239.900 ;
        RECT 56.830 238.900 57.830 239.900 ;
        RECT 71.630 240.100 72.630 241.100 ;
        RECT 72.730 240.100 73.730 241.100 ;
        RECT 73.880 240.100 75.480 241.100 ;
        RECT 75.680 240.100 76.680 241.100 ;
        RECT 76.830 240.100 77.830 241.100 ;
        RECT 71.630 238.900 72.630 239.900 ;
        RECT 72.780 238.900 73.780 239.900 ;
        RECT 73.930 238.900 75.530 239.900 ;
        RECT 75.680 238.900 76.680 239.900 ;
        RECT 76.830 238.900 77.830 239.900 ;
        RECT 91.630 240.100 92.630 241.100 ;
        RECT 92.730 240.100 93.730 241.100 ;
        RECT 93.880 240.100 95.480 241.100 ;
        RECT 95.680 240.100 96.680 241.100 ;
        RECT 96.830 240.100 97.830 241.100 ;
        RECT 91.630 238.900 92.630 239.900 ;
        RECT 92.780 238.900 93.780 239.900 ;
        RECT 93.930 238.900 95.530 239.900 ;
        RECT 95.680 238.900 96.680 239.900 ;
        RECT 96.830 238.900 97.830 239.900 ;
        RECT 111.630 240.100 112.630 241.100 ;
        RECT 112.730 240.100 113.730 241.100 ;
        RECT 113.880 240.100 115.480 241.100 ;
        RECT 115.680 240.100 116.680 241.100 ;
        RECT 116.830 240.100 117.830 241.100 ;
        RECT 111.630 238.900 112.630 239.900 ;
        RECT 112.780 238.900 113.780 239.900 ;
        RECT 113.930 238.900 115.530 239.900 ;
        RECT 115.680 238.900 116.680 239.900 ;
        RECT 116.830 238.900 117.830 239.900 ;
        RECT 4.830 232.400 5.530 233.100 ;
        RECT 4.830 231.550 5.530 232.250 ;
        RECT 4.830 230.700 5.530 231.400 ;
        RECT 23.930 232.400 24.630 233.100 ;
        RECT 24.830 232.400 25.530 233.100 ;
        RECT 23.930 231.550 24.630 232.250 ;
        RECT 24.830 231.550 25.530 232.250 ;
        RECT 23.930 230.700 24.630 231.400 ;
        RECT 24.830 230.700 25.530 231.400 ;
        RECT 4.830 228.600 5.530 229.300 ;
        RECT 4.830 227.750 5.530 228.450 ;
        RECT 4.830 226.900 5.530 227.600 ;
        RECT 43.930 232.400 44.630 233.100 ;
        RECT 44.830 232.400 45.530 233.100 ;
        RECT 43.930 231.550 44.630 232.250 ;
        RECT 44.830 231.550 45.530 232.250 ;
        RECT 43.930 230.700 44.630 231.400 ;
        RECT 44.830 230.700 45.530 231.400 ;
        RECT 23.930 228.600 24.630 229.300 ;
        RECT 24.830 228.600 25.530 229.300 ;
        RECT 23.930 227.750 24.630 228.450 ;
        RECT 24.830 227.750 25.530 228.450 ;
        RECT 23.930 226.900 24.630 227.600 ;
        RECT 24.830 226.900 25.530 227.600 ;
        RECT 63.930 232.400 64.630 233.100 ;
        RECT 64.830 232.400 65.530 233.100 ;
        RECT 63.930 231.550 64.630 232.250 ;
        RECT 64.830 231.550 65.530 232.250 ;
        RECT 63.930 230.700 64.630 231.400 ;
        RECT 64.830 230.700 65.530 231.400 ;
        RECT 43.930 228.600 44.630 229.300 ;
        RECT 44.830 228.600 45.530 229.300 ;
        RECT 43.930 227.750 44.630 228.450 ;
        RECT 44.830 227.750 45.530 228.450 ;
        RECT 43.930 226.900 44.630 227.600 ;
        RECT 44.830 226.900 45.530 227.600 ;
        RECT 83.930 232.400 84.630 233.100 ;
        RECT 84.830 232.400 85.530 233.100 ;
        RECT 83.930 231.550 84.630 232.250 ;
        RECT 84.830 231.550 85.530 232.250 ;
        RECT 83.930 230.700 84.630 231.400 ;
        RECT 84.830 230.700 85.530 231.400 ;
        RECT 63.930 228.600 64.630 229.300 ;
        RECT 64.830 228.600 65.530 229.300 ;
        RECT 63.930 227.750 64.630 228.450 ;
        RECT 64.830 227.750 65.530 228.450 ;
        RECT 63.930 226.900 64.630 227.600 ;
        RECT 64.830 226.900 65.530 227.600 ;
        RECT 103.930 232.400 104.630 233.100 ;
        RECT 104.830 232.400 105.530 233.100 ;
        RECT 103.930 231.550 104.630 232.250 ;
        RECT 104.830 231.550 105.530 232.250 ;
        RECT 103.930 230.700 104.630 231.400 ;
        RECT 104.830 230.700 105.530 231.400 ;
        RECT 83.930 228.600 84.630 229.300 ;
        RECT 84.830 228.600 85.530 229.300 ;
        RECT 83.930 227.750 84.630 228.450 ;
        RECT 84.830 227.750 85.530 228.450 ;
        RECT 83.930 226.900 84.630 227.600 ;
        RECT 84.830 226.900 85.530 227.600 ;
        RECT 123.930 232.400 124.630 233.100 ;
        RECT 123.930 231.550 124.630 232.250 ;
        RECT 123.930 230.700 124.630 231.400 ;
        RECT 103.930 228.600 104.630 229.300 ;
        RECT 104.830 228.600 105.530 229.300 ;
        RECT 103.930 227.750 104.630 228.450 ;
        RECT 104.830 227.750 105.530 228.450 ;
        RECT 103.930 226.900 104.630 227.600 ;
        RECT 104.830 226.900 105.530 227.600 ;
        RECT 130.050 230.410 130.410 230.790 ;
        RECT 130.680 230.410 131.040 230.790 ;
        RECT 131.280 230.410 131.640 230.790 ;
        RECT 130.050 229.820 130.410 230.200 ;
        RECT 130.680 229.820 131.040 230.200 ;
        RECT 131.280 229.820 131.640 230.200 ;
        RECT 123.930 228.600 124.630 229.300 ;
        RECT 123.930 227.750 124.630 228.450 ;
        RECT 123.930 226.900 124.630 227.600 ;
        RECT 11.630 220.100 12.630 221.100 ;
        RECT 12.730 220.100 13.730 221.100 ;
        RECT 13.880 220.100 15.480 221.100 ;
        RECT 15.680 220.100 16.680 221.100 ;
        RECT 16.830 220.100 17.830 221.100 ;
        RECT 11.630 218.900 12.630 219.900 ;
        RECT 12.780 218.900 13.780 219.900 ;
        RECT 13.930 218.900 15.530 219.900 ;
        RECT 15.680 218.900 16.680 219.900 ;
        RECT 16.830 218.900 17.830 219.900 ;
        RECT 31.630 220.100 32.630 221.100 ;
        RECT 32.730 220.100 33.730 221.100 ;
        RECT 33.880 220.100 35.480 221.100 ;
        RECT 35.680 220.100 36.680 221.100 ;
        RECT 36.830 220.100 37.830 221.100 ;
        RECT 31.630 218.900 32.630 219.900 ;
        RECT 32.780 218.900 33.780 219.900 ;
        RECT 33.930 218.900 35.530 219.900 ;
        RECT 35.680 218.900 36.680 219.900 ;
        RECT 36.830 218.900 37.830 219.900 ;
        RECT 51.630 220.100 52.630 221.100 ;
        RECT 52.730 220.100 53.730 221.100 ;
        RECT 53.880 220.100 55.480 221.100 ;
        RECT 55.680 220.100 56.680 221.100 ;
        RECT 56.830 220.100 57.830 221.100 ;
        RECT 51.630 218.900 52.630 219.900 ;
        RECT 52.780 218.900 53.780 219.900 ;
        RECT 53.930 218.900 55.530 219.900 ;
        RECT 55.680 218.900 56.680 219.900 ;
        RECT 56.830 218.900 57.830 219.900 ;
        RECT 71.630 220.100 72.630 221.100 ;
        RECT 72.730 220.100 73.730 221.100 ;
        RECT 73.880 220.100 75.480 221.100 ;
        RECT 75.680 220.100 76.680 221.100 ;
        RECT 76.830 220.100 77.830 221.100 ;
        RECT 71.630 218.900 72.630 219.900 ;
        RECT 72.780 218.900 73.780 219.900 ;
        RECT 73.930 218.900 75.530 219.900 ;
        RECT 75.680 218.900 76.680 219.900 ;
        RECT 76.830 218.900 77.830 219.900 ;
        RECT 91.630 220.100 92.630 221.100 ;
        RECT 92.730 220.100 93.730 221.100 ;
        RECT 93.880 220.100 95.480 221.100 ;
        RECT 95.680 220.100 96.680 221.100 ;
        RECT 96.830 220.100 97.830 221.100 ;
        RECT 91.630 218.900 92.630 219.900 ;
        RECT 92.780 218.900 93.780 219.900 ;
        RECT 93.930 218.900 95.530 219.900 ;
        RECT 95.680 218.900 96.680 219.900 ;
        RECT 96.830 218.900 97.830 219.900 ;
        RECT 111.630 220.100 112.630 221.100 ;
        RECT 112.730 220.100 113.730 221.100 ;
        RECT 113.880 220.100 115.480 221.100 ;
        RECT 115.680 220.100 116.680 221.100 ;
        RECT 116.830 220.100 117.830 221.100 ;
        RECT 111.630 218.900 112.630 219.900 ;
        RECT 112.780 218.900 113.780 219.900 ;
        RECT 113.930 218.900 115.530 219.900 ;
        RECT 115.680 218.900 116.680 219.900 ;
        RECT 116.830 218.900 117.830 219.900 ;
        RECT 4.830 212.400 5.530 213.100 ;
        RECT 4.830 211.550 5.530 212.250 ;
        RECT 4.830 210.700 5.530 211.400 ;
        RECT 23.930 212.400 24.630 213.100 ;
        RECT 24.830 212.400 25.530 213.100 ;
        RECT 23.930 211.550 24.630 212.250 ;
        RECT 24.830 211.550 25.530 212.250 ;
        RECT 23.930 210.700 24.630 211.400 ;
        RECT 24.830 210.700 25.530 211.400 ;
        RECT 4.830 208.600 5.530 209.300 ;
        RECT 4.830 207.750 5.530 208.450 ;
        RECT 4.830 206.900 5.530 207.600 ;
        RECT 43.930 212.400 44.630 213.100 ;
        RECT 44.830 212.400 45.530 213.100 ;
        RECT 43.930 211.550 44.630 212.250 ;
        RECT 44.830 211.550 45.530 212.250 ;
        RECT 43.930 210.700 44.630 211.400 ;
        RECT 44.830 210.700 45.530 211.400 ;
        RECT 23.930 208.600 24.630 209.300 ;
        RECT 24.830 208.600 25.530 209.300 ;
        RECT 23.930 207.750 24.630 208.450 ;
        RECT 24.830 207.750 25.530 208.450 ;
        RECT 23.930 206.900 24.630 207.600 ;
        RECT 24.830 206.900 25.530 207.600 ;
        RECT 63.930 212.400 64.630 213.100 ;
        RECT 64.830 212.400 65.530 213.100 ;
        RECT 63.930 211.550 64.630 212.250 ;
        RECT 64.830 211.550 65.530 212.250 ;
        RECT 63.930 210.700 64.630 211.400 ;
        RECT 64.830 210.700 65.530 211.400 ;
        RECT 43.930 208.600 44.630 209.300 ;
        RECT 44.830 208.600 45.530 209.300 ;
        RECT 43.930 207.750 44.630 208.450 ;
        RECT 44.830 207.750 45.530 208.450 ;
        RECT 43.930 206.900 44.630 207.600 ;
        RECT 44.830 206.900 45.530 207.600 ;
        RECT 83.930 212.400 84.630 213.100 ;
        RECT 84.830 212.400 85.530 213.100 ;
        RECT 83.930 211.550 84.630 212.250 ;
        RECT 84.830 211.550 85.530 212.250 ;
        RECT 83.930 210.700 84.630 211.400 ;
        RECT 84.830 210.700 85.530 211.400 ;
        RECT 63.930 208.600 64.630 209.300 ;
        RECT 64.830 208.600 65.530 209.300 ;
        RECT 63.930 207.750 64.630 208.450 ;
        RECT 64.830 207.750 65.530 208.450 ;
        RECT 63.930 206.900 64.630 207.600 ;
        RECT 64.830 206.900 65.530 207.600 ;
        RECT 103.930 212.400 104.630 213.100 ;
        RECT 104.830 212.400 105.530 213.100 ;
        RECT 103.930 211.550 104.630 212.250 ;
        RECT 104.830 211.550 105.530 212.250 ;
        RECT 103.930 210.700 104.630 211.400 ;
        RECT 104.830 210.700 105.530 211.400 ;
        RECT 83.930 208.600 84.630 209.300 ;
        RECT 84.830 208.600 85.530 209.300 ;
        RECT 83.930 207.750 84.630 208.450 ;
        RECT 84.830 207.750 85.530 208.450 ;
        RECT 83.930 206.900 84.630 207.600 ;
        RECT 84.830 206.900 85.530 207.600 ;
        RECT 123.930 212.400 124.630 213.100 ;
        RECT 123.930 211.550 124.630 212.250 ;
        RECT 123.930 210.700 124.630 211.400 ;
        RECT 103.930 208.600 104.630 209.300 ;
        RECT 104.830 208.600 105.530 209.300 ;
        RECT 103.930 207.750 104.630 208.450 ;
        RECT 104.830 207.750 105.530 208.450 ;
        RECT 103.930 206.900 104.630 207.600 ;
        RECT 104.830 206.900 105.530 207.600 ;
        RECT 123.930 208.600 124.630 209.300 ;
        RECT 130.050 209.120 130.410 209.500 ;
        RECT 130.680 209.120 131.040 209.500 ;
        RECT 131.280 209.120 131.640 209.500 ;
        RECT 130.050 208.530 130.410 208.910 ;
        RECT 130.680 208.530 131.040 208.910 ;
        RECT 131.280 208.530 131.640 208.910 ;
        RECT 123.930 207.750 124.630 208.450 ;
        RECT 123.930 206.900 124.630 207.600 ;
        RECT 11.630 200.100 12.630 201.100 ;
        RECT 12.730 200.100 13.730 201.100 ;
        RECT 13.880 200.100 15.480 201.100 ;
        RECT 15.680 200.100 16.680 201.100 ;
        RECT 16.830 200.100 17.830 201.100 ;
        RECT 31.630 200.100 32.630 201.100 ;
        RECT 32.730 200.100 33.730 201.100 ;
        RECT 33.880 200.100 35.480 201.100 ;
        RECT 35.680 200.100 36.680 201.100 ;
        RECT 36.830 200.100 37.830 201.100 ;
        RECT 51.630 200.100 52.630 201.100 ;
        RECT 52.730 200.100 53.730 201.100 ;
        RECT 53.880 200.100 55.480 201.100 ;
        RECT 55.680 200.100 56.680 201.100 ;
        RECT 56.830 200.100 57.830 201.100 ;
        RECT 71.630 200.100 72.630 201.100 ;
        RECT 72.730 200.100 73.730 201.100 ;
        RECT 73.880 200.100 75.480 201.100 ;
        RECT 75.680 200.100 76.680 201.100 ;
        RECT 76.830 200.100 77.830 201.100 ;
        RECT 91.630 200.100 92.630 201.100 ;
        RECT 92.730 200.100 93.730 201.100 ;
        RECT 93.880 200.100 95.480 201.100 ;
        RECT 95.680 200.100 96.680 201.100 ;
        RECT 96.830 200.100 97.830 201.100 ;
        RECT 111.630 200.100 112.630 201.100 ;
        RECT 112.730 200.100 113.730 201.100 ;
        RECT 113.880 200.100 115.480 201.100 ;
        RECT 115.680 200.100 116.680 201.100 ;
        RECT 116.830 200.100 117.830 201.100 ;
        RECT 9.425 176.405 10.015 176.975 ;
        RECT 10.205 176.405 10.795 176.975 ;
        RECT 10.985 176.405 11.575 176.975 ;
        RECT 11.630 138.900 12.630 139.900 ;
        RECT 12.780 138.900 13.780 139.900 ;
        RECT 13.930 138.900 15.530 139.900 ;
        RECT 15.680 138.900 16.680 139.900 ;
        RECT 16.830 138.900 17.830 139.900 ;
        RECT 31.630 138.900 32.630 139.900 ;
        RECT 32.780 138.900 33.780 139.900 ;
        RECT 33.930 138.900 35.530 139.900 ;
        RECT 35.680 138.900 36.680 139.900 ;
        RECT 36.830 138.900 37.830 139.900 ;
        RECT 51.630 138.900 52.630 139.900 ;
        RECT 52.780 138.900 53.780 139.900 ;
        RECT 53.930 138.900 55.530 139.900 ;
        RECT 55.680 138.900 56.680 139.900 ;
        RECT 56.830 138.900 57.830 139.900 ;
        RECT 71.630 138.900 72.630 139.900 ;
        RECT 72.780 138.900 73.780 139.900 ;
        RECT 73.930 138.900 75.530 139.900 ;
        RECT 75.680 138.900 76.680 139.900 ;
        RECT 76.830 138.900 77.830 139.900 ;
        RECT 91.630 138.900 92.630 139.900 ;
        RECT 92.780 138.900 93.780 139.900 ;
        RECT 93.930 138.900 95.530 139.900 ;
        RECT 95.680 138.900 96.680 139.900 ;
        RECT 96.830 138.900 97.830 139.900 ;
        RECT 111.630 138.900 112.630 139.900 ;
        RECT 112.780 138.900 113.780 139.900 ;
        RECT 113.930 138.900 115.530 139.900 ;
        RECT 115.680 138.900 116.680 139.900 ;
        RECT 116.830 138.900 117.830 139.900 ;
        RECT 4.830 132.400 5.530 133.100 ;
        RECT 4.830 131.550 5.530 132.250 ;
        RECT 4.830 130.700 5.530 131.400 ;
        RECT 23.930 132.400 24.630 133.100 ;
        RECT 24.830 132.400 25.530 133.100 ;
        RECT 23.930 131.550 24.630 132.250 ;
        RECT 24.830 131.550 25.530 132.250 ;
        RECT 23.930 130.700 24.630 131.400 ;
        RECT 24.830 130.700 25.530 131.400 ;
        RECT 4.830 128.600 5.530 129.300 ;
        RECT 4.830 127.750 5.530 128.450 ;
        RECT 4.830 126.900 5.530 127.600 ;
        RECT 43.930 132.400 44.630 133.100 ;
        RECT 44.830 132.400 45.530 133.100 ;
        RECT 43.930 131.550 44.630 132.250 ;
        RECT 44.830 131.550 45.530 132.250 ;
        RECT 43.930 130.700 44.630 131.400 ;
        RECT 44.830 130.700 45.530 131.400 ;
        RECT 23.930 128.600 24.630 129.300 ;
        RECT 24.830 128.600 25.530 129.300 ;
        RECT 23.930 127.750 24.630 128.450 ;
        RECT 24.830 127.750 25.530 128.450 ;
        RECT 23.930 126.900 24.630 127.600 ;
        RECT 24.830 126.900 25.530 127.600 ;
        RECT 63.930 132.400 64.630 133.100 ;
        RECT 64.830 132.400 65.530 133.100 ;
        RECT 63.930 131.550 64.630 132.250 ;
        RECT 64.830 131.550 65.530 132.250 ;
        RECT 63.930 130.700 64.630 131.400 ;
        RECT 64.830 130.700 65.530 131.400 ;
        RECT 43.930 128.600 44.630 129.300 ;
        RECT 44.830 128.600 45.530 129.300 ;
        RECT 43.930 127.750 44.630 128.450 ;
        RECT 44.830 127.750 45.530 128.450 ;
        RECT 43.930 126.900 44.630 127.600 ;
        RECT 44.830 126.900 45.530 127.600 ;
        RECT 83.930 132.400 84.630 133.100 ;
        RECT 84.830 132.400 85.530 133.100 ;
        RECT 83.930 131.550 84.630 132.250 ;
        RECT 84.830 131.550 85.530 132.250 ;
        RECT 83.930 130.700 84.630 131.400 ;
        RECT 84.830 130.700 85.530 131.400 ;
        RECT 63.930 128.600 64.630 129.300 ;
        RECT 64.830 128.600 65.530 129.300 ;
        RECT 63.930 127.750 64.630 128.450 ;
        RECT 64.830 127.750 65.530 128.450 ;
        RECT 63.930 126.900 64.630 127.600 ;
        RECT 64.830 126.900 65.530 127.600 ;
        RECT 103.930 132.400 104.630 133.100 ;
        RECT 104.830 132.400 105.530 133.100 ;
        RECT 103.930 131.550 104.630 132.250 ;
        RECT 104.830 131.550 105.530 132.250 ;
        RECT 103.930 130.700 104.630 131.400 ;
        RECT 104.830 130.700 105.530 131.400 ;
        RECT 83.930 128.600 84.630 129.300 ;
        RECT 84.830 128.600 85.530 129.300 ;
        RECT 83.930 127.750 84.630 128.450 ;
        RECT 84.830 127.750 85.530 128.450 ;
        RECT 83.930 126.900 84.630 127.600 ;
        RECT 84.830 126.900 85.530 127.600 ;
        RECT 123.930 132.400 124.630 133.100 ;
        RECT 123.930 131.550 124.630 132.250 ;
        RECT 123.930 130.700 124.630 131.400 ;
        RECT 103.930 128.600 104.630 129.300 ;
        RECT 104.830 128.600 105.530 129.300 ;
        RECT 103.930 127.750 104.630 128.450 ;
        RECT 104.830 127.750 105.530 128.450 ;
        RECT 103.930 126.900 104.630 127.600 ;
        RECT 104.830 126.900 105.530 127.600 ;
        RECT 130.050 130.270 130.410 130.650 ;
        RECT 130.680 130.270 131.040 130.650 ;
        RECT 131.280 130.270 131.640 130.650 ;
        RECT 130.050 129.680 130.410 130.060 ;
        RECT 130.680 129.680 131.040 130.060 ;
        RECT 131.280 129.680 131.640 130.060 ;
        RECT 123.930 128.600 124.630 129.300 ;
        RECT 123.930 127.750 124.630 128.450 ;
        RECT 123.930 126.900 124.630 127.600 ;
        RECT 11.630 120.100 12.630 121.100 ;
        RECT 12.730 120.100 13.730 121.100 ;
        RECT 13.880 120.100 15.480 121.100 ;
        RECT 15.680 120.100 16.680 121.100 ;
        RECT 16.830 120.100 17.830 121.100 ;
        RECT 11.630 118.900 12.630 119.900 ;
        RECT 12.780 118.900 13.780 119.900 ;
        RECT 13.930 118.900 15.530 119.900 ;
        RECT 15.680 118.900 16.680 119.900 ;
        RECT 16.830 118.900 17.830 119.900 ;
        RECT 31.630 120.100 32.630 121.100 ;
        RECT 32.730 120.100 33.730 121.100 ;
        RECT 33.880 120.100 35.480 121.100 ;
        RECT 35.680 120.100 36.680 121.100 ;
        RECT 36.830 120.100 37.830 121.100 ;
        RECT 31.630 118.900 32.630 119.900 ;
        RECT 32.780 118.900 33.780 119.900 ;
        RECT 33.930 118.900 35.530 119.900 ;
        RECT 35.680 118.900 36.680 119.900 ;
        RECT 36.830 118.900 37.830 119.900 ;
        RECT 51.630 120.100 52.630 121.100 ;
        RECT 52.730 120.100 53.730 121.100 ;
        RECT 53.880 120.100 55.480 121.100 ;
        RECT 55.680 120.100 56.680 121.100 ;
        RECT 56.830 120.100 57.830 121.100 ;
        RECT 51.630 118.900 52.630 119.900 ;
        RECT 52.780 118.900 53.780 119.900 ;
        RECT 53.930 118.900 55.530 119.900 ;
        RECT 55.680 118.900 56.680 119.900 ;
        RECT 56.830 118.900 57.830 119.900 ;
        RECT 71.630 120.100 72.630 121.100 ;
        RECT 72.730 120.100 73.730 121.100 ;
        RECT 73.880 120.100 75.480 121.100 ;
        RECT 75.680 120.100 76.680 121.100 ;
        RECT 76.830 120.100 77.830 121.100 ;
        RECT 71.630 118.900 72.630 119.900 ;
        RECT 72.780 118.900 73.780 119.900 ;
        RECT 73.930 118.900 75.530 119.900 ;
        RECT 75.680 118.900 76.680 119.900 ;
        RECT 76.830 118.900 77.830 119.900 ;
        RECT 91.630 120.100 92.630 121.100 ;
        RECT 92.730 120.100 93.730 121.100 ;
        RECT 93.880 120.100 95.480 121.100 ;
        RECT 95.680 120.100 96.680 121.100 ;
        RECT 96.830 120.100 97.830 121.100 ;
        RECT 91.630 118.900 92.630 119.900 ;
        RECT 92.780 118.900 93.780 119.900 ;
        RECT 93.930 118.900 95.530 119.900 ;
        RECT 95.680 118.900 96.680 119.900 ;
        RECT 96.830 118.900 97.830 119.900 ;
        RECT 111.630 120.100 112.630 121.100 ;
        RECT 112.730 120.100 113.730 121.100 ;
        RECT 113.880 120.100 115.480 121.100 ;
        RECT 115.680 120.100 116.680 121.100 ;
        RECT 116.830 120.100 117.830 121.100 ;
        RECT 111.630 118.900 112.630 119.900 ;
        RECT 112.780 118.900 113.780 119.900 ;
        RECT 113.930 118.900 115.530 119.900 ;
        RECT 115.680 118.900 116.680 119.900 ;
        RECT 116.830 118.900 117.830 119.900 ;
        RECT 4.830 112.400 5.530 113.100 ;
        RECT 4.830 111.550 5.530 112.250 ;
        RECT 4.830 110.700 5.530 111.400 ;
        RECT 23.930 112.400 24.630 113.100 ;
        RECT 24.830 112.400 25.530 113.100 ;
        RECT 23.930 111.550 24.630 112.250 ;
        RECT 24.830 111.550 25.530 112.250 ;
        RECT 23.930 110.700 24.630 111.400 ;
        RECT 24.830 110.700 25.530 111.400 ;
        RECT 4.830 108.600 5.530 109.300 ;
        RECT 4.830 107.750 5.530 108.450 ;
        RECT 4.830 106.900 5.530 107.600 ;
        RECT 43.930 112.400 44.630 113.100 ;
        RECT 44.830 112.400 45.530 113.100 ;
        RECT 43.930 111.550 44.630 112.250 ;
        RECT 44.830 111.550 45.530 112.250 ;
        RECT 43.930 110.700 44.630 111.400 ;
        RECT 44.830 110.700 45.530 111.400 ;
        RECT 23.930 108.600 24.630 109.300 ;
        RECT 24.830 108.600 25.530 109.300 ;
        RECT 23.930 107.750 24.630 108.450 ;
        RECT 24.830 107.750 25.530 108.450 ;
        RECT 23.930 106.900 24.630 107.600 ;
        RECT 24.830 106.900 25.530 107.600 ;
        RECT 63.930 112.400 64.630 113.100 ;
        RECT 64.830 112.400 65.530 113.100 ;
        RECT 63.930 111.550 64.630 112.250 ;
        RECT 64.830 111.550 65.530 112.250 ;
        RECT 63.930 110.700 64.630 111.400 ;
        RECT 64.830 110.700 65.530 111.400 ;
        RECT 43.930 108.600 44.630 109.300 ;
        RECT 44.830 108.600 45.530 109.300 ;
        RECT 43.930 107.750 44.630 108.450 ;
        RECT 44.830 107.750 45.530 108.450 ;
        RECT 43.930 106.900 44.630 107.600 ;
        RECT 44.830 106.900 45.530 107.600 ;
        RECT 83.930 112.400 84.630 113.100 ;
        RECT 84.830 112.400 85.530 113.100 ;
        RECT 83.930 111.550 84.630 112.250 ;
        RECT 84.830 111.550 85.530 112.250 ;
        RECT 83.930 110.700 84.630 111.400 ;
        RECT 84.830 110.700 85.530 111.400 ;
        RECT 63.930 108.600 64.630 109.300 ;
        RECT 64.830 108.600 65.530 109.300 ;
        RECT 63.930 107.750 64.630 108.450 ;
        RECT 64.830 107.750 65.530 108.450 ;
        RECT 63.930 106.900 64.630 107.600 ;
        RECT 64.830 106.900 65.530 107.600 ;
        RECT 103.930 112.400 104.630 113.100 ;
        RECT 104.830 112.400 105.530 113.100 ;
        RECT 103.930 111.550 104.630 112.250 ;
        RECT 104.830 111.550 105.530 112.250 ;
        RECT 103.930 110.700 104.630 111.400 ;
        RECT 104.830 110.700 105.530 111.400 ;
        RECT 83.930 108.600 84.630 109.300 ;
        RECT 84.830 108.600 85.530 109.300 ;
        RECT 83.930 107.750 84.630 108.450 ;
        RECT 84.830 107.750 85.530 108.450 ;
        RECT 83.930 106.900 84.630 107.600 ;
        RECT 84.830 106.900 85.530 107.600 ;
        RECT 123.930 112.400 124.630 113.100 ;
        RECT 123.930 111.550 124.630 112.250 ;
        RECT 123.930 110.700 124.630 111.400 ;
        RECT 103.930 108.600 104.630 109.300 ;
        RECT 104.830 108.600 105.530 109.300 ;
        RECT 103.930 107.750 104.630 108.450 ;
        RECT 104.830 107.750 105.530 108.450 ;
        RECT 103.930 106.900 104.630 107.600 ;
        RECT 104.830 106.900 105.530 107.600 ;
        RECT 130.050 109.475 130.410 109.855 ;
        RECT 130.680 109.475 131.040 109.855 ;
        RECT 131.280 109.475 131.640 109.855 ;
        RECT 123.930 108.600 124.630 109.300 ;
        RECT 130.050 108.885 130.410 109.265 ;
        RECT 130.680 108.885 131.040 109.265 ;
        RECT 131.280 108.885 131.640 109.265 ;
        RECT 123.930 107.750 124.630 108.450 ;
        RECT 123.930 106.900 124.630 107.600 ;
        RECT 11.630 100.100 12.630 101.100 ;
        RECT 12.730 100.100 13.730 101.100 ;
        RECT 13.880 100.100 15.480 101.100 ;
        RECT 15.680 100.100 16.680 101.100 ;
        RECT 16.830 100.100 17.830 101.100 ;
        RECT 11.630 98.900 12.630 99.900 ;
        RECT 12.780 98.900 13.780 99.900 ;
        RECT 13.930 98.900 15.530 99.900 ;
        RECT 15.680 98.900 16.680 99.900 ;
        RECT 16.830 98.900 17.830 99.900 ;
        RECT 31.630 100.100 32.630 101.100 ;
        RECT 32.730 100.100 33.730 101.100 ;
        RECT 33.880 100.100 35.480 101.100 ;
        RECT 35.680 100.100 36.680 101.100 ;
        RECT 36.830 100.100 37.830 101.100 ;
        RECT 31.630 98.900 32.630 99.900 ;
        RECT 32.780 98.900 33.780 99.900 ;
        RECT 33.930 98.900 35.530 99.900 ;
        RECT 35.680 98.900 36.680 99.900 ;
        RECT 36.830 98.900 37.830 99.900 ;
        RECT 51.630 100.100 52.630 101.100 ;
        RECT 52.730 100.100 53.730 101.100 ;
        RECT 53.880 100.100 55.480 101.100 ;
        RECT 55.680 100.100 56.680 101.100 ;
        RECT 56.830 100.100 57.830 101.100 ;
        RECT 51.630 98.900 52.630 99.900 ;
        RECT 52.780 98.900 53.780 99.900 ;
        RECT 53.930 98.900 55.530 99.900 ;
        RECT 55.680 98.900 56.680 99.900 ;
        RECT 56.830 98.900 57.830 99.900 ;
        RECT 71.630 100.100 72.630 101.100 ;
        RECT 72.730 100.100 73.730 101.100 ;
        RECT 73.880 100.100 75.480 101.100 ;
        RECT 75.680 100.100 76.680 101.100 ;
        RECT 76.830 100.100 77.830 101.100 ;
        RECT 71.630 98.900 72.630 99.900 ;
        RECT 72.780 98.900 73.780 99.900 ;
        RECT 73.930 98.900 75.530 99.900 ;
        RECT 75.680 98.900 76.680 99.900 ;
        RECT 76.830 98.900 77.830 99.900 ;
        RECT 91.630 100.100 92.630 101.100 ;
        RECT 92.730 100.100 93.730 101.100 ;
        RECT 93.880 100.100 95.480 101.100 ;
        RECT 95.680 100.100 96.680 101.100 ;
        RECT 96.830 100.100 97.830 101.100 ;
        RECT 91.630 98.900 92.630 99.900 ;
        RECT 92.780 98.900 93.780 99.900 ;
        RECT 93.930 98.900 95.530 99.900 ;
        RECT 95.680 98.900 96.680 99.900 ;
        RECT 96.830 98.900 97.830 99.900 ;
        RECT 111.630 100.100 112.630 101.100 ;
        RECT 112.730 100.100 113.730 101.100 ;
        RECT 113.880 100.100 115.480 101.100 ;
        RECT 115.680 100.100 116.680 101.100 ;
        RECT 116.830 100.100 117.830 101.100 ;
        RECT 111.630 98.900 112.630 99.900 ;
        RECT 112.780 98.900 113.780 99.900 ;
        RECT 113.930 98.900 115.530 99.900 ;
        RECT 115.680 98.900 116.680 99.900 ;
        RECT 116.830 98.900 117.830 99.900 ;
        RECT 4.830 92.400 5.530 93.100 ;
        RECT 4.830 91.550 5.530 92.250 ;
        RECT 4.830 90.700 5.530 91.400 ;
        RECT 23.930 92.400 24.630 93.100 ;
        RECT 24.830 92.400 25.530 93.100 ;
        RECT 23.930 91.550 24.630 92.250 ;
        RECT 24.830 91.550 25.530 92.250 ;
        RECT 23.930 90.700 24.630 91.400 ;
        RECT 24.830 90.700 25.530 91.400 ;
        RECT 4.830 88.600 5.530 89.300 ;
        RECT 4.830 87.750 5.530 88.450 ;
        RECT 4.830 86.900 5.530 87.600 ;
        RECT 43.930 92.400 44.630 93.100 ;
        RECT 44.830 92.400 45.530 93.100 ;
        RECT 43.930 91.550 44.630 92.250 ;
        RECT 44.830 91.550 45.530 92.250 ;
        RECT 43.930 90.700 44.630 91.400 ;
        RECT 44.830 90.700 45.530 91.400 ;
        RECT 23.930 88.600 24.630 89.300 ;
        RECT 24.830 88.600 25.530 89.300 ;
        RECT 23.930 87.750 24.630 88.450 ;
        RECT 24.830 87.750 25.530 88.450 ;
        RECT 23.930 86.900 24.630 87.600 ;
        RECT 24.830 86.900 25.530 87.600 ;
        RECT 63.930 92.400 64.630 93.100 ;
        RECT 64.830 92.400 65.530 93.100 ;
        RECT 63.930 91.550 64.630 92.250 ;
        RECT 64.830 91.550 65.530 92.250 ;
        RECT 63.930 90.700 64.630 91.400 ;
        RECT 64.830 90.700 65.530 91.400 ;
        RECT 43.930 88.600 44.630 89.300 ;
        RECT 44.830 88.600 45.530 89.300 ;
        RECT 43.930 87.750 44.630 88.450 ;
        RECT 44.830 87.750 45.530 88.450 ;
        RECT 43.930 86.900 44.630 87.600 ;
        RECT 44.830 86.900 45.530 87.600 ;
        RECT 83.930 92.400 84.630 93.100 ;
        RECT 84.830 92.400 85.530 93.100 ;
        RECT 83.930 91.550 84.630 92.250 ;
        RECT 84.830 91.550 85.530 92.250 ;
        RECT 83.930 90.700 84.630 91.400 ;
        RECT 84.830 90.700 85.530 91.400 ;
        RECT 63.930 88.600 64.630 89.300 ;
        RECT 64.830 88.600 65.530 89.300 ;
        RECT 63.930 87.750 64.630 88.450 ;
        RECT 64.830 87.750 65.530 88.450 ;
        RECT 63.930 86.900 64.630 87.600 ;
        RECT 64.830 86.900 65.530 87.600 ;
        RECT 103.930 92.400 104.630 93.100 ;
        RECT 104.830 92.400 105.530 93.100 ;
        RECT 103.930 91.550 104.630 92.250 ;
        RECT 104.830 91.550 105.530 92.250 ;
        RECT 103.930 90.700 104.630 91.400 ;
        RECT 104.830 90.700 105.530 91.400 ;
        RECT 83.930 88.600 84.630 89.300 ;
        RECT 84.830 88.600 85.530 89.300 ;
        RECT 83.930 87.750 84.630 88.450 ;
        RECT 84.830 87.750 85.530 88.450 ;
        RECT 83.930 86.900 84.630 87.600 ;
        RECT 84.830 86.900 85.530 87.600 ;
        RECT 123.930 92.400 124.630 93.100 ;
        RECT 123.930 91.550 124.630 92.250 ;
        RECT 123.930 90.700 124.630 91.400 ;
        RECT 130.050 90.525 130.410 90.905 ;
        RECT 130.680 90.525 131.040 90.905 ;
        RECT 131.280 90.525 131.640 90.905 ;
        RECT 103.930 88.600 104.630 89.300 ;
        RECT 104.830 88.600 105.530 89.300 ;
        RECT 103.930 87.750 104.630 88.450 ;
        RECT 104.830 87.750 105.530 88.450 ;
        RECT 103.930 86.900 104.630 87.600 ;
        RECT 104.830 86.900 105.530 87.600 ;
        RECT 130.050 89.935 130.410 90.315 ;
        RECT 130.680 89.935 131.040 90.315 ;
        RECT 131.280 89.935 131.640 90.315 ;
        RECT 123.930 88.600 124.630 89.300 ;
        RECT 123.930 87.750 124.630 88.450 ;
        RECT 123.930 86.900 124.630 87.600 ;
        RECT 11.630 80.100 12.630 81.100 ;
        RECT 12.730 80.100 13.730 81.100 ;
        RECT 13.880 80.100 15.480 81.100 ;
        RECT 15.680 80.100 16.680 81.100 ;
        RECT 16.830 80.100 17.830 81.100 ;
        RECT 11.630 78.900 12.630 79.900 ;
        RECT 12.780 78.900 13.780 79.900 ;
        RECT 13.930 78.900 15.530 79.900 ;
        RECT 15.680 78.900 16.680 79.900 ;
        RECT 16.830 78.900 17.830 79.900 ;
        RECT 31.630 80.100 32.630 81.100 ;
        RECT 32.730 80.100 33.730 81.100 ;
        RECT 33.880 80.100 35.480 81.100 ;
        RECT 35.680 80.100 36.680 81.100 ;
        RECT 36.830 80.100 37.830 81.100 ;
        RECT 31.630 78.900 32.630 79.900 ;
        RECT 32.780 78.900 33.780 79.900 ;
        RECT 33.930 78.900 35.530 79.900 ;
        RECT 35.680 78.900 36.680 79.900 ;
        RECT 36.830 78.900 37.830 79.900 ;
        RECT 51.630 80.100 52.630 81.100 ;
        RECT 52.730 80.100 53.730 81.100 ;
        RECT 53.880 80.100 55.480 81.100 ;
        RECT 55.680 80.100 56.680 81.100 ;
        RECT 56.830 80.100 57.830 81.100 ;
        RECT 51.630 78.900 52.630 79.900 ;
        RECT 52.780 78.900 53.780 79.900 ;
        RECT 53.930 78.900 55.530 79.900 ;
        RECT 55.680 78.900 56.680 79.900 ;
        RECT 56.830 78.900 57.830 79.900 ;
        RECT 71.630 80.100 72.630 81.100 ;
        RECT 72.730 80.100 73.730 81.100 ;
        RECT 73.880 80.100 75.480 81.100 ;
        RECT 75.680 80.100 76.680 81.100 ;
        RECT 76.830 80.100 77.830 81.100 ;
        RECT 71.630 78.900 72.630 79.900 ;
        RECT 72.780 78.900 73.780 79.900 ;
        RECT 73.930 78.900 75.530 79.900 ;
        RECT 75.680 78.900 76.680 79.900 ;
        RECT 76.830 78.900 77.830 79.900 ;
        RECT 91.630 80.100 92.630 81.100 ;
        RECT 92.730 80.100 93.730 81.100 ;
        RECT 93.880 80.100 95.480 81.100 ;
        RECT 95.680 80.100 96.680 81.100 ;
        RECT 96.830 80.100 97.830 81.100 ;
        RECT 91.630 78.900 92.630 79.900 ;
        RECT 92.780 78.900 93.780 79.900 ;
        RECT 93.930 78.900 95.530 79.900 ;
        RECT 95.680 78.900 96.680 79.900 ;
        RECT 96.830 78.900 97.830 79.900 ;
        RECT 111.630 80.100 112.630 81.100 ;
        RECT 112.730 80.100 113.730 81.100 ;
        RECT 113.880 80.100 115.480 81.100 ;
        RECT 115.680 80.100 116.680 81.100 ;
        RECT 116.830 80.100 117.830 81.100 ;
        RECT 111.630 78.900 112.630 79.900 ;
        RECT 112.780 78.900 113.780 79.900 ;
        RECT 113.930 78.900 115.530 79.900 ;
        RECT 115.680 78.900 116.680 79.900 ;
        RECT 116.830 78.900 117.830 79.900 ;
        RECT 4.830 72.400 5.530 73.100 ;
        RECT 4.830 71.550 5.530 72.250 ;
        RECT 4.830 70.700 5.530 71.400 ;
        RECT 23.930 72.400 24.630 73.100 ;
        RECT 24.830 72.400 25.530 73.100 ;
        RECT 23.930 71.550 24.630 72.250 ;
        RECT 24.830 71.550 25.530 72.250 ;
        RECT 23.930 70.700 24.630 71.400 ;
        RECT 24.830 70.700 25.530 71.400 ;
        RECT 4.830 68.600 5.530 69.300 ;
        RECT 4.830 67.750 5.530 68.450 ;
        RECT 4.830 66.900 5.530 67.600 ;
        RECT 43.930 72.400 44.630 73.100 ;
        RECT 44.830 72.400 45.530 73.100 ;
        RECT 43.930 71.550 44.630 72.250 ;
        RECT 44.830 71.550 45.530 72.250 ;
        RECT 43.930 70.700 44.630 71.400 ;
        RECT 44.830 70.700 45.530 71.400 ;
        RECT 23.930 68.600 24.630 69.300 ;
        RECT 24.830 68.600 25.530 69.300 ;
        RECT 23.930 67.750 24.630 68.450 ;
        RECT 24.830 67.750 25.530 68.450 ;
        RECT 23.930 66.900 24.630 67.600 ;
        RECT 24.830 66.900 25.530 67.600 ;
        RECT 63.930 72.400 64.630 73.100 ;
        RECT 64.830 72.400 65.530 73.100 ;
        RECT 63.930 71.550 64.630 72.250 ;
        RECT 64.830 71.550 65.530 72.250 ;
        RECT 63.930 70.700 64.630 71.400 ;
        RECT 64.830 70.700 65.530 71.400 ;
        RECT 43.930 68.600 44.630 69.300 ;
        RECT 44.830 68.600 45.530 69.300 ;
        RECT 43.930 67.750 44.630 68.450 ;
        RECT 44.830 67.750 45.530 68.450 ;
        RECT 43.930 66.900 44.630 67.600 ;
        RECT 44.830 66.900 45.530 67.600 ;
        RECT 83.930 72.400 84.630 73.100 ;
        RECT 84.830 72.400 85.530 73.100 ;
        RECT 83.930 71.550 84.630 72.250 ;
        RECT 84.830 71.550 85.530 72.250 ;
        RECT 83.930 70.700 84.630 71.400 ;
        RECT 84.830 70.700 85.530 71.400 ;
        RECT 63.930 68.600 64.630 69.300 ;
        RECT 64.830 68.600 65.530 69.300 ;
        RECT 63.930 67.750 64.630 68.450 ;
        RECT 64.830 67.750 65.530 68.450 ;
        RECT 63.930 66.900 64.630 67.600 ;
        RECT 64.830 66.900 65.530 67.600 ;
        RECT 103.930 72.400 104.630 73.100 ;
        RECT 104.830 72.400 105.530 73.100 ;
        RECT 103.930 71.550 104.630 72.250 ;
        RECT 104.830 71.550 105.530 72.250 ;
        RECT 103.930 70.700 104.630 71.400 ;
        RECT 104.830 70.700 105.530 71.400 ;
        RECT 83.930 68.600 84.630 69.300 ;
        RECT 84.830 68.600 85.530 69.300 ;
        RECT 83.930 67.750 84.630 68.450 ;
        RECT 84.830 67.750 85.530 68.450 ;
        RECT 83.930 66.900 84.630 67.600 ;
        RECT 84.830 66.900 85.530 67.600 ;
        RECT 123.930 72.400 124.630 73.100 ;
        RECT 123.930 71.550 124.630 72.250 ;
        RECT 123.930 70.700 124.630 71.400 ;
        RECT 103.930 68.600 104.630 69.300 ;
        RECT 104.830 68.600 105.530 69.300 ;
        RECT 103.930 67.750 104.630 68.450 ;
        RECT 104.830 67.750 105.530 68.450 ;
        RECT 103.930 66.900 104.630 67.600 ;
        RECT 104.830 66.900 105.530 67.600 ;
        RECT 130.050 69.990 130.410 70.370 ;
        RECT 130.680 69.990 131.040 70.370 ;
        RECT 131.280 69.990 131.640 70.370 ;
        RECT 130.050 69.400 130.410 69.780 ;
        RECT 130.680 69.400 131.040 69.780 ;
        RECT 131.280 69.400 131.640 69.780 ;
        RECT 123.930 68.600 124.630 69.300 ;
        RECT 123.930 67.750 124.630 68.450 ;
        RECT 123.930 66.900 124.630 67.600 ;
        RECT 11.630 60.100 12.630 61.100 ;
        RECT 12.730 60.100 13.730 61.100 ;
        RECT 13.880 60.100 15.480 61.100 ;
        RECT 15.680 60.100 16.680 61.100 ;
        RECT 16.830 60.100 17.830 61.100 ;
        RECT 11.630 58.900 12.630 59.900 ;
        RECT 12.780 58.900 13.780 59.900 ;
        RECT 13.930 58.900 15.530 59.900 ;
        RECT 15.680 58.900 16.680 59.900 ;
        RECT 16.830 58.900 17.830 59.900 ;
        RECT 31.630 60.100 32.630 61.100 ;
        RECT 32.730 60.100 33.730 61.100 ;
        RECT 33.880 60.100 35.480 61.100 ;
        RECT 35.680 60.100 36.680 61.100 ;
        RECT 36.830 60.100 37.830 61.100 ;
        RECT 31.630 58.900 32.630 59.900 ;
        RECT 32.780 58.900 33.780 59.900 ;
        RECT 33.930 58.900 35.530 59.900 ;
        RECT 35.680 58.900 36.680 59.900 ;
        RECT 36.830 58.900 37.830 59.900 ;
        RECT 51.630 60.100 52.630 61.100 ;
        RECT 52.730 60.100 53.730 61.100 ;
        RECT 53.880 60.100 55.480 61.100 ;
        RECT 55.680 60.100 56.680 61.100 ;
        RECT 56.830 60.100 57.830 61.100 ;
        RECT 51.630 58.900 52.630 59.900 ;
        RECT 52.780 58.900 53.780 59.900 ;
        RECT 53.930 58.900 55.530 59.900 ;
        RECT 55.680 58.900 56.680 59.900 ;
        RECT 56.830 58.900 57.830 59.900 ;
        RECT 71.630 60.100 72.630 61.100 ;
        RECT 72.730 60.100 73.730 61.100 ;
        RECT 73.880 60.100 75.480 61.100 ;
        RECT 75.680 60.100 76.680 61.100 ;
        RECT 76.830 60.100 77.830 61.100 ;
        RECT 71.630 58.900 72.630 59.900 ;
        RECT 72.780 58.900 73.780 59.900 ;
        RECT 73.930 58.900 75.530 59.900 ;
        RECT 75.680 58.900 76.680 59.900 ;
        RECT 76.830 58.900 77.830 59.900 ;
        RECT 91.630 60.100 92.630 61.100 ;
        RECT 92.730 60.100 93.730 61.100 ;
        RECT 93.880 60.100 95.480 61.100 ;
        RECT 95.680 60.100 96.680 61.100 ;
        RECT 96.830 60.100 97.830 61.100 ;
        RECT 91.630 58.900 92.630 59.900 ;
        RECT 92.780 58.900 93.780 59.900 ;
        RECT 93.930 58.900 95.530 59.900 ;
        RECT 95.680 58.900 96.680 59.900 ;
        RECT 96.830 58.900 97.830 59.900 ;
        RECT 111.630 60.100 112.630 61.100 ;
        RECT 112.730 60.100 113.730 61.100 ;
        RECT 113.880 60.100 115.480 61.100 ;
        RECT 115.680 60.100 116.680 61.100 ;
        RECT 116.830 60.100 117.830 61.100 ;
        RECT 111.630 58.900 112.630 59.900 ;
        RECT 112.780 58.900 113.780 59.900 ;
        RECT 113.930 58.900 115.530 59.900 ;
        RECT 115.680 58.900 116.680 59.900 ;
        RECT 116.830 58.900 117.830 59.900 ;
        RECT 4.830 52.400 5.530 53.100 ;
        RECT 4.830 51.550 5.530 52.250 ;
        RECT 4.830 50.700 5.530 51.400 ;
        RECT 23.930 52.400 24.630 53.100 ;
        RECT 24.830 52.400 25.530 53.100 ;
        RECT 23.930 51.550 24.630 52.250 ;
        RECT 24.830 51.550 25.530 52.250 ;
        RECT 23.930 50.700 24.630 51.400 ;
        RECT 24.830 50.700 25.530 51.400 ;
        RECT 4.830 48.600 5.530 49.300 ;
        RECT 4.830 47.750 5.530 48.450 ;
        RECT 4.830 46.900 5.530 47.600 ;
        RECT 43.930 52.400 44.630 53.100 ;
        RECT 44.830 52.400 45.530 53.100 ;
        RECT 43.930 51.550 44.630 52.250 ;
        RECT 44.830 51.550 45.530 52.250 ;
        RECT 43.930 50.700 44.630 51.400 ;
        RECT 44.830 50.700 45.530 51.400 ;
        RECT 23.930 48.600 24.630 49.300 ;
        RECT 24.830 48.600 25.530 49.300 ;
        RECT 23.930 47.750 24.630 48.450 ;
        RECT 24.830 47.750 25.530 48.450 ;
        RECT 23.930 46.900 24.630 47.600 ;
        RECT 24.830 46.900 25.530 47.600 ;
        RECT 63.930 52.400 64.630 53.100 ;
        RECT 64.830 52.400 65.530 53.100 ;
        RECT 63.930 51.550 64.630 52.250 ;
        RECT 64.830 51.550 65.530 52.250 ;
        RECT 63.930 50.700 64.630 51.400 ;
        RECT 64.830 50.700 65.530 51.400 ;
        RECT 43.930 48.600 44.630 49.300 ;
        RECT 44.830 48.600 45.530 49.300 ;
        RECT 43.930 47.750 44.630 48.450 ;
        RECT 44.830 47.750 45.530 48.450 ;
        RECT 43.930 46.900 44.630 47.600 ;
        RECT 44.830 46.900 45.530 47.600 ;
        RECT 83.930 52.400 84.630 53.100 ;
        RECT 84.830 52.400 85.530 53.100 ;
        RECT 83.930 51.550 84.630 52.250 ;
        RECT 84.830 51.550 85.530 52.250 ;
        RECT 83.930 50.700 84.630 51.400 ;
        RECT 84.830 50.700 85.530 51.400 ;
        RECT 63.930 48.600 64.630 49.300 ;
        RECT 64.830 48.600 65.530 49.300 ;
        RECT 63.930 47.750 64.630 48.450 ;
        RECT 64.830 47.750 65.530 48.450 ;
        RECT 63.930 46.900 64.630 47.600 ;
        RECT 64.830 46.900 65.530 47.600 ;
        RECT 103.930 52.400 104.630 53.100 ;
        RECT 104.830 52.400 105.530 53.100 ;
        RECT 103.930 51.550 104.630 52.250 ;
        RECT 104.830 51.550 105.530 52.250 ;
        RECT 103.930 50.700 104.630 51.400 ;
        RECT 104.830 50.700 105.530 51.400 ;
        RECT 83.930 48.600 84.630 49.300 ;
        RECT 84.830 48.600 85.530 49.300 ;
        RECT 83.930 47.750 84.630 48.450 ;
        RECT 84.830 47.750 85.530 48.450 ;
        RECT 83.930 46.900 84.630 47.600 ;
        RECT 84.830 46.900 85.530 47.600 ;
        RECT 123.930 52.400 124.630 53.100 ;
        RECT 123.930 51.550 124.630 52.250 ;
        RECT 123.930 50.700 124.630 51.400 ;
        RECT 130.050 50.900 130.410 51.280 ;
        RECT 130.680 50.900 131.040 51.280 ;
        RECT 131.280 50.900 131.640 51.280 ;
        RECT 103.930 48.600 104.630 49.300 ;
        RECT 104.830 48.600 105.530 49.300 ;
        RECT 103.930 47.750 104.630 48.450 ;
        RECT 104.830 47.750 105.530 48.450 ;
        RECT 103.930 46.900 104.630 47.600 ;
        RECT 104.830 46.900 105.530 47.600 ;
        RECT 130.050 50.310 130.410 50.690 ;
        RECT 130.680 50.310 131.040 50.690 ;
        RECT 131.280 50.310 131.640 50.690 ;
        RECT 123.930 48.600 124.630 49.300 ;
        RECT 123.930 47.750 124.630 48.450 ;
        RECT 123.930 46.900 124.630 47.600 ;
        RECT 11.630 40.100 12.630 41.100 ;
        RECT 12.730 40.100 13.730 41.100 ;
        RECT 13.880 40.100 15.480 41.100 ;
        RECT 15.680 40.100 16.680 41.100 ;
        RECT 16.830 40.100 17.830 41.100 ;
        RECT 11.630 38.900 12.630 39.900 ;
        RECT 12.780 38.900 13.780 39.900 ;
        RECT 13.930 38.900 15.530 39.900 ;
        RECT 15.680 38.900 16.680 39.900 ;
        RECT 16.830 38.900 17.830 39.900 ;
        RECT 31.630 40.100 32.630 41.100 ;
        RECT 32.730 40.100 33.730 41.100 ;
        RECT 33.880 40.100 35.480 41.100 ;
        RECT 35.680 40.100 36.680 41.100 ;
        RECT 36.830 40.100 37.830 41.100 ;
        RECT 31.630 38.900 32.630 39.900 ;
        RECT 32.780 38.900 33.780 39.900 ;
        RECT 33.930 38.900 35.530 39.900 ;
        RECT 35.680 38.900 36.680 39.900 ;
        RECT 36.830 38.900 37.830 39.900 ;
        RECT 51.630 40.100 52.630 41.100 ;
        RECT 52.730 40.100 53.730 41.100 ;
        RECT 53.880 40.100 55.480 41.100 ;
        RECT 55.680 40.100 56.680 41.100 ;
        RECT 56.830 40.100 57.830 41.100 ;
        RECT 51.630 38.900 52.630 39.900 ;
        RECT 52.780 38.900 53.780 39.900 ;
        RECT 53.930 38.900 55.530 39.900 ;
        RECT 55.680 38.900 56.680 39.900 ;
        RECT 56.830 38.900 57.830 39.900 ;
        RECT 71.630 40.100 72.630 41.100 ;
        RECT 72.730 40.100 73.730 41.100 ;
        RECT 73.880 40.100 75.480 41.100 ;
        RECT 75.680 40.100 76.680 41.100 ;
        RECT 76.830 40.100 77.830 41.100 ;
        RECT 71.630 38.900 72.630 39.900 ;
        RECT 72.780 38.900 73.780 39.900 ;
        RECT 73.930 38.900 75.530 39.900 ;
        RECT 75.680 38.900 76.680 39.900 ;
        RECT 76.830 38.900 77.830 39.900 ;
        RECT 91.630 40.100 92.630 41.100 ;
        RECT 92.730 40.100 93.730 41.100 ;
        RECT 93.880 40.100 95.480 41.100 ;
        RECT 95.680 40.100 96.680 41.100 ;
        RECT 96.830 40.100 97.830 41.100 ;
        RECT 91.630 38.900 92.630 39.900 ;
        RECT 92.780 38.900 93.780 39.900 ;
        RECT 93.930 38.900 95.530 39.900 ;
        RECT 95.680 38.900 96.680 39.900 ;
        RECT 96.830 38.900 97.830 39.900 ;
        RECT 111.630 40.100 112.630 41.100 ;
        RECT 112.730 40.100 113.730 41.100 ;
        RECT 113.880 40.100 115.480 41.100 ;
        RECT 115.680 40.100 116.680 41.100 ;
        RECT 116.830 40.100 117.830 41.100 ;
        RECT 111.630 38.900 112.630 39.900 ;
        RECT 112.780 38.900 113.780 39.900 ;
        RECT 113.930 38.900 115.530 39.900 ;
        RECT 115.680 38.900 116.680 39.900 ;
        RECT 116.830 38.900 117.830 39.900 ;
        RECT 4.830 32.400 5.530 33.100 ;
        RECT 4.830 31.550 5.530 32.250 ;
        RECT 4.830 30.700 5.530 31.400 ;
        RECT 23.930 32.400 24.630 33.100 ;
        RECT 24.830 32.400 25.530 33.100 ;
        RECT 23.930 31.550 24.630 32.250 ;
        RECT 24.830 31.550 25.530 32.250 ;
        RECT 23.930 30.700 24.630 31.400 ;
        RECT 24.830 30.700 25.530 31.400 ;
        RECT 4.830 28.600 5.530 29.300 ;
        RECT 4.830 27.750 5.530 28.450 ;
        RECT 4.830 26.900 5.530 27.600 ;
        RECT 43.930 32.400 44.630 33.100 ;
        RECT 44.830 32.400 45.530 33.100 ;
        RECT 43.930 31.550 44.630 32.250 ;
        RECT 44.830 31.550 45.530 32.250 ;
        RECT 43.930 30.700 44.630 31.400 ;
        RECT 44.830 30.700 45.530 31.400 ;
        RECT 23.930 28.600 24.630 29.300 ;
        RECT 24.830 28.600 25.530 29.300 ;
        RECT 23.930 27.750 24.630 28.450 ;
        RECT 24.830 27.750 25.530 28.450 ;
        RECT 23.930 26.900 24.630 27.600 ;
        RECT 24.830 26.900 25.530 27.600 ;
        RECT 63.930 32.400 64.630 33.100 ;
        RECT 64.830 32.400 65.530 33.100 ;
        RECT 63.930 31.550 64.630 32.250 ;
        RECT 64.830 31.550 65.530 32.250 ;
        RECT 63.930 30.700 64.630 31.400 ;
        RECT 64.830 30.700 65.530 31.400 ;
        RECT 43.930 28.600 44.630 29.300 ;
        RECT 44.830 28.600 45.530 29.300 ;
        RECT 43.930 27.750 44.630 28.450 ;
        RECT 44.830 27.750 45.530 28.450 ;
        RECT 43.930 26.900 44.630 27.600 ;
        RECT 44.830 26.900 45.530 27.600 ;
        RECT 83.930 32.400 84.630 33.100 ;
        RECT 84.830 32.400 85.530 33.100 ;
        RECT 83.930 31.550 84.630 32.250 ;
        RECT 84.830 31.550 85.530 32.250 ;
        RECT 83.930 30.700 84.630 31.400 ;
        RECT 84.830 30.700 85.530 31.400 ;
        RECT 63.930 28.600 64.630 29.300 ;
        RECT 64.830 28.600 65.530 29.300 ;
        RECT 63.930 27.750 64.630 28.450 ;
        RECT 64.830 27.750 65.530 28.450 ;
        RECT 63.930 26.900 64.630 27.600 ;
        RECT 64.830 26.900 65.530 27.600 ;
        RECT 103.930 32.400 104.630 33.100 ;
        RECT 104.830 32.400 105.530 33.100 ;
        RECT 103.930 31.550 104.630 32.250 ;
        RECT 104.830 31.550 105.530 32.250 ;
        RECT 103.930 30.700 104.630 31.400 ;
        RECT 104.830 30.700 105.530 31.400 ;
        RECT 83.930 28.600 84.630 29.300 ;
        RECT 84.830 28.600 85.530 29.300 ;
        RECT 83.930 27.750 84.630 28.450 ;
        RECT 84.830 27.750 85.530 28.450 ;
        RECT 83.930 26.900 84.630 27.600 ;
        RECT 84.830 26.900 85.530 27.600 ;
        RECT 123.930 32.400 124.630 33.100 ;
        RECT 123.930 31.550 124.630 32.250 ;
        RECT 123.930 30.700 124.630 31.400 ;
        RECT 130.050 31.080 130.410 31.460 ;
        RECT 130.680 31.080 131.040 31.460 ;
        RECT 131.280 31.080 131.640 31.460 ;
        RECT 130.050 30.490 130.410 30.870 ;
        RECT 130.680 30.490 131.040 30.870 ;
        RECT 131.280 30.490 131.640 30.870 ;
        RECT 103.930 28.600 104.630 29.300 ;
        RECT 104.830 28.600 105.530 29.300 ;
        RECT 103.930 27.750 104.630 28.450 ;
        RECT 104.830 27.750 105.530 28.450 ;
        RECT 103.930 26.900 104.630 27.600 ;
        RECT 104.830 26.900 105.530 27.600 ;
        RECT 123.930 28.600 124.630 29.300 ;
        RECT 123.930 27.750 124.630 28.450 ;
        RECT 123.930 26.900 124.630 27.600 ;
        RECT 11.630 20.100 12.630 21.100 ;
        RECT 12.730 20.100 13.730 21.100 ;
        RECT 13.880 20.100 15.480 21.100 ;
        RECT 15.680 20.100 16.680 21.100 ;
        RECT 16.830 20.100 17.830 21.100 ;
        RECT 11.630 18.900 12.630 19.900 ;
        RECT 12.780 18.900 13.780 19.900 ;
        RECT 13.930 18.900 15.530 19.900 ;
        RECT 15.680 18.900 16.680 19.900 ;
        RECT 16.830 18.900 17.830 19.900 ;
        RECT 31.630 20.100 32.630 21.100 ;
        RECT 32.730 20.100 33.730 21.100 ;
        RECT 33.880 20.100 35.480 21.100 ;
        RECT 35.680 20.100 36.680 21.100 ;
        RECT 36.830 20.100 37.830 21.100 ;
        RECT 31.630 18.900 32.630 19.900 ;
        RECT 32.780 18.900 33.780 19.900 ;
        RECT 33.930 18.900 35.530 19.900 ;
        RECT 35.680 18.900 36.680 19.900 ;
        RECT 36.830 18.900 37.830 19.900 ;
        RECT 51.630 20.100 52.630 21.100 ;
        RECT 52.730 20.100 53.730 21.100 ;
        RECT 53.880 20.100 55.480 21.100 ;
        RECT 55.680 20.100 56.680 21.100 ;
        RECT 56.830 20.100 57.830 21.100 ;
        RECT 51.630 18.900 52.630 19.900 ;
        RECT 52.780 18.900 53.780 19.900 ;
        RECT 53.930 18.900 55.530 19.900 ;
        RECT 55.680 18.900 56.680 19.900 ;
        RECT 56.830 18.900 57.830 19.900 ;
        RECT 71.630 20.100 72.630 21.100 ;
        RECT 72.730 20.100 73.730 21.100 ;
        RECT 73.880 20.100 75.480 21.100 ;
        RECT 75.680 20.100 76.680 21.100 ;
        RECT 76.830 20.100 77.830 21.100 ;
        RECT 71.630 18.900 72.630 19.900 ;
        RECT 72.780 18.900 73.780 19.900 ;
        RECT 73.930 18.900 75.530 19.900 ;
        RECT 75.680 18.900 76.680 19.900 ;
        RECT 76.830 18.900 77.830 19.900 ;
        RECT 91.630 20.100 92.630 21.100 ;
        RECT 92.730 20.100 93.730 21.100 ;
        RECT 93.880 20.100 95.480 21.100 ;
        RECT 95.680 20.100 96.680 21.100 ;
        RECT 96.830 20.100 97.830 21.100 ;
        RECT 91.630 18.900 92.630 19.900 ;
        RECT 92.780 18.900 93.780 19.900 ;
        RECT 93.930 18.900 95.530 19.900 ;
        RECT 95.680 18.900 96.680 19.900 ;
        RECT 96.830 18.900 97.830 19.900 ;
        RECT 111.630 20.100 112.630 21.100 ;
        RECT 112.730 20.100 113.730 21.100 ;
        RECT 113.880 20.100 115.480 21.100 ;
        RECT 115.680 20.100 116.680 21.100 ;
        RECT 116.830 20.100 117.830 21.100 ;
        RECT 111.630 18.900 112.630 19.900 ;
        RECT 112.780 18.900 113.780 19.900 ;
        RECT 113.930 18.900 115.530 19.900 ;
        RECT 115.680 18.900 116.680 19.900 ;
        RECT 116.830 18.900 117.830 19.900 ;
        RECT 4.830 12.400 5.530 13.100 ;
        RECT 4.830 11.550 5.530 12.250 ;
        RECT 4.830 10.700 5.530 11.400 ;
        RECT 23.930 12.400 24.630 13.100 ;
        RECT 24.830 12.400 25.530 13.100 ;
        RECT 23.930 11.550 24.630 12.250 ;
        RECT 24.830 11.550 25.530 12.250 ;
        RECT 23.930 10.700 24.630 11.400 ;
        RECT 24.830 10.700 25.530 11.400 ;
        RECT 4.830 8.600 5.530 9.300 ;
        RECT 4.830 7.750 5.530 8.450 ;
        RECT 4.830 6.900 5.530 7.600 ;
        RECT 43.930 12.400 44.630 13.100 ;
        RECT 44.830 12.400 45.530 13.100 ;
        RECT 43.930 11.550 44.630 12.250 ;
        RECT 44.830 11.550 45.530 12.250 ;
        RECT 43.930 10.700 44.630 11.400 ;
        RECT 44.830 10.700 45.530 11.400 ;
        RECT 23.930 8.600 24.630 9.300 ;
        RECT 24.830 8.600 25.530 9.300 ;
        RECT 23.930 7.750 24.630 8.450 ;
        RECT 24.830 7.750 25.530 8.450 ;
        RECT 23.930 6.900 24.630 7.600 ;
        RECT 24.830 6.900 25.530 7.600 ;
        RECT 63.930 12.400 64.630 13.100 ;
        RECT 64.830 12.400 65.530 13.100 ;
        RECT 63.930 11.550 64.630 12.250 ;
        RECT 64.830 11.550 65.530 12.250 ;
        RECT 63.930 10.700 64.630 11.400 ;
        RECT 64.830 10.700 65.530 11.400 ;
        RECT 43.930 8.600 44.630 9.300 ;
        RECT 44.830 8.600 45.530 9.300 ;
        RECT 43.930 7.750 44.630 8.450 ;
        RECT 44.830 7.750 45.530 8.450 ;
        RECT 43.930 6.900 44.630 7.600 ;
        RECT 44.830 6.900 45.530 7.600 ;
        RECT 83.930 12.400 84.630 13.100 ;
        RECT 84.830 12.400 85.530 13.100 ;
        RECT 83.930 11.550 84.630 12.250 ;
        RECT 84.830 11.550 85.530 12.250 ;
        RECT 83.930 10.700 84.630 11.400 ;
        RECT 84.830 10.700 85.530 11.400 ;
        RECT 63.930 8.600 64.630 9.300 ;
        RECT 64.830 8.600 65.530 9.300 ;
        RECT 63.930 7.750 64.630 8.450 ;
        RECT 64.830 7.750 65.530 8.450 ;
        RECT 63.930 6.900 64.630 7.600 ;
        RECT 64.830 6.900 65.530 7.600 ;
        RECT 103.930 12.400 104.630 13.100 ;
        RECT 104.830 12.400 105.530 13.100 ;
        RECT 103.930 11.550 104.630 12.250 ;
        RECT 104.830 11.550 105.530 12.250 ;
        RECT 103.930 10.700 104.630 11.400 ;
        RECT 104.830 10.700 105.530 11.400 ;
        RECT 83.930 8.600 84.630 9.300 ;
        RECT 84.830 8.600 85.530 9.300 ;
        RECT 83.930 7.750 84.630 8.450 ;
        RECT 84.830 7.750 85.530 8.450 ;
        RECT 83.930 6.900 84.630 7.600 ;
        RECT 84.830 6.900 85.530 7.600 ;
        RECT 123.930 12.400 124.630 13.100 ;
        RECT 123.930 11.550 124.630 12.250 ;
        RECT 123.930 10.700 124.630 11.400 ;
        RECT 130.050 11.020 130.410 11.400 ;
        RECT 130.680 11.020 131.040 11.400 ;
        RECT 131.280 11.020 131.640 11.400 ;
        RECT 103.930 8.600 104.630 9.300 ;
        RECT 104.830 8.600 105.530 9.300 ;
        RECT 103.930 7.750 104.630 8.450 ;
        RECT 104.830 7.750 105.530 8.450 ;
        RECT 103.930 6.900 104.630 7.600 ;
        RECT 104.830 6.900 105.530 7.600 ;
        RECT 130.050 10.430 130.410 10.810 ;
        RECT 130.680 10.430 131.040 10.810 ;
        RECT 131.280 10.430 131.640 10.810 ;
        RECT 123.930 8.600 124.630 9.300 ;
        RECT 123.930 7.750 124.630 8.450 ;
        RECT 123.930 6.900 124.630 7.600 ;
        RECT 11.630 0.100 12.630 1.100 ;
        RECT 12.730 0.100 13.730 1.100 ;
        RECT 13.880 0.100 15.480 1.100 ;
        RECT 15.680 0.100 16.680 1.100 ;
        RECT 16.830 0.100 17.830 1.100 ;
        RECT 31.630 0.100 32.630 1.100 ;
        RECT 32.730 0.100 33.730 1.100 ;
        RECT 33.880 0.100 35.480 1.100 ;
        RECT 35.680 0.100 36.680 1.100 ;
        RECT 36.830 0.100 37.830 1.100 ;
        RECT 51.630 0.100 52.630 1.100 ;
        RECT 52.730 0.100 53.730 1.100 ;
        RECT 53.880 0.100 55.480 1.100 ;
        RECT 55.680 0.100 56.680 1.100 ;
        RECT 56.830 0.100 57.830 1.100 ;
        RECT 71.630 0.100 72.630 1.100 ;
        RECT 72.730 0.100 73.730 1.100 ;
        RECT 73.880 0.100 75.480 1.100 ;
        RECT 75.680 0.100 76.680 1.100 ;
        RECT 76.830 0.100 77.830 1.100 ;
        RECT 91.630 0.100 92.630 1.100 ;
        RECT 92.730 0.100 93.730 1.100 ;
        RECT 93.880 0.100 95.480 1.100 ;
        RECT 95.680 0.100 96.680 1.100 ;
        RECT 96.830 0.100 97.830 1.100 ;
        RECT 111.630 0.100 112.630 1.100 ;
        RECT 112.730 0.100 113.730 1.100 ;
        RECT 113.880 0.100 115.480 1.100 ;
        RECT 115.680 0.100 116.680 1.100 ;
        RECT 116.830 0.100 117.830 1.100 ;
      LAYER met2 ;
        RECT 11.530 339.100 17.930 340.000 ;
        RECT 31.530 339.100 37.930 340.000 ;
        RECT 51.530 339.100 57.930 340.000 ;
        RECT 71.530 339.100 77.930 340.000 ;
        RECT 91.530 339.100 97.930 340.000 ;
        RECT 111.530 339.100 117.930 340.000 ;
        RECT 9.630 338.600 19.830 339.100 ;
        RECT 29.630 338.600 39.830 339.100 ;
        RECT 49.630 338.600 59.830 339.100 ;
        RECT 69.630 338.600 79.830 339.100 ;
        RECT 89.630 338.600 99.830 339.100 ;
        RECT 109.630 338.600 119.830 339.100 ;
        RECT 6.530 338.550 22.930 338.600 ;
        RECT 6.530 338.000 10.330 338.550 ;
        RECT 10.030 337.550 10.330 338.000 ;
        RECT 6.480 337.400 10.330 337.550 ;
        RECT 10.030 336.950 10.330 337.400 ;
        RECT 6.480 336.800 10.330 336.950 ;
        RECT 10.030 336.350 10.330 336.800 ;
        RECT 6.480 336.200 10.330 336.350 ;
        RECT 10.030 335.750 10.330 336.200 ;
        RECT 6.480 335.600 10.330 335.750 ;
        RECT 10.030 335.150 10.330 335.600 ;
        RECT 6.480 335.000 10.330 335.150 ;
        RECT 10.030 334.550 10.330 335.000 ;
        RECT 6.480 334.400 10.330 334.550 ;
        RECT 10.030 333.950 10.330 334.400 ;
        RECT 6.480 333.800 10.330 333.950 ;
        RECT 10.030 333.350 10.330 333.800 ;
        RECT 6.480 333.200 10.330 333.350 ;
        RECT 4.730 326.800 5.630 333.200 ;
        RECT 10.030 332.750 10.330 333.200 ;
        RECT 6.480 332.600 10.330 332.750 ;
        RECT 10.030 332.150 10.330 332.600 ;
        RECT 6.480 332.000 10.330 332.150 ;
        RECT 10.030 331.550 10.330 332.000 ;
        RECT 6.480 331.400 10.330 331.550 ;
        RECT 10.030 330.950 10.330 331.400 ;
        RECT 6.480 330.800 10.330 330.950 ;
        RECT 10.030 330.350 10.330 330.800 ;
        RECT 10.780 330.350 10.930 338.550 ;
        RECT 11.380 330.350 11.530 338.550 ;
        RECT 11.980 330.350 12.130 338.550 ;
        RECT 12.580 330.350 12.730 338.550 ;
        RECT 13.180 330.350 13.330 338.550 ;
        RECT 13.780 330.350 13.930 338.550 ;
        RECT 10.030 329.200 10.330 329.650 ;
        RECT 6.480 329.050 10.330 329.200 ;
        RECT 10.030 328.600 10.330 329.050 ;
        RECT 6.480 328.450 10.330 328.600 ;
        RECT 10.030 328.000 10.330 328.450 ;
        RECT 6.480 327.850 10.330 328.000 ;
        RECT 10.030 327.400 10.330 327.850 ;
        RECT 6.480 327.250 10.330 327.400 ;
        RECT 10.030 326.800 10.330 327.250 ;
        RECT 6.480 326.650 10.330 326.800 ;
        RECT 10.030 326.200 10.330 326.650 ;
        RECT 6.480 326.050 10.330 326.200 ;
        RECT 10.030 325.600 10.330 326.050 ;
        RECT 6.480 325.450 10.330 325.600 ;
        RECT 10.030 325.000 10.330 325.450 ;
        RECT 6.480 324.850 10.330 325.000 ;
        RECT 10.030 324.400 10.330 324.850 ;
        RECT 6.480 324.250 10.330 324.400 ;
        RECT 10.030 323.800 10.330 324.250 ;
        RECT 6.480 323.650 10.330 323.800 ;
        RECT 10.030 323.200 10.330 323.650 ;
        RECT 6.480 323.050 10.330 323.200 ;
        RECT 10.030 322.600 10.330 323.050 ;
        RECT 6.480 322.450 10.330 322.600 ;
        RECT 10.030 322.000 10.330 322.450 ;
        RECT 6.530 321.450 10.330 322.000 ;
        RECT 10.780 321.450 10.930 329.650 ;
        RECT 11.380 321.450 11.530 329.650 ;
        RECT 11.980 321.450 12.130 329.650 ;
        RECT 12.580 321.450 12.730 329.650 ;
        RECT 13.180 321.450 13.330 329.650 ;
        RECT 13.780 321.450 13.930 329.650 ;
        RECT 14.380 321.450 15.080 338.550 ;
        RECT 15.530 330.350 15.680 338.550 ;
        RECT 16.130 330.350 16.280 338.550 ;
        RECT 16.730 330.350 16.880 338.550 ;
        RECT 17.330 330.350 17.480 338.550 ;
        RECT 17.930 330.350 18.080 338.550 ;
        RECT 18.530 330.350 18.680 338.550 ;
        RECT 19.130 338.000 22.930 338.550 ;
        RECT 26.530 338.550 42.930 338.600 ;
        RECT 26.530 338.000 30.330 338.550 ;
        RECT 19.130 337.550 19.430 338.000 ;
        RECT 30.030 337.550 30.330 338.000 ;
        RECT 19.130 337.400 22.980 337.550 ;
        RECT 26.480 337.400 30.330 337.550 ;
        RECT 19.130 336.950 19.430 337.400 ;
        RECT 30.030 336.950 30.330 337.400 ;
        RECT 19.130 336.800 22.980 336.950 ;
        RECT 26.480 336.800 30.330 336.950 ;
        RECT 19.130 336.350 19.430 336.800 ;
        RECT 30.030 336.350 30.330 336.800 ;
        RECT 19.130 336.200 22.980 336.350 ;
        RECT 26.480 336.200 30.330 336.350 ;
        RECT 19.130 335.750 19.430 336.200 ;
        RECT 30.030 335.750 30.330 336.200 ;
        RECT 19.130 335.600 22.980 335.750 ;
        RECT 26.480 335.600 30.330 335.750 ;
        RECT 19.130 335.150 19.430 335.600 ;
        RECT 30.030 335.150 30.330 335.600 ;
        RECT 19.130 335.000 22.980 335.150 ;
        RECT 26.480 335.000 30.330 335.150 ;
        RECT 19.130 334.550 19.430 335.000 ;
        RECT 30.030 334.550 30.330 335.000 ;
        RECT 19.130 334.400 22.980 334.550 ;
        RECT 26.480 334.400 30.330 334.550 ;
        RECT 19.130 333.950 19.430 334.400 ;
        RECT 30.030 333.950 30.330 334.400 ;
        RECT 19.130 333.800 22.980 333.950 ;
        RECT 26.480 333.800 30.330 333.950 ;
        RECT 19.130 333.350 19.430 333.800 ;
        RECT 30.030 333.350 30.330 333.800 ;
        RECT 19.130 333.200 22.980 333.350 ;
        RECT 26.480 333.200 30.330 333.350 ;
        RECT 19.130 332.750 19.430 333.200 ;
        RECT 19.130 332.600 22.980 332.750 ;
        RECT 19.130 332.150 19.430 332.600 ;
        RECT 19.130 332.000 22.980 332.150 ;
        RECT 19.130 331.550 19.430 332.000 ;
        RECT 19.130 331.400 22.980 331.550 ;
        RECT 19.130 330.950 19.430 331.400 ;
        RECT 19.130 330.800 22.980 330.950 ;
        RECT 19.130 330.350 19.430 330.800 ;
        RECT 15.530 321.450 15.680 329.650 ;
        RECT 16.130 321.450 16.280 329.650 ;
        RECT 16.730 321.450 16.880 329.650 ;
        RECT 17.330 321.450 17.480 329.650 ;
        RECT 17.930 321.450 18.080 329.650 ;
        RECT 18.530 321.450 18.680 329.650 ;
        RECT 19.130 329.200 19.430 329.650 ;
        RECT 19.130 329.050 22.980 329.200 ;
        RECT 19.130 328.600 19.430 329.050 ;
        RECT 19.130 328.450 22.980 328.600 ;
        RECT 19.130 328.000 19.430 328.450 ;
        RECT 19.130 327.850 22.980 328.000 ;
        RECT 19.130 327.400 19.430 327.850 ;
        RECT 19.130 327.250 22.980 327.400 ;
        RECT 19.130 326.800 19.430 327.250 ;
        RECT 23.830 326.800 25.630 333.200 ;
        RECT 30.030 332.750 30.330 333.200 ;
        RECT 26.480 332.600 30.330 332.750 ;
        RECT 30.030 332.150 30.330 332.600 ;
        RECT 26.480 332.000 30.330 332.150 ;
        RECT 30.030 331.550 30.330 332.000 ;
        RECT 26.480 331.400 30.330 331.550 ;
        RECT 30.030 330.950 30.330 331.400 ;
        RECT 26.480 330.800 30.330 330.950 ;
        RECT 30.030 330.350 30.330 330.800 ;
        RECT 30.780 330.350 30.930 338.550 ;
        RECT 31.380 330.350 31.530 338.550 ;
        RECT 31.980 330.350 32.130 338.550 ;
        RECT 32.580 330.350 32.730 338.550 ;
        RECT 33.180 330.350 33.330 338.550 ;
        RECT 33.780 330.350 33.930 338.550 ;
        RECT 30.030 329.200 30.330 329.650 ;
        RECT 26.480 329.050 30.330 329.200 ;
        RECT 30.030 328.600 30.330 329.050 ;
        RECT 26.480 328.450 30.330 328.600 ;
        RECT 30.030 328.000 30.330 328.450 ;
        RECT 26.480 327.850 30.330 328.000 ;
        RECT 30.030 327.400 30.330 327.850 ;
        RECT 26.480 327.250 30.330 327.400 ;
        RECT 30.030 326.800 30.330 327.250 ;
        RECT 19.130 326.650 22.980 326.800 ;
        RECT 26.480 326.650 30.330 326.800 ;
        RECT 19.130 326.200 19.430 326.650 ;
        RECT 30.030 326.200 30.330 326.650 ;
        RECT 19.130 326.050 22.980 326.200 ;
        RECT 26.480 326.050 30.330 326.200 ;
        RECT 19.130 325.600 19.430 326.050 ;
        RECT 30.030 325.600 30.330 326.050 ;
        RECT 19.130 325.450 22.980 325.600 ;
        RECT 26.480 325.450 30.330 325.600 ;
        RECT 19.130 325.000 19.430 325.450 ;
        RECT 30.030 325.000 30.330 325.450 ;
        RECT 19.130 324.850 22.980 325.000 ;
        RECT 26.480 324.850 30.330 325.000 ;
        RECT 19.130 324.400 19.430 324.850 ;
        RECT 30.030 324.400 30.330 324.850 ;
        RECT 19.130 324.250 22.980 324.400 ;
        RECT 26.480 324.250 30.330 324.400 ;
        RECT 19.130 323.800 19.430 324.250 ;
        RECT 30.030 323.800 30.330 324.250 ;
        RECT 19.130 323.650 22.980 323.800 ;
        RECT 26.480 323.650 30.330 323.800 ;
        RECT 19.130 323.200 19.430 323.650 ;
        RECT 30.030 323.200 30.330 323.650 ;
        RECT 19.130 323.050 22.980 323.200 ;
        RECT 26.480 323.050 30.330 323.200 ;
        RECT 19.130 322.600 19.430 323.050 ;
        RECT 30.030 322.600 30.330 323.050 ;
        RECT 19.130 322.450 22.980 322.600 ;
        RECT 26.480 322.450 30.330 322.600 ;
        RECT 19.130 322.000 19.430 322.450 ;
        RECT 30.030 322.000 30.330 322.450 ;
        RECT 19.130 321.450 22.930 322.000 ;
        RECT 6.530 321.400 22.930 321.450 ;
        RECT 26.530 321.450 30.330 322.000 ;
        RECT 30.780 321.450 30.930 329.650 ;
        RECT 31.380 321.450 31.530 329.650 ;
        RECT 31.980 321.450 32.130 329.650 ;
        RECT 32.580 321.450 32.730 329.650 ;
        RECT 33.180 321.450 33.330 329.650 ;
        RECT 33.780 321.450 33.930 329.650 ;
        RECT 34.380 321.450 35.080 338.550 ;
        RECT 35.530 330.350 35.680 338.550 ;
        RECT 36.130 330.350 36.280 338.550 ;
        RECT 36.730 330.350 36.880 338.550 ;
        RECT 37.330 330.350 37.480 338.550 ;
        RECT 37.930 330.350 38.080 338.550 ;
        RECT 38.530 330.350 38.680 338.550 ;
        RECT 39.130 338.000 42.930 338.550 ;
        RECT 46.530 338.550 62.930 338.600 ;
        RECT 46.530 338.000 50.330 338.550 ;
        RECT 39.130 337.550 39.430 338.000 ;
        RECT 50.030 337.550 50.330 338.000 ;
        RECT 39.130 337.400 42.980 337.550 ;
        RECT 46.480 337.400 50.330 337.550 ;
        RECT 39.130 336.950 39.430 337.400 ;
        RECT 50.030 336.950 50.330 337.400 ;
        RECT 39.130 336.800 42.980 336.950 ;
        RECT 46.480 336.800 50.330 336.950 ;
        RECT 39.130 336.350 39.430 336.800 ;
        RECT 50.030 336.350 50.330 336.800 ;
        RECT 39.130 336.200 42.980 336.350 ;
        RECT 46.480 336.200 50.330 336.350 ;
        RECT 39.130 335.750 39.430 336.200 ;
        RECT 50.030 335.750 50.330 336.200 ;
        RECT 39.130 335.600 42.980 335.750 ;
        RECT 46.480 335.600 50.330 335.750 ;
        RECT 39.130 335.150 39.430 335.600 ;
        RECT 50.030 335.150 50.330 335.600 ;
        RECT 39.130 335.000 42.980 335.150 ;
        RECT 46.480 335.000 50.330 335.150 ;
        RECT 39.130 334.550 39.430 335.000 ;
        RECT 50.030 334.550 50.330 335.000 ;
        RECT 39.130 334.400 42.980 334.550 ;
        RECT 46.480 334.400 50.330 334.550 ;
        RECT 39.130 333.950 39.430 334.400 ;
        RECT 50.030 333.950 50.330 334.400 ;
        RECT 39.130 333.800 42.980 333.950 ;
        RECT 46.480 333.800 50.330 333.950 ;
        RECT 39.130 333.350 39.430 333.800 ;
        RECT 50.030 333.350 50.330 333.800 ;
        RECT 39.130 333.200 42.980 333.350 ;
        RECT 46.480 333.200 50.330 333.350 ;
        RECT 39.130 332.750 39.430 333.200 ;
        RECT 39.130 332.600 42.980 332.750 ;
        RECT 39.130 332.150 39.430 332.600 ;
        RECT 39.130 332.000 42.980 332.150 ;
        RECT 39.130 331.550 39.430 332.000 ;
        RECT 39.130 331.400 42.980 331.550 ;
        RECT 39.130 330.950 39.430 331.400 ;
        RECT 39.130 330.800 42.980 330.950 ;
        RECT 39.130 330.350 39.430 330.800 ;
        RECT 35.530 321.450 35.680 329.650 ;
        RECT 36.130 321.450 36.280 329.650 ;
        RECT 36.730 321.450 36.880 329.650 ;
        RECT 37.330 321.450 37.480 329.650 ;
        RECT 37.930 321.450 38.080 329.650 ;
        RECT 38.530 321.450 38.680 329.650 ;
        RECT 39.130 329.200 39.430 329.650 ;
        RECT 39.130 329.050 42.980 329.200 ;
        RECT 39.130 328.600 39.430 329.050 ;
        RECT 39.130 328.450 42.980 328.600 ;
        RECT 39.130 328.000 39.430 328.450 ;
        RECT 39.130 327.850 42.980 328.000 ;
        RECT 39.130 327.400 39.430 327.850 ;
        RECT 39.130 327.250 42.980 327.400 ;
        RECT 39.130 326.800 39.430 327.250 ;
        RECT 43.830 326.800 45.630 333.200 ;
        RECT 50.030 332.750 50.330 333.200 ;
        RECT 46.480 332.600 50.330 332.750 ;
        RECT 50.030 332.150 50.330 332.600 ;
        RECT 46.480 332.000 50.330 332.150 ;
        RECT 50.030 331.550 50.330 332.000 ;
        RECT 46.480 331.400 50.330 331.550 ;
        RECT 50.030 330.950 50.330 331.400 ;
        RECT 46.480 330.800 50.330 330.950 ;
        RECT 50.030 330.350 50.330 330.800 ;
        RECT 50.780 330.350 50.930 338.550 ;
        RECT 51.380 330.350 51.530 338.550 ;
        RECT 51.980 330.350 52.130 338.550 ;
        RECT 52.580 330.350 52.730 338.550 ;
        RECT 53.180 330.350 53.330 338.550 ;
        RECT 53.780 330.350 53.930 338.550 ;
        RECT 50.030 329.200 50.330 329.650 ;
        RECT 46.480 329.050 50.330 329.200 ;
        RECT 50.030 328.600 50.330 329.050 ;
        RECT 46.480 328.450 50.330 328.600 ;
        RECT 50.030 328.000 50.330 328.450 ;
        RECT 46.480 327.850 50.330 328.000 ;
        RECT 50.030 327.400 50.330 327.850 ;
        RECT 46.480 327.250 50.330 327.400 ;
        RECT 50.030 326.800 50.330 327.250 ;
        RECT 39.130 326.650 42.980 326.800 ;
        RECT 46.480 326.650 50.330 326.800 ;
        RECT 39.130 326.200 39.430 326.650 ;
        RECT 50.030 326.200 50.330 326.650 ;
        RECT 39.130 326.050 42.980 326.200 ;
        RECT 46.480 326.050 50.330 326.200 ;
        RECT 39.130 325.600 39.430 326.050 ;
        RECT 50.030 325.600 50.330 326.050 ;
        RECT 39.130 325.450 42.980 325.600 ;
        RECT 46.480 325.450 50.330 325.600 ;
        RECT 39.130 325.000 39.430 325.450 ;
        RECT 50.030 325.000 50.330 325.450 ;
        RECT 39.130 324.850 42.980 325.000 ;
        RECT 46.480 324.850 50.330 325.000 ;
        RECT 39.130 324.400 39.430 324.850 ;
        RECT 50.030 324.400 50.330 324.850 ;
        RECT 39.130 324.250 42.980 324.400 ;
        RECT 46.480 324.250 50.330 324.400 ;
        RECT 39.130 323.800 39.430 324.250 ;
        RECT 50.030 323.800 50.330 324.250 ;
        RECT 39.130 323.650 42.980 323.800 ;
        RECT 46.480 323.650 50.330 323.800 ;
        RECT 39.130 323.200 39.430 323.650 ;
        RECT 50.030 323.200 50.330 323.650 ;
        RECT 39.130 323.050 42.980 323.200 ;
        RECT 46.480 323.050 50.330 323.200 ;
        RECT 39.130 322.600 39.430 323.050 ;
        RECT 50.030 322.600 50.330 323.050 ;
        RECT 39.130 322.450 42.980 322.600 ;
        RECT 46.480 322.450 50.330 322.600 ;
        RECT 39.130 322.000 39.430 322.450 ;
        RECT 50.030 322.000 50.330 322.450 ;
        RECT 39.130 321.450 42.930 322.000 ;
        RECT 26.530 321.400 42.930 321.450 ;
        RECT 46.530 321.450 50.330 322.000 ;
        RECT 50.780 321.450 50.930 329.650 ;
        RECT 51.380 321.450 51.530 329.650 ;
        RECT 51.980 321.450 52.130 329.650 ;
        RECT 52.580 321.450 52.730 329.650 ;
        RECT 53.180 321.450 53.330 329.650 ;
        RECT 53.780 321.450 53.930 329.650 ;
        RECT 54.380 321.450 55.080 338.550 ;
        RECT 55.530 330.350 55.680 338.550 ;
        RECT 56.130 330.350 56.280 338.550 ;
        RECT 56.730 330.350 56.880 338.550 ;
        RECT 57.330 330.350 57.480 338.550 ;
        RECT 57.930 330.350 58.080 338.550 ;
        RECT 58.530 330.350 58.680 338.550 ;
        RECT 59.130 338.000 62.930 338.550 ;
        RECT 66.530 338.550 82.930 338.600 ;
        RECT 66.530 338.000 70.330 338.550 ;
        RECT 59.130 337.550 59.430 338.000 ;
        RECT 70.030 337.550 70.330 338.000 ;
        RECT 59.130 337.400 62.980 337.550 ;
        RECT 66.480 337.400 70.330 337.550 ;
        RECT 59.130 336.950 59.430 337.400 ;
        RECT 70.030 336.950 70.330 337.400 ;
        RECT 59.130 336.800 62.980 336.950 ;
        RECT 66.480 336.800 70.330 336.950 ;
        RECT 59.130 336.350 59.430 336.800 ;
        RECT 70.030 336.350 70.330 336.800 ;
        RECT 59.130 336.200 62.980 336.350 ;
        RECT 66.480 336.200 70.330 336.350 ;
        RECT 59.130 335.750 59.430 336.200 ;
        RECT 70.030 335.750 70.330 336.200 ;
        RECT 59.130 335.600 62.980 335.750 ;
        RECT 66.480 335.600 70.330 335.750 ;
        RECT 59.130 335.150 59.430 335.600 ;
        RECT 70.030 335.150 70.330 335.600 ;
        RECT 59.130 335.000 62.980 335.150 ;
        RECT 66.480 335.000 70.330 335.150 ;
        RECT 59.130 334.550 59.430 335.000 ;
        RECT 70.030 334.550 70.330 335.000 ;
        RECT 59.130 334.400 62.980 334.550 ;
        RECT 66.480 334.400 70.330 334.550 ;
        RECT 59.130 333.950 59.430 334.400 ;
        RECT 70.030 333.950 70.330 334.400 ;
        RECT 59.130 333.800 62.980 333.950 ;
        RECT 66.480 333.800 70.330 333.950 ;
        RECT 59.130 333.350 59.430 333.800 ;
        RECT 70.030 333.350 70.330 333.800 ;
        RECT 59.130 333.200 62.980 333.350 ;
        RECT 66.480 333.200 70.330 333.350 ;
        RECT 59.130 332.750 59.430 333.200 ;
        RECT 59.130 332.600 62.980 332.750 ;
        RECT 59.130 332.150 59.430 332.600 ;
        RECT 59.130 332.000 62.980 332.150 ;
        RECT 59.130 331.550 59.430 332.000 ;
        RECT 59.130 331.400 62.980 331.550 ;
        RECT 59.130 330.950 59.430 331.400 ;
        RECT 59.130 330.800 62.980 330.950 ;
        RECT 59.130 330.350 59.430 330.800 ;
        RECT 55.530 321.450 55.680 329.650 ;
        RECT 56.130 321.450 56.280 329.650 ;
        RECT 56.730 321.450 56.880 329.650 ;
        RECT 57.330 321.450 57.480 329.650 ;
        RECT 57.930 321.450 58.080 329.650 ;
        RECT 58.530 321.450 58.680 329.650 ;
        RECT 59.130 329.200 59.430 329.650 ;
        RECT 59.130 329.050 62.980 329.200 ;
        RECT 59.130 328.600 59.430 329.050 ;
        RECT 59.130 328.450 62.980 328.600 ;
        RECT 59.130 328.000 59.430 328.450 ;
        RECT 59.130 327.850 62.980 328.000 ;
        RECT 59.130 327.400 59.430 327.850 ;
        RECT 59.130 327.250 62.980 327.400 ;
        RECT 59.130 326.800 59.430 327.250 ;
        RECT 63.830 326.800 65.630 333.200 ;
        RECT 70.030 332.750 70.330 333.200 ;
        RECT 66.480 332.600 70.330 332.750 ;
        RECT 70.030 332.150 70.330 332.600 ;
        RECT 66.480 332.000 70.330 332.150 ;
        RECT 70.030 331.550 70.330 332.000 ;
        RECT 66.480 331.400 70.330 331.550 ;
        RECT 70.030 330.950 70.330 331.400 ;
        RECT 66.480 330.800 70.330 330.950 ;
        RECT 70.030 330.350 70.330 330.800 ;
        RECT 70.780 330.350 70.930 338.550 ;
        RECT 71.380 330.350 71.530 338.550 ;
        RECT 71.980 330.350 72.130 338.550 ;
        RECT 72.580 330.350 72.730 338.550 ;
        RECT 73.180 330.350 73.330 338.550 ;
        RECT 73.780 330.350 73.930 338.550 ;
        RECT 70.030 329.200 70.330 329.650 ;
        RECT 66.480 329.050 70.330 329.200 ;
        RECT 70.030 328.600 70.330 329.050 ;
        RECT 66.480 328.450 70.330 328.600 ;
        RECT 70.030 328.000 70.330 328.450 ;
        RECT 66.480 327.850 70.330 328.000 ;
        RECT 70.030 327.400 70.330 327.850 ;
        RECT 66.480 327.250 70.330 327.400 ;
        RECT 70.030 326.800 70.330 327.250 ;
        RECT 59.130 326.650 62.980 326.800 ;
        RECT 66.480 326.650 70.330 326.800 ;
        RECT 59.130 326.200 59.430 326.650 ;
        RECT 70.030 326.200 70.330 326.650 ;
        RECT 59.130 326.050 62.980 326.200 ;
        RECT 66.480 326.050 70.330 326.200 ;
        RECT 59.130 325.600 59.430 326.050 ;
        RECT 70.030 325.600 70.330 326.050 ;
        RECT 59.130 325.450 62.980 325.600 ;
        RECT 66.480 325.450 70.330 325.600 ;
        RECT 59.130 325.000 59.430 325.450 ;
        RECT 70.030 325.000 70.330 325.450 ;
        RECT 59.130 324.850 62.980 325.000 ;
        RECT 66.480 324.850 70.330 325.000 ;
        RECT 59.130 324.400 59.430 324.850 ;
        RECT 70.030 324.400 70.330 324.850 ;
        RECT 59.130 324.250 62.980 324.400 ;
        RECT 66.480 324.250 70.330 324.400 ;
        RECT 59.130 323.800 59.430 324.250 ;
        RECT 70.030 323.800 70.330 324.250 ;
        RECT 59.130 323.650 62.980 323.800 ;
        RECT 66.480 323.650 70.330 323.800 ;
        RECT 59.130 323.200 59.430 323.650 ;
        RECT 70.030 323.200 70.330 323.650 ;
        RECT 59.130 323.050 62.980 323.200 ;
        RECT 66.480 323.050 70.330 323.200 ;
        RECT 59.130 322.600 59.430 323.050 ;
        RECT 70.030 322.600 70.330 323.050 ;
        RECT 59.130 322.450 62.980 322.600 ;
        RECT 66.480 322.450 70.330 322.600 ;
        RECT 59.130 322.000 59.430 322.450 ;
        RECT 70.030 322.000 70.330 322.450 ;
        RECT 59.130 321.450 62.930 322.000 ;
        RECT 46.530 321.400 62.930 321.450 ;
        RECT 66.530 321.450 70.330 322.000 ;
        RECT 70.780 321.450 70.930 329.650 ;
        RECT 71.380 321.450 71.530 329.650 ;
        RECT 71.980 321.450 72.130 329.650 ;
        RECT 72.580 321.450 72.730 329.650 ;
        RECT 73.180 321.450 73.330 329.650 ;
        RECT 73.780 321.450 73.930 329.650 ;
        RECT 74.380 321.450 75.080 338.550 ;
        RECT 75.530 330.350 75.680 338.550 ;
        RECT 76.130 330.350 76.280 338.550 ;
        RECT 76.730 330.350 76.880 338.550 ;
        RECT 77.330 330.350 77.480 338.550 ;
        RECT 77.930 330.350 78.080 338.550 ;
        RECT 78.530 330.350 78.680 338.550 ;
        RECT 79.130 338.000 82.930 338.550 ;
        RECT 86.530 338.550 102.930 338.600 ;
        RECT 86.530 338.000 90.330 338.550 ;
        RECT 79.130 337.550 79.430 338.000 ;
        RECT 90.030 337.550 90.330 338.000 ;
        RECT 79.130 337.400 82.980 337.550 ;
        RECT 86.480 337.400 90.330 337.550 ;
        RECT 79.130 336.950 79.430 337.400 ;
        RECT 90.030 336.950 90.330 337.400 ;
        RECT 79.130 336.800 82.980 336.950 ;
        RECT 86.480 336.800 90.330 336.950 ;
        RECT 79.130 336.350 79.430 336.800 ;
        RECT 90.030 336.350 90.330 336.800 ;
        RECT 79.130 336.200 82.980 336.350 ;
        RECT 86.480 336.200 90.330 336.350 ;
        RECT 79.130 335.750 79.430 336.200 ;
        RECT 90.030 335.750 90.330 336.200 ;
        RECT 79.130 335.600 82.980 335.750 ;
        RECT 86.480 335.600 90.330 335.750 ;
        RECT 79.130 335.150 79.430 335.600 ;
        RECT 90.030 335.150 90.330 335.600 ;
        RECT 79.130 335.000 82.980 335.150 ;
        RECT 86.480 335.000 90.330 335.150 ;
        RECT 79.130 334.550 79.430 335.000 ;
        RECT 90.030 334.550 90.330 335.000 ;
        RECT 79.130 334.400 82.980 334.550 ;
        RECT 86.480 334.400 90.330 334.550 ;
        RECT 79.130 333.950 79.430 334.400 ;
        RECT 90.030 333.950 90.330 334.400 ;
        RECT 79.130 333.800 82.980 333.950 ;
        RECT 86.480 333.800 90.330 333.950 ;
        RECT 79.130 333.350 79.430 333.800 ;
        RECT 90.030 333.350 90.330 333.800 ;
        RECT 79.130 333.200 82.980 333.350 ;
        RECT 86.480 333.200 90.330 333.350 ;
        RECT 79.130 332.750 79.430 333.200 ;
        RECT 79.130 332.600 82.980 332.750 ;
        RECT 79.130 332.150 79.430 332.600 ;
        RECT 79.130 332.000 82.980 332.150 ;
        RECT 79.130 331.550 79.430 332.000 ;
        RECT 79.130 331.400 82.980 331.550 ;
        RECT 79.130 330.950 79.430 331.400 ;
        RECT 79.130 330.800 82.980 330.950 ;
        RECT 79.130 330.350 79.430 330.800 ;
        RECT 75.530 321.450 75.680 329.650 ;
        RECT 76.130 321.450 76.280 329.650 ;
        RECT 76.730 321.450 76.880 329.650 ;
        RECT 77.330 321.450 77.480 329.650 ;
        RECT 77.930 321.450 78.080 329.650 ;
        RECT 78.530 321.450 78.680 329.650 ;
        RECT 79.130 329.200 79.430 329.650 ;
        RECT 79.130 329.050 82.980 329.200 ;
        RECT 79.130 328.600 79.430 329.050 ;
        RECT 79.130 328.450 82.980 328.600 ;
        RECT 79.130 328.000 79.430 328.450 ;
        RECT 79.130 327.850 82.980 328.000 ;
        RECT 79.130 327.400 79.430 327.850 ;
        RECT 79.130 327.250 82.980 327.400 ;
        RECT 79.130 326.800 79.430 327.250 ;
        RECT 83.830 326.800 85.630 333.200 ;
        RECT 90.030 332.750 90.330 333.200 ;
        RECT 86.480 332.600 90.330 332.750 ;
        RECT 90.030 332.150 90.330 332.600 ;
        RECT 86.480 332.000 90.330 332.150 ;
        RECT 90.030 331.550 90.330 332.000 ;
        RECT 86.480 331.400 90.330 331.550 ;
        RECT 90.030 330.950 90.330 331.400 ;
        RECT 86.480 330.800 90.330 330.950 ;
        RECT 90.030 330.350 90.330 330.800 ;
        RECT 90.780 330.350 90.930 338.550 ;
        RECT 91.380 330.350 91.530 338.550 ;
        RECT 91.980 330.350 92.130 338.550 ;
        RECT 92.580 330.350 92.730 338.550 ;
        RECT 93.180 330.350 93.330 338.550 ;
        RECT 93.780 330.350 93.930 338.550 ;
        RECT 90.030 329.200 90.330 329.650 ;
        RECT 86.480 329.050 90.330 329.200 ;
        RECT 90.030 328.600 90.330 329.050 ;
        RECT 86.480 328.450 90.330 328.600 ;
        RECT 90.030 328.000 90.330 328.450 ;
        RECT 86.480 327.850 90.330 328.000 ;
        RECT 90.030 327.400 90.330 327.850 ;
        RECT 86.480 327.250 90.330 327.400 ;
        RECT 90.030 326.800 90.330 327.250 ;
        RECT 79.130 326.650 82.980 326.800 ;
        RECT 86.480 326.650 90.330 326.800 ;
        RECT 79.130 326.200 79.430 326.650 ;
        RECT 90.030 326.200 90.330 326.650 ;
        RECT 79.130 326.050 82.980 326.200 ;
        RECT 86.480 326.050 90.330 326.200 ;
        RECT 79.130 325.600 79.430 326.050 ;
        RECT 90.030 325.600 90.330 326.050 ;
        RECT 79.130 325.450 82.980 325.600 ;
        RECT 86.480 325.450 90.330 325.600 ;
        RECT 79.130 325.000 79.430 325.450 ;
        RECT 90.030 325.000 90.330 325.450 ;
        RECT 79.130 324.850 82.980 325.000 ;
        RECT 86.480 324.850 90.330 325.000 ;
        RECT 79.130 324.400 79.430 324.850 ;
        RECT 90.030 324.400 90.330 324.850 ;
        RECT 79.130 324.250 82.980 324.400 ;
        RECT 86.480 324.250 90.330 324.400 ;
        RECT 79.130 323.800 79.430 324.250 ;
        RECT 90.030 323.800 90.330 324.250 ;
        RECT 79.130 323.650 82.980 323.800 ;
        RECT 86.480 323.650 90.330 323.800 ;
        RECT 79.130 323.200 79.430 323.650 ;
        RECT 90.030 323.200 90.330 323.650 ;
        RECT 79.130 323.050 82.980 323.200 ;
        RECT 86.480 323.050 90.330 323.200 ;
        RECT 79.130 322.600 79.430 323.050 ;
        RECT 90.030 322.600 90.330 323.050 ;
        RECT 79.130 322.450 82.980 322.600 ;
        RECT 86.480 322.450 90.330 322.600 ;
        RECT 79.130 322.000 79.430 322.450 ;
        RECT 90.030 322.000 90.330 322.450 ;
        RECT 79.130 321.450 82.930 322.000 ;
        RECT 66.530 321.400 82.930 321.450 ;
        RECT 86.530 321.450 90.330 322.000 ;
        RECT 90.780 321.450 90.930 329.650 ;
        RECT 91.380 321.450 91.530 329.650 ;
        RECT 91.980 321.450 92.130 329.650 ;
        RECT 92.580 321.450 92.730 329.650 ;
        RECT 93.180 321.450 93.330 329.650 ;
        RECT 93.780 321.450 93.930 329.650 ;
        RECT 94.380 321.450 95.080 338.550 ;
        RECT 95.530 330.350 95.680 338.550 ;
        RECT 96.130 330.350 96.280 338.550 ;
        RECT 96.730 330.350 96.880 338.550 ;
        RECT 97.330 330.350 97.480 338.550 ;
        RECT 97.930 330.350 98.080 338.550 ;
        RECT 98.530 330.350 98.680 338.550 ;
        RECT 99.130 338.000 102.930 338.550 ;
        RECT 106.530 338.550 122.930 338.600 ;
        RECT 106.530 338.000 110.330 338.550 ;
        RECT 99.130 337.550 99.430 338.000 ;
        RECT 110.030 337.550 110.330 338.000 ;
        RECT 99.130 337.400 102.980 337.550 ;
        RECT 106.480 337.400 110.330 337.550 ;
        RECT 99.130 336.950 99.430 337.400 ;
        RECT 110.030 336.950 110.330 337.400 ;
        RECT 99.130 336.800 102.980 336.950 ;
        RECT 106.480 336.800 110.330 336.950 ;
        RECT 99.130 336.350 99.430 336.800 ;
        RECT 110.030 336.350 110.330 336.800 ;
        RECT 99.130 336.200 102.980 336.350 ;
        RECT 106.480 336.200 110.330 336.350 ;
        RECT 99.130 335.750 99.430 336.200 ;
        RECT 110.030 335.750 110.330 336.200 ;
        RECT 99.130 335.600 102.980 335.750 ;
        RECT 106.480 335.600 110.330 335.750 ;
        RECT 99.130 335.150 99.430 335.600 ;
        RECT 110.030 335.150 110.330 335.600 ;
        RECT 99.130 335.000 102.980 335.150 ;
        RECT 106.480 335.000 110.330 335.150 ;
        RECT 99.130 334.550 99.430 335.000 ;
        RECT 110.030 334.550 110.330 335.000 ;
        RECT 99.130 334.400 102.980 334.550 ;
        RECT 106.480 334.400 110.330 334.550 ;
        RECT 99.130 333.950 99.430 334.400 ;
        RECT 110.030 333.950 110.330 334.400 ;
        RECT 99.130 333.800 102.980 333.950 ;
        RECT 106.480 333.800 110.330 333.950 ;
        RECT 99.130 333.350 99.430 333.800 ;
        RECT 110.030 333.350 110.330 333.800 ;
        RECT 99.130 333.200 102.980 333.350 ;
        RECT 106.480 333.200 110.330 333.350 ;
        RECT 99.130 332.750 99.430 333.200 ;
        RECT 99.130 332.600 102.980 332.750 ;
        RECT 99.130 332.150 99.430 332.600 ;
        RECT 99.130 332.000 102.980 332.150 ;
        RECT 99.130 331.550 99.430 332.000 ;
        RECT 99.130 331.400 102.980 331.550 ;
        RECT 99.130 330.950 99.430 331.400 ;
        RECT 99.130 330.800 102.980 330.950 ;
        RECT 99.130 330.350 99.430 330.800 ;
        RECT 95.530 321.450 95.680 329.650 ;
        RECT 96.130 321.450 96.280 329.650 ;
        RECT 96.730 321.450 96.880 329.650 ;
        RECT 97.330 321.450 97.480 329.650 ;
        RECT 97.930 321.450 98.080 329.650 ;
        RECT 98.530 321.450 98.680 329.650 ;
        RECT 99.130 329.200 99.430 329.650 ;
        RECT 99.130 329.050 102.980 329.200 ;
        RECT 99.130 328.600 99.430 329.050 ;
        RECT 99.130 328.450 102.980 328.600 ;
        RECT 99.130 328.000 99.430 328.450 ;
        RECT 99.130 327.850 102.980 328.000 ;
        RECT 99.130 327.400 99.430 327.850 ;
        RECT 99.130 327.250 102.980 327.400 ;
        RECT 99.130 326.800 99.430 327.250 ;
        RECT 103.830 326.800 105.630 333.200 ;
        RECT 110.030 332.750 110.330 333.200 ;
        RECT 106.480 332.600 110.330 332.750 ;
        RECT 110.030 332.150 110.330 332.600 ;
        RECT 106.480 332.000 110.330 332.150 ;
        RECT 110.030 331.550 110.330 332.000 ;
        RECT 106.480 331.400 110.330 331.550 ;
        RECT 110.030 330.950 110.330 331.400 ;
        RECT 106.480 330.800 110.330 330.950 ;
        RECT 110.030 330.350 110.330 330.800 ;
        RECT 110.780 330.350 110.930 338.550 ;
        RECT 111.380 330.350 111.530 338.550 ;
        RECT 111.980 330.350 112.130 338.550 ;
        RECT 112.580 330.350 112.730 338.550 ;
        RECT 113.180 330.350 113.330 338.550 ;
        RECT 113.780 330.350 113.930 338.550 ;
        RECT 110.030 329.200 110.330 329.650 ;
        RECT 106.480 329.050 110.330 329.200 ;
        RECT 110.030 328.600 110.330 329.050 ;
        RECT 106.480 328.450 110.330 328.600 ;
        RECT 110.030 328.000 110.330 328.450 ;
        RECT 106.480 327.850 110.330 328.000 ;
        RECT 110.030 327.400 110.330 327.850 ;
        RECT 106.480 327.250 110.330 327.400 ;
        RECT 110.030 326.800 110.330 327.250 ;
        RECT 99.130 326.650 102.980 326.800 ;
        RECT 106.480 326.650 110.330 326.800 ;
        RECT 99.130 326.200 99.430 326.650 ;
        RECT 110.030 326.200 110.330 326.650 ;
        RECT 99.130 326.050 102.980 326.200 ;
        RECT 106.480 326.050 110.330 326.200 ;
        RECT 99.130 325.600 99.430 326.050 ;
        RECT 110.030 325.600 110.330 326.050 ;
        RECT 99.130 325.450 102.980 325.600 ;
        RECT 106.480 325.450 110.330 325.600 ;
        RECT 99.130 325.000 99.430 325.450 ;
        RECT 110.030 325.000 110.330 325.450 ;
        RECT 99.130 324.850 102.980 325.000 ;
        RECT 106.480 324.850 110.330 325.000 ;
        RECT 99.130 324.400 99.430 324.850 ;
        RECT 110.030 324.400 110.330 324.850 ;
        RECT 99.130 324.250 102.980 324.400 ;
        RECT 106.480 324.250 110.330 324.400 ;
        RECT 99.130 323.800 99.430 324.250 ;
        RECT 110.030 323.800 110.330 324.250 ;
        RECT 99.130 323.650 102.980 323.800 ;
        RECT 106.480 323.650 110.330 323.800 ;
        RECT 99.130 323.200 99.430 323.650 ;
        RECT 110.030 323.200 110.330 323.650 ;
        RECT 99.130 323.050 102.980 323.200 ;
        RECT 106.480 323.050 110.330 323.200 ;
        RECT 99.130 322.600 99.430 323.050 ;
        RECT 110.030 322.600 110.330 323.050 ;
        RECT 99.130 322.450 102.980 322.600 ;
        RECT 106.480 322.450 110.330 322.600 ;
        RECT 99.130 322.000 99.430 322.450 ;
        RECT 110.030 322.000 110.330 322.450 ;
        RECT 99.130 321.450 102.930 322.000 ;
        RECT 86.530 321.400 102.930 321.450 ;
        RECT 106.530 321.450 110.330 322.000 ;
        RECT 110.780 321.450 110.930 329.650 ;
        RECT 111.380 321.450 111.530 329.650 ;
        RECT 111.980 321.450 112.130 329.650 ;
        RECT 112.580 321.450 112.730 329.650 ;
        RECT 113.180 321.450 113.330 329.650 ;
        RECT 113.780 321.450 113.930 329.650 ;
        RECT 114.380 321.450 115.080 338.550 ;
        RECT 115.530 330.350 115.680 338.550 ;
        RECT 116.130 330.350 116.280 338.550 ;
        RECT 116.730 330.350 116.880 338.550 ;
        RECT 117.330 330.350 117.480 338.550 ;
        RECT 117.930 330.350 118.080 338.550 ;
        RECT 118.530 330.350 118.680 338.550 ;
        RECT 119.130 338.000 122.930 338.550 ;
        RECT 119.130 337.550 119.430 338.000 ;
        RECT 119.130 337.400 122.980 337.550 ;
        RECT 119.130 336.950 119.430 337.400 ;
        RECT 119.130 336.800 122.980 336.950 ;
        RECT 119.130 336.350 119.430 336.800 ;
        RECT 119.130 336.200 122.980 336.350 ;
        RECT 119.130 335.750 119.430 336.200 ;
        RECT 119.130 335.600 122.980 335.750 ;
        RECT 119.130 335.150 119.430 335.600 ;
        RECT 119.130 335.000 122.980 335.150 ;
        RECT 119.130 334.550 119.430 335.000 ;
        RECT 119.130 334.400 122.980 334.550 ;
        RECT 119.130 333.950 119.430 334.400 ;
        RECT 119.130 333.800 122.980 333.950 ;
        RECT 119.130 333.350 119.430 333.800 ;
        RECT 119.130 333.200 122.980 333.350 ;
        RECT 119.130 332.750 119.430 333.200 ;
        RECT 119.130 332.600 122.980 332.750 ;
        RECT 119.130 332.150 119.430 332.600 ;
        RECT 119.130 332.000 122.980 332.150 ;
        RECT 119.130 331.550 119.430 332.000 ;
        RECT 119.130 331.400 122.980 331.550 ;
        RECT 119.130 330.950 119.430 331.400 ;
        RECT 119.130 330.800 122.980 330.950 ;
        RECT 119.130 330.350 119.430 330.800 ;
        RECT 115.530 321.450 115.680 329.650 ;
        RECT 116.130 321.450 116.280 329.650 ;
        RECT 116.730 321.450 116.880 329.650 ;
        RECT 117.330 321.450 117.480 329.650 ;
        RECT 117.930 321.450 118.080 329.650 ;
        RECT 118.530 321.450 118.680 329.650 ;
        RECT 119.130 329.200 119.430 329.650 ;
        RECT 119.130 329.050 122.980 329.200 ;
        RECT 119.130 328.600 119.430 329.050 ;
        RECT 119.130 328.450 122.980 328.600 ;
        RECT 119.130 328.000 119.430 328.450 ;
        RECT 119.130 327.850 122.980 328.000 ;
        RECT 119.130 327.400 119.430 327.850 ;
        RECT 119.130 327.250 122.980 327.400 ;
        RECT 119.130 326.800 119.430 327.250 ;
        RECT 123.830 326.800 124.730 333.200 ;
        RECT 129.850 329.205 131.850 330.480 ;
        RECT 119.130 326.650 122.980 326.800 ;
        RECT 119.130 326.200 119.430 326.650 ;
        RECT 119.130 326.050 122.980 326.200 ;
        RECT 119.130 325.600 119.430 326.050 ;
        RECT 119.130 325.450 122.980 325.600 ;
        RECT 119.130 325.000 119.430 325.450 ;
        RECT 119.130 324.850 122.980 325.000 ;
        RECT 119.130 324.400 119.430 324.850 ;
        RECT 119.130 324.250 122.980 324.400 ;
        RECT 119.130 323.800 119.430 324.250 ;
        RECT 119.130 323.650 122.980 323.800 ;
        RECT 119.130 323.200 119.430 323.650 ;
        RECT 119.130 323.050 122.980 323.200 ;
        RECT 119.130 322.600 119.430 323.050 ;
        RECT 119.130 322.450 122.980 322.600 ;
        RECT 119.130 322.000 119.430 322.450 ;
        RECT 119.130 321.450 122.930 322.000 ;
        RECT 106.530 321.400 122.930 321.450 ;
        RECT 9.630 320.900 19.830 321.400 ;
        RECT 29.630 320.900 39.830 321.400 ;
        RECT 49.630 320.900 59.830 321.400 ;
        RECT 69.630 320.900 79.830 321.400 ;
        RECT 89.630 320.900 99.830 321.400 ;
        RECT 109.630 320.900 119.830 321.400 ;
        RECT 11.530 319.100 17.930 320.900 ;
        RECT 31.530 319.100 37.930 320.900 ;
        RECT 51.530 319.100 57.930 320.900 ;
        RECT 71.530 319.100 77.930 320.900 ;
        RECT 91.530 319.100 97.930 320.900 ;
        RECT 111.530 319.100 117.930 320.900 ;
        RECT 9.630 318.600 19.830 319.100 ;
        RECT 29.630 318.600 39.830 319.100 ;
        RECT 49.630 318.600 59.830 319.100 ;
        RECT 69.630 318.600 79.830 319.100 ;
        RECT 89.630 318.600 99.830 319.100 ;
        RECT 109.630 318.600 119.830 319.100 ;
        RECT 6.530 318.550 22.930 318.600 ;
        RECT 6.530 318.000 10.330 318.550 ;
        RECT 10.030 317.550 10.330 318.000 ;
        RECT 6.480 317.400 10.330 317.550 ;
        RECT 10.030 316.950 10.330 317.400 ;
        RECT 6.480 316.800 10.330 316.950 ;
        RECT 10.030 316.350 10.330 316.800 ;
        RECT 6.480 316.200 10.330 316.350 ;
        RECT 10.030 315.750 10.330 316.200 ;
        RECT 6.480 315.600 10.330 315.750 ;
        RECT 10.030 315.150 10.330 315.600 ;
        RECT 6.480 315.000 10.330 315.150 ;
        RECT 10.030 314.550 10.330 315.000 ;
        RECT 6.480 314.400 10.330 314.550 ;
        RECT 10.030 313.950 10.330 314.400 ;
        RECT 6.480 313.800 10.330 313.950 ;
        RECT 10.030 313.350 10.330 313.800 ;
        RECT 6.480 313.200 10.330 313.350 ;
        RECT 4.730 306.800 5.630 313.200 ;
        RECT 10.030 312.750 10.330 313.200 ;
        RECT 6.480 312.600 10.330 312.750 ;
        RECT 10.030 312.150 10.330 312.600 ;
        RECT 6.480 312.000 10.330 312.150 ;
        RECT 10.030 311.550 10.330 312.000 ;
        RECT 6.480 311.400 10.330 311.550 ;
        RECT 10.030 310.950 10.330 311.400 ;
        RECT 6.480 310.800 10.330 310.950 ;
        RECT 10.030 310.350 10.330 310.800 ;
        RECT 10.780 310.350 10.930 318.550 ;
        RECT 11.380 310.350 11.530 318.550 ;
        RECT 11.980 310.350 12.130 318.550 ;
        RECT 12.580 310.350 12.730 318.550 ;
        RECT 13.180 310.350 13.330 318.550 ;
        RECT 13.780 310.350 13.930 318.550 ;
        RECT 10.030 309.200 10.330 309.650 ;
        RECT 6.480 309.050 10.330 309.200 ;
        RECT 10.030 308.600 10.330 309.050 ;
        RECT 6.480 308.450 10.330 308.600 ;
        RECT 10.030 308.000 10.330 308.450 ;
        RECT 6.480 307.850 10.330 308.000 ;
        RECT 10.030 307.400 10.330 307.850 ;
        RECT 6.480 307.250 10.330 307.400 ;
        RECT 10.030 306.800 10.330 307.250 ;
        RECT 6.480 306.650 10.330 306.800 ;
        RECT 10.030 306.200 10.330 306.650 ;
        RECT 6.480 306.050 10.330 306.200 ;
        RECT 10.030 305.600 10.330 306.050 ;
        RECT 6.480 305.450 10.330 305.600 ;
        RECT 10.030 305.000 10.330 305.450 ;
        RECT 6.480 304.850 10.330 305.000 ;
        RECT 10.030 304.400 10.330 304.850 ;
        RECT 6.480 304.250 10.330 304.400 ;
        RECT 10.030 303.800 10.330 304.250 ;
        RECT 6.480 303.650 10.330 303.800 ;
        RECT 10.030 303.200 10.330 303.650 ;
        RECT 6.480 303.050 10.330 303.200 ;
        RECT 10.030 302.600 10.330 303.050 ;
        RECT 6.480 302.450 10.330 302.600 ;
        RECT 10.030 302.000 10.330 302.450 ;
        RECT 6.530 301.450 10.330 302.000 ;
        RECT 10.780 301.450 10.930 309.650 ;
        RECT 11.380 301.450 11.530 309.650 ;
        RECT 11.980 301.450 12.130 309.650 ;
        RECT 12.580 301.450 12.730 309.650 ;
        RECT 13.180 301.450 13.330 309.650 ;
        RECT 13.780 301.450 13.930 309.650 ;
        RECT 14.380 301.450 15.080 318.550 ;
        RECT 15.530 310.350 15.680 318.550 ;
        RECT 16.130 310.350 16.280 318.550 ;
        RECT 16.730 310.350 16.880 318.550 ;
        RECT 17.330 310.350 17.480 318.550 ;
        RECT 17.930 310.350 18.080 318.550 ;
        RECT 18.530 310.350 18.680 318.550 ;
        RECT 19.130 318.000 22.930 318.550 ;
        RECT 26.530 318.550 42.930 318.600 ;
        RECT 26.530 318.000 30.330 318.550 ;
        RECT 19.130 317.550 19.430 318.000 ;
        RECT 30.030 317.550 30.330 318.000 ;
        RECT 19.130 317.400 22.980 317.550 ;
        RECT 26.480 317.400 30.330 317.550 ;
        RECT 19.130 316.950 19.430 317.400 ;
        RECT 30.030 316.950 30.330 317.400 ;
        RECT 19.130 316.800 22.980 316.950 ;
        RECT 26.480 316.800 30.330 316.950 ;
        RECT 19.130 316.350 19.430 316.800 ;
        RECT 30.030 316.350 30.330 316.800 ;
        RECT 19.130 316.200 22.980 316.350 ;
        RECT 26.480 316.200 30.330 316.350 ;
        RECT 19.130 315.750 19.430 316.200 ;
        RECT 30.030 315.750 30.330 316.200 ;
        RECT 19.130 315.600 22.980 315.750 ;
        RECT 26.480 315.600 30.330 315.750 ;
        RECT 19.130 315.150 19.430 315.600 ;
        RECT 30.030 315.150 30.330 315.600 ;
        RECT 19.130 315.000 22.980 315.150 ;
        RECT 26.480 315.000 30.330 315.150 ;
        RECT 19.130 314.550 19.430 315.000 ;
        RECT 30.030 314.550 30.330 315.000 ;
        RECT 19.130 314.400 22.980 314.550 ;
        RECT 26.480 314.400 30.330 314.550 ;
        RECT 19.130 313.950 19.430 314.400 ;
        RECT 30.030 313.950 30.330 314.400 ;
        RECT 19.130 313.800 22.980 313.950 ;
        RECT 26.480 313.800 30.330 313.950 ;
        RECT 19.130 313.350 19.430 313.800 ;
        RECT 30.030 313.350 30.330 313.800 ;
        RECT 19.130 313.200 22.980 313.350 ;
        RECT 26.480 313.200 30.330 313.350 ;
        RECT 19.130 312.750 19.430 313.200 ;
        RECT 19.130 312.600 22.980 312.750 ;
        RECT 19.130 312.150 19.430 312.600 ;
        RECT 19.130 312.000 22.980 312.150 ;
        RECT 19.130 311.550 19.430 312.000 ;
        RECT 19.130 311.400 22.980 311.550 ;
        RECT 19.130 310.950 19.430 311.400 ;
        RECT 19.130 310.800 22.980 310.950 ;
        RECT 19.130 310.350 19.430 310.800 ;
        RECT 15.530 301.450 15.680 309.650 ;
        RECT 16.130 301.450 16.280 309.650 ;
        RECT 16.730 301.450 16.880 309.650 ;
        RECT 17.330 301.450 17.480 309.650 ;
        RECT 17.930 301.450 18.080 309.650 ;
        RECT 18.530 301.450 18.680 309.650 ;
        RECT 19.130 309.200 19.430 309.650 ;
        RECT 19.130 309.050 22.980 309.200 ;
        RECT 19.130 308.600 19.430 309.050 ;
        RECT 19.130 308.450 22.980 308.600 ;
        RECT 19.130 308.000 19.430 308.450 ;
        RECT 19.130 307.850 22.980 308.000 ;
        RECT 19.130 307.400 19.430 307.850 ;
        RECT 19.130 307.250 22.980 307.400 ;
        RECT 19.130 306.800 19.430 307.250 ;
        RECT 23.830 306.800 25.630 313.200 ;
        RECT 30.030 312.750 30.330 313.200 ;
        RECT 26.480 312.600 30.330 312.750 ;
        RECT 30.030 312.150 30.330 312.600 ;
        RECT 26.480 312.000 30.330 312.150 ;
        RECT 30.030 311.550 30.330 312.000 ;
        RECT 26.480 311.400 30.330 311.550 ;
        RECT 30.030 310.950 30.330 311.400 ;
        RECT 26.480 310.800 30.330 310.950 ;
        RECT 30.030 310.350 30.330 310.800 ;
        RECT 30.780 310.350 30.930 318.550 ;
        RECT 31.380 310.350 31.530 318.550 ;
        RECT 31.980 310.350 32.130 318.550 ;
        RECT 32.580 310.350 32.730 318.550 ;
        RECT 33.180 310.350 33.330 318.550 ;
        RECT 33.780 310.350 33.930 318.550 ;
        RECT 30.030 309.200 30.330 309.650 ;
        RECT 26.480 309.050 30.330 309.200 ;
        RECT 30.030 308.600 30.330 309.050 ;
        RECT 26.480 308.450 30.330 308.600 ;
        RECT 30.030 308.000 30.330 308.450 ;
        RECT 26.480 307.850 30.330 308.000 ;
        RECT 30.030 307.400 30.330 307.850 ;
        RECT 26.480 307.250 30.330 307.400 ;
        RECT 30.030 306.800 30.330 307.250 ;
        RECT 19.130 306.650 22.980 306.800 ;
        RECT 26.480 306.650 30.330 306.800 ;
        RECT 19.130 306.200 19.430 306.650 ;
        RECT 30.030 306.200 30.330 306.650 ;
        RECT 19.130 306.050 22.980 306.200 ;
        RECT 26.480 306.050 30.330 306.200 ;
        RECT 19.130 305.600 19.430 306.050 ;
        RECT 30.030 305.600 30.330 306.050 ;
        RECT 19.130 305.450 22.980 305.600 ;
        RECT 26.480 305.450 30.330 305.600 ;
        RECT 19.130 305.000 19.430 305.450 ;
        RECT 30.030 305.000 30.330 305.450 ;
        RECT 19.130 304.850 22.980 305.000 ;
        RECT 26.480 304.850 30.330 305.000 ;
        RECT 19.130 304.400 19.430 304.850 ;
        RECT 30.030 304.400 30.330 304.850 ;
        RECT 19.130 304.250 22.980 304.400 ;
        RECT 26.480 304.250 30.330 304.400 ;
        RECT 19.130 303.800 19.430 304.250 ;
        RECT 30.030 303.800 30.330 304.250 ;
        RECT 19.130 303.650 22.980 303.800 ;
        RECT 26.480 303.650 30.330 303.800 ;
        RECT 19.130 303.200 19.430 303.650 ;
        RECT 30.030 303.200 30.330 303.650 ;
        RECT 19.130 303.050 22.980 303.200 ;
        RECT 26.480 303.050 30.330 303.200 ;
        RECT 19.130 302.600 19.430 303.050 ;
        RECT 30.030 302.600 30.330 303.050 ;
        RECT 19.130 302.450 22.980 302.600 ;
        RECT 26.480 302.450 30.330 302.600 ;
        RECT 19.130 302.000 19.430 302.450 ;
        RECT 30.030 302.000 30.330 302.450 ;
        RECT 19.130 301.450 22.930 302.000 ;
        RECT 6.530 301.400 22.930 301.450 ;
        RECT 26.530 301.450 30.330 302.000 ;
        RECT 30.780 301.450 30.930 309.650 ;
        RECT 31.380 301.450 31.530 309.650 ;
        RECT 31.980 301.450 32.130 309.650 ;
        RECT 32.580 301.450 32.730 309.650 ;
        RECT 33.180 301.450 33.330 309.650 ;
        RECT 33.780 301.450 33.930 309.650 ;
        RECT 34.380 301.450 35.080 318.550 ;
        RECT 35.530 310.350 35.680 318.550 ;
        RECT 36.130 310.350 36.280 318.550 ;
        RECT 36.730 310.350 36.880 318.550 ;
        RECT 37.330 310.350 37.480 318.550 ;
        RECT 37.930 310.350 38.080 318.550 ;
        RECT 38.530 310.350 38.680 318.550 ;
        RECT 39.130 318.000 42.930 318.550 ;
        RECT 46.530 318.550 62.930 318.600 ;
        RECT 46.530 318.000 50.330 318.550 ;
        RECT 39.130 317.550 39.430 318.000 ;
        RECT 50.030 317.550 50.330 318.000 ;
        RECT 39.130 317.400 42.980 317.550 ;
        RECT 46.480 317.400 50.330 317.550 ;
        RECT 39.130 316.950 39.430 317.400 ;
        RECT 50.030 316.950 50.330 317.400 ;
        RECT 39.130 316.800 42.980 316.950 ;
        RECT 46.480 316.800 50.330 316.950 ;
        RECT 39.130 316.350 39.430 316.800 ;
        RECT 50.030 316.350 50.330 316.800 ;
        RECT 39.130 316.200 42.980 316.350 ;
        RECT 46.480 316.200 50.330 316.350 ;
        RECT 39.130 315.750 39.430 316.200 ;
        RECT 50.030 315.750 50.330 316.200 ;
        RECT 39.130 315.600 42.980 315.750 ;
        RECT 46.480 315.600 50.330 315.750 ;
        RECT 39.130 315.150 39.430 315.600 ;
        RECT 50.030 315.150 50.330 315.600 ;
        RECT 39.130 315.000 42.980 315.150 ;
        RECT 46.480 315.000 50.330 315.150 ;
        RECT 39.130 314.550 39.430 315.000 ;
        RECT 50.030 314.550 50.330 315.000 ;
        RECT 39.130 314.400 42.980 314.550 ;
        RECT 46.480 314.400 50.330 314.550 ;
        RECT 39.130 313.950 39.430 314.400 ;
        RECT 50.030 313.950 50.330 314.400 ;
        RECT 39.130 313.800 42.980 313.950 ;
        RECT 46.480 313.800 50.330 313.950 ;
        RECT 39.130 313.350 39.430 313.800 ;
        RECT 50.030 313.350 50.330 313.800 ;
        RECT 39.130 313.200 42.980 313.350 ;
        RECT 46.480 313.200 50.330 313.350 ;
        RECT 39.130 312.750 39.430 313.200 ;
        RECT 39.130 312.600 42.980 312.750 ;
        RECT 39.130 312.150 39.430 312.600 ;
        RECT 39.130 312.000 42.980 312.150 ;
        RECT 39.130 311.550 39.430 312.000 ;
        RECT 39.130 311.400 42.980 311.550 ;
        RECT 39.130 310.950 39.430 311.400 ;
        RECT 39.130 310.800 42.980 310.950 ;
        RECT 39.130 310.350 39.430 310.800 ;
        RECT 35.530 301.450 35.680 309.650 ;
        RECT 36.130 301.450 36.280 309.650 ;
        RECT 36.730 301.450 36.880 309.650 ;
        RECT 37.330 301.450 37.480 309.650 ;
        RECT 37.930 301.450 38.080 309.650 ;
        RECT 38.530 301.450 38.680 309.650 ;
        RECT 39.130 309.200 39.430 309.650 ;
        RECT 39.130 309.050 42.980 309.200 ;
        RECT 39.130 308.600 39.430 309.050 ;
        RECT 39.130 308.450 42.980 308.600 ;
        RECT 39.130 308.000 39.430 308.450 ;
        RECT 39.130 307.850 42.980 308.000 ;
        RECT 39.130 307.400 39.430 307.850 ;
        RECT 39.130 307.250 42.980 307.400 ;
        RECT 39.130 306.800 39.430 307.250 ;
        RECT 43.830 306.800 45.630 313.200 ;
        RECT 50.030 312.750 50.330 313.200 ;
        RECT 46.480 312.600 50.330 312.750 ;
        RECT 50.030 312.150 50.330 312.600 ;
        RECT 46.480 312.000 50.330 312.150 ;
        RECT 50.030 311.550 50.330 312.000 ;
        RECT 46.480 311.400 50.330 311.550 ;
        RECT 50.030 310.950 50.330 311.400 ;
        RECT 46.480 310.800 50.330 310.950 ;
        RECT 50.030 310.350 50.330 310.800 ;
        RECT 50.780 310.350 50.930 318.550 ;
        RECT 51.380 310.350 51.530 318.550 ;
        RECT 51.980 310.350 52.130 318.550 ;
        RECT 52.580 310.350 52.730 318.550 ;
        RECT 53.180 310.350 53.330 318.550 ;
        RECT 53.780 310.350 53.930 318.550 ;
        RECT 50.030 309.200 50.330 309.650 ;
        RECT 46.480 309.050 50.330 309.200 ;
        RECT 50.030 308.600 50.330 309.050 ;
        RECT 46.480 308.450 50.330 308.600 ;
        RECT 50.030 308.000 50.330 308.450 ;
        RECT 46.480 307.850 50.330 308.000 ;
        RECT 50.030 307.400 50.330 307.850 ;
        RECT 46.480 307.250 50.330 307.400 ;
        RECT 50.030 306.800 50.330 307.250 ;
        RECT 39.130 306.650 42.980 306.800 ;
        RECT 46.480 306.650 50.330 306.800 ;
        RECT 39.130 306.200 39.430 306.650 ;
        RECT 50.030 306.200 50.330 306.650 ;
        RECT 39.130 306.050 42.980 306.200 ;
        RECT 46.480 306.050 50.330 306.200 ;
        RECT 39.130 305.600 39.430 306.050 ;
        RECT 50.030 305.600 50.330 306.050 ;
        RECT 39.130 305.450 42.980 305.600 ;
        RECT 46.480 305.450 50.330 305.600 ;
        RECT 39.130 305.000 39.430 305.450 ;
        RECT 50.030 305.000 50.330 305.450 ;
        RECT 39.130 304.850 42.980 305.000 ;
        RECT 46.480 304.850 50.330 305.000 ;
        RECT 39.130 304.400 39.430 304.850 ;
        RECT 50.030 304.400 50.330 304.850 ;
        RECT 39.130 304.250 42.980 304.400 ;
        RECT 46.480 304.250 50.330 304.400 ;
        RECT 39.130 303.800 39.430 304.250 ;
        RECT 50.030 303.800 50.330 304.250 ;
        RECT 39.130 303.650 42.980 303.800 ;
        RECT 46.480 303.650 50.330 303.800 ;
        RECT 39.130 303.200 39.430 303.650 ;
        RECT 50.030 303.200 50.330 303.650 ;
        RECT 39.130 303.050 42.980 303.200 ;
        RECT 46.480 303.050 50.330 303.200 ;
        RECT 39.130 302.600 39.430 303.050 ;
        RECT 50.030 302.600 50.330 303.050 ;
        RECT 39.130 302.450 42.980 302.600 ;
        RECT 46.480 302.450 50.330 302.600 ;
        RECT 39.130 302.000 39.430 302.450 ;
        RECT 50.030 302.000 50.330 302.450 ;
        RECT 39.130 301.450 42.930 302.000 ;
        RECT 26.530 301.400 42.930 301.450 ;
        RECT 46.530 301.450 50.330 302.000 ;
        RECT 50.780 301.450 50.930 309.650 ;
        RECT 51.380 301.450 51.530 309.650 ;
        RECT 51.980 301.450 52.130 309.650 ;
        RECT 52.580 301.450 52.730 309.650 ;
        RECT 53.180 301.450 53.330 309.650 ;
        RECT 53.780 301.450 53.930 309.650 ;
        RECT 54.380 301.450 55.080 318.550 ;
        RECT 55.530 310.350 55.680 318.550 ;
        RECT 56.130 310.350 56.280 318.550 ;
        RECT 56.730 310.350 56.880 318.550 ;
        RECT 57.330 310.350 57.480 318.550 ;
        RECT 57.930 310.350 58.080 318.550 ;
        RECT 58.530 310.350 58.680 318.550 ;
        RECT 59.130 318.000 62.930 318.550 ;
        RECT 66.530 318.550 82.930 318.600 ;
        RECT 66.530 318.000 70.330 318.550 ;
        RECT 59.130 317.550 59.430 318.000 ;
        RECT 70.030 317.550 70.330 318.000 ;
        RECT 59.130 317.400 62.980 317.550 ;
        RECT 66.480 317.400 70.330 317.550 ;
        RECT 59.130 316.950 59.430 317.400 ;
        RECT 70.030 316.950 70.330 317.400 ;
        RECT 59.130 316.800 62.980 316.950 ;
        RECT 66.480 316.800 70.330 316.950 ;
        RECT 59.130 316.350 59.430 316.800 ;
        RECT 70.030 316.350 70.330 316.800 ;
        RECT 59.130 316.200 62.980 316.350 ;
        RECT 66.480 316.200 70.330 316.350 ;
        RECT 59.130 315.750 59.430 316.200 ;
        RECT 70.030 315.750 70.330 316.200 ;
        RECT 59.130 315.600 62.980 315.750 ;
        RECT 66.480 315.600 70.330 315.750 ;
        RECT 59.130 315.150 59.430 315.600 ;
        RECT 70.030 315.150 70.330 315.600 ;
        RECT 59.130 315.000 62.980 315.150 ;
        RECT 66.480 315.000 70.330 315.150 ;
        RECT 59.130 314.550 59.430 315.000 ;
        RECT 70.030 314.550 70.330 315.000 ;
        RECT 59.130 314.400 62.980 314.550 ;
        RECT 66.480 314.400 70.330 314.550 ;
        RECT 59.130 313.950 59.430 314.400 ;
        RECT 70.030 313.950 70.330 314.400 ;
        RECT 59.130 313.800 62.980 313.950 ;
        RECT 66.480 313.800 70.330 313.950 ;
        RECT 59.130 313.350 59.430 313.800 ;
        RECT 70.030 313.350 70.330 313.800 ;
        RECT 59.130 313.200 62.980 313.350 ;
        RECT 66.480 313.200 70.330 313.350 ;
        RECT 59.130 312.750 59.430 313.200 ;
        RECT 59.130 312.600 62.980 312.750 ;
        RECT 59.130 312.150 59.430 312.600 ;
        RECT 59.130 312.000 62.980 312.150 ;
        RECT 59.130 311.550 59.430 312.000 ;
        RECT 59.130 311.400 62.980 311.550 ;
        RECT 59.130 310.950 59.430 311.400 ;
        RECT 59.130 310.800 62.980 310.950 ;
        RECT 59.130 310.350 59.430 310.800 ;
        RECT 55.530 301.450 55.680 309.650 ;
        RECT 56.130 301.450 56.280 309.650 ;
        RECT 56.730 301.450 56.880 309.650 ;
        RECT 57.330 301.450 57.480 309.650 ;
        RECT 57.930 301.450 58.080 309.650 ;
        RECT 58.530 301.450 58.680 309.650 ;
        RECT 59.130 309.200 59.430 309.650 ;
        RECT 59.130 309.050 62.980 309.200 ;
        RECT 59.130 308.600 59.430 309.050 ;
        RECT 59.130 308.450 62.980 308.600 ;
        RECT 59.130 308.000 59.430 308.450 ;
        RECT 59.130 307.850 62.980 308.000 ;
        RECT 59.130 307.400 59.430 307.850 ;
        RECT 59.130 307.250 62.980 307.400 ;
        RECT 59.130 306.800 59.430 307.250 ;
        RECT 63.830 306.800 65.630 313.200 ;
        RECT 70.030 312.750 70.330 313.200 ;
        RECT 66.480 312.600 70.330 312.750 ;
        RECT 70.030 312.150 70.330 312.600 ;
        RECT 66.480 312.000 70.330 312.150 ;
        RECT 70.030 311.550 70.330 312.000 ;
        RECT 66.480 311.400 70.330 311.550 ;
        RECT 70.030 310.950 70.330 311.400 ;
        RECT 66.480 310.800 70.330 310.950 ;
        RECT 70.030 310.350 70.330 310.800 ;
        RECT 70.780 310.350 70.930 318.550 ;
        RECT 71.380 310.350 71.530 318.550 ;
        RECT 71.980 310.350 72.130 318.550 ;
        RECT 72.580 310.350 72.730 318.550 ;
        RECT 73.180 310.350 73.330 318.550 ;
        RECT 73.780 310.350 73.930 318.550 ;
        RECT 70.030 309.200 70.330 309.650 ;
        RECT 66.480 309.050 70.330 309.200 ;
        RECT 70.030 308.600 70.330 309.050 ;
        RECT 66.480 308.450 70.330 308.600 ;
        RECT 70.030 308.000 70.330 308.450 ;
        RECT 66.480 307.850 70.330 308.000 ;
        RECT 70.030 307.400 70.330 307.850 ;
        RECT 66.480 307.250 70.330 307.400 ;
        RECT 70.030 306.800 70.330 307.250 ;
        RECT 59.130 306.650 62.980 306.800 ;
        RECT 66.480 306.650 70.330 306.800 ;
        RECT 59.130 306.200 59.430 306.650 ;
        RECT 70.030 306.200 70.330 306.650 ;
        RECT 59.130 306.050 62.980 306.200 ;
        RECT 66.480 306.050 70.330 306.200 ;
        RECT 59.130 305.600 59.430 306.050 ;
        RECT 70.030 305.600 70.330 306.050 ;
        RECT 59.130 305.450 62.980 305.600 ;
        RECT 66.480 305.450 70.330 305.600 ;
        RECT 59.130 305.000 59.430 305.450 ;
        RECT 70.030 305.000 70.330 305.450 ;
        RECT 59.130 304.850 62.980 305.000 ;
        RECT 66.480 304.850 70.330 305.000 ;
        RECT 59.130 304.400 59.430 304.850 ;
        RECT 70.030 304.400 70.330 304.850 ;
        RECT 59.130 304.250 62.980 304.400 ;
        RECT 66.480 304.250 70.330 304.400 ;
        RECT 59.130 303.800 59.430 304.250 ;
        RECT 70.030 303.800 70.330 304.250 ;
        RECT 59.130 303.650 62.980 303.800 ;
        RECT 66.480 303.650 70.330 303.800 ;
        RECT 59.130 303.200 59.430 303.650 ;
        RECT 70.030 303.200 70.330 303.650 ;
        RECT 59.130 303.050 62.980 303.200 ;
        RECT 66.480 303.050 70.330 303.200 ;
        RECT 59.130 302.600 59.430 303.050 ;
        RECT 70.030 302.600 70.330 303.050 ;
        RECT 59.130 302.450 62.980 302.600 ;
        RECT 66.480 302.450 70.330 302.600 ;
        RECT 59.130 302.000 59.430 302.450 ;
        RECT 70.030 302.000 70.330 302.450 ;
        RECT 59.130 301.450 62.930 302.000 ;
        RECT 46.530 301.400 62.930 301.450 ;
        RECT 66.530 301.450 70.330 302.000 ;
        RECT 70.780 301.450 70.930 309.650 ;
        RECT 71.380 301.450 71.530 309.650 ;
        RECT 71.980 301.450 72.130 309.650 ;
        RECT 72.580 301.450 72.730 309.650 ;
        RECT 73.180 301.450 73.330 309.650 ;
        RECT 73.780 301.450 73.930 309.650 ;
        RECT 74.380 301.450 75.080 318.550 ;
        RECT 75.530 310.350 75.680 318.550 ;
        RECT 76.130 310.350 76.280 318.550 ;
        RECT 76.730 310.350 76.880 318.550 ;
        RECT 77.330 310.350 77.480 318.550 ;
        RECT 77.930 310.350 78.080 318.550 ;
        RECT 78.530 310.350 78.680 318.550 ;
        RECT 79.130 318.000 82.930 318.550 ;
        RECT 86.530 318.550 102.930 318.600 ;
        RECT 86.530 318.000 90.330 318.550 ;
        RECT 79.130 317.550 79.430 318.000 ;
        RECT 90.030 317.550 90.330 318.000 ;
        RECT 79.130 317.400 82.980 317.550 ;
        RECT 86.480 317.400 90.330 317.550 ;
        RECT 79.130 316.950 79.430 317.400 ;
        RECT 90.030 316.950 90.330 317.400 ;
        RECT 79.130 316.800 82.980 316.950 ;
        RECT 86.480 316.800 90.330 316.950 ;
        RECT 79.130 316.350 79.430 316.800 ;
        RECT 90.030 316.350 90.330 316.800 ;
        RECT 79.130 316.200 82.980 316.350 ;
        RECT 86.480 316.200 90.330 316.350 ;
        RECT 79.130 315.750 79.430 316.200 ;
        RECT 90.030 315.750 90.330 316.200 ;
        RECT 79.130 315.600 82.980 315.750 ;
        RECT 86.480 315.600 90.330 315.750 ;
        RECT 79.130 315.150 79.430 315.600 ;
        RECT 90.030 315.150 90.330 315.600 ;
        RECT 79.130 315.000 82.980 315.150 ;
        RECT 86.480 315.000 90.330 315.150 ;
        RECT 79.130 314.550 79.430 315.000 ;
        RECT 90.030 314.550 90.330 315.000 ;
        RECT 79.130 314.400 82.980 314.550 ;
        RECT 86.480 314.400 90.330 314.550 ;
        RECT 79.130 313.950 79.430 314.400 ;
        RECT 90.030 313.950 90.330 314.400 ;
        RECT 79.130 313.800 82.980 313.950 ;
        RECT 86.480 313.800 90.330 313.950 ;
        RECT 79.130 313.350 79.430 313.800 ;
        RECT 90.030 313.350 90.330 313.800 ;
        RECT 79.130 313.200 82.980 313.350 ;
        RECT 86.480 313.200 90.330 313.350 ;
        RECT 79.130 312.750 79.430 313.200 ;
        RECT 79.130 312.600 82.980 312.750 ;
        RECT 79.130 312.150 79.430 312.600 ;
        RECT 79.130 312.000 82.980 312.150 ;
        RECT 79.130 311.550 79.430 312.000 ;
        RECT 79.130 311.400 82.980 311.550 ;
        RECT 79.130 310.950 79.430 311.400 ;
        RECT 79.130 310.800 82.980 310.950 ;
        RECT 79.130 310.350 79.430 310.800 ;
        RECT 75.530 301.450 75.680 309.650 ;
        RECT 76.130 301.450 76.280 309.650 ;
        RECT 76.730 301.450 76.880 309.650 ;
        RECT 77.330 301.450 77.480 309.650 ;
        RECT 77.930 301.450 78.080 309.650 ;
        RECT 78.530 301.450 78.680 309.650 ;
        RECT 79.130 309.200 79.430 309.650 ;
        RECT 79.130 309.050 82.980 309.200 ;
        RECT 79.130 308.600 79.430 309.050 ;
        RECT 79.130 308.450 82.980 308.600 ;
        RECT 79.130 308.000 79.430 308.450 ;
        RECT 79.130 307.850 82.980 308.000 ;
        RECT 79.130 307.400 79.430 307.850 ;
        RECT 79.130 307.250 82.980 307.400 ;
        RECT 79.130 306.800 79.430 307.250 ;
        RECT 83.830 306.800 85.630 313.200 ;
        RECT 90.030 312.750 90.330 313.200 ;
        RECT 86.480 312.600 90.330 312.750 ;
        RECT 90.030 312.150 90.330 312.600 ;
        RECT 86.480 312.000 90.330 312.150 ;
        RECT 90.030 311.550 90.330 312.000 ;
        RECT 86.480 311.400 90.330 311.550 ;
        RECT 90.030 310.950 90.330 311.400 ;
        RECT 86.480 310.800 90.330 310.950 ;
        RECT 90.030 310.350 90.330 310.800 ;
        RECT 90.780 310.350 90.930 318.550 ;
        RECT 91.380 310.350 91.530 318.550 ;
        RECT 91.980 310.350 92.130 318.550 ;
        RECT 92.580 310.350 92.730 318.550 ;
        RECT 93.180 310.350 93.330 318.550 ;
        RECT 93.780 310.350 93.930 318.550 ;
        RECT 90.030 309.200 90.330 309.650 ;
        RECT 86.480 309.050 90.330 309.200 ;
        RECT 90.030 308.600 90.330 309.050 ;
        RECT 86.480 308.450 90.330 308.600 ;
        RECT 90.030 308.000 90.330 308.450 ;
        RECT 86.480 307.850 90.330 308.000 ;
        RECT 90.030 307.400 90.330 307.850 ;
        RECT 86.480 307.250 90.330 307.400 ;
        RECT 90.030 306.800 90.330 307.250 ;
        RECT 79.130 306.650 82.980 306.800 ;
        RECT 86.480 306.650 90.330 306.800 ;
        RECT 79.130 306.200 79.430 306.650 ;
        RECT 90.030 306.200 90.330 306.650 ;
        RECT 79.130 306.050 82.980 306.200 ;
        RECT 86.480 306.050 90.330 306.200 ;
        RECT 79.130 305.600 79.430 306.050 ;
        RECT 90.030 305.600 90.330 306.050 ;
        RECT 79.130 305.450 82.980 305.600 ;
        RECT 86.480 305.450 90.330 305.600 ;
        RECT 79.130 305.000 79.430 305.450 ;
        RECT 90.030 305.000 90.330 305.450 ;
        RECT 79.130 304.850 82.980 305.000 ;
        RECT 86.480 304.850 90.330 305.000 ;
        RECT 79.130 304.400 79.430 304.850 ;
        RECT 90.030 304.400 90.330 304.850 ;
        RECT 79.130 304.250 82.980 304.400 ;
        RECT 86.480 304.250 90.330 304.400 ;
        RECT 79.130 303.800 79.430 304.250 ;
        RECT 90.030 303.800 90.330 304.250 ;
        RECT 79.130 303.650 82.980 303.800 ;
        RECT 86.480 303.650 90.330 303.800 ;
        RECT 79.130 303.200 79.430 303.650 ;
        RECT 90.030 303.200 90.330 303.650 ;
        RECT 79.130 303.050 82.980 303.200 ;
        RECT 86.480 303.050 90.330 303.200 ;
        RECT 79.130 302.600 79.430 303.050 ;
        RECT 90.030 302.600 90.330 303.050 ;
        RECT 79.130 302.450 82.980 302.600 ;
        RECT 86.480 302.450 90.330 302.600 ;
        RECT 79.130 302.000 79.430 302.450 ;
        RECT 90.030 302.000 90.330 302.450 ;
        RECT 79.130 301.450 82.930 302.000 ;
        RECT 66.530 301.400 82.930 301.450 ;
        RECT 86.530 301.450 90.330 302.000 ;
        RECT 90.780 301.450 90.930 309.650 ;
        RECT 91.380 301.450 91.530 309.650 ;
        RECT 91.980 301.450 92.130 309.650 ;
        RECT 92.580 301.450 92.730 309.650 ;
        RECT 93.180 301.450 93.330 309.650 ;
        RECT 93.780 301.450 93.930 309.650 ;
        RECT 94.380 301.450 95.080 318.550 ;
        RECT 95.530 310.350 95.680 318.550 ;
        RECT 96.130 310.350 96.280 318.550 ;
        RECT 96.730 310.350 96.880 318.550 ;
        RECT 97.330 310.350 97.480 318.550 ;
        RECT 97.930 310.350 98.080 318.550 ;
        RECT 98.530 310.350 98.680 318.550 ;
        RECT 99.130 318.000 102.930 318.550 ;
        RECT 106.530 318.550 122.930 318.600 ;
        RECT 106.530 318.000 110.330 318.550 ;
        RECT 99.130 317.550 99.430 318.000 ;
        RECT 110.030 317.550 110.330 318.000 ;
        RECT 99.130 317.400 102.980 317.550 ;
        RECT 106.480 317.400 110.330 317.550 ;
        RECT 99.130 316.950 99.430 317.400 ;
        RECT 110.030 316.950 110.330 317.400 ;
        RECT 99.130 316.800 102.980 316.950 ;
        RECT 106.480 316.800 110.330 316.950 ;
        RECT 99.130 316.350 99.430 316.800 ;
        RECT 110.030 316.350 110.330 316.800 ;
        RECT 99.130 316.200 102.980 316.350 ;
        RECT 106.480 316.200 110.330 316.350 ;
        RECT 99.130 315.750 99.430 316.200 ;
        RECT 110.030 315.750 110.330 316.200 ;
        RECT 99.130 315.600 102.980 315.750 ;
        RECT 106.480 315.600 110.330 315.750 ;
        RECT 99.130 315.150 99.430 315.600 ;
        RECT 110.030 315.150 110.330 315.600 ;
        RECT 99.130 315.000 102.980 315.150 ;
        RECT 106.480 315.000 110.330 315.150 ;
        RECT 99.130 314.550 99.430 315.000 ;
        RECT 110.030 314.550 110.330 315.000 ;
        RECT 99.130 314.400 102.980 314.550 ;
        RECT 106.480 314.400 110.330 314.550 ;
        RECT 99.130 313.950 99.430 314.400 ;
        RECT 110.030 313.950 110.330 314.400 ;
        RECT 99.130 313.800 102.980 313.950 ;
        RECT 106.480 313.800 110.330 313.950 ;
        RECT 99.130 313.350 99.430 313.800 ;
        RECT 110.030 313.350 110.330 313.800 ;
        RECT 99.130 313.200 102.980 313.350 ;
        RECT 106.480 313.200 110.330 313.350 ;
        RECT 99.130 312.750 99.430 313.200 ;
        RECT 99.130 312.600 102.980 312.750 ;
        RECT 99.130 312.150 99.430 312.600 ;
        RECT 99.130 312.000 102.980 312.150 ;
        RECT 99.130 311.550 99.430 312.000 ;
        RECT 99.130 311.400 102.980 311.550 ;
        RECT 99.130 310.950 99.430 311.400 ;
        RECT 99.130 310.800 102.980 310.950 ;
        RECT 99.130 310.350 99.430 310.800 ;
        RECT 95.530 301.450 95.680 309.650 ;
        RECT 96.130 301.450 96.280 309.650 ;
        RECT 96.730 301.450 96.880 309.650 ;
        RECT 97.330 301.450 97.480 309.650 ;
        RECT 97.930 301.450 98.080 309.650 ;
        RECT 98.530 301.450 98.680 309.650 ;
        RECT 99.130 309.200 99.430 309.650 ;
        RECT 99.130 309.050 102.980 309.200 ;
        RECT 99.130 308.600 99.430 309.050 ;
        RECT 99.130 308.450 102.980 308.600 ;
        RECT 99.130 308.000 99.430 308.450 ;
        RECT 99.130 307.850 102.980 308.000 ;
        RECT 99.130 307.400 99.430 307.850 ;
        RECT 99.130 307.250 102.980 307.400 ;
        RECT 99.130 306.800 99.430 307.250 ;
        RECT 103.830 306.800 105.630 313.200 ;
        RECT 110.030 312.750 110.330 313.200 ;
        RECT 106.480 312.600 110.330 312.750 ;
        RECT 110.030 312.150 110.330 312.600 ;
        RECT 106.480 312.000 110.330 312.150 ;
        RECT 110.030 311.550 110.330 312.000 ;
        RECT 106.480 311.400 110.330 311.550 ;
        RECT 110.030 310.950 110.330 311.400 ;
        RECT 106.480 310.800 110.330 310.950 ;
        RECT 110.030 310.350 110.330 310.800 ;
        RECT 110.780 310.350 110.930 318.550 ;
        RECT 111.380 310.350 111.530 318.550 ;
        RECT 111.980 310.350 112.130 318.550 ;
        RECT 112.580 310.350 112.730 318.550 ;
        RECT 113.180 310.350 113.330 318.550 ;
        RECT 113.780 310.350 113.930 318.550 ;
        RECT 110.030 309.200 110.330 309.650 ;
        RECT 106.480 309.050 110.330 309.200 ;
        RECT 110.030 308.600 110.330 309.050 ;
        RECT 106.480 308.450 110.330 308.600 ;
        RECT 110.030 308.000 110.330 308.450 ;
        RECT 106.480 307.850 110.330 308.000 ;
        RECT 110.030 307.400 110.330 307.850 ;
        RECT 106.480 307.250 110.330 307.400 ;
        RECT 110.030 306.800 110.330 307.250 ;
        RECT 99.130 306.650 102.980 306.800 ;
        RECT 106.480 306.650 110.330 306.800 ;
        RECT 99.130 306.200 99.430 306.650 ;
        RECT 110.030 306.200 110.330 306.650 ;
        RECT 99.130 306.050 102.980 306.200 ;
        RECT 106.480 306.050 110.330 306.200 ;
        RECT 99.130 305.600 99.430 306.050 ;
        RECT 110.030 305.600 110.330 306.050 ;
        RECT 99.130 305.450 102.980 305.600 ;
        RECT 106.480 305.450 110.330 305.600 ;
        RECT 99.130 305.000 99.430 305.450 ;
        RECT 110.030 305.000 110.330 305.450 ;
        RECT 99.130 304.850 102.980 305.000 ;
        RECT 106.480 304.850 110.330 305.000 ;
        RECT 99.130 304.400 99.430 304.850 ;
        RECT 110.030 304.400 110.330 304.850 ;
        RECT 99.130 304.250 102.980 304.400 ;
        RECT 106.480 304.250 110.330 304.400 ;
        RECT 99.130 303.800 99.430 304.250 ;
        RECT 110.030 303.800 110.330 304.250 ;
        RECT 99.130 303.650 102.980 303.800 ;
        RECT 106.480 303.650 110.330 303.800 ;
        RECT 99.130 303.200 99.430 303.650 ;
        RECT 110.030 303.200 110.330 303.650 ;
        RECT 99.130 303.050 102.980 303.200 ;
        RECT 106.480 303.050 110.330 303.200 ;
        RECT 99.130 302.600 99.430 303.050 ;
        RECT 110.030 302.600 110.330 303.050 ;
        RECT 99.130 302.450 102.980 302.600 ;
        RECT 106.480 302.450 110.330 302.600 ;
        RECT 99.130 302.000 99.430 302.450 ;
        RECT 110.030 302.000 110.330 302.450 ;
        RECT 99.130 301.450 102.930 302.000 ;
        RECT 86.530 301.400 102.930 301.450 ;
        RECT 106.530 301.450 110.330 302.000 ;
        RECT 110.780 301.450 110.930 309.650 ;
        RECT 111.380 301.450 111.530 309.650 ;
        RECT 111.980 301.450 112.130 309.650 ;
        RECT 112.580 301.450 112.730 309.650 ;
        RECT 113.180 301.450 113.330 309.650 ;
        RECT 113.780 301.450 113.930 309.650 ;
        RECT 114.380 301.450 115.080 318.550 ;
        RECT 115.530 310.350 115.680 318.550 ;
        RECT 116.130 310.350 116.280 318.550 ;
        RECT 116.730 310.350 116.880 318.550 ;
        RECT 117.330 310.350 117.480 318.550 ;
        RECT 117.930 310.350 118.080 318.550 ;
        RECT 118.530 310.350 118.680 318.550 ;
        RECT 119.130 318.000 122.930 318.550 ;
        RECT 119.130 317.550 119.430 318.000 ;
        RECT 119.130 317.400 122.980 317.550 ;
        RECT 119.130 316.950 119.430 317.400 ;
        RECT 119.130 316.800 122.980 316.950 ;
        RECT 119.130 316.350 119.430 316.800 ;
        RECT 119.130 316.200 122.980 316.350 ;
        RECT 119.130 315.750 119.430 316.200 ;
        RECT 119.130 315.600 122.980 315.750 ;
        RECT 119.130 315.150 119.430 315.600 ;
        RECT 119.130 315.000 122.980 315.150 ;
        RECT 119.130 314.550 119.430 315.000 ;
        RECT 119.130 314.400 122.980 314.550 ;
        RECT 119.130 313.950 119.430 314.400 ;
        RECT 119.130 313.800 122.980 313.950 ;
        RECT 119.130 313.350 119.430 313.800 ;
        RECT 119.130 313.200 122.980 313.350 ;
        RECT 119.130 312.750 119.430 313.200 ;
        RECT 119.130 312.600 122.980 312.750 ;
        RECT 119.130 312.150 119.430 312.600 ;
        RECT 119.130 312.000 122.980 312.150 ;
        RECT 119.130 311.550 119.430 312.000 ;
        RECT 119.130 311.400 122.980 311.550 ;
        RECT 119.130 310.950 119.430 311.400 ;
        RECT 119.130 310.800 122.980 310.950 ;
        RECT 119.130 310.350 119.430 310.800 ;
        RECT 115.530 301.450 115.680 309.650 ;
        RECT 116.130 301.450 116.280 309.650 ;
        RECT 116.730 301.450 116.880 309.650 ;
        RECT 117.330 301.450 117.480 309.650 ;
        RECT 117.930 301.450 118.080 309.650 ;
        RECT 118.530 301.450 118.680 309.650 ;
        RECT 119.130 309.200 119.430 309.650 ;
        RECT 119.130 309.050 122.980 309.200 ;
        RECT 119.130 308.600 119.430 309.050 ;
        RECT 119.130 308.450 122.980 308.600 ;
        RECT 119.130 308.000 119.430 308.450 ;
        RECT 119.130 307.850 122.980 308.000 ;
        RECT 119.130 307.400 119.430 307.850 ;
        RECT 119.130 307.250 122.980 307.400 ;
        RECT 119.130 306.800 119.430 307.250 ;
        RECT 123.830 306.800 124.730 313.200 ;
        RECT 129.850 309.140 131.850 310.415 ;
        RECT 119.130 306.650 122.980 306.800 ;
        RECT 119.130 306.200 119.430 306.650 ;
        RECT 119.130 306.050 122.980 306.200 ;
        RECT 119.130 305.600 119.430 306.050 ;
        RECT 119.130 305.450 122.980 305.600 ;
        RECT 119.130 305.000 119.430 305.450 ;
        RECT 119.130 304.850 122.980 305.000 ;
        RECT 119.130 304.400 119.430 304.850 ;
        RECT 119.130 304.250 122.980 304.400 ;
        RECT 119.130 303.800 119.430 304.250 ;
        RECT 119.130 303.650 122.980 303.800 ;
        RECT 119.130 303.200 119.430 303.650 ;
        RECT 119.130 303.050 122.980 303.200 ;
        RECT 119.130 302.600 119.430 303.050 ;
        RECT 119.130 302.450 122.980 302.600 ;
        RECT 119.130 302.000 119.430 302.450 ;
        RECT 119.130 301.450 122.930 302.000 ;
        RECT 106.530 301.400 122.930 301.450 ;
        RECT 9.630 300.900 19.830 301.400 ;
        RECT 29.630 300.900 39.830 301.400 ;
        RECT 49.630 300.900 59.830 301.400 ;
        RECT 69.630 300.900 79.830 301.400 ;
        RECT 89.630 300.900 99.830 301.400 ;
        RECT 109.630 300.900 119.830 301.400 ;
        RECT 11.530 299.100 17.930 300.900 ;
        RECT 31.530 299.100 37.930 300.900 ;
        RECT 51.530 299.100 57.930 300.900 ;
        RECT 71.530 299.100 77.930 300.900 ;
        RECT 91.530 299.100 97.930 300.900 ;
        RECT 111.530 299.100 117.930 300.900 ;
        RECT 9.630 298.600 19.830 299.100 ;
        RECT 29.630 298.600 39.830 299.100 ;
        RECT 49.630 298.600 59.830 299.100 ;
        RECT 69.630 298.600 79.830 299.100 ;
        RECT 89.630 298.600 99.830 299.100 ;
        RECT 109.630 298.600 119.830 299.100 ;
        RECT 6.530 298.550 22.930 298.600 ;
        RECT 6.530 298.000 10.330 298.550 ;
        RECT 10.030 297.550 10.330 298.000 ;
        RECT 6.480 297.400 10.330 297.550 ;
        RECT 10.030 296.950 10.330 297.400 ;
        RECT 6.480 296.800 10.330 296.950 ;
        RECT 10.030 296.350 10.330 296.800 ;
        RECT 6.480 296.200 10.330 296.350 ;
        RECT 10.030 295.750 10.330 296.200 ;
        RECT 6.480 295.600 10.330 295.750 ;
        RECT 10.030 295.150 10.330 295.600 ;
        RECT 6.480 295.000 10.330 295.150 ;
        RECT 10.030 294.550 10.330 295.000 ;
        RECT 6.480 294.400 10.330 294.550 ;
        RECT 10.030 293.950 10.330 294.400 ;
        RECT 6.480 293.800 10.330 293.950 ;
        RECT 10.030 293.350 10.330 293.800 ;
        RECT 6.480 293.200 10.330 293.350 ;
        RECT 4.730 286.800 5.630 293.200 ;
        RECT 10.030 292.750 10.330 293.200 ;
        RECT 6.480 292.600 10.330 292.750 ;
        RECT 10.030 292.150 10.330 292.600 ;
        RECT 6.480 292.000 10.330 292.150 ;
        RECT 10.030 291.550 10.330 292.000 ;
        RECT 6.480 291.400 10.330 291.550 ;
        RECT 10.030 290.950 10.330 291.400 ;
        RECT 6.480 290.800 10.330 290.950 ;
        RECT 10.030 290.350 10.330 290.800 ;
        RECT 10.780 290.350 10.930 298.550 ;
        RECT 11.380 290.350 11.530 298.550 ;
        RECT 11.980 290.350 12.130 298.550 ;
        RECT 12.580 290.350 12.730 298.550 ;
        RECT 13.180 290.350 13.330 298.550 ;
        RECT 13.780 290.350 13.930 298.550 ;
        RECT 10.030 289.200 10.330 289.650 ;
        RECT 6.480 289.050 10.330 289.200 ;
        RECT 10.030 288.600 10.330 289.050 ;
        RECT 6.480 288.450 10.330 288.600 ;
        RECT 10.030 288.000 10.330 288.450 ;
        RECT 6.480 287.850 10.330 288.000 ;
        RECT 10.030 287.400 10.330 287.850 ;
        RECT 6.480 287.250 10.330 287.400 ;
        RECT 10.030 286.800 10.330 287.250 ;
        RECT 6.480 286.650 10.330 286.800 ;
        RECT 10.030 286.200 10.330 286.650 ;
        RECT 6.480 286.050 10.330 286.200 ;
        RECT 10.030 285.600 10.330 286.050 ;
        RECT 6.480 285.450 10.330 285.600 ;
        RECT 10.030 285.000 10.330 285.450 ;
        RECT 6.480 284.850 10.330 285.000 ;
        RECT 10.030 284.400 10.330 284.850 ;
        RECT 6.480 284.250 10.330 284.400 ;
        RECT 10.030 283.800 10.330 284.250 ;
        RECT 6.480 283.650 10.330 283.800 ;
        RECT 10.030 283.200 10.330 283.650 ;
        RECT 6.480 283.050 10.330 283.200 ;
        RECT 10.030 282.600 10.330 283.050 ;
        RECT 6.480 282.450 10.330 282.600 ;
        RECT 10.030 282.000 10.330 282.450 ;
        RECT 6.530 281.450 10.330 282.000 ;
        RECT 10.780 281.450 10.930 289.650 ;
        RECT 11.380 281.450 11.530 289.650 ;
        RECT 11.980 281.450 12.130 289.650 ;
        RECT 12.580 281.450 12.730 289.650 ;
        RECT 13.180 281.450 13.330 289.650 ;
        RECT 13.780 281.450 13.930 289.650 ;
        RECT 14.380 281.450 15.080 298.550 ;
        RECT 15.530 290.350 15.680 298.550 ;
        RECT 16.130 290.350 16.280 298.550 ;
        RECT 16.730 290.350 16.880 298.550 ;
        RECT 17.330 290.350 17.480 298.550 ;
        RECT 17.930 290.350 18.080 298.550 ;
        RECT 18.530 290.350 18.680 298.550 ;
        RECT 19.130 298.000 22.930 298.550 ;
        RECT 26.530 298.550 42.930 298.600 ;
        RECT 26.530 298.000 30.330 298.550 ;
        RECT 19.130 297.550 19.430 298.000 ;
        RECT 30.030 297.550 30.330 298.000 ;
        RECT 19.130 297.400 22.980 297.550 ;
        RECT 26.480 297.400 30.330 297.550 ;
        RECT 19.130 296.950 19.430 297.400 ;
        RECT 30.030 296.950 30.330 297.400 ;
        RECT 19.130 296.800 22.980 296.950 ;
        RECT 26.480 296.800 30.330 296.950 ;
        RECT 19.130 296.350 19.430 296.800 ;
        RECT 30.030 296.350 30.330 296.800 ;
        RECT 19.130 296.200 22.980 296.350 ;
        RECT 26.480 296.200 30.330 296.350 ;
        RECT 19.130 295.750 19.430 296.200 ;
        RECT 30.030 295.750 30.330 296.200 ;
        RECT 19.130 295.600 22.980 295.750 ;
        RECT 26.480 295.600 30.330 295.750 ;
        RECT 19.130 295.150 19.430 295.600 ;
        RECT 30.030 295.150 30.330 295.600 ;
        RECT 19.130 295.000 22.980 295.150 ;
        RECT 26.480 295.000 30.330 295.150 ;
        RECT 19.130 294.550 19.430 295.000 ;
        RECT 30.030 294.550 30.330 295.000 ;
        RECT 19.130 294.400 22.980 294.550 ;
        RECT 26.480 294.400 30.330 294.550 ;
        RECT 19.130 293.950 19.430 294.400 ;
        RECT 30.030 293.950 30.330 294.400 ;
        RECT 19.130 293.800 22.980 293.950 ;
        RECT 26.480 293.800 30.330 293.950 ;
        RECT 19.130 293.350 19.430 293.800 ;
        RECT 30.030 293.350 30.330 293.800 ;
        RECT 19.130 293.200 22.980 293.350 ;
        RECT 26.480 293.200 30.330 293.350 ;
        RECT 19.130 292.750 19.430 293.200 ;
        RECT 19.130 292.600 22.980 292.750 ;
        RECT 19.130 292.150 19.430 292.600 ;
        RECT 19.130 292.000 22.980 292.150 ;
        RECT 19.130 291.550 19.430 292.000 ;
        RECT 19.130 291.400 22.980 291.550 ;
        RECT 19.130 290.950 19.430 291.400 ;
        RECT 19.130 290.800 22.980 290.950 ;
        RECT 19.130 290.350 19.430 290.800 ;
        RECT 15.530 281.450 15.680 289.650 ;
        RECT 16.130 281.450 16.280 289.650 ;
        RECT 16.730 281.450 16.880 289.650 ;
        RECT 17.330 281.450 17.480 289.650 ;
        RECT 17.930 281.450 18.080 289.650 ;
        RECT 18.530 281.450 18.680 289.650 ;
        RECT 19.130 289.200 19.430 289.650 ;
        RECT 19.130 289.050 22.980 289.200 ;
        RECT 19.130 288.600 19.430 289.050 ;
        RECT 19.130 288.450 22.980 288.600 ;
        RECT 19.130 288.000 19.430 288.450 ;
        RECT 19.130 287.850 22.980 288.000 ;
        RECT 19.130 287.400 19.430 287.850 ;
        RECT 19.130 287.250 22.980 287.400 ;
        RECT 19.130 286.800 19.430 287.250 ;
        RECT 23.830 286.800 25.630 293.200 ;
        RECT 30.030 292.750 30.330 293.200 ;
        RECT 26.480 292.600 30.330 292.750 ;
        RECT 30.030 292.150 30.330 292.600 ;
        RECT 26.480 292.000 30.330 292.150 ;
        RECT 30.030 291.550 30.330 292.000 ;
        RECT 26.480 291.400 30.330 291.550 ;
        RECT 30.030 290.950 30.330 291.400 ;
        RECT 26.480 290.800 30.330 290.950 ;
        RECT 30.030 290.350 30.330 290.800 ;
        RECT 30.780 290.350 30.930 298.550 ;
        RECT 31.380 290.350 31.530 298.550 ;
        RECT 31.980 290.350 32.130 298.550 ;
        RECT 32.580 290.350 32.730 298.550 ;
        RECT 33.180 290.350 33.330 298.550 ;
        RECT 33.780 290.350 33.930 298.550 ;
        RECT 30.030 289.200 30.330 289.650 ;
        RECT 26.480 289.050 30.330 289.200 ;
        RECT 30.030 288.600 30.330 289.050 ;
        RECT 26.480 288.450 30.330 288.600 ;
        RECT 30.030 288.000 30.330 288.450 ;
        RECT 26.480 287.850 30.330 288.000 ;
        RECT 30.030 287.400 30.330 287.850 ;
        RECT 26.480 287.250 30.330 287.400 ;
        RECT 30.030 286.800 30.330 287.250 ;
        RECT 19.130 286.650 22.980 286.800 ;
        RECT 26.480 286.650 30.330 286.800 ;
        RECT 19.130 286.200 19.430 286.650 ;
        RECT 30.030 286.200 30.330 286.650 ;
        RECT 19.130 286.050 22.980 286.200 ;
        RECT 26.480 286.050 30.330 286.200 ;
        RECT 19.130 285.600 19.430 286.050 ;
        RECT 30.030 285.600 30.330 286.050 ;
        RECT 19.130 285.450 22.980 285.600 ;
        RECT 26.480 285.450 30.330 285.600 ;
        RECT 19.130 285.000 19.430 285.450 ;
        RECT 30.030 285.000 30.330 285.450 ;
        RECT 19.130 284.850 22.980 285.000 ;
        RECT 26.480 284.850 30.330 285.000 ;
        RECT 19.130 284.400 19.430 284.850 ;
        RECT 30.030 284.400 30.330 284.850 ;
        RECT 19.130 284.250 22.980 284.400 ;
        RECT 26.480 284.250 30.330 284.400 ;
        RECT 19.130 283.800 19.430 284.250 ;
        RECT 30.030 283.800 30.330 284.250 ;
        RECT 19.130 283.650 22.980 283.800 ;
        RECT 26.480 283.650 30.330 283.800 ;
        RECT 19.130 283.200 19.430 283.650 ;
        RECT 30.030 283.200 30.330 283.650 ;
        RECT 19.130 283.050 22.980 283.200 ;
        RECT 26.480 283.050 30.330 283.200 ;
        RECT 19.130 282.600 19.430 283.050 ;
        RECT 30.030 282.600 30.330 283.050 ;
        RECT 19.130 282.450 22.980 282.600 ;
        RECT 26.480 282.450 30.330 282.600 ;
        RECT 19.130 282.000 19.430 282.450 ;
        RECT 30.030 282.000 30.330 282.450 ;
        RECT 19.130 281.450 22.930 282.000 ;
        RECT 6.530 281.400 22.930 281.450 ;
        RECT 26.530 281.450 30.330 282.000 ;
        RECT 30.780 281.450 30.930 289.650 ;
        RECT 31.380 281.450 31.530 289.650 ;
        RECT 31.980 281.450 32.130 289.650 ;
        RECT 32.580 281.450 32.730 289.650 ;
        RECT 33.180 281.450 33.330 289.650 ;
        RECT 33.780 281.450 33.930 289.650 ;
        RECT 34.380 281.450 35.080 298.550 ;
        RECT 35.530 290.350 35.680 298.550 ;
        RECT 36.130 290.350 36.280 298.550 ;
        RECT 36.730 290.350 36.880 298.550 ;
        RECT 37.330 290.350 37.480 298.550 ;
        RECT 37.930 290.350 38.080 298.550 ;
        RECT 38.530 290.350 38.680 298.550 ;
        RECT 39.130 298.000 42.930 298.550 ;
        RECT 46.530 298.550 62.930 298.600 ;
        RECT 46.530 298.000 50.330 298.550 ;
        RECT 39.130 297.550 39.430 298.000 ;
        RECT 50.030 297.550 50.330 298.000 ;
        RECT 39.130 297.400 42.980 297.550 ;
        RECT 46.480 297.400 50.330 297.550 ;
        RECT 39.130 296.950 39.430 297.400 ;
        RECT 50.030 296.950 50.330 297.400 ;
        RECT 39.130 296.800 42.980 296.950 ;
        RECT 46.480 296.800 50.330 296.950 ;
        RECT 39.130 296.350 39.430 296.800 ;
        RECT 50.030 296.350 50.330 296.800 ;
        RECT 39.130 296.200 42.980 296.350 ;
        RECT 46.480 296.200 50.330 296.350 ;
        RECT 39.130 295.750 39.430 296.200 ;
        RECT 50.030 295.750 50.330 296.200 ;
        RECT 39.130 295.600 42.980 295.750 ;
        RECT 46.480 295.600 50.330 295.750 ;
        RECT 39.130 295.150 39.430 295.600 ;
        RECT 50.030 295.150 50.330 295.600 ;
        RECT 39.130 295.000 42.980 295.150 ;
        RECT 46.480 295.000 50.330 295.150 ;
        RECT 39.130 294.550 39.430 295.000 ;
        RECT 50.030 294.550 50.330 295.000 ;
        RECT 39.130 294.400 42.980 294.550 ;
        RECT 46.480 294.400 50.330 294.550 ;
        RECT 39.130 293.950 39.430 294.400 ;
        RECT 50.030 293.950 50.330 294.400 ;
        RECT 39.130 293.800 42.980 293.950 ;
        RECT 46.480 293.800 50.330 293.950 ;
        RECT 39.130 293.350 39.430 293.800 ;
        RECT 50.030 293.350 50.330 293.800 ;
        RECT 39.130 293.200 42.980 293.350 ;
        RECT 46.480 293.200 50.330 293.350 ;
        RECT 39.130 292.750 39.430 293.200 ;
        RECT 39.130 292.600 42.980 292.750 ;
        RECT 39.130 292.150 39.430 292.600 ;
        RECT 39.130 292.000 42.980 292.150 ;
        RECT 39.130 291.550 39.430 292.000 ;
        RECT 39.130 291.400 42.980 291.550 ;
        RECT 39.130 290.950 39.430 291.400 ;
        RECT 39.130 290.800 42.980 290.950 ;
        RECT 39.130 290.350 39.430 290.800 ;
        RECT 35.530 281.450 35.680 289.650 ;
        RECT 36.130 281.450 36.280 289.650 ;
        RECT 36.730 281.450 36.880 289.650 ;
        RECT 37.330 281.450 37.480 289.650 ;
        RECT 37.930 281.450 38.080 289.650 ;
        RECT 38.530 281.450 38.680 289.650 ;
        RECT 39.130 289.200 39.430 289.650 ;
        RECT 39.130 289.050 42.980 289.200 ;
        RECT 39.130 288.600 39.430 289.050 ;
        RECT 39.130 288.450 42.980 288.600 ;
        RECT 39.130 288.000 39.430 288.450 ;
        RECT 39.130 287.850 42.980 288.000 ;
        RECT 39.130 287.400 39.430 287.850 ;
        RECT 39.130 287.250 42.980 287.400 ;
        RECT 39.130 286.800 39.430 287.250 ;
        RECT 43.830 286.800 45.630 293.200 ;
        RECT 50.030 292.750 50.330 293.200 ;
        RECT 46.480 292.600 50.330 292.750 ;
        RECT 50.030 292.150 50.330 292.600 ;
        RECT 46.480 292.000 50.330 292.150 ;
        RECT 50.030 291.550 50.330 292.000 ;
        RECT 46.480 291.400 50.330 291.550 ;
        RECT 50.030 290.950 50.330 291.400 ;
        RECT 46.480 290.800 50.330 290.950 ;
        RECT 50.030 290.350 50.330 290.800 ;
        RECT 50.780 290.350 50.930 298.550 ;
        RECT 51.380 290.350 51.530 298.550 ;
        RECT 51.980 290.350 52.130 298.550 ;
        RECT 52.580 290.350 52.730 298.550 ;
        RECT 53.180 290.350 53.330 298.550 ;
        RECT 53.780 290.350 53.930 298.550 ;
        RECT 50.030 289.200 50.330 289.650 ;
        RECT 46.480 289.050 50.330 289.200 ;
        RECT 50.030 288.600 50.330 289.050 ;
        RECT 46.480 288.450 50.330 288.600 ;
        RECT 50.030 288.000 50.330 288.450 ;
        RECT 46.480 287.850 50.330 288.000 ;
        RECT 50.030 287.400 50.330 287.850 ;
        RECT 46.480 287.250 50.330 287.400 ;
        RECT 50.030 286.800 50.330 287.250 ;
        RECT 39.130 286.650 42.980 286.800 ;
        RECT 46.480 286.650 50.330 286.800 ;
        RECT 39.130 286.200 39.430 286.650 ;
        RECT 50.030 286.200 50.330 286.650 ;
        RECT 39.130 286.050 42.980 286.200 ;
        RECT 46.480 286.050 50.330 286.200 ;
        RECT 39.130 285.600 39.430 286.050 ;
        RECT 50.030 285.600 50.330 286.050 ;
        RECT 39.130 285.450 42.980 285.600 ;
        RECT 46.480 285.450 50.330 285.600 ;
        RECT 39.130 285.000 39.430 285.450 ;
        RECT 50.030 285.000 50.330 285.450 ;
        RECT 39.130 284.850 42.980 285.000 ;
        RECT 46.480 284.850 50.330 285.000 ;
        RECT 39.130 284.400 39.430 284.850 ;
        RECT 50.030 284.400 50.330 284.850 ;
        RECT 39.130 284.250 42.980 284.400 ;
        RECT 46.480 284.250 50.330 284.400 ;
        RECT 39.130 283.800 39.430 284.250 ;
        RECT 50.030 283.800 50.330 284.250 ;
        RECT 39.130 283.650 42.980 283.800 ;
        RECT 46.480 283.650 50.330 283.800 ;
        RECT 39.130 283.200 39.430 283.650 ;
        RECT 50.030 283.200 50.330 283.650 ;
        RECT 39.130 283.050 42.980 283.200 ;
        RECT 46.480 283.050 50.330 283.200 ;
        RECT 39.130 282.600 39.430 283.050 ;
        RECT 50.030 282.600 50.330 283.050 ;
        RECT 39.130 282.450 42.980 282.600 ;
        RECT 46.480 282.450 50.330 282.600 ;
        RECT 39.130 282.000 39.430 282.450 ;
        RECT 50.030 282.000 50.330 282.450 ;
        RECT 39.130 281.450 42.930 282.000 ;
        RECT 26.530 281.400 42.930 281.450 ;
        RECT 46.530 281.450 50.330 282.000 ;
        RECT 50.780 281.450 50.930 289.650 ;
        RECT 51.380 281.450 51.530 289.650 ;
        RECT 51.980 281.450 52.130 289.650 ;
        RECT 52.580 281.450 52.730 289.650 ;
        RECT 53.180 281.450 53.330 289.650 ;
        RECT 53.780 281.450 53.930 289.650 ;
        RECT 54.380 281.450 55.080 298.550 ;
        RECT 55.530 290.350 55.680 298.550 ;
        RECT 56.130 290.350 56.280 298.550 ;
        RECT 56.730 290.350 56.880 298.550 ;
        RECT 57.330 290.350 57.480 298.550 ;
        RECT 57.930 290.350 58.080 298.550 ;
        RECT 58.530 290.350 58.680 298.550 ;
        RECT 59.130 298.000 62.930 298.550 ;
        RECT 66.530 298.550 82.930 298.600 ;
        RECT 66.530 298.000 70.330 298.550 ;
        RECT 59.130 297.550 59.430 298.000 ;
        RECT 70.030 297.550 70.330 298.000 ;
        RECT 59.130 297.400 62.980 297.550 ;
        RECT 66.480 297.400 70.330 297.550 ;
        RECT 59.130 296.950 59.430 297.400 ;
        RECT 70.030 296.950 70.330 297.400 ;
        RECT 59.130 296.800 62.980 296.950 ;
        RECT 66.480 296.800 70.330 296.950 ;
        RECT 59.130 296.350 59.430 296.800 ;
        RECT 70.030 296.350 70.330 296.800 ;
        RECT 59.130 296.200 62.980 296.350 ;
        RECT 66.480 296.200 70.330 296.350 ;
        RECT 59.130 295.750 59.430 296.200 ;
        RECT 70.030 295.750 70.330 296.200 ;
        RECT 59.130 295.600 62.980 295.750 ;
        RECT 66.480 295.600 70.330 295.750 ;
        RECT 59.130 295.150 59.430 295.600 ;
        RECT 70.030 295.150 70.330 295.600 ;
        RECT 59.130 295.000 62.980 295.150 ;
        RECT 66.480 295.000 70.330 295.150 ;
        RECT 59.130 294.550 59.430 295.000 ;
        RECT 70.030 294.550 70.330 295.000 ;
        RECT 59.130 294.400 62.980 294.550 ;
        RECT 66.480 294.400 70.330 294.550 ;
        RECT 59.130 293.950 59.430 294.400 ;
        RECT 70.030 293.950 70.330 294.400 ;
        RECT 59.130 293.800 62.980 293.950 ;
        RECT 66.480 293.800 70.330 293.950 ;
        RECT 59.130 293.350 59.430 293.800 ;
        RECT 70.030 293.350 70.330 293.800 ;
        RECT 59.130 293.200 62.980 293.350 ;
        RECT 66.480 293.200 70.330 293.350 ;
        RECT 59.130 292.750 59.430 293.200 ;
        RECT 59.130 292.600 62.980 292.750 ;
        RECT 59.130 292.150 59.430 292.600 ;
        RECT 59.130 292.000 62.980 292.150 ;
        RECT 59.130 291.550 59.430 292.000 ;
        RECT 59.130 291.400 62.980 291.550 ;
        RECT 59.130 290.950 59.430 291.400 ;
        RECT 59.130 290.800 62.980 290.950 ;
        RECT 59.130 290.350 59.430 290.800 ;
        RECT 55.530 281.450 55.680 289.650 ;
        RECT 56.130 281.450 56.280 289.650 ;
        RECT 56.730 281.450 56.880 289.650 ;
        RECT 57.330 281.450 57.480 289.650 ;
        RECT 57.930 281.450 58.080 289.650 ;
        RECT 58.530 281.450 58.680 289.650 ;
        RECT 59.130 289.200 59.430 289.650 ;
        RECT 59.130 289.050 62.980 289.200 ;
        RECT 59.130 288.600 59.430 289.050 ;
        RECT 59.130 288.450 62.980 288.600 ;
        RECT 59.130 288.000 59.430 288.450 ;
        RECT 59.130 287.850 62.980 288.000 ;
        RECT 59.130 287.400 59.430 287.850 ;
        RECT 59.130 287.250 62.980 287.400 ;
        RECT 59.130 286.800 59.430 287.250 ;
        RECT 63.830 286.800 65.630 293.200 ;
        RECT 70.030 292.750 70.330 293.200 ;
        RECT 66.480 292.600 70.330 292.750 ;
        RECT 70.030 292.150 70.330 292.600 ;
        RECT 66.480 292.000 70.330 292.150 ;
        RECT 70.030 291.550 70.330 292.000 ;
        RECT 66.480 291.400 70.330 291.550 ;
        RECT 70.030 290.950 70.330 291.400 ;
        RECT 66.480 290.800 70.330 290.950 ;
        RECT 70.030 290.350 70.330 290.800 ;
        RECT 70.780 290.350 70.930 298.550 ;
        RECT 71.380 290.350 71.530 298.550 ;
        RECT 71.980 290.350 72.130 298.550 ;
        RECT 72.580 290.350 72.730 298.550 ;
        RECT 73.180 290.350 73.330 298.550 ;
        RECT 73.780 290.350 73.930 298.550 ;
        RECT 70.030 289.200 70.330 289.650 ;
        RECT 66.480 289.050 70.330 289.200 ;
        RECT 70.030 288.600 70.330 289.050 ;
        RECT 66.480 288.450 70.330 288.600 ;
        RECT 70.030 288.000 70.330 288.450 ;
        RECT 66.480 287.850 70.330 288.000 ;
        RECT 70.030 287.400 70.330 287.850 ;
        RECT 66.480 287.250 70.330 287.400 ;
        RECT 70.030 286.800 70.330 287.250 ;
        RECT 59.130 286.650 62.980 286.800 ;
        RECT 66.480 286.650 70.330 286.800 ;
        RECT 59.130 286.200 59.430 286.650 ;
        RECT 70.030 286.200 70.330 286.650 ;
        RECT 59.130 286.050 62.980 286.200 ;
        RECT 66.480 286.050 70.330 286.200 ;
        RECT 59.130 285.600 59.430 286.050 ;
        RECT 70.030 285.600 70.330 286.050 ;
        RECT 59.130 285.450 62.980 285.600 ;
        RECT 66.480 285.450 70.330 285.600 ;
        RECT 59.130 285.000 59.430 285.450 ;
        RECT 70.030 285.000 70.330 285.450 ;
        RECT 59.130 284.850 62.980 285.000 ;
        RECT 66.480 284.850 70.330 285.000 ;
        RECT 59.130 284.400 59.430 284.850 ;
        RECT 70.030 284.400 70.330 284.850 ;
        RECT 59.130 284.250 62.980 284.400 ;
        RECT 66.480 284.250 70.330 284.400 ;
        RECT 59.130 283.800 59.430 284.250 ;
        RECT 70.030 283.800 70.330 284.250 ;
        RECT 59.130 283.650 62.980 283.800 ;
        RECT 66.480 283.650 70.330 283.800 ;
        RECT 59.130 283.200 59.430 283.650 ;
        RECT 70.030 283.200 70.330 283.650 ;
        RECT 59.130 283.050 62.980 283.200 ;
        RECT 66.480 283.050 70.330 283.200 ;
        RECT 59.130 282.600 59.430 283.050 ;
        RECT 70.030 282.600 70.330 283.050 ;
        RECT 59.130 282.450 62.980 282.600 ;
        RECT 66.480 282.450 70.330 282.600 ;
        RECT 59.130 282.000 59.430 282.450 ;
        RECT 70.030 282.000 70.330 282.450 ;
        RECT 59.130 281.450 62.930 282.000 ;
        RECT 46.530 281.400 62.930 281.450 ;
        RECT 66.530 281.450 70.330 282.000 ;
        RECT 70.780 281.450 70.930 289.650 ;
        RECT 71.380 281.450 71.530 289.650 ;
        RECT 71.980 281.450 72.130 289.650 ;
        RECT 72.580 281.450 72.730 289.650 ;
        RECT 73.180 281.450 73.330 289.650 ;
        RECT 73.780 281.450 73.930 289.650 ;
        RECT 74.380 281.450 75.080 298.550 ;
        RECT 75.530 290.350 75.680 298.550 ;
        RECT 76.130 290.350 76.280 298.550 ;
        RECT 76.730 290.350 76.880 298.550 ;
        RECT 77.330 290.350 77.480 298.550 ;
        RECT 77.930 290.350 78.080 298.550 ;
        RECT 78.530 290.350 78.680 298.550 ;
        RECT 79.130 298.000 82.930 298.550 ;
        RECT 86.530 298.550 102.930 298.600 ;
        RECT 86.530 298.000 90.330 298.550 ;
        RECT 79.130 297.550 79.430 298.000 ;
        RECT 90.030 297.550 90.330 298.000 ;
        RECT 79.130 297.400 82.980 297.550 ;
        RECT 86.480 297.400 90.330 297.550 ;
        RECT 79.130 296.950 79.430 297.400 ;
        RECT 90.030 296.950 90.330 297.400 ;
        RECT 79.130 296.800 82.980 296.950 ;
        RECT 86.480 296.800 90.330 296.950 ;
        RECT 79.130 296.350 79.430 296.800 ;
        RECT 90.030 296.350 90.330 296.800 ;
        RECT 79.130 296.200 82.980 296.350 ;
        RECT 86.480 296.200 90.330 296.350 ;
        RECT 79.130 295.750 79.430 296.200 ;
        RECT 90.030 295.750 90.330 296.200 ;
        RECT 79.130 295.600 82.980 295.750 ;
        RECT 86.480 295.600 90.330 295.750 ;
        RECT 79.130 295.150 79.430 295.600 ;
        RECT 90.030 295.150 90.330 295.600 ;
        RECT 79.130 295.000 82.980 295.150 ;
        RECT 86.480 295.000 90.330 295.150 ;
        RECT 79.130 294.550 79.430 295.000 ;
        RECT 90.030 294.550 90.330 295.000 ;
        RECT 79.130 294.400 82.980 294.550 ;
        RECT 86.480 294.400 90.330 294.550 ;
        RECT 79.130 293.950 79.430 294.400 ;
        RECT 90.030 293.950 90.330 294.400 ;
        RECT 79.130 293.800 82.980 293.950 ;
        RECT 86.480 293.800 90.330 293.950 ;
        RECT 79.130 293.350 79.430 293.800 ;
        RECT 90.030 293.350 90.330 293.800 ;
        RECT 79.130 293.200 82.980 293.350 ;
        RECT 86.480 293.200 90.330 293.350 ;
        RECT 79.130 292.750 79.430 293.200 ;
        RECT 79.130 292.600 82.980 292.750 ;
        RECT 79.130 292.150 79.430 292.600 ;
        RECT 79.130 292.000 82.980 292.150 ;
        RECT 79.130 291.550 79.430 292.000 ;
        RECT 79.130 291.400 82.980 291.550 ;
        RECT 79.130 290.950 79.430 291.400 ;
        RECT 79.130 290.800 82.980 290.950 ;
        RECT 79.130 290.350 79.430 290.800 ;
        RECT 75.530 281.450 75.680 289.650 ;
        RECT 76.130 281.450 76.280 289.650 ;
        RECT 76.730 281.450 76.880 289.650 ;
        RECT 77.330 281.450 77.480 289.650 ;
        RECT 77.930 281.450 78.080 289.650 ;
        RECT 78.530 281.450 78.680 289.650 ;
        RECT 79.130 289.200 79.430 289.650 ;
        RECT 79.130 289.050 82.980 289.200 ;
        RECT 79.130 288.600 79.430 289.050 ;
        RECT 79.130 288.450 82.980 288.600 ;
        RECT 79.130 288.000 79.430 288.450 ;
        RECT 79.130 287.850 82.980 288.000 ;
        RECT 79.130 287.400 79.430 287.850 ;
        RECT 79.130 287.250 82.980 287.400 ;
        RECT 79.130 286.800 79.430 287.250 ;
        RECT 83.830 286.800 85.630 293.200 ;
        RECT 90.030 292.750 90.330 293.200 ;
        RECT 86.480 292.600 90.330 292.750 ;
        RECT 90.030 292.150 90.330 292.600 ;
        RECT 86.480 292.000 90.330 292.150 ;
        RECT 90.030 291.550 90.330 292.000 ;
        RECT 86.480 291.400 90.330 291.550 ;
        RECT 90.030 290.950 90.330 291.400 ;
        RECT 86.480 290.800 90.330 290.950 ;
        RECT 90.030 290.350 90.330 290.800 ;
        RECT 90.780 290.350 90.930 298.550 ;
        RECT 91.380 290.350 91.530 298.550 ;
        RECT 91.980 290.350 92.130 298.550 ;
        RECT 92.580 290.350 92.730 298.550 ;
        RECT 93.180 290.350 93.330 298.550 ;
        RECT 93.780 290.350 93.930 298.550 ;
        RECT 90.030 289.200 90.330 289.650 ;
        RECT 86.480 289.050 90.330 289.200 ;
        RECT 90.030 288.600 90.330 289.050 ;
        RECT 86.480 288.450 90.330 288.600 ;
        RECT 90.030 288.000 90.330 288.450 ;
        RECT 86.480 287.850 90.330 288.000 ;
        RECT 90.030 287.400 90.330 287.850 ;
        RECT 86.480 287.250 90.330 287.400 ;
        RECT 90.030 286.800 90.330 287.250 ;
        RECT 79.130 286.650 82.980 286.800 ;
        RECT 86.480 286.650 90.330 286.800 ;
        RECT 79.130 286.200 79.430 286.650 ;
        RECT 90.030 286.200 90.330 286.650 ;
        RECT 79.130 286.050 82.980 286.200 ;
        RECT 86.480 286.050 90.330 286.200 ;
        RECT 79.130 285.600 79.430 286.050 ;
        RECT 90.030 285.600 90.330 286.050 ;
        RECT 79.130 285.450 82.980 285.600 ;
        RECT 86.480 285.450 90.330 285.600 ;
        RECT 79.130 285.000 79.430 285.450 ;
        RECT 90.030 285.000 90.330 285.450 ;
        RECT 79.130 284.850 82.980 285.000 ;
        RECT 86.480 284.850 90.330 285.000 ;
        RECT 79.130 284.400 79.430 284.850 ;
        RECT 90.030 284.400 90.330 284.850 ;
        RECT 79.130 284.250 82.980 284.400 ;
        RECT 86.480 284.250 90.330 284.400 ;
        RECT 79.130 283.800 79.430 284.250 ;
        RECT 90.030 283.800 90.330 284.250 ;
        RECT 79.130 283.650 82.980 283.800 ;
        RECT 86.480 283.650 90.330 283.800 ;
        RECT 79.130 283.200 79.430 283.650 ;
        RECT 90.030 283.200 90.330 283.650 ;
        RECT 79.130 283.050 82.980 283.200 ;
        RECT 86.480 283.050 90.330 283.200 ;
        RECT 79.130 282.600 79.430 283.050 ;
        RECT 90.030 282.600 90.330 283.050 ;
        RECT 79.130 282.450 82.980 282.600 ;
        RECT 86.480 282.450 90.330 282.600 ;
        RECT 79.130 282.000 79.430 282.450 ;
        RECT 90.030 282.000 90.330 282.450 ;
        RECT 79.130 281.450 82.930 282.000 ;
        RECT 66.530 281.400 82.930 281.450 ;
        RECT 86.530 281.450 90.330 282.000 ;
        RECT 90.780 281.450 90.930 289.650 ;
        RECT 91.380 281.450 91.530 289.650 ;
        RECT 91.980 281.450 92.130 289.650 ;
        RECT 92.580 281.450 92.730 289.650 ;
        RECT 93.180 281.450 93.330 289.650 ;
        RECT 93.780 281.450 93.930 289.650 ;
        RECT 94.380 281.450 95.080 298.550 ;
        RECT 95.530 290.350 95.680 298.550 ;
        RECT 96.130 290.350 96.280 298.550 ;
        RECT 96.730 290.350 96.880 298.550 ;
        RECT 97.330 290.350 97.480 298.550 ;
        RECT 97.930 290.350 98.080 298.550 ;
        RECT 98.530 290.350 98.680 298.550 ;
        RECT 99.130 298.000 102.930 298.550 ;
        RECT 106.530 298.550 122.930 298.600 ;
        RECT 106.530 298.000 110.330 298.550 ;
        RECT 99.130 297.550 99.430 298.000 ;
        RECT 110.030 297.550 110.330 298.000 ;
        RECT 99.130 297.400 102.980 297.550 ;
        RECT 106.480 297.400 110.330 297.550 ;
        RECT 99.130 296.950 99.430 297.400 ;
        RECT 110.030 296.950 110.330 297.400 ;
        RECT 99.130 296.800 102.980 296.950 ;
        RECT 106.480 296.800 110.330 296.950 ;
        RECT 99.130 296.350 99.430 296.800 ;
        RECT 110.030 296.350 110.330 296.800 ;
        RECT 99.130 296.200 102.980 296.350 ;
        RECT 106.480 296.200 110.330 296.350 ;
        RECT 99.130 295.750 99.430 296.200 ;
        RECT 110.030 295.750 110.330 296.200 ;
        RECT 99.130 295.600 102.980 295.750 ;
        RECT 106.480 295.600 110.330 295.750 ;
        RECT 99.130 295.150 99.430 295.600 ;
        RECT 110.030 295.150 110.330 295.600 ;
        RECT 99.130 295.000 102.980 295.150 ;
        RECT 106.480 295.000 110.330 295.150 ;
        RECT 99.130 294.550 99.430 295.000 ;
        RECT 110.030 294.550 110.330 295.000 ;
        RECT 99.130 294.400 102.980 294.550 ;
        RECT 106.480 294.400 110.330 294.550 ;
        RECT 99.130 293.950 99.430 294.400 ;
        RECT 110.030 293.950 110.330 294.400 ;
        RECT 99.130 293.800 102.980 293.950 ;
        RECT 106.480 293.800 110.330 293.950 ;
        RECT 99.130 293.350 99.430 293.800 ;
        RECT 110.030 293.350 110.330 293.800 ;
        RECT 99.130 293.200 102.980 293.350 ;
        RECT 106.480 293.200 110.330 293.350 ;
        RECT 99.130 292.750 99.430 293.200 ;
        RECT 99.130 292.600 102.980 292.750 ;
        RECT 99.130 292.150 99.430 292.600 ;
        RECT 99.130 292.000 102.980 292.150 ;
        RECT 99.130 291.550 99.430 292.000 ;
        RECT 99.130 291.400 102.980 291.550 ;
        RECT 99.130 290.950 99.430 291.400 ;
        RECT 99.130 290.800 102.980 290.950 ;
        RECT 99.130 290.350 99.430 290.800 ;
        RECT 95.530 281.450 95.680 289.650 ;
        RECT 96.130 281.450 96.280 289.650 ;
        RECT 96.730 281.450 96.880 289.650 ;
        RECT 97.330 281.450 97.480 289.650 ;
        RECT 97.930 281.450 98.080 289.650 ;
        RECT 98.530 281.450 98.680 289.650 ;
        RECT 99.130 289.200 99.430 289.650 ;
        RECT 99.130 289.050 102.980 289.200 ;
        RECT 99.130 288.600 99.430 289.050 ;
        RECT 99.130 288.450 102.980 288.600 ;
        RECT 99.130 288.000 99.430 288.450 ;
        RECT 99.130 287.850 102.980 288.000 ;
        RECT 99.130 287.400 99.430 287.850 ;
        RECT 99.130 287.250 102.980 287.400 ;
        RECT 99.130 286.800 99.430 287.250 ;
        RECT 103.830 286.800 105.630 293.200 ;
        RECT 110.030 292.750 110.330 293.200 ;
        RECT 106.480 292.600 110.330 292.750 ;
        RECT 110.030 292.150 110.330 292.600 ;
        RECT 106.480 292.000 110.330 292.150 ;
        RECT 110.030 291.550 110.330 292.000 ;
        RECT 106.480 291.400 110.330 291.550 ;
        RECT 110.030 290.950 110.330 291.400 ;
        RECT 106.480 290.800 110.330 290.950 ;
        RECT 110.030 290.350 110.330 290.800 ;
        RECT 110.780 290.350 110.930 298.550 ;
        RECT 111.380 290.350 111.530 298.550 ;
        RECT 111.980 290.350 112.130 298.550 ;
        RECT 112.580 290.350 112.730 298.550 ;
        RECT 113.180 290.350 113.330 298.550 ;
        RECT 113.780 290.350 113.930 298.550 ;
        RECT 110.030 289.200 110.330 289.650 ;
        RECT 106.480 289.050 110.330 289.200 ;
        RECT 110.030 288.600 110.330 289.050 ;
        RECT 106.480 288.450 110.330 288.600 ;
        RECT 110.030 288.000 110.330 288.450 ;
        RECT 106.480 287.850 110.330 288.000 ;
        RECT 110.030 287.400 110.330 287.850 ;
        RECT 106.480 287.250 110.330 287.400 ;
        RECT 110.030 286.800 110.330 287.250 ;
        RECT 99.130 286.650 102.980 286.800 ;
        RECT 106.480 286.650 110.330 286.800 ;
        RECT 99.130 286.200 99.430 286.650 ;
        RECT 110.030 286.200 110.330 286.650 ;
        RECT 99.130 286.050 102.980 286.200 ;
        RECT 106.480 286.050 110.330 286.200 ;
        RECT 99.130 285.600 99.430 286.050 ;
        RECT 110.030 285.600 110.330 286.050 ;
        RECT 99.130 285.450 102.980 285.600 ;
        RECT 106.480 285.450 110.330 285.600 ;
        RECT 99.130 285.000 99.430 285.450 ;
        RECT 110.030 285.000 110.330 285.450 ;
        RECT 99.130 284.850 102.980 285.000 ;
        RECT 106.480 284.850 110.330 285.000 ;
        RECT 99.130 284.400 99.430 284.850 ;
        RECT 110.030 284.400 110.330 284.850 ;
        RECT 99.130 284.250 102.980 284.400 ;
        RECT 106.480 284.250 110.330 284.400 ;
        RECT 99.130 283.800 99.430 284.250 ;
        RECT 110.030 283.800 110.330 284.250 ;
        RECT 99.130 283.650 102.980 283.800 ;
        RECT 106.480 283.650 110.330 283.800 ;
        RECT 99.130 283.200 99.430 283.650 ;
        RECT 110.030 283.200 110.330 283.650 ;
        RECT 99.130 283.050 102.980 283.200 ;
        RECT 106.480 283.050 110.330 283.200 ;
        RECT 99.130 282.600 99.430 283.050 ;
        RECT 110.030 282.600 110.330 283.050 ;
        RECT 99.130 282.450 102.980 282.600 ;
        RECT 106.480 282.450 110.330 282.600 ;
        RECT 99.130 282.000 99.430 282.450 ;
        RECT 110.030 282.000 110.330 282.450 ;
        RECT 99.130 281.450 102.930 282.000 ;
        RECT 86.530 281.400 102.930 281.450 ;
        RECT 106.530 281.450 110.330 282.000 ;
        RECT 110.780 281.450 110.930 289.650 ;
        RECT 111.380 281.450 111.530 289.650 ;
        RECT 111.980 281.450 112.130 289.650 ;
        RECT 112.580 281.450 112.730 289.650 ;
        RECT 113.180 281.450 113.330 289.650 ;
        RECT 113.780 281.450 113.930 289.650 ;
        RECT 114.380 281.450 115.080 298.550 ;
        RECT 115.530 290.350 115.680 298.550 ;
        RECT 116.130 290.350 116.280 298.550 ;
        RECT 116.730 290.350 116.880 298.550 ;
        RECT 117.330 290.350 117.480 298.550 ;
        RECT 117.930 290.350 118.080 298.550 ;
        RECT 118.530 290.350 118.680 298.550 ;
        RECT 119.130 298.000 122.930 298.550 ;
        RECT 119.130 297.550 119.430 298.000 ;
        RECT 119.130 297.400 122.980 297.550 ;
        RECT 119.130 296.950 119.430 297.400 ;
        RECT 119.130 296.800 122.980 296.950 ;
        RECT 119.130 296.350 119.430 296.800 ;
        RECT 119.130 296.200 122.980 296.350 ;
        RECT 119.130 295.750 119.430 296.200 ;
        RECT 119.130 295.600 122.980 295.750 ;
        RECT 119.130 295.150 119.430 295.600 ;
        RECT 119.130 295.000 122.980 295.150 ;
        RECT 119.130 294.550 119.430 295.000 ;
        RECT 119.130 294.400 122.980 294.550 ;
        RECT 119.130 293.950 119.430 294.400 ;
        RECT 119.130 293.800 122.980 293.950 ;
        RECT 119.130 293.350 119.430 293.800 ;
        RECT 119.130 293.200 122.980 293.350 ;
        RECT 119.130 292.750 119.430 293.200 ;
        RECT 119.130 292.600 122.980 292.750 ;
        RECT 119.130 292.150 119.430 292.600 ;
        RECT 119.130 292.000 122.980 292.150 ;
        RECT 119.130 291.550 119.430 292.000 ;
        RECT 119.130 291.400 122.980 291.550 ;
        RECT 119.130 290.950 119.430 291.400 ;
        RECT 119.130 290.800 122.980 290.950 ;
        RECT 119.130 290.350 119.430 290.800 ;
        RECT 115.530 281.450 115.680 289.650 ;
        RECT 116.130 281.450 116.280 289.650 ;
        RECT 116.730 281.450 116.880 289.650 ;
        RECT 117.330 281.450 117.480 289.650 ;
        RECT 117.930 281.450 118.080 289.650 ;
        RECT 118.530 281.450 118.680 289.650 ;
        RECT 119.130 289.200 119.430 289.650 ;
        RECT 119.130 289.050 122.980 289.200 ;
        RECT 119.130 288.600 119.430 289.050 ;
        RECT 119.130 288.450 122.980 288.600 ;
        RECT 119.130 288.000 119.430 288.450 ;
        RECT 119.130 287.850 122.980 288.000 ;
        RECT 119.130 287.400 119.430 287.850 ;
        RECT 119.130 287.250 122.980 287.400 ;
        RECT 119.130 286.800 119.430 287.250 ;
        RECT 123.830 286.800 124.730 293.200 ;
        RECT 129.850 289.135 131.850 290.410 ;
        RECT 119.130 286.650 122.980 286.800 ;
        RECT 119.130 286.200 119.430 286.650 ;
        RECT 119.130 286.050 122.980 286.200 ;
        RECT 119.130 285.600 119.430 286.050 ;
        RECT 119.130 285.450 122.980 285.600 ;
        RECT 119.130 285.000 119.430 285.450 ;
        RECT 119.130 284.850 122.980 285.000 ;
        RECT 119.130 284.400 119.430 284.850 ;
        RECT 119.130 284.250 122.980 284.400 ;
        RECT 119.130 283.800 119.430 284.250 ;
        RECT 119.130 283.650 122.980 283.800 ;
        RECT 119.130 283.200 119.430 283.650 ;
        RECT 119.130 283.050 122.980 283.200 ;
        RECT 119.130 282.600 119.430 283.050 ;
        RECT 119.130 282.450 122.980 282.600 ;
        RECT 119.130 282.000 119.430 282.450 ;
        RECT 119.130 281.450 122.930 282.000 ;
        RECT 106.530 281.400 122.930 281.450 ;
        RECT 9.630 280.900 19.830 281.400 ;
        RECT 29.630 280.900 39.830 281.400 ;
        RECT 49.630 280.900 59.830 281.400 ;
        RECT 69.630 280.900 79.830 281.400 ;
        RECT 89.630 280.900 99.830 281.400 ;
        RECT 109.630 280.900 119.830 281.400 ;
        RECT 11.530 279.100 17.930 280.900 ;
        RECT 31.530 279.100 37.930 280.900 ;
        RECT 51.530 279.100 57.930 280.900 ;
        RECT 71.530 279.100 77.930 280.900 ;
        RECT 91.530 279.100 97.930 280.900 ;
        RECT 111.530 279.100 117.930 280.900 ;
        RECT 9.630 278.600 19.830 279.100 ;
        RECT 29.630 278.600 39.830 279.100 ;
        RECT 49.630 278.600 59.830 279.100 ;
        RECT 69.630 278.600 79.830 279.100 ;
        RECT 89.630 278.600 99.830 279.100 ;
        RECT 109.630 278.600 119.830 279.100 ;
        RECT 6.530 278.550 22.930 278.600 ;
        RECT 6.530 278.000 10.330 278.550 ;
        RECT 10.030 277.550 10.330 278.000 ;
        RECT 6.480 277.400 10.330 277.550 ;
        RECT 10.030 276.950 10.330 277.400 ;
        RECT 6.480 276.800 10.330 276.950 ;
        RECT 10.030 276.350 10.330 276.800 ;
        RECT 6.480 276.200 10.330 276.350 ;
        RECT 10.030 275.750 10.330 276.200 ;
        RECT 6.480 275.600 10.330 275.750 ;
        RECT 10.030 275.150 10.330 275.600 ;
        RECT 6.480 275.000 10.330 275.150 ;
        RECT 10.030 274.550 10.330 275.000 ;
        RECT 6.480 274.400 10.330 274.550 ;
        RECT 10.030 273.950 10.330 274.400 ;
        RECT 6.480 273.800 10.330 273.950 ;
        RECT 10.030 273.350 10.330 273.800 ;
        RECT 6.480 273.200 10.330 273.350 ;
        RECT 4.730 266.800 5.630 273.200 ;
        RECT 10.030 272.750 10.330 273.200 ;
        RECT 6.480 272.600 10.330 272.750 ;
        RECT 10.030 272.150 10.330 272.600 ;
        RECT 6.480 272.000 10.330 272.150 ;
        RECT 10.030 271.550 10.330 272.000 ;
        RECT 6.480 271.400 10.330 271.550 ;
        RECT 10.030 270.950 10.330 271.400 ;
        RECT 6.480 270.800 10.330 270.950 ;
        RECT 10.030 270.350 10.330 270.800 ;
        RECT 10.780 270.350 10.930 278.550 ;
        RECT 11.380 270.350 11.530 278.550 ;
        RECT 11.980 270.350 12.130 278.550 ;
        RECT 12.580 270.350 12.730 278.550 ;
        RECT 13.180 270.350 13.330 278.550 ;
        RECT 13.780 270.350 13.930 278.550 ;
        RECT 10.030 269.200 10.330 269.650 ;
        RECT 6.480 269.050 10.330 269.200 ;
        RECT 10.030 268.600 10.330 269.050 ;
        RECT 6.480 268.450 10.330 268.600 ;
        RECT 10.030 268.000 10.330 268.450 ;
        RECT 6.480 267.850 10.330 268.000 ;
        RECT 10.030 267.400 10.330 267.850 ;
        RECT 6.480 267.250 10.330 267.400 ;
        RECT 10.030 266.800 10.330 267.250 ;
        RECT 6.480 266.650 10.330 266.800 ;
        RECT 10.030 266.200 10.330 266.650 ;
        RECT 6.480 266.050 10.330 266.200 ;
        RECT 10.030 265.600 10.330 266.050 ;
        RECT 6.480 265.450 10.330 265.600 ;
        RECT 10.030 265.000 10.330 265.450 ;
        RECT 6.480 264.850 10.330 265.000 ;
        RECT 10.030 264.400 10.330 264.850 ;
        RECT 6.480 264.250 10.330 264.400 ;
        RECT 10.030 263.800 10.330 264.250 ;
        RECT 6.480 263.650 10.330 263.800 ;
        RECT 10.030 263.200 10.330 263.650 ;
        RECT 6.480 263.050 10.330 263.200 ;
        RECT 10.030 262.600 10.330 263.050 ;
        RECT 6.480 262.450 10.330 262.600 ;
        RECT 10.030 262.000 10.330 262.450 ;
        RECT 6.530 261.450 10.330 262.000 ;
        RECT 10.780 261.450 10.930 269.650 ;
        RECT 11.380 261.450 11.530 269.650 ;
        RECT 11.980 261.450 12.130 269.650 ;
        RECT 12.580 261.450 12.730 269.650 ;
        RECT 13.180 261.450 13.330 269.650 ;
        RECT 13.780 261.450 13.930 269.650 ;
        RECT 14.380 261.450 15.080 278.550 ;
        RECT 15.530 270.350 15.680 278.550 ;
        RECT 16.130 270.350 16.280 278.550 ;
        RECT 16.730 270.350 16.880 278.550 ;
        RECT 17.330 270.350 17.480 278.550 ;
        RECT 17.930 270.350 18.080 278.550 ;
        RECT 18.530 270.350 18.680 278.550 ;
        RECT 19.130 278.000 22.930 278.550 ;
        RECT 26.530 278.550 42.930 278.600 ;
        RECT 26.530 278.000 30.330 278.550 ;
        RECT 19.130 277.550 19.430 278.000 ;
        RECT 30.030 277.550 30.330 278.000 ;
        RECT 19.130 277.400 22.980 277.550 ;
        RECT 26.480 277.400 30.330 277.550 ;
        RECT 19.130 276.950 19.430 277.400 ;
        RECT 30.030 276.950 30.330 277.400 ;
        RECT 19.130 276.800 22.980 276.950 ;
        RECT 26.480 276.800 30.330 276.950 ;
        RECT 19.130 276.350 19.430 276.800 ;
        RECT 30.030 276.350 30.330 276.800 ;
        RECT 19.130 276.200 22.980 276.350 ;
        RECT 26.480 276.200 30.330 276.350 ;
        RECT 19.130 275.750 19.430 276.200 ;
        RECT 30.030 275.750 30.330 276.200 ;
        RECT 19.130 275.600 22.980 275.750 ;
        RECT 26.480 275.600 30.330 275.750 ;
        RECT 19.130 275.150 19.430 275.600 ;
        RECT 30.030 275.150 30.330 275.600 ;
        RECT 19.130 275.000 22.980 275.150 ;
        RECT 26.480 275.000 30.330 275.150 ;
        RECT 19.130 274.550 19.430 275.000 ;
        RECT 30.030 274.550 30.330 275.000 ;
        RECT 19.130 274.400 22.980 274.550 ;
        RECT 26.480 274.400 30.330 274.550 ;
        RECT 19.130 273.950 19.430 274.400 ;
        RECT 30.030 273.950 30.330 274.400 ;
        RECT 19.130 273.800 22.980 273.950 ;
        RECT 26.480 273.800 30.330 273.950 ;
        RECT 19.130 273.350 19.430 273.800 ;
        RECT 30.030 273.350 30.330 273.800 ;
        RECT 19.130 273.200 22.980 273.350 ;
        RECT 26.480 273.200 30.330 273.350 ;
        RECT 19.130 272.750 19.430 273.200 ;
        RECT 19.130 272.600 22.980 272.750 ;
        RECT 19.130 272.150 19.430 272.600 ;
        RECT 19.130 272.000 22.980 272.150 ;
        RECT 19.130 271.550 19.430 272.000 ;
        RECT 19.130 271.400 22.980 271.550 ;
        RECT 19.130 270.950 19.430 271.400 ;
        RECT 19.130 270.800 22.980 270.950 ;
        RECT 19.130 270.350 19.430 270.800 ;
        RECT 15.530 261.450 15.680 269.650 ;
        RECT 16.130 261.450 16.280 269.650 ;
        RECT 16.730 261.450 16.880 269.650 ;
        RECT 17.330 261.450 17.480 269.650 ;
        RECT 17.930 261.450 18.080 269.650 ;
        RECT 18.530 261.450 18.680 269.650 ;
        RECT 19.130 269.200 19.430 269.650 ;
        RECT 19.130 269.050 22.980 269.200 ;
        RECT 19.130 268.600 19.430 269.050 ;
        RECT 19.130 268.450 22.980 268.600 ;
        RECT 19.130 268.000 19.430 268.450 ;
        RECT 19.130 267.850 22.980 268.000 ;
        RECT 19.130 267.400 19.430 267.850 ;
        RECT 19.130 267.250 22.980 267.400 ;
        RECT 19.130 266.800 19.430 267.250 ;
        RECT 23.830 266.800 25.630 273.200 ;
        RECT 30.030 272.750 30.330 273.200 ;
        RECT 26.480 272.600 30.330 272.750 ;
        RECT 30.030 272.150 30.330 272.600 ;
        RECT 26.480 272.000 30.330 272.150 ;
        RECT 30.030 271.550 30.330 272.000 ;
        RECT 26.480 271.400 30.330 271.550 ;
        RECT 30.030 270.950 30.330 271.400 ;
        RECT 26.480 270.800 30.330 270.950 ;
        RECT 30.030 270.350 30.330 270.800 ;
        RECT 30.780 270.350 30.930 278.550 ;
        RECT 31.380 270.350 31.530 278.550 ;
        RECT 31.980 270.350 32.130 278.550 ;
        RECT 32.580 270.350 32.730 278.550 ;
        RECT 33.180 270.350 33.330 278.550 ;
        RECT 33.780 270.350 33.930 278.550 ;
        RECT 30.030 269.200 30.330 269.650 ;
        RECT 26.480 269.050 30.330 269.200 ;
        RECT 30.030 268.600 30.330 269.050 ;
        RECT 26.480 268.450 30.330 268.600 ;
        RECT 30.030 268.000 30.330 268.450 ;
        RECT 26.480 267.850 30.330 268.000 ;
        RECT 30.030 267.400 30.330 267.850 ;
        RECT 26.480 267.250 30.330 267.400 ;
        RECT 30.030 266.800 30.330 267.250 ;
        RECT 19.130 266.650 22.980 266.800 ;
        RECT 26.480 266.650 30.330 266.800 ;
        RECT 19.130 266.200 19.430 266.650 ;
        RECT 30.030 266.200 30.330 266.650 ;
        RECT 19.130 266.050 22.980 266.200 ;
        RECT 26.480 266.050 30.330 266.200 ;
        RECT 19.130 265.600 19.430 266.050 ;
        RECT 30.030 265.600 30.330 266.050 ;
        RECT 19.130 265.450 22.980 265.600 ;
        RECT 26.480 265.450 30.330 265.600 ;
        RECT 19.130 265.000 19.430 265.450 ;
        RECT 30.030 265.000 30.330 265.450 ;
        RECT 19.130 264.850 22.980 265.000 ;
        RECT 26.480 264.850 30.330 265.000 ;
        RECT 19.130 264.400 19.430 264.850 ;
        RECT 30.030 264.400 30.330 264.850 ;
        RECT 19.130 264.250 22.980 264.400 ;
        RECT 26.480 264.250 30.330 264.400 ;
        RECT 19.130 263.800 19.430 264.250 ;
        RECT 30.030 263.800 30.330 264.250 ;
        RECT 19.130 263.650 22.980 263.800 ;
        RECT 26.480 263.650 30.330 263.800 ;
        RECT 19.130 263.200 19.430 263.650 ;
        RECT 30.030 263.200 30.330 263.650 ;
        RECT 19.130 263.050 22.980 263.200 ;
        RECT 26.480 263.050 30.330 263.200 ;
        RECT 19.130 262.600 19.430 263.050 ;
        RECT 30.030 262.600 30.330 263.050 ;
        RECT 19.130 262.450 22.980 262.600 ;
        RECT 26.480 262.450 30.330 262.600 ;
        RECT 19.130 262.000 19.430 262.450 ;
        RECT 30.030 262.000 30.330 262.450 ;
        RECT 19.130 261.450 22.930 262.000 ;
        RECT 6.530 261.400 22.930 261.450 ;
        RECT 26.530 261.450 30.330 262.000 ;
        RECT 30.780 261.450 30.930 269.650 ;
        RECT 31.380 261.450 31.530 269.650 ;
        RECT 31.980 261.450 32.130 269.650 ;
        RECT 32.580 261.450 32.730 269.650 ;
        RECT 33.180 261.450 33.330 269.650 ;
        RECT 33.780 261.450 33.930 269.650 ;
        RECT 34.380 261.450 35.080 278.550 ;
        RECT 35.530 270.350 35.680 278.550 ;
        RECT 36.130 270.350 36.280 278.550 ;
        RECT 36.730 270.350 36.880 278.550 ;
        RECT 37.330 270.350 37.480 278.550 ;
        RECT 37.930 270.350 38.080 278.550 ;
        RECT 38.530 270.350 38.680 278.550 ;
        RECT 39.130 278.000 42.930 278.550 ;
        RECT 46.530 278.550 62.930 278.600 ;
        RECT 46.530 278.000 50.330 278.550 ;
        RECT 39.130 277.550 39.430 278.000 ;
        RECT 50.030 277.550 50.330 278.000 ;
        RECT 39.130 277.400 42.980 277.550 ;
        RECT 46.480 277.400 50.330 277.550 ;
        RECT 39.130 276.950 39.430 277.400 ;
        RECT 50.030 276.950 50.330 277.400 ;
        RECT 39.130 276.800 42.980 276.950 ;
        RECT 46.480 276.800 50.330 276.950 ;
        RECT 39.130 276.350 39.430 276.800 ;
        RECT 50.030 276.350 50.330 276.800 ;
        RECT 39.130 276.200 42.980 276.350 ;
        RECT 46.480 276.200 50.330 276.350 ;
        RECT 39.130 275.750 39.430 276.200 ;
        RECT 50.030 275.750 50.330 276.200 ;
        RECT 39.130 275.600 42.980 275.750 ;
        RECT 46.480 275.600 50.330 275.750 ;
        RECT 39.130 275.150 39.430 275.600 ;
        RECT 50.030 275.150 50.330 275.600 ;
        RECT 39.130 275.000 42.980 275.150 ;
        RECT 46.480 275.000 50.330 275.150 ;
        RECT 39.130 274.550 39.430 275.000 ;
        RECT 50.030 274.550 50.330 275.000 ;
        RECT 39.130 274.400 42.980 274.550 ;
        RECT 46.480 274.400 50.330 274.550 ;
        RECT 39.130 273.950 39.430 274.400 ;
        RECT 50.030 273.950 50.330 274.400 ;
        RECT 39.130 273.800 42.980 273.950 ;
        RECT 46.480 273.800 50.330 273.950 ;
        RECT 39.130 273.350 39.430 273.800 ;
        RECT 50.030 273.350 50.330 273.800 ;
        RECT 39.130 273.200 42.980 273.350 ;
        RECT 46.480 273.200 50.330 273.350 ;
        RECT 39.130 272.750 39.430 273.200 ;
        RECT 39.130 272.600 42.980 272.750 ;
        RECT 39.130 272.150 39.430 272.600 ;
        RECT 39.130 272.000 42.980 272.150 ;
        RECT 39.130 271.550 39.430 272.000 ;
        RECT 39.130 271.400 42.980 271.550 ;
        RECT 39.130 270.950 39.430 271.400 ;
        RECT 39.130 270.800 42.980 270.950 ;
        RECT 39.130 270.350 39.430 270.800 ;
        RECT 35.530 261.450 35.680 269.650 ;
        RECT 36.130 261.450 36.280 269.650 ;
        RECT 36.730 261.450 36.880 269.650 ;
        RECT 37.330 261.450 37.480 269.650 ;
        RECT 37.930 261.450 38.080 269.650 ;
        RECT 38.530 261.450 38.680 269.650 ;
        RECT 39.130 269.200 39.430 269.650 ;
        RECT 39.130 269.050 42.980 269.200 ;
        RECT 39.130 268.600 39.430 269.050 ;
        RECT 39.130 268.450 42.980 268.600 ;
        RECT 39.130 268.000 39.430 268.450 ;
        RECT 39.130 267.850 42.980 268.000 ;
        RECT 39.130 267.400 39.430 267.850 ;
        RECT 39.130 267.250 42.980 267.400 ;
        RECT 39.130 266.800 39.430 267.250 ;
        RECT 43.830 266.800 45.630 273.200 ;
        RECT 50.030 272.750 50.330 273.200 ;
        RECT 46.480 272.600 50.330 272.750 ;
        RECT 50.030 272.150 50.330 272.600 ;
        RECT 46.480 272.000 50.330 272.150 ;
        RECT 50.030 271.550 50.330 272.000 ;
        RECT 46.480 271.400 50.330 271.550 ;
        RECT 50.030 270.950 50.330 271.400 ;
        RECT 46.480 270.800 50.330 270.950 ;
        RECT 50.030 270.350 50.330 270.800 ;
        RECT 50.780 270.350 50.930 278.550 ;
        RECT 51.380 270.350 51.530 278.550 ;
        RECT 51.980 270.350 52.130 278.550 ;
        RECT 52.580 270.350 52.730 278.550 ;
        RECT 53.180 270.350 53.330 278.550 ;
        RECT 53.780 270.350 53.930 278.550 ;
        RECT 50.030 269.200 50.330 269.650 ;
        RECT 46.480 269.050 50.330 269.200 ;
        RECT 50.030 268.600 50.330 269.050 ;
        RECT 46.480 268.450 50.330 268.600 ;
        RECT 50.030 268.000 50.330 268.450 ;
        RECT 46.480 267.850 50.330 268.000 ;
        RECT 50.030 267.400 50.330 267.850 ;
        RECT 46.480 267.250 50.330 267.400 ;
        RECT 50.030 266.800 50.330 267.250 ;
        RECT 39.130 266.650 42.980 266.800 ;
        RECT 46.480 266.650 50.330 266.800 ;
        RECT 39.130 266.200 39.430 266.650 ;
        RECT 50.030 266.200 50.330 266.650 ;
        RECT 39.130 266.050 42.980 266.200 ;
        RECT 46.480 266.050 50.330 266.200 ;
        RECT 39.130 265.600 39.430 266.050 ;
        RECT 50.030 265.600 50.330 266.050 ;
        RECT 39.130 265.450 42.980 265.600 ;
        RECT 46.480 265.450 50.330 265.600 ;
        RECT 39.130 265.000 39.430 265.450 ;
        RECT 50.030 265.000 50.330 265.450 ;
        RECT 39.130 264.850 42.980 265.000 ;
        RECT 46.480 264.850 50.330 265.000 ;
        RECT 39.130 264.400 39.430 264.850 ;
        RECT 50.030 264.400 50.330 264.850 ;
        RECT 39.130 264.250 42.980 264.400 ;
        RECT 46.480 264.250 50.330 264.400 ;
        RECT 39.130 263.800 39.430 264.250 ;
        RECT 50.030 263.800 50.330 264.250 ;
        RECT 39.130 263.650 42.980 263.800 ;
        RECT 46.480 263.650 50.330 263.800 ;
        RECT 39.130 263.200 39.430 263.650 ;
        RECT 50.030 263.200 50.330 263.650 ;
        RECT 39.130 263.050 42.980 263.200 ;
        RECT 46.480 263.050 50.330 263.200 ;
        RECT 39.130 262.600 39.430 263.050 ;
        RECT 50.030 262.600 50.330 263.050 ;
        RECT 39.130 262.450 42.980 262.600 ;
        RECT 46.480 262.450 50.330 262.600 ;
        RECT 39.130 262.000 39.430 262.450 ;
        RECT 50.030 262.000 50.330 262.450 ;
        RECT 39.130 261.450 42.930 262.000 ;
        RECT 26.530 261.400 42.930 261.450 ;
        RECT 46.530 261.450 50.330 262.000 ;
        RECT 50.780 261.450 50.930 269.650 ;
        RECT 51.380 261.450 51.530 269.650 ;
        RECT 51.980 261.450 52.130 269.650 ;
        RECT 52.580 261.450 52.730 269.650 ;
        RECT 53.180 261.450 53.330 269.650 ;
        RECT 53.780 261.450 53.930 269.650 ;
        RECT 54.380 261.450 55.080 278.550 ;
        RECT 55.530 270.350 55.680 278.550 ;
        RECT 56.130 270.350 56.280 278.550 ;
        RECT 56.730 270.350 56.880 278.550 ;
        RECT 57.330 270.350 57.480 278.550 ;
        RECT 57.930 270.350 58.080 278.550 ;
        RECT 58.530 270.350 58.680 278.550 ;
        RECT 59.130 278.000 62.930 278.550 ;
        RECT 66.530 278.550 82.930 278.600 ;
        RECT 66.530 278.000 70.330 278.550 ;
        RECT 59.130 277.550 59.430 278.000 ;
        RECT 70.030 277.550 70.330 278.000 ;
        RECT 59.130 277.400 62.980 277.550 ;
        RECT 66.480 277.400 70.330 277.550 ;
        RECT 59.130 276.950 59.430 277.400 ;
        RECT 70.030 276.950 70.330 277.400 ;
        RECT 59.130 276.800 62.980 276.950 ;
        RECT 66.480 276.800 70.330 276.950 ;
        RECT 59.130 276.350 59.430 276.800 ;
        RECT 70.030 276.350 70.330 276.800 ;
        RECT 59.130 276.200 62.980 276.350 ;
        RECT 66.480 276.200 70.330 276.350 ;
        RECT 59.130 275.750 59.430 276.200 ;
        RECT 70.030 275.750 70.330 276.200 ;
        RECT 59.130 275.600 62.980 275.750 ;
        RECT 66.480 275.600 70.330 275.750 ;
        RECT 59.130 275.150 59.430 275.600 ;
        RECT 70.030 275.150 70.330 275.600 ;
        RECT 59.130 275.000 62.980 275.150 ;
        RECT 66.480 275.000 70.330 275.150 ;
        RECT 59.130 274.550 59.430 275.000 ;
        RECT 70.030 274.550 70.330 275.000 ;
        RECT 59.130 274.400 62.980 274.550 ;
        RECT 66.480 274.400 70.330 274.550 ;
        RECT 59.130 273.950 59.430 274.400 ;
        RECT 70.030 273.950 70.330 274.400 ;
        RECT 59.130 273.800 62.980 273.950 ;
        RECT 66.480 273.800 70.330 273.950 ;
        RECT 59.130 273.350 59.430 273.800 ;
        RECT 70.030 273.350 70.330 273.800 ;
        RECT 59.130 273.200 62.980 273.350 ;
        RECT 66.480 273.200 70.330 273.350 ;
        RECT 59.130 272.750 59.430 273.200 ;
        RECT 59.130 272.600 62.980 272.750 ;
        RECT 59.130 272.150 59.430 272.600 ;
        RECT 59.130 272.000 62.980 272.150 ;
        RECT 59.130 271.550 59.430 272.000 ;
        RECT 59.130 271.400 62.980 271.550 ;
        RECT 59.130 270.950 59.430 271.400 ;
        RECT 59.130 270.800 62.980 270.950 ;
        RECT 59.130 270.350 59.430 270.800 ;
        RECT 55.530 261.450 55.680 269.650 ;
        RECT 56.130 261.450 56.280 269.650 ;
        RECT 56.730 261.450 56.880 269.650 ;
        RECT 57.330 261.450 57.480 269.650 ;
        RECT 57.930 261.450 58.080 269.650 ;
        RECT 58.530 261.450 58.680 269.650 ;
        RECT 59.130 269.200 59.430 269.650 ;
        RECT 59.130 269.050 62.980 269.200 ;
        RECT 59.130 268.600 59.430 269.050 ;
        RECT 59.130 268.450 62.980 268.600 ;
        RECT 59.130 268.000 59.430 268.450 ;
        RECT 59.130 267.850 62.980 268.000 ;
        RECT 59.130 267.400 59.430 267.850 ;
        RECT 59.130 267.250 62.980 267.400 ;
        RECT 59.130 266.800 59.430 267.250 ;
        RECT 63.830 266.800 65.630 273.200 ;
        RECT 70.030 272.750 70.330 273.200 ;
        RECT 66.480 272.600 70.330 272.750 ;
        RECT 70.030 272.150 70.330 272.600 ;
        RECT 66.480 272.000 70.330 272.150 ;
        RECT 70.030 271.550 70.330 272.000 ;
        RECT 66.480 271.400 70.330 271.550 ;
        RECT 70.030 270.950 70.330 271.400 ;
        RECT 66.480 270.800 70.330 270.950 ;
        RECT 70.030 270.350 70.330 270.800 ;
        RECT 70.780 270.350 70.930 278.550 ;
        RECT 71.380 270.350 71.530 278.550 ;
        RECT 71.980 270.350 72.130 278.550 ;
        RECT 72.580 270.350 72.730 278.550 ;
        RECT 73.180 270.350 73.330 278.550 ;
        RECT 73.780 270.350 73.930 278.550 ;
        RECT 70.030 269.200 70.330 269.650 ;
        RECT 66.480 269.050 70.330 269.200 ;
        RECT 70.030 268.600 70.330 269.050 ;
        RECT 66.480 268.450 70.330 268.600 ;
        RECT 70.030 268.000 70.330 268.450 ;
        RECT 66.480 267.850 70.330 268.000 ;
        RECT 70.030 267.400 70.330 267.850 ;
        RECT 66.480 267.250 70.330 267.400 ;
        RECT 70.030 266.800 70.330 267.250 ;
        RECT 59.130 266.650 62.980 266.800 ;
        RECT 66.480 266.650 70.330 266.800 ;
        RECT 59.130 266.200 59.430 266.650 ;
        RECT 70.030 266.200 70.330 266.650 ;
        RECT 59.130 266.050 62.980 266.200 ;
        RECT 66.480 266.050 70.330 266.200 ;
        RECT 59.130 265.600 59.430 266.050 ;
        RECT 70.030 265.600 70.330 266.050 ;
        RECT 59.130 265.450 62.980 265.600 ;
        RECT 66.480 265.450 70.330 265.600 ;
        RECT 59.130 265.000 59.430 265.450 ;
        RECT 70.030 265.000 70.330 265.450 ;
        RECT 59.130 264.850 62.980 265.000 ;
        RECT 66.480 264.850 70.330 265.000 ;
        RECT 59.130 264.400 59.430 264.850 ;
        RECT 70.030 264.400 70.330 264.850 ;
        RECT 59.130 264.250 62.980 264.400 ;
        RECT 66.480 264.250 70.330 264.400 ;
        RECT 59.130 263.800 59.430 264.250 ;
        RECT 70.030 263.800 70.330 264.250 ;
        RECT 59.130 263.650 62.980 263.800 ;
        RECT 66.480 263.650 70.330 263.800 ;
        RECT 59.130 263.200 59.430 263.650 ;
        RECT 70.030 263.200 70.330 263.650 ;
        RECT 59.130 263.050 62.980 263.200 ;
        RECT 66.480 263.050 70.330 263.200 ;
        RECT 59.130 262.600 59.430 263.050 ;
        RECT 70.030 262.600 70.330 263.050 ;
        RECT 59.130 262.450 62.980 262.600 ;
        RECT 66.480 262.450 70.330 262.600 ;
        RECT 59.130 262.000 59.430 262.450 ;
        RECT 70.030 262.000 70.330 262.450 ;
        RECT 59.130 261.450 62.930 262.000 ;
        RECT 46.530 261.400 62.930 261.450 ;
        RECT 66.530 261.450 70.330 262.000 ;
        RECT 70.780 261.450 70.930 269.650 ;
        RECT 71.380 261.450 71.530 269.650 ;
        RECT 71.980 261.450 72.130 269.650 ;
        RECT 72.580 261.450 72.730 269.650 ;
        RECT 73.180 261.450 73.330 269.650 ;
        RECT 73.780 261.450 73.930 269.650 ;
        RECT 74.380 261.450 75.080 278.550 ;
        RECT 75.530 270.350 75.680 278.550 ;
        RECT 76.130 270.350 76.280 278.550 ;
        RECT 76.730 270.350 76.880 278.550 ;
        RECT 77.330 270.350 77.480 278.550 ;
        RECT 77.930 270.350 78.080 278.550 ;
        RECT 78.530 270.350 78.680 278.550 ;
        RECT 79.130 278.000 82.930 278.550 ;
        RECT 86.530 278.550 102.930 278.600 ;
        RECT 86.530 278.000 90.330 278.550 ;
        RECT 79.130 277.550 79.430 278.000 ;
        RECT 90.030 277.550 90.330 278.000 ;
        RECT 79.130 277.400 82.980 277.550 ;
        RECT 86.480 277.400 90.330 277.550 ;
        RECT 79.130 276.950 79.430 277.400 ;
        RECT 90.030 276.950 90.330 277.400 ;
        RECT 79.130 276.800 82.980 276.950 ;
        RECT 86.480 276.800 90.330 276.950 ;
        RECT 79.130 276.350 79.430 276.800 ;
        RECT 90.030 276.350 90.330 276.800 ;
        RECT 79.130 276.200 82.980 276.350 ;
        RECT 86.480 276.200 90.330 276.350 ;
        RECT 79.130 275.750 79.430 276.200 ;
        RECT 90.030 275.750 90.330 276.200 ;
        RECT 79.130 275.600 82.980 275.750 ;
        RECT 86.480 275.600 90.330 275.750 ;
        RECT 79.130 275.150 79.430 275.600 ;
        RECT 90.030 275.150 90.330 275.600 ;
        RECT 79.130 275.000 82.980 275.150 ;
        RECT 86.480 275.000 90.330 275.150 ;
        RECT 79.130 274.550 79.430 275.000 ;
        RECT 90.030 274.550 90.330 275.000 ;
        RECT 79.130 274.400 82.980 274.550 ;
        RECT 86.480 274.400 90.330 274.550 ;
        RECT 79.130 273.950 79.430 274.400 ;
        RECT 90.030 273.950 90.330 274.400 ;
        RECT 79.130 273.800 82.980 273.950 ;
        RECT 86.480 273.800 90.330 273.950 ;
        RECT 79.130 273.350 79.430 273.800 ;
        RECT 90.030 273.350 90.330 273.800 ;
        RECT 79.130 273.200 82.980 273.350 ;
        RECT 86.480 273.200 90.330 273.350 ;
        RECT 79.130 272.750 79.430 273.200 ;
        RECT 79.130 272.600 82.980 272.750 ;
        RECT 79.130 272.150 79.430 272.600 ;
        RECT 79.130 272.000 82.980 272.150 ;
        RECT 79.130 271.550 79.430 272.000 ;
        RECT 79.130 271.400 82.980 271.550 ;
        RECT 79.130 270.950 79.430 271.400 ;
        RECT 79.130 270.800 82.980 270.950 ;
        RECT 79.130 270.350 79.430 270.800 ;
        RECT 75.530 261.450 75.680 269.650 ;
        RECT 76.130 261.450 76.280 269.650 ;
        RECT 76.730 261.450 76.880 269.650 ;
        RECT 77.330 261.450 77.480 269.650 ;
        RECT 77.930 261.450 78.080 269.650 ;
        RECT 78.530 261.450 78.680 269.650 ;
        RECT 79.130 269.200 79.430 269.650 ;
        RECT 79.130 269.050 82.980 269.200 ;
        RECT 79.130 268.600 79.430 269.050 ;
        RECT 79.130 268.450 82.980 268.600 ;
        RECT 79.130 268.000 79.430 268.450 ;
        RECT 79.130 267.850 82.980 268.000 ;
        RECT 79.130 267.400 79.430 267.850 ;
        RECT 79.130 267.250 82.980 267.400 ;
        RECT 79.130 266.800 79.430 267.250 ;
        RECT 83.830 266.800 85.630 273.200 ;
        RECT 90.030 272.750 90.330 273.200 ;
        RECT 86.480 272.600 90.330 272.750 ;
        RECT 90.030 272.150 90.330 272.600 ;
        RECT 86.480 272.000 90.330 272.150 ;
        RECT 90.030 271.550 90.330 272.000 ;
        RECT 86.480 271.400 90.330 271.550 ;
        RECT 90.030 270.950 90.330 271.400 ;
        RECT 86.480 270.800 90.330 270.950 ;
        RECT 90.030 270.350 90.330 270.800 ;
        RECT 90.780 270.350 90.930 278.550 ;
        RECT 91.380 270.350 91.530 278.550 ;
        RECT 91.980 270.350 92.130 278.550 ;
        RECT 92.580 270.350 92.730 278.550 ;
        RECT 93.180 270.350 93.330 278.550 ;
        RECT 93.780 270.350 93.930 278.550 ;
        RECT 90.030 269.200 90.330 269.650 ;
        RECT 86.480 269.050 90.330 269.200 ;
        RECT 90.030 268.600 90.330 269.050 ;
        RECT 86.480 268.450 90.330 268.600 ;
        RECT 90.030 268.000 90.330 268.450 ;
        RECT 86.480 267.850 90.330 268.000 ;
        RECT 90.030 267.400 90.330 267.850 ;
        RECT 86.480 267.250 90.330 267.400 ;
        RECT 90.030 266.800 90.330 267.250 ;
        RECT 79.130 266.650 82.980 266.800 ;
        RECT 86.480 266.650 90.330 266.800 ;
        RECT 79.130 266.200 79.430 266.650 ;
        RECT 90.030 266.200 90.330 266.650 ;
        RECT 79.130 266.050 82.980 266.200 ;
        RECT 86.480 266.050 90.330 266.200 ;
        RECT 79.130 265.600 79.430 266.050 ;
        RECT 90.030 265.600 90.330 266.050 ;
        RECT 79.130 265.450 82.980 265.600 ;
        RECT 86.480 265.450 90.330 265.600 ;
        RECT 79.130 265.000 79.430 265.450 ;
        RECT 90.030 265.000 90.330 265.450 ;
        RECT 79.130 264.850 82.980 265.000 ;
        RECT 86.480 264.850 90.330 265.000 ;
        RECT 79.130 264.400 79.430 264.850 ;
        RECT 90.030 264.400 90.330 264.850 ;
        RECT 79.130 264.250 82.980 264.400 ;
        RECT 86.480 264.250 90.330 264.400 ;
        RECT 79.130 263.800 79.430 264.250 ;
        RECT 90.030 263.800 90.330 264.250 ;
        RECT 79.130 263.650 82.980 263.800 ;
        RECT 86.480 263.650 90.330 263.800 ;
        RECT 79.130 263.200 79.430 263.650 ;
        RECT 90.030 263.200 90.330 263.650 ;
        RECT 79.130 263.050 82.980 263.200 ;
        RECT 86.480 263.050 90.330 263.200 ;
        RECT 79.130 262.600 79.430 263.050 ;
        RECT 90.030 262.600 90.330 263.050 ;
        RECT 79.130 262.450 82.980 262.600 ;
        RECT 86.480 262.450 90.330 262.600 ;
        RECT 79.130 262.000 79.430 262.450 ;
        RECT 90.030 262.000 90.330 262.450 ;
        RECT 79.130 261.450 82.930 262.000 ;
        RECT 66.530 261.400 82.930 261.450 ;
        RECT 86.530 261.450 90.330 262.000 ;
        RECT 90.780 261.450 90.930 269.650 ;
        RECT 91.380 261.450 91.530 269.650 ;
        RECT 91.980 261.450 92.130 269.650 ;
        RECT 92.580 261.450 92.730 269.650 ;
        RECT 93.180 261.450 93.330 269.650 ;
        RECT 93.780 261.450 93.930 269.650 ;
        RECT 94.380 261.450 95.080 278.550 ;
        RECT 95.530 270.350 95.680 278.550 ;
        RECT 96.130 270.350 96.280 278.550 ;
        RECT 96.730 270.350 96.880 278.550 ;
        RECT 97.330 270.350 97.480 278.550 ;
        RECT 97.930 270.350 98.080 278.550 ;
        RECT 98.530 270.350 98.680 278.550 ;
        RECT 99.130 278.000 102.930 278.550 ;
        RECT 106.530 278.550 122.930 278.600 ;
        RECT 106.530 278.000 110.330 278.550 ;
        RECT 99.130 277.550 99.430 278.000 ;
        RECT 110.030 277.550 110.330 278.000 ;
        RECT 99.130 277.400 102.980 277.550 ;
        RECT 106.480 277.400 110.330 277.550 ;
        RECT 99.130 276.950 99.430 277.400 ;
        RECT 110.030 276.950 110.330 277.400 ;
        RECT 99.130 276.800 102.980 276.950 ;
        RECT 106.480 276.800 110.330 276.950 ;
        RECT 99.130 276.350 99.430 276.800 ;
        RECT 110.030 276.350 110.330 276.800 ;
        RECT 99.130 276.200 102.980 276.350 ;
        RECT 106.480 276.200 110.330 276.350 ;
        RECT 99.130 275.750 99.430 276.200 ;
        RECT 110.030 275.750 110.330 276.200 ;
        RECT 99.130 275.600 102.980 275.750 ;
        RECT 106.480 275.600 110.330 275.750 ;
        RECT 99.130 275.150 99.430 275.600 ;
        RECT 110.030 275.150 110.330 275.600 ;
        RECT 99.130 275.000 102.980 275.150 ;
        RECT 106.480 275.000 110.330 275.150 ;
        RECT 99.130 274.550 99.430 275.000 ;
        RECT 110.030 274.550 110.330 275.000 ;
        RECT 99.130 274.400 102.980 274.550 ;
        RECT 106.480 274.400 110.330 274.550 ;
        RECT 99.130 273.950 99.430 274.400 ;
        RECT 110.030 273.950 110.330 274.400 ;
        RECT 99.130 273.800 102.980 273.950 ;
        RECT 106.480 273.800 110.330 273.950 ;
        RECT 99.130 273.350 99.430 273.800 ;
        RECT 110.030 273.350 110.330 273.800 ;
        RECT 99.130 273.200 102.980 273.350 ;
        RECT 106.480 273.200 110.330 273.350 ;
        RECT 99.130 272.750 99.430 273.200 ;
        RECT 99.130 272.600 102.980 272.750 ;
        RECT 99.130 272.150 99.430 272.600 ;
        RECT 99.130 272.000 102.980 272.150 ;
        RECT 99.130 271.550 99.430 272.000 ;
        RECT 99.130 271.400 102.980 271.550 ;
        RECT 99.130 270.950 99.430 271.400 ;
        RECT 99.130 270.800 102.980 270.950 ;
        RECT 99.130 270.350 99.430 270.800 ;
        RECT 95.530 261.450 95.680 269.650 ;
        RECT 96.130 261.450 96.280 269.650 ;
        RECT 96.730 261.450 96.880 269.650 ;
        RECT 97.330 261.450 97.480 269.650 ;
        RECT 97.930 261.450 98.080 269.650 ;
        RECT 98.530 261.450 98.680 269.650 ;
        RECT 99.130 269.200 99.430 269.650 ;
        RECT 99.130 269.050 102.980 269.200 ;
        RECT 99.130 268.600 99.430 269.050 ;
        RECT 99.130 268.450 102.980 268.600 ;
        RECT 99.130 268.000 99.430 268.450 ;
        RECT 99.130 267.850 102.980 268.000 ;
        RECT 99.130 267.400 99.430 267.850 ;
        RECT 99.130 267.250 102.980 267.400 ;
        RECT 99.130 266.800 99.430 267.250 ;
        RECT 103.830 266.800 105.630 273.200 ;
        RECT 110.030 272.750 110.330 273.200 ;
        RECT 106.480 272.600 110.330 272.750 ;
        RECT 110.030 272.150 110.330 272.600 ;
        RECT 106.480 272.000 110.330 272.150 ;
        RECT 110.030 271.550 110.330 272.000 ;
        RECT 106.480 271.400 110.330 271.550 ;
        RECT 110.030 270.950 110.330 271.400 ;
        RECT 106.480 270.800 110.330 270.950 ;
        RECT 110.030 270.350 110.330 270.800 ;
        RECT 110.780 270.350 110.930 278.550 ;
        RECT 111.380 270.350 111.530 278.550 ;
        RECT 111.980 270.350 112.130 278.550 ;
        RECT 112.580 270.350 112.730 278.550 ;
        RECT 113.180 270.350 113.330 278.550 ;
        RECT 113.780 270.350 113.930 278.550 ;
        RECT 110.030 269.200 110.330 269.650 ;
        RECT 106.480 269.050 110.330 269.200 ;
        RECT 110.030 268.600 110.330 269.050 ;
        RECT 106.480 268.450 110.330 268.600 ;
        RECT 110.030 268.000 110.330 268.450 ;
        RECT 106.480 267.850 110.330 268.000 ;
        RECT 110.030 267.400 110.330 267.850 ;
        RECT 106.480 267.250 110.330 267.400 ;
        RECT 110.030 266.800 110.330 267.250 ;
        RECT 99.130 266.650 102.980 266.800 ;
        RECT 106.480 266.650 110.330 266.800 ;
        RECT 99.130 266.200 99.430 266.650 ;
        RECT 110.030 266.200 110.330 266.650 ;
        RECT 99.130 266.050 102.980 266.200 ;
        RECT 106.480 266.050 110.330 266.200 ;
        RECT 99.130 265.600 99.430 266.050 ;
        RECT 110.030 265.600 110.330 266.050 ;
        RECT 99.130 265.450 102.980 265.600 ;
        RECT 106.480 265.450 110.330 265.600 ;
        RECT 99.130 265.000 99.430 265.450 ;
        RECT 110.030 265.000 110.330 265.450 ;
        RECT 99.130 264.850 102.980 265.000 ;
        RECT 106.480 264.850 110.330 265.000 ;
        RECT 99.130 264.400 99.430 264.850 ;
        RECT 110.030 264.400 110.330 264.850 ;
        RECT 99.130 264.250 102.980 264.400 ;
        RECT 106.480 264.250 110.330 264.400 ;
        RECT 99.130 263.800 99.430 264.250 ;
        RECT 110.030 263.800 110.330 264.250 ;
        RECT 99.130 263.650 102.980 263.800 ;
        RECT 106.480 263.650 110.330 263.800 ;
        RECT 99.130 263.200 99.430 263.650 ;
        RECT 110.030 263.200 110.330 263.650 ;
        RECT 99.130 263.050 102.980 263.200 ;
        RECT 106.480 263.050 110.330 263.200 ;
        RECT 99.130 262.600 99.430 263.050 ;
        RECT 110.030 262.600 110.330 263.050 ;
        RECT 99.130 262.450 102.980 262.600 ;
        RECT 106.480 262.450 110.330 262.600 ;
        RECT 99.130 262.000 99.430 262.450 ;
        RECT 110.030 262.000 110.330 262.450 ;
        RECT 99.130 261.450 102.930 262.000 ;
        RECT 86.530 261.400 102.930 261.450 ;
        RECT 106.530 261.450 110.330 262.000 ;
        RECT 110.780 261.450 110.930 269.650 ;
        RECT 111.380 261.450 111.530 269.650 ;
        RECT 111.980 261.450 112.130 269.650 ;
        RECT 112.580 261.450 112.730 269.650 ;
        RECT 113.180 261.450 113.330 269.650 ;
        RECT 113.780 261.450 113.930 269.650 ;
        RECT 114.380 261.450 115.080 278.550 ;
        RECT 115.530 270.350 115.680 278.550 ;
        RECT 116.130 270.350 116.280 278.550 ;
        RECT 116.730 270.350 116.880 278.550 ;
        RECT 117.330 270.350 117.480 278.550 ;
        RECT 117.930 270.350 118.080 278.550 ;
        RECT 118.530 270.350 118.680 278.550 ;
        RECT 119.130 278.000 122.930 278.550 ;
        RECT 119.130 277.550 119.430 278.000 ;
        RECT 119.130 277.400 122.980 277.550 ;
        RECT 119.130 276.950 119.430 277.400 ;
        RECT 119.130 276.800 122.980 276.950 ;
        RECT 119.130 276.350 119.430 276.800 ;
        RECT 119.130 276.200 122.980 276.350 ;
        RECT 119.130 275.750 119.430 276.200 ;
        RECT 119.130 275.600 122.980 275.750 ;
        RECT 119.130 275.150 119.430 275.600 ;
        RECT 119.130 275.000 122.980 275.150 ;
        RECT 119.130 274.550 119.430 275.000 ;
        RECT 119.130 274.400 122.980 274.550 ;
        RECT 119.130 273.950 119.430 274.400 ;
        RECT 119.130 273.800 122.980 273.950 ;
        RECT 119.130 273.350 119.430 273.800 ;
        RECT 119.130 273.200 122.980 273.350 ;
        RECT 119.130 272.750 119.430 273.200 ;
        RECT 119.130 272.600 122.980 272.750 ;
        RECT 119.130 272.150 119.430 272.600 ;
        RECT 119.130 272.000 122.980 272.150 ;
        RECT 119.130 271.550 119.430 272.000 ;
        RECT 119.130 271.400 122.980 271.550 ;
        RECT 119.130 270.950 119.430 271.400 ;
        RECT 119.130 270.800 122.980 270.950 ;
        RECT 119.130 270.350 119.430 270.800 ;
        RECT 115.530 261.450 115.680 269.650 ;
        RECT 116.130 261.450 116.280 269.650 ;
        RECT 116.730 261.450 116.880 269.650 ;
        RECT 117.330 261.450 117.480 269.650 ;
        RECT 117.930 261.450 118.080 269.650 ;
        RECT 118.530 261.450 118.680 269.650 ;
        RECT 119.130 269.200 119.430 269.650 ;
        RECT 119.130 269.050 122.980 269.200 ;
        RECT 119.130 268.600 119.430 269.050 ;
        RECT 119.130 268.450 122.980 268.600 ;
        RECT 119.130 268.000 119.430 268.450 ;
        RECT 119.130 267.850 122.980 268.000 ;
        RECT 119.130 267.400 119.430 267.850 ;
        RECT 119.130 267.250 122.980 267.400 ;
        RECT 119.130 266.800 119.430 267.250 ;
        RECT 123.830 266.800 124.730 273.200 ;
        RECT 129.850 269.330 131.850 270.605 ;
        RECT 119.130 266.650 122.980 266.800 ;
        RECT 119.130 266.200 119.430 266.650 ;
        RECT 119.130 266.050 122.980 266.200 ;
        RECT 119.130 265.600 119.430 266.050 ;
        RECT 119.130 265.450 122.980 265.600 ;
        RECT 119.130 265.000 119.430 265.450 ;
        RECT 119.130 264.850 122.980 265.000 ;
        RECT 119.130 264.400 119.430 264.850 ;
        RECT 119.130 264.250 122.980 264.400 ;
        RECT 119.130 263.800 119.430 264.250 ;
        RECT 119.130 263.650 122.980 263.800 ;
        RECT 119.130 263.200 119.430 263.650 ;
        RECT 119.130 263.050 122.980 263.200 ;
        RECT 119.130 262.600 119.430 263.050 ;
        RECT 119.130 262.450 122.980 262.600 ;
        RECT 119.130 262.000 119.430 262.450 ;
        RECT 119.130 261.450 122.930 262.000 ;
        RECT 106.530 261.400 122.930 261.450 ;
        RECT 9.630 260.900 19.830 261.400 ;
        RECT 29.630 260.900 39.830 261.400 ;
        RECT 49.630 260.900 59.830 261.400 ;
        RECT 69.630 260.900 79.830 261.400 ;
        RECT 89.630 260.900 99.830 261.400 ;
        RECT 109.630 260.900 119.830 261.400 ;
        RECT 11.530 259.100 17.930 260.900 ;
        RECT 31.530 259.100 37.930 260.900 ;
        RECT 51.530 259.100 57.930 260.900 ;
        RECT 71.530 259.100 77.930 260.900 ;
        RECT 91.530 259.100 97.930 260.900 ;
        RECT 111.530 259.100 117.930 260.900 ;
        RECT 9.630 258.600 19.830 259.100 ;
        RECT 29.630 258.600 39.830 259.100 ;
        RECT 49.630 258.600 59.830 259.100 ;
        RECT 69.630 258.600 79.830 259.100 ;
        RECT 89.630 258.600 99.830 259.100 ;
        RECT 109.630 258.600 119.830 259.100 ;
        RECT 6.530 258.550 22.930 258.600 ;
        RECT 6.530 258.000 10.330 258.550 ;
        RECT 10.030 257.550 10.330 258.000 ;
        RECT 6.480 257.400 10.330 257.550 ;
        RECT 10.030 256.950 10.330 257.400 ;
        RECT 6.480 256.800 10.330 256.950 ;
        RECT 10.030 256.350 10.330 256.800 ;
        RECT 6.480 256.200 10.330 256.350 ;
        RECT 10.030 255.750 10.330 256.200 ;
        RECT 6.480 255.600 10.330 255.750 ;
        RECT 10.030 255.150 10.330 255.600 ;
        RECT 6.480 255.000 10.330 255.150 ;
        RECT 10.030 254.550 10.330 255.000 ;
        RECT 6.480 254.400 10.330 254.550 ;
        RECT 10.030 253.950 10.330 254.400 ;
        RECT 6.480 253.800 10.330 253.950 ;
        RECT 10.030 253.350 10.330 253.800 ;
        RECT 6.480 253.200 10.330 253.350 ;
        RECT 4.730 246.800 5.630 253.200 ;
        RECT 10.030 252.750 10.330 253.200 ;
        RECT 6.480 252.600 10.330 252.750 ;
        RECT 10.030 252.150 10.330 252.600 ;
        RECT 6.480 252.000 10.330 252.150 ;
        RECT 10.030 251.550 10.330 252.000 ;
        RECT 6.480 251.400 10.330 251.550 ;
        RECT 10.030 250.950 10.330 251.400 ;
        RECT 6.480 250.800 10.330 250.950 ;
        RECT 10.030 250.350 10.330 250.800 ;
        RECT 10.780 250.350 10.930 258.550 ;
        RECT 11.380 250.350 11.530 258.550 ;
        RECT 11.980 250.350 12.130 258.550 ;
        RECT 12.580 250.350 12.730 258.550 ;
        RECT 13.180 250.350 13.330 258.550 ;
        RECT 13.780 250.350 13.930 258.550 ;
        RECT 10.030 249.200 10.330 249.650 ;
        RECT 6.480 249.050 10.330 249.200 ;
        RECT 10.030 248.600 10.330 249.050 ;
        RECT 6.480 248.450 10.330 248.600 ;
        RECT 10.030 248.000 10.330 248.450 ;
        RECT 6.480 247.850 10.330 248.000 ;
        RECT 10.030 247.400 10.330 247.850 ;
        RECT 6.480 247.250 10.330 247.400 ;
        RECT 10.030 246.800 10.330 247.250 ;
        RECT 6.480 246.650 10.330 246.800 ;
        RECT 10.030 246.200 10.330 246.650 ;
        RECT 6.480 246.050 10.330 246.200 ;
        RECT 10.030 245.600 10.330 246.050 ;
        RECT 6.480 245.450 10.330 245.600 ;
        RECT 10.030 245.000 10.330 245.450 ;
        RECT 6.480 244.850 10.330 245.000 ;
        RECT 10.030 244.400 10.330 244.850 ;
        RECT 6.480 244.250 10.330 244.400 ;
        RECT 10.030 243.800 10.330 244.250 ;
        RECT 6.480 243.650 10.330 243.800 ;
        RECT 10.030 243.200 10.330 243.650 ;
        RECT 6.480 243.050 10.330 243.200 ;
        RECT 10.030 242.600 10.330 243.050 ;
        RECT 6.480 242.450 10.330 242.600 ;
        RECT 10.030 242.000 10.330 242.450 ;
        RECT 6.530 241.450 10.330 242.000 ;
        RECT 10.780 241.450 10.930 249.650 ;
        RECT 11.380 241.450 11.530 249.650 ;
        RECT 11.980 241.450 12.130 249.650 ;
        RECT 12.580 241.450 12.730 249.650 ;
        RECT 13.180 241.450 13.330 249.650 ;
        RECT 13.780 241.450 13.930 249.650 ;
        RECT 14.380 241.450 15.080 258.550 ;
        RECT 15.530 250.350 15.680 258.550 ;
        RECT 16.130 250.350 16.280 258.550 ;
        RECT 16.730 250.350 16.880 258.550 ;
        RECT 17.330 250.350 17.480 258.550 ;
        RECT 17.930 250.350 18.080 258.550 ;
        RECT 18.530 250.350 18.680 258.550 ;
        RECT 19.130 258.000 22.930 258.550 ;
        RECT 26.530 258.550 42.930 258.600 ;
        RECT 26.530 258.000 30.330 258.550 ;
        RECT 19.130 257.550 19.430 258.000 ;
        RECT 30.030 257.550 30.330 258.000 ;
        RECT 19.130 257.400 22.980 257.550 ;
        RECT 26.480 257.400 30.330 257.550 ;
        RECT 19.130 256.950 19.430 257.400 ;
        RECT 30.030 256.950 30.330 257.400 ;
        RECT 19.130 256.800 22.980 256.950 ;
        RECT 26.480 256.800 30.330 256.950 ;
        RECT 19.130 256.350 19.430 256.800 ;
        RECT 30.030 256.350 30.330 256.800 ;
        RECT 19.130 256.200 22.980 256.350 ;
        RECT 26.480 256.200 30.330 256.350 ;
        RECT 19.130 255.750 19.430 256.200 ;
        RECT 30.030 255.750 30.330 256.200 ;
        RECT 19.130 255.600 22.980 255.750 ;
        RECT 26.480 255.600 30.330 255.750 ;
        RECT 19.130 255.150 19.430 255.600 ;
        RECT 30.030 255.150 30.330 255.600 ;
        RECT 19.130 255.000 22.980 255.150 ;
        RECT 26.480 255.000 30.330 255.150 ;
        RECT 19.130 254.550 19.430 255.000 ;
        RECT 30.030 254.550 30.330 255.000 ;
        RECT 19.130 254.400 22.980 254.550 ;
        RECT 26.480 254.400 30.330 254.550 ;
        RECT 19.130 253.950 19.430 254.400 ;
        RECT 30.030 253.950 30.330 254.400 ;
        RECT 19.130 253.800 22.980 253.950 ;
        RECT 26.480 253.800 30.330 253.950 ;
        RECT 19.130 253.350 19.430 253.800 ;
        RECT 30.030 253.350 30.330 253.800 ;
        RECT 19.130 253.200 22.980 253.350 ;
        RECT 26.480 253.200 30.330 253.350 ;
        RECT 19.130 252.750 19.430 253.200 ;
        RECT 19.130 252.600 22.980 252.750 ;
        RECT 19.130 252.150 19.430 252.600 ;
        RECT 19.130 252.000 22.980 252.150 ;
        RECT 19.130 251.550 19.430 252.000 ;
        RECT 19.130 251.400 22.980 251.550 ;
        RECT 19.130 250.950 19.430 251.400 ;
        RECT 19.130 250.800 22.980 250.950 ;
        RECT 19.130 250.350 19.430 250.800 ;
        RECT 15.530 241.450 15.680 249.650 ;
        RECT 16.130 241.450 16.280 249.650 ;
        RECT 16.730 241.450 16.880 249.650 ;
        RECT 17.330 241.450 17.480 249.650 ;
        RECT 17.930 241.450 18.080 249.650 ;
        RECT 18.530 241.450 18.680 249.650 ;
        RECT 19.130 249.200 19.430 249.650 ;
        RECT 19.130 249.050 22.980 249.200 ;
        RECT 19.130 248.600 19.430 249.050 ;
        RECT 19.130 248.450 22.980 248.600 ;
        RECT 19.130 248.000 19.430 248.450 ;
        RECT 19.130 247.850 22.980 248.000 ;
        RECT 19.130 247.400 19.430 247.850 ;
        RECT 19.130 247.250 22.980 247.400 ;
        RECT 19.130 246.800 19.430 247.250 ;
        RECT 23.830 246.800 25.630 253.200 ;
        RECT 30.030 252.750 30.330 253.200 ;
        RECT 26.480 252.600 30.330 252.750 ;
        RECT 30.030 252.150 30.330 252.600 ;
        RECT 26.480 252.000 30.330 252.150 ;
        RECT 30.030 251.550 30.330 252.000 ;
        RECT 26.480 251.400 30.330 251.550 ;
        RECT 30.030 250.950 30.330 251.400 ;
        RECT 26.480 250.800 30.330 250.950 ;
        RECT 30.030 250.350 30.330 250.800 ;
        RECT 30.780 250.350 30.930 258.550 ;
        RECT 31.380 250.350 31.530 258.550 ;
        RECT 31.980 250.350 32.130 258.550 ;
        RECT 32.580 250.350 32.730 258.550 ;
        RECT 33.180 250.350 33.330 258.550 ;
        RECT 33.780 250.350 33.930 258.550 ;
        RECT 30.030 249.200 30.330 249.650 ;
        RECT 26.480 249.050 30.330 249.200 ;
        RECT 30.030 248.600 30.330 249.050 ;
        RECT 26.480 248.450 30.330 248.600 ;
        RECT 30.030 248.000 30.330 248.450 ;
        RECT 26.480 247.850 30.330 248.000 ;
        RECT 30.030 247.400 30.330 247.850 ;
        RECT 26.480 247.250 30.330 247.400 ;
        RECT 30.030 246.800 30.330 247.250 ;
        RECT 19.130 246.650 22.980 246.800 ;
        RECT 26.480 246.650 30.330 246.800 ;
        RECT 19.130 246.200 19.430 246.650 ;
        RECT 30.030 246.200 30.330 246.650 ;
        RECT 19.130 246.050 22.980 246.200 ;
        RECT 26.480 246.050 30.330 246.200 ;
        RECT 19.130 245.600 19.430 246.050 ;
        RECT 30.030 245.600 30.330 246.050 ;
        RECT 19.130 245.450 22.980 245.600 ;
        RECT 26.480 245.450 30.330 245.600 ;
        RECT 19.130 245.000 19.430 245.450 ;
        RECT 30.030 245.000 30.330 245.450 ;
        RECT 19.130 244.850 22.980 245.000 ;
        RECT 26.480 244.850 30.330 245.000 ;
        RECT 19.130 244.400 19.430 244.850 ;
        RECT 30.030 244.400 30.330 244.850 ;
        RECT 19.130 244.250 22.980 244.400 ;
        RECT 26.480 244.250 30.330 244.400 ;
        RECT 19.130 243.800 19.430 244.250 ;
        RECT 30.030 243.800 30.330 244.250 ;
        RECT 19.130 243.650 22.980 243.800 ;
        RECT 26.480 243.650 30.330 243.800 ;
        RECT 19.130 243.200 19.430 243.650 ;
        RECT 30.030 243.200 30.330 243.650 ;
        RECT 19.130 243.050 22.980 243.200 ;
        RECT 26.480 243.050 30.330 243.200 ;
        RECT 19.130 242.600 19.430 243.050 ;
        RECT 30.030 242.600 30.330 243.050 ;
        RECT 19.130 242.450 22.980 242.600 ;
        RECT 26.480 242.450 30.330 242.600 ;
        RECT 19.130 242.000 19.430 242.450 ;
        RECT 30.030 242.000 30.330 242.450 ;
        RECT 19.130 241.450 22.930 242.000 ;
        RECT 6.530 241.400 22.930 241.450 ;
        RECT 26.530 241.450 30.330 242.000 ;
        RECT 30.780 241.450 30.930 249.650 ;
        RECT 31.380 241.450 31.530 249.650 ;
        RECT 31.980 241.450 32.130 249.650 ;
        RECT 32.580 241.450 32.730 249.650 ;
        RECT 33.180 241.450 33.330 249.650 ;
        RECT 33.780 241.450 33.930 249.650 ;
        RECT 34.380 241.450 35.080 258.550 ;
        RECT 35.530 250.350 35.680 258.550 ;
        RECT 36.130 250.350 36.280 258.550 ;
        RECT 36.730 250.350 36.880 258.550 ;
        RECT 37.330 250.350 37.480 258.550 ;
        RECT 37.930 250.350 38.080 258.550 ;
        RECT 38.530 250.350 38.680 258.550 ;
        RECT 39.130 258.000 42.930 258.550 ;
        RECT 46.530 258.550 62.930 258.600 ;
        RECT 46.530 258.000 50.330 258.550 ;
        RECT 39.130 257.550 39.430 258.000 ;
        RECT 50.030 257.550 50.330 258.000 ;
        RECT 39.130 257.400 42.980 257.550 ;
        RECT 46.480 257.400 50.330 257.550 ;
        RECT 39.130 256.950 39.430 257.400 ;
        RECT 50.030 256.950 50.330 257.400 ;
        RECT 39.130 256.800 42.980 256.950 ;
        RECT 46.480 256.800 50.330 256.950 ;
        RECT 39.130 256.350 39.430 256.800 ;
        RECT 50.030 256.350 50.330 256.800 ;
        RECT 39.130 256.200 42.980 256.350 ;
        RECT 46.480 256.200 50.330 256.350 ;
        RECT 39.130 255.750 39.430 256.200 ;
        RECT 50.030 255.750 50.330 256.200 ;
        RECT 39.130 255.600 42.980 255.750 ;
        RECT 46.480 255.600 50.330 255.750 ;
        RECT 39.130 255.150 39.430 255.600 ;
        RECT 50.030 255.150 50.330 255.600 ;
        RECT 39.130 255.000 42.980 255.150 ;
        RECT 46.480 255.000 50.330 255.150 ;
        RECT 39.130 254.550 39.430 255.000 ;
        RECT 50.030 254.550 50.330 255.000 ;
        RECT 39.130 254.400 42.980 254.550 ;
        RECT 46.480 254.400 50.330 254.550 ;
        RECT 39.130 253.950 39.430 254.400 ;
        RECT 50.030 253.950 50.330 254.400 ;
        RECT 39.130 253.800 42.980 253.950 ;
        RECT 46.480 253.800 50.330 253.950 ;
        RECT 39.130 253.350 39.430 253.800 ;
        RECT 50.030 253.350 50.330 253.800 ;
        RECT 39.130 253.200 42.980 253.350 ;
        RECT 46.480 253.200 50.330 253.350 ;
        RECT 39.130 252.750 39.430 253.200 ;
        RECT 39.130 252.600 42.980 252.750 ;
        RECT 39.130 252.150 39.430 252.600 ;
        RECT 39.130 252.000 42.980 252.150 ;
        RECT 39.130 251.550 39.430 252.000 ;
        RECT 39.130 251.400 42.980 251.550 ;
        RECT 39.130 250.950 39.430 251.400 ;
        RECT 39.130 250.800 42.980 250.950 ;
        RECT 39.130 250.350 39.430 250.800 ;
        RECT 35.530 241.450 35.680 249.650 ;
        RECT 36.130 241.450 36.280 249.650 ;
        RECT 36.730 241.450 36.880 249.650 ;
        RECT 37.330 241.450 37.480 249.650 ;
        RECT 37.930 241.450 38.080 249.650 ;
        RECT 38.530 241.450 38.680 249.650 ;
        RECT 39.130 249.200 39.430 249.650 ;
        RECT 39.130 249.050 42.980 249.200 ;
        RECT 39.130 248.600 39.430 249.050 ;
        RECT 39.130 248.450 42.980 248.600 ;
        RECT 39.130 248.000 39.430 248.450 ;
        RECT 39.130 247.850 42.980 248.000 ;
        RECT 39.130 247.400 39.430 247.850 ;
        RECT 39.130 247.250 42.980 247.400 ;
        RECT 39.130 246.800 39.430 247.250 ;
        RECT 43.830 246.800 45.630 253.200 ;
        RECT 50.030 252.750 50.330 253.200 ;
        RECT 46.480 252.600 50.330 252.750 ;
        RECT 50.030 252.150 50.330 252.600 ;
        RECT 46.480 252.000 50.330 252.150 ;
        RECT 50.030 251.550 50.330 252.000 ;
        RECT 46.480 251.400 50.330 251.550 ;
        RECT 50.030 250.950 50.330 251.400 ;
        RECT 46.480 250.800 50.330 250.950 ;
        RECT 50.030 250.350 50.330 250.800 ;
        RECT 50.780 250.350 50.930 258.550 ;
        RECT 51.380 250.350 51.530 258.550 ;
        RECT 51.980 250.350 52.130 258.550 ;
        RECT 52.580 250.350 52.730 258.550 ;
        RECT 53.180 250.350 53.330 258.550 ;
        RECT 53.780 250.350 53.930 258.550 ;
        RECT 50.030 249.200 50.330 249.650 ;
        RECT 46.480 249.050 50.330 249.200 ;
        RECT 50.030 248.600 50.330 249.050 ;
        RECT 46.480 248.450 50.330 248.600 ;
        RECT 50.030 248.000 50.330 248.450 ;
        RECT 46.480 247.850 50.330 248.000 ;
        RECT 50.030 247.400 50.330 247.850 ;
        RECT 46.480 247.250 50.330 247.400 ;
        RECT 50.030 246.800 50.330 247.250 ;
        RECT 39.130 246.650 42.980 246.800 ;
        RECT 46.480 246.650 50.330 246.800 ;
        RECT 39.130 246.200 39.430 246.650 ;
        RECT 50.030 246.200 50.330 246.650 ;
        RECT 39.130 246.050 42.980 246.200 ;
        RECT 46.480 246.050 50.330 246.200 ;
        RECT 39.130 245.600 39.430 246.050 ;
        RECT 50.030 245.600 50.330 246.050 ;
        RECT 39.130 245.450 42.980 245.600 ;
        RECT 46.480 245.450 50.330 245.600 ;
        RECT 39.130 245.000 39.430 245.450 ;
        RECT 50.030 245.000 50.330 245.450 ;
        RECT 39.130 244.850 42.980 245.000 ;
        RECT 46.480 244.850 50.330 245.000 ;
        RECT 39.130 244.400 39.430 244.850 ;
        RECT 50.030 244.400 50.330 244.850 ;
        RECT 39.130 244.250 42.980 244.400 ;
        RECT 46.480 244.250 50.330 244.400 ;
        RECT 39.130 243.800 39.430 244.250 ;
        RECT 50.030 243.800 50.330 244.250 ;
        RECT 39.130 243.650 42.980 243.800 ;
        RECT 46.480 243.650 50.330 243.800 ;
        RECT 39.130 243.200 39.430 243.650 ;
        RECT 50.030 243.200 50.330 243.650 ;
        RECT 39.130 243.050 42.980 243.200 ;
        RECT 46.480 243.050 50.330 243.200 ;
        RECT 39.130 242.600 39.430 243.050 ;
        RECT 50.030 242.600 50.330 243.050 ;
        RECT 39.130 242.450 42.980 242.600 ;
        RECT 46.480 242.450 50.330 242.600 ;
        RECT 39.130 242.000 39.430 242.450 ;
        RECT 50.030 242.000 50.330 242.450 ;
        RECT 39.130 241.450 42.930 242.000 ;
        RECT 26.530 241.400 42.930 241.450 ;
        RECT 46.530 241.450 50.330 242.000 ;
        RECT 50.780 241.450 50.930 249.650 ;
        RECT 51.380 241.450 51.530 249.650 ;
        RECT 51.980 241.450 52.130 249.650 ;
        RECT 52.580 241.450 52.730 249.650 ;
        RECT 53.180 241.450 53.330 249.650 ;
        RECT 53.780 241.450 53.930 249.650 ;
        RECT 54.380 241.450 55.080 258.550 ;
        RECT 55.530 250.350 55.680 258.550 ;
        RECT 56.130 250.350 56.280 258.550 ;
        RECT 56.730 250.350 56.880 258.550 ;
        RECT 57.330 250.350 57.480 258.550 ;
        RECT 57.930 250.350 58.080 258.550 ;
        RECT 58.530 250.350 58.680 258.550 ;
        RECT 59.130 258.000 62.930 258.550 ;
        RECT 66.530 258.550 82.930 258.600 ;
        RECT 66.530 258.000 70.330 258.550 ;
        RECT 59.130 257.550 59.430 258.000 ;
        RECT 70.030 257.550 70.330 258.000 ;
        RECT 59.130 257.400 62.980 257.550 ;
        RECT 66.480 257.400 70.330 257.550 ;
        RECT 59.130 256.950 59.430 257.400 ;
        RECT 70.030 256.950 70.330 257.400 ;
        RECT 59.130 256.800 62.980 256.950 ;
        RECT 66.480 256.800 70.330 256.950 ;
        RECT 59.130 256.350 59.430 256.800 ;
        RECT 70.030 256.350 70.330 256.800 ;
        RECT 59.130 256.200 62.980 256.350 ;
        RECT 66.480 256.200 70.330 256.350 ;
        RECT 59.130 255.750 59.430 256.200 ;
        RECT 70.030 255.750 70.330 256.200 ;
        RECT 59.130 255.600 62.980 255.750 ;
        RECT 66.480 255.600 70.330 255.750 ;
        RECT 59.130 255.150 59.430 255.600 ;
        RECT 70.030 255.150 70.330 255.600 ;
        RECT 59.130 255.000 62.980 255.150 ;
        RECT 66.480 255.000 70.330 255.150 ;
        RECT 59.130 254.550 59.430 255.000 ;
        RECT 70.030 254.550 70.330 255.000 ;
        RECT 59.130 254.400 62.980 254.550 ;
        RECT 66.480 254.400 70.330 254.550 ;
        RECT 59.130 253.950 59.430 254.400 ;
        RECT 70.030 253.950 70.330 254.400 ;
        RECT 59.130 253.800 62.980 253.950 ;
        RECT 66.480 253.800 70.330 253.950 ;
        RECT 59.130 253.350 59.430 253.800 ;
        RECT 70.030 253.350 70.330 253.800 ;
        RECT 59.130 253.200 62.980 253.350 ;
        RECT 66.480 253.200 70.330 253.350 ;
        RECT 59.130 252.750 59.430 253.200 ;
        RECT 59.130 252.600 62.980 252.750 ;
        RECT 59.130 252.150 59.430 252.600 ;
        RECT 59.130 252.000 62.980 252.150 ;
        RECT 59.130 251.550 59.430 252.000 ;
        RECT 59.130 251.400 62.980 251.550 ;
        RECT 59.130 250.950 59.430 251.400 ;
        RECT 59.130 250.800 62.980 250.950 ;
        RECT 59.130 250.350 59.430 250.800 ;
        RECT 55.530 241.450 55.680 249.650 ;
        RECT 56.130 241.450 56.280 249.650 ;
        RECT 56.730 241.450 56.880 249.650 ;
        RECT 57.330 241.450 57.480 249.650 ;
        RECT 57.930 241.450 58.080 249.650 ;
        RECT 58.530 241.450 58.680 249.650 ;
        RECT 59.130 249.200 59.430 249.650 ;
        RECT 59.130 249.050 62.980 249.200 ;
        RECT 59.130 248.600 59.430 249.050 ;
        RECT 59.130 248.450 62.980 248.600 ;
        RECT 59.130 248.000 59.430 248.450 ;
        RECT 59.130 247.850 62.980 248.000 ;
        RECT 59.130 247.400 59.430 247.850 ;
        RECT 59.130 247.250 62.980 247.400 ;
        RECT 59.130 246.800 59.430 247.250 ;
        RECT 63.830 246.800 65.630 253.200 ;
        RECT 70.030 252.750 70.330 253.200 ;
        RECT 66.480 252.600 70.330 252.750 ;
        RECT 70.030 252.150 70.330 252.600 ;
        RECT 66.480 252.000 70.330 252.150 ;
        RECT 70.030 251.550 70.330 252.000 ;
        RECT 66.480 251.400 70.330 251.550 ;
        RECT 70.030 250.950 70.330 251.400 ;
        RECT 66.480 250.800 70.330 250.950 ;
        RECT 70.030 250.350 70.330 250.800 ;
        RECT 70.780 250.350 70.930 258.550 ;
        RECT 71.380 250.350 71.530 258.550 ;
        RECT 71.980 250.350 72.130 258.550 ;
        RECT 72.580 250.350 72.730 258.550 ;
        RECT 73.180 250.350 73.330 258.550 ;
        RECT 73.780 250.350 73.930 258.550 ;
        RECT 70.030 249.200 70.330 249.650 ;
        RECT 66.480 249.050 70.330 249.200 ;
        RECT 70.030 248.600 70.330 249.050 ;
        RECT 66.480 248.450 70.330 248.600 ;
        RECT 70.030 248.000 70.330 248.450 ;
        RECT 66.480 247.850 70.330 248.000 ;
        RECT 70.030 247.400 70.330 247.850 ;
        RECT 66.480 247.250 70.330 247.400 ;
        RECT 70.030 246.800 70.330 247.250 ;
        RECT 59.130 246.650 62.980 246.800 ;
        RECT 66.480 246.650 70.330 246.800 ;
        RECT 59.130 246.200 59.430 246.650 ;
        RECT 70.030 246.200 70.330 246.650 ;
        RECT 59.130 246.050 62.980 246.200 ;
        RECT 66.480 246.050 70.330 246.200 ;
        RECT 59.130 245.600 59.430 246.050 ;
        RECT 70.030 245.600 70.330 246.050 ;
        RECT 59.130 245.450 62.980 245.600 ;
        RECT 66.480 245.450 70.330 245.600 ;
        RECT 59.130 245.000 59.430 245.450 ;
        RECT 70.030 245.000 70.330 245.450 ;
        RECT 59.130 244.850 62.980 245.000 ;
        RECT 66.480 244.850 70.330 245.000 ;
        RECT 59.130 244.400 59.430 244.850 ;
        RECT 70.030 244.400 70.330 244.850 ;
        RECT 59.130 244.250 62.980 244.400 ;
        RECT 66.480 244.250 70.330 244.400 ;
        RECT 59.130 243.800 59.430 244.250 ;
        RECT 70.030 243.800 70.330 244.250 ;
        RECT 59.130 243.650 62.980 243.800 ;
        RECT 66.480 243.650 70.330 243.800 ;
        RECT 59.130 243.200 59.430 243.650 ;
        RECT 70.030 243.200 70.330 243.650 ;
        RECT 59.130 243.050 62.980 243.200 ;
        RECT 66.480 243.050 70.330 243.200 ;
        RECT 59.130 242.600 59.430 243.050 ;
        RECT 70.030 242.600 70.330 243.050 ;
        RECT 59.130 242.450 62.980 242.600 ;
        RECT 66.480 242.450 70.330 242.600 ;
        RECT 59.130 242.000 59.430 242.450 ;
        RECT 70.030 242.000 70.330 242.450 ;
        RECT 59.130 241.450 62.930 242.000 ;
        RECT 46.530 241.400 62.930 241.450 ;
        RECT 66.530 241.450 70.330 242.000 ;
        RECT 70.780 241.450 70.930 249.650 ;
        RECT 71.380 241.450 71.530 249.650 ;
        RECT 71.980 241.450 72.130 249.650 ;
        RECT 72.580 241.450 72.730 249.650 ;
        RECT 73.180 241.450 73.330 249.650 ;
        RECT 73.780 241.450 73.930 249.650 ;
        RECT 74.380 241.450 75.080 258.550 ;
        RECT 75.530 250.350 75.680 258.550 ;
        RECT 76.130 250.350 76.280 258.550 ;
        RECT 76.730 250.350 76.880 258.550 ;
        RECT 77.330 250.350 77.480 258.550 ;
        RECT 77.930 250.350 78.080 258.550 ;
        RECT 78.530 250.350 78.680 258.550 ;
        RECT 79.130 258.000 82.930 258.550 ;
        RECT 86.530 258.550 102.930 258.600 ;
        RECT 86.530 258.000 90.330 258.550 ;
        RECT 79.130 257.550 79.430 258.000 ;
        RECT 90.030 257.550 90.330 258.000 ;
        RECT 79.130 257.400 82.980 257.550 ;
        RECT 86.480 257.400 90.330 257.550 ;
        RECT 79.130 256.950 79.430 257.400 ;
        RECT 90.030 256.950 90.330 257.400 ;
        RECT 79.130 256.800 82.980 256.950 ;
        RECT 86.480 256.800 90.330 256.950 ;
        RECT 79.130 256.350 79.430 256.800 ;
        RECT 90.030 256.350 90.330 256.800 ;
        RECT 79.130 256.200 82.980 256.350 ;
        RECT 86.480 256.200 90.330 256.350 ;
        RECT 79.130 255.750 79.430 256.200 ;
        RECT 90.030 255.750 90.330 256.200 ;
        RECT 79.130 255.600 82.980 255.750 ;
        RECT 86.480 255.600 90.330 255.750 ;
        RECT 79.130 255.150 79.430 255.600 ;
        RECT 90.030 255.150 90.330 255.600 ;
        RECT 79.130 255.000 82.980 255.150 ;
        RECT 86.480 255.000 90.330 255.150 ;
        RECT 79.130 254.550 79.430 255.000 ;
        RECT 90.030 254.550 90.330 255.000 ;
        RECT 79.130 254.400 82.980 254.550 ;
        RECT 86.480 254.400 90.330 254.550 ;
        RECT 79.130 253.950 79.430 254.400 ;
        RECT 90.030 253.950 90.330 254.400 ;
        RECT 79.130 253.800 82.980 253.950 ;
        RECT 86.480 253.800 90.330 253.950 ;
        RECT 79.130 253.350 79.430 253.800 ;
        RECT 90.030 253.350 90.330 253.800 ;
        RECT 79.130 253.200 82.980 253.350 ;
        RECT 86.480 253.200 90.330 253.350 ;
        RECT 79.130 252.750 79.430 253.200 ;
        RECT 79.130 252.600 82.980 252.750 ;
        RECT 79.130 252.150 79.430 252.600 ;
        RECT 79.130 252.000 82.980 252.150 ;
        RECT 79.130 251.550 79.430 252.000 ;
        RECT 79.130 251.400 82.980 251.550 ;
        RECT 79.130 250.950 79.430 251.400 ;
        RECT 79.130 250.800 82.980 250.950 ;
        RECT 79.130 250.350 79.430 250.800 ;
        RECT 75.530 241.450 75.680 249.650 ;
        RECT 76.130 241.450 76.280 249.650 ;
        RECT 76.730 241.450 76.880 249.650 ;
        RECT 77.330 241.450 77.480 249.650 ;
        RECT 77.930 241.450 78.080 249.650 ;
        RECT 78.530 241.450 78.680 249.650 ;
        RECT 79.130 249.200 79.430 249.650 ;
        RECT 79.130 249.050 82.980 249.200 ;
        RECT 79.130 248.600 79.430 249.050 ;
        RECT 79.130 248.450 82.980 248.600 ;
        RECT 79.130 248.000 79.430 248.450 ;
        RECT 79.130 247.850 82.980 248.000 ;
        RECT 79.130 247.400 79.430 247.850 ;
        RECT 79.130 247.250 82.980 247.400 ;
        RECT 79.130 246.800 79.430 247.250 ;
        RECT 83.830 246.800 85.630 253.200 ;
        RECT 90.030 252.750 90.330 253.200 ;
        RECT 86.480 252.600 90.330 252.750 ;
        RECT 90.030 252.150 90.330 252.600 ;
        RECT 86.480 252.000 90.330 252.150 ;
        RECT 90.030 251.550 90.330 252.000 ;
        RECT 86.480 251.400 90.330 251.550 ;
        RECT 90.030 250.950 90.330 251.400 ;
        RECT 86.480 250.800 90.330 250.950 ;
        RECT 90.030 250.350 90.330 250.800 ;
        RECT 90.780 250.350 90.930 258.550 ;
        RECT 91.380 250.350 91.530 258.550 ;
        RECT 91.980 250.350 92.130 258.550 ;
        RECT 92.580 250.350 92.730 258.550 ;
        RECT 93.180 250.350 93.330 258.550 ;
        RECT 93.780 250.350 93.930 258.550 ;
        RECT 90.030 249.200 90.330 249.650 ;
        RECT 86.480 249.050 90.330 249.200 ;
        RECT 90.030 248.600 90.330 249.050 ;
        RECT 86.480 248.450 90.330 248.600 ;
        RECT 90.030 248.000 90.330 248.450 ;
        RECT 86.480 247.850 90.330 248.000 ;
        RECT 90.030 247.400 90.330 247.850 ;
        RECT 86.480 247.250 90.330 247.400 ;
        RECT 90.030 246.800 90.330 247.250 ;
        RECT 79.130 246.650 82.980 246.800 ;
        RECT 86.480 246.650 90.330 246.800 ;
        RECT 79.130 246.200 79.430 246.650 ;
        RECT 90.030 246.200 90.330 246.650 ;
        RECT 79.130 246.050 82.980 246.200 ;
        RECT 86.480 246.050 90.330 246.200 ;
        RECT 79.130 245.600 79.430 246.050 ;
        RECT 90.030 245.600 90.330 246.050 ;
        RECT 79.130 245.450 82.980 245.600 ;
        RECT 86.480 245.450 90.330 245.600 ;
        RECT 79.130 245.000 79.430 245.450 ;
        RECT 90.030 245.000 90.330 245.450 ;
        RECT 79.130 244.850 82.980 245.000 ;
        RECT 86.480 244.850 90.330 245.000 ;
        RECT 79.130 244.400 79.430 244.850 ;
        RECT 90.030 244.400 90.330 244.850 ;
        RECT 79.130 244.250 82.980 244.400 ;
        RECT 86.480 244.250 90.330 244.400 ;
        RECT 79.130 243.800 79.430 244.250 ;
        RECT 90.030 243.800 90.330 244.250 ;
        RECT 79.130 243.650 82.980 243.800 ;
        RECT 86.480 243.650 90.330 243.800 ;
        RECT 79.130 243.200 79.430 243.650 ;
        RECT 90.030 243.200 90.330 243.650 ;
        RECT 79.130 243.050 82.980 243.200 ;
        RECT 86.480 243.050 90.330 243.200 ;
        RECT 79.130 242.600 79.430 243.050 ;
        RECT 90.030 242.600 90.330 243.050 ;
        RECT 79.130 242.450 82.980 242.600 ;
        RECT 86.480 242.450 90.330 242.600 ;
        RECT 79.130 242.000 79.430 242.450 ;
        RECT 90.030 242.000 90.330 242.450 ;
        RECT 79.130 241.450 82.930 242.000 ;
        RECT 66.530 241.400 82.930 241.450 ;
        RECT 86.530 241.450 90.330 242.000 ;
        RECT 90.780 241.450 90.930 249.650 ;
        RECT 91.380 241.450 91.530 249.650 ;
        RECT 91.980 241.450 92.130 249.650 ;
        RECT 92.580 241.450 92.730 249.650 ;
        RECT 93.180 241.450 93.330 249.650 ;
        RECT 93.780 241.450 93.930 249.650 ;
        RECT 94.380 241.450 95.080 258.550 ;
        RECT 95.530 250.350 95.680 258.550 ;
        RECT 96.130 250.350 96.280 258.550 ;
        RECT 96.730 250.350 96.880 258.550 ;
        RECT 97.330 250.350 97.480 258.550 ;
        RECT 97.930 250.350 98.080 258.550 ;
        RECT 98.530 250.350 98.680 258.550 ;
        RECT 99.130 258.000 102.930 258.550 ;
        RECT 106.530 258.550 122.930 258.600 ;
        RECT 106.530 258.000 110.330 258.550 ;
        RECT 99.130 257.550 99.430 258.000 ;
        RECT 110.030 257.550 110.330 258.000 ;
        RECT 99.130 257.400 102.980 257.550 ;
        RECT 106.480 257.400 110.330 257.550 ;
        RECT 99.130 256.950 99.430 257.400 ;
        RECT 110.030 256.950 110.330 257.400 ;
        RECT 99.130 256.800 102.980 256.950 ;
        RECT 106.480 256.800 110.330 256.950 ;
        RECT 99.130 256.350 99.430 256.800 ;
        RECT 110.030 256.350 110.330 256.800 ;
        RECT 99.130 256.200 102.980 256.350 ;
        RECT 106.480 256.200 110.330 256.350 ;
        RECT 99.130 255.750 99.430 256.200 ;
        RECT 110.030 255.750 110.330 256.200 ;
        RECT 99.130 255.600 102.980 255.750 ;
        RECT 106.480 255.600 110.330 255.750 ;
        RECT 99.130 255.150 99.430 255.600 ;
        RECT 110.030 255.150 110.330 255.600 ;
        RECT 99.130 255.000 102.980 255.150 ;
        RECT 106.480 255.000 110.330 255.150 ;
        RECT 99.130 254.550 99.430 255.000 ;
        RECT 110.030 254.550 110.330 255.000 ;
        RECT 99.130 254.400 102.980 254.550 ;
        RECT 106.480 254.400 110.330 254.550 ;
        RECT 99.130 253.950 99.430 254.400 ;
        RECT 110.030 253.950 110.330 254.400 ;
        RECT 99.130 253.800 102.980 253.950 ;
        RECT 106.480 253.800 110.330 253.950 ;
        RECT 99.130 253.350 99.430 253.800 ;
        RECT 110.030 253.350 110.330 253.800 ;
        RECT 99.130 253.200 102.980 253.350 ;
        RECT 106.480 253.200 110.330 253.350 ;
        RECT 99.130 252.750 99.430 253.200 ;
        RECT 99.130 252.600 102.980 252.750 ;
        RECT 99.130 252.150 99.430 252.600 ;
        RECT 99.130 252.000 102.980 252.150 ;
        RECT 99.130 251.550 99.430 252.000 ;
        RECT 99.130 251.400 102.980 251.550 ;
        RECT 99.130 250.950 99.430 251.400 ;
        RECT 99.130 250.800 102.980 250.950 ;
        RECT 99.130 250.350 99.430 250.800 ;
        RECT 95.530 241.450 95.680 249.650 ;
        RECT 96.130 241.450 96.280 249.650 ;
        RECT 96.730 241.450 96.880 249.650 ;
        RECT 97.330 241.450 97.480 249.650 ;
        RECT 97.930 241.450 98.080 249.650 ;
        RECT 98.530 241.450 98.680 249.650 ;
        RECT 99.130 249.200 99.430 249.650 ;
        RECT 99.130 249.050 102.980 249.200 ;
        RECT 99.130 248.600 99.430 249.050 ;
        RECT 99.130 248.450 102.980 248.600 ;
        RECT 99.130 248.000 99.430 248.450 ;
        RECT 99.130 247.850 102.980 248.000 ;
        RECT 99.130 247.400 99.430 247.850 ;
        RECT 99.130 247.250 102.980 247.400 ;
        RECT 99.130 246.800 99.430 247.250 ;
        RECT 103.830 246.800 105.630 253.200 ;
        RECT 110.030 252.750 110.330 253.200 ;
        RECT 106.480 252.600 110.330 252.750 ;
        RECT 110.030 252.150 110.330 252.600 ;
        RECT 106.480 252.000 110.330 252.150 ;
        RECT 110.030 251.550 110.330 252.000 ;
        RECT 106.480 251.400 110.330 251.550 ;
        RECT 110.030 250.950 110.330 251.400 ;
        RECT 106.480 250.800 110.330 250.950 ;
        RECT 110.030 250.350 110.330 250.800 ;
        RECT 110.780 250.350 110.930 258.550 ;
        RECT 111.380 250.350 111.530 258.550 ;
        RECT 111.980 250.350 112.130 258.550 ;
        RECT 112.580 250.350 112.730 258.550 ;
        RECT 113.180 250.350 113.330 258.550 ;
        RECT 113.780 250.350 113.930 258.550 ;
        RECT 110.030 249.200 110.330 249.650 ;
        RECT 106.480 249.050 110.330 249.200 ;
        RECT 110.030 248.600 110.330 249.050 ;
        RECT 106.480 248.450 110.330 248.600 ;
        RECT 110.030 248.000 110.330 248.450 ;
        RECT 106.480 247.850 110.330 248.000 ;
        RECT 110.030 247.400 110.330 247.850 ;
        RECT 106.480 247.250 110.330 247.400 ;
        RECT 110.030 246.800 110.330 247.250 ;
        RECT 99.130 246.650 102.980 246.800 ;
        RECT 106.480 246.650 110.330 246.800 ;
        RECT 99.130 246.200 99.430 246.650 ;
        RECT 110.030 246.200 110.330 246.650 ;
        RECT 99.130 246.050 102.980 246.200 ;
        RECT 106.480 246.050 110.330 246.200 ;
        RECT 99.130 245.600 99.430 246.050 ;
        RECT 110.030 245.600 110.330 246.050 ;
        RECT 99.130 245.450 102.980 245.600 ;
        RECT 106.480 245.450 110.330 245.600 ;
        RECT 99.130 245.000 99.430 245.450 ;
        RECT 110.030 245.000 110.330 245.450 ;
        RECT 99.130 244.850 102.980 245.000 ;
        RECT 106.480 244.850 110.330 245.000 ;
        RECT 99.130 244.400 99.430 244.850 ;
        RECT 110.030 244.400 110.330 244.850 ;
        RECT 99.130 244.250 102.980 244.400 ;
        RECT 106.480 244.250 110.330 244.400 ;
        RECT 99.130 243.800 99.430 244.250 ;
        RECT 110.030 243.800 110.330 244.250 ;
        RECT 99.130 243.650 102.980 243.800 ;
        RECT 106.480 243.650 110.330 243.800 ;
        RECT 99.130 243.200 99.430 243.650 ;
        RECT 110.030 243.200 110.330 243.650 ;
        RECT 99.130 243.050 102.980 243.200 ;
        RECT 106.480 243.050 110.330 243.200 ;
        RECT 99.130 242.600 99.430 243.050 ;
        RECT 110.030 242.600 110.330 243.050 ;
        RECT 99.130 242.450 102.980 242.600 ;
        RECT 106.480 242.450 110.330 242.600 ;
        RECT 99.130 242.000 99.430 242.450 ;
        RECT 110.030 242.000 110.330 242.450 ;
        RECT 99.130 241.450 102.930 242.000 ;
        RECT 86.530 241.400 102.930 241.450 ;
        RECT 106.530 241.450 110.330 242.000 ;
        RECT 110.780 241.450 110.930 249.650 ;
        RECT 111.380 241.450 111.530 249.650 ;
        RECT 111.980 241.450 112.130 249.650 ;
        RECT 112.580 241.450 112.730 249.650 ;
        RECT 113.180 241.450 113.330 249.650 ;
        RECT 113.780 241.450 113.930 249.650 ;
        RECT 114.380 241.450 115.080 258.550 ;
        RECT 115.530 250.350 115.680 258.550 ;
        RECT 116.130 250.350 116.280 258.550 ;
        RECT 116.730 250.350 116.880 258.550 ;
        RECT 117.330 250.350 117.480 258.550 ;
        RECT 117.930 250.350 118.080 258.550 ;
        RECT 118.530 250.350 118.680 258.550 ;
        RECT 119.130 258.000 122.930 258.550 ;
        RECT 119.130 257.550 119.430 258.000 ;
        RECT 119.130 257.400 122.980 257.550 ;
        RECT 119.130 256.950 119.430 257.400 ;
        RECT 119.130 256.800 122.980 256.950 ;
        RECT 119.130 256.350 119.430 256.800 ;
        RECT 119.130 256.200 122.980 256.350 ;
        RECT 119.130 255.750 119.430 256.200 ;
        RECT 119.130 255.600 122.980 255.750 ;
        RECT 119.130 255.150 119.430 255.600 ;
        RECT 119.130 255.000 122.980 255.150 ;
        RECT 119.130 254.550 119.430 255.000 ;
        RECT 119.130 254.400 122.980 254.550 ;
        RECT 119.130 253.950 119.430 254.400 ;
        RECT 119.130 253.800 122.980 253.950 ;
        RECT 119.130 253.350 119.430 253.800 ;
        RECT 119.130 253.200 122.980 253.350 ;
        RECT 119.130 252.750 119.430 253.200 ;
        RECT 119.130 252.600 122.980 252.750 ;
        RECT 119.130 252.150 119.430 252.600 ;
        RECT 119.130 252.000 122.980 252.150 ;
        RECT 119.130 251.550 119.430 252.000 ;
        RECT 119.130 251.400 122.980 251.550 ;
        RECT 119.130 250.950 119.430 251.400 ;
        RECT 119.130 250.800 122.980 250.950 ;
        RECT 119.130 250.350 119.430 250.800 ;
        RECT 115.530 241.450 115.680 249.650 ;
        RECT 116.130 241.450 116.280 249.650 ;
        RECT 116.730 241.450 116.880 249.650 ;
        RECT 117.330 241.450 117.480 249.650 ;
        RECT 117.930 241.450 118.080 249.650 ;
        RECT 118.530 241.450 118.680 249.650 ;
        RECT 119.130 249.200 119.430 249.650 ;
        RECT 119.130 249.050 122.980 249.200 ;
        RECT 119.130 248.600 119.430 249.050 ;
        RECT 119.130 248.450 122.980 248.600 ;
        RECT 119.130 248.000 119.430 248.450 ;
        RECT 119.130 247.850 122.980 248.000 ;
        RECT 119.130 247.400 119.430 247.850 ;
        RECT 119.130 247.250 122.980 247.400 ;
        RECT 119.130 246.800 119.430 247.250 ;
        RECT 123.830 246.800 124.730 253.200 ;
        RECT 129.850 249.245 131.850 250.520 ;
        RECT 119.130 246.650 122.980 246.800 ;
        RECT 119.130 246.200 119.430 246.650 ;
        RECT 119.130 246.050 122.980 246.200 ;
        RECT 119.130 245.600 119.430 246.050 ;
        RECT 119.130 245.450 122.980 245.600 ;
        RECT 119.130 245.000 119.430 245.450 ;
        RECT 119.130 244.850 122.980 245.000 ;
        RECT 119.130 244.400 119.430 244.850 ;
        RECT 119.130 244.250 122.980 244.400 ;
        RECT 119.130 243.800 119.430 244.250 ;
        RECT 119.130 243.650 122.980 243.800 ;
        RECT 119.130 243.200 119.430 243.650 ;
        RECT 119.130 243.050 122.980 243.200 ;
        RECT 119.130 242.600 119.430 243.050 ;
        RECT 119.130 242.450 122.980 242.600 ;
        RECT 119.130 242.000 119.430 242.450 ;
        RECT 119.130 241.450 122.930 242.000 ;
        RECT 106.530 241.400 122.930 241.450 ;
        RECT 9.630 240.900 19.830 241.400 ;
        RECT 29.630 240.900 39.830 241.400 ;
        RECT 49.630 240.900 59.830 241.400 ;
        RECT 69.630 240.900 79.830 241.400 ;
        RECT 89.630 240.900 99.830 241.400 ;
        RECT 109.630 240.900 119.830 241.400 ;
        RECT 11.530 239.100 17.930 240.900 ;
        RECT 31.530 239.100 37.930 240.900 ;
        RECT 51.530 239.100 57.930 240.900 ;
        RECT 71.530 239.100 77.930 240.900 ;
        RECT 91.530 239.100 97.930 240.900 ;
        RECT 111.530 239.100 117.930 240.900 ;
        RECT 9.630 238.600 19.830 239.100 ;
        RECT 29.630 238.600 39.830 239.100 ;
        RECT 49.630 238.600 59.830 239.100 ;
        RECT 69.630 238.600 79.830 239.100 ;
        RECT 89.630 238.600 99.830 239.100 ;
        RECT 109.630 238.600 119.830 239.100 ;
        RECT 6.530 238.550 22.930 238.600 ;
        RECT 6.530 238.000 10.330 238.550 ;
        RECT 10.030 237.550 10.330 238.000 ;
        RECT 6.480 237.400 10.330 237.550 ;
        RECT 10.030 236.950 10.330 237.400 ;
        RECT 6.480 236.800 10.330 236.950 ;
        RECT 10.030 236.350 10.330 236.800 ;
        RECT 6.480 236.200 10.330 236.350 ;
        RECT 10.030 235.750 10.330 236.200 ;
        RECT 6.480 235.600 10.330 235.750 ;
        RECT 10.030 235.150 10.330 235.600 ;
        RECT 6.480 235.000 10.330 235.150 ;
        RECT 10.030 234.550 10.330 235.000 ;
        RECT 6.480 234.400 10.330 234.550 ;
        RECT 10.030 233.950 10.330 234.400 ;
        RECT 6.480 233.800 10.330 233.950 ;
        RECT 10.030 233.350 10.330 233.800 ;
        RECT 6.480 233.200 10.330 233.350 ;
        RECT 4.730 226.800 5.630 233.200 ;
        RECT 10.030 232.750 10.330 233.200 ;
        RECT 6.480 232.600 10.330 232.750 ;
        RECT 10.030 232.150 10.330 232.600 ;
        RECT 6.480 232.000 10.330 232.150 ;
        RECT 10.030 231.550 10.330 232.000 ;
        RECT 6.480 231.400 10.330 231.550 ;
        RECT 10.030 230.950 10.330 231.400 ;
        RECT 6.480 230.800 10.330 230.950 ;
        RECT 10.030 230.350 10.330 230.800 ;
        RECT 10.780 230.350 10.930 238.550 ;
        RECT 11.380 230.350 11.530 238.550 ;
        RECT 11.980 230.350 12.130 238.550 ;
        RECT 12.580 230.350 12.730 238.550 ;
        RECT 13.180 230.350 13.330 238.550 ;
        RECT 13.780 230.350 13.930 238.550 ;
        RECT 10.030 229.200 10.330 229.650 ;
        RECT 6.480 229.050 10.330 229.200 ;
        RECT 10.030 228.600 10.330 229.050 ;
        RECT 6.480 228.450 10.330 228.600 ;
        RECT 10.030 228.000 10.330 228.450 ;
        RECT 6.480 227.850 10.330 228.000 ;
        RECT 10.030 227.400 10.330 227.850 ;
        RECT 6.480 227.250 10.330 227.400 ;
        RECT 10.030 226.800 10.330 227.250 ;
        RECT 6.480 226.650 10.330 226.800 ;
        RECT 10.030 226.200 10.330 226.650 ;
        RECT 6.480 226.050 10.330 226.200 ;
        RECT 10.030 225.600 10.330 226.050 ;
        RECT 6.480 225.450 10.330 225.600 ;
        RECT 10.030 225.000 10.330 225.450 ;
        RECT 6.480 224.850 10.330 225.000 ;
        RECT 10.030 224.400 10.330 224.850 ;
        RECT 6.480 224.250 10.330 224.400 ;
        RECT 10.030 223.800 10.330 224.250 ;
        RECT 6.480 223.650 10.330 223.800 ;
        RECT 10.030 223.200 10.330 223.650 ;
        RECT 6.480 223.050 10.330 223.200 ;
        RECT 10.030 222.600 10.330 223.050 ;
        RECT 6.480 222.450 10.330 222.600 ;
        RECT 10.030 222.000 10.330 222.450 ;
        RECT 6.530 221.450 10.330 222.000 ;
        RECT 10.780 221.450 10.930 229.650 ;
        RECT 11.380 221.450 11.530 229.650 ;
        RECT 11.980 221.450 12.130 229.650 ;
        RECT 12.580 221.450 12.730 229.650 ;
        RECT 13.180 221.450 13.330 229.650 ;
        RECT 13.780 221.450 13.930 229.650 ;
        RECT 14.380 221.450 15.080 238.550 ;
        RECT 15.530 230.350 15.680 238.550 ;
        RECT 16.130 230.350 16.280 238.550 ;
        RECT 16.730 230.350 16.880 238.550 ;
        RECT 17.330 230.350 17.480 238.550 ;
        RECT 17.930 230.350 18.080 238.550 ;
        RECT 18.530 230.350 18.680 238.550 ;
        RECT 19.130 238.000 22.930 238.550 ;
        RECT 26.530 238.550 42.930 238.600 ;
        RECT 26.530 238.000 30.330 238.550 ;
        RECT 19.130 237.550 19.430 238.000 ;
        RECT 30.030 237.550 30.330 238.000 ;
        RECT 19.130 237.400 22.980 237.550 ;
        RECT 26.480 237.400 30.330 237.550 ;
        RECT 19.130 236.950 19.430 237.400 ;
        RECT 30.030 236.950 30.330 237.400 ;
        RECT 19.130 236.800 22.980 236.950 ;
        RECT 26.480 236.800 30.330 236.950 ;
        RECT 19.130 236.350 19.430 236.800 ;
        RECT 30.030 236.350 30.330 236.800 ;
        RECT 19.130 236.200 22.980 236.350 ;
        RECT 26.480 236.200 30.330 236.350 ;
        RECT 19.130 235.750 19.430 236.200 ;
        RECT 30.030 235.750 30.330 236.200 ;
        RECT 19.130 235.600 22.980 235.750 ;
        RECT 26.480 235.600 30.330 235.750 ;
        RECT 19.130 235.150 19.430 235.600 ;
        RECT 30.030 235.150 30.330 235.600 ;
        RECT 19.130 235.000 22.980 235.150 ;
        RECT 26.480 235.000 30.330 235.150 ;
        RECT 19.130 234.550 19.430 235.000 ;
        RECT 30.030 234.550 30.330 235.000 ;
        RECT 19.130 234.400 22.980 234.550 ;
        RECT 26.480 234.400 30.330 234.550 ;
        RECT 19.130 233.950 19.430 234.400 ;
        RECT 30.030 233.950 30.330 234.400 ;
        RECT 19.130 233.800 22.980 233.950 ;
        RECT 26.480 233.800 30.330 233.950 ;
        RECT 19.130 233.350 19.430 233.800 ;
        RECT 30.030 233.350 30.330 233.800 ;
        RECT 19.130 233.200 22.980 233.350 ;
        RECT 26.480 233.200 30.330 233.350 ;
        RECT 19.130 232.750 19.430 233.200 ;
        RECT 19.130 232.600 22.980 232.750 ;
        RECT 19.130 232.150 19.430 232.600 ;
        RECT 19.130 232.000 22.980 232.150 ;
        RECT 19.130 231.550 19.430 232.000 ;
        RECT 19.130 231.400 22.980 231.550 ;
        RECT 19.130 230.950 19.430 231.400 ;
        RECT 19.130 230.800 22.980 230.950 ;
        RECT 19.130 230.350 19.430 230.800 ;
        RECT 15.530 221.450 15.680 229.650 ;
        RECT 16.130 221.450 16.280 229.650 ;
        RECT 16.730 221.450 16.880 229.650 ;
        RECT 17.330 221.450 17.480 229.650 ;
        RECT 17.930 221.450 18.080 229.650 ;
        RECT 18.530 221.450 18.680 229.650 ;
        RECT 19.130 229.200 19.430 229.650 ;
        RECT 19.130 229.050 22.980 229.200 ;
        RECT 19.130 228.600 19.430 229.050 ;
        RECT 19.130 228.450 22.980 228.600 ;
        RECT 19.130 228.000 19.430 228.450 ;
        RECT 19.130 227.850 22.980 228.000 ;
        RECT 19.130 227.400 19.430 227.850 ;
        RECT 19.130 227.250 22.980 227.400 ;
        RECT 19.130 226.800 19.430 227.250 ;
        RECT 23.830 226.800 25.630 233.200 ;
        RECT 30.030 232.750 30.330 233.200 ;
        RECT 26.480 232.600 30.330 232.750 ;
        RECT 30.030 232.150 30.330 232.600 ;
        RECT 26.480 232.000 30.330 232.150 ;
        RECT 30.030 231.550 30.330 232.000 ;
        RECT 26.480 231.400 30.330 231.550 ;
        RECT 30.030 230.950 30.330 231.400 ;
        RECT 26.480 230.800 30.330 230.950 ;
        RECT 30.030 230.350 30.330 230.800 ;
        RECT 30.780 230.350 30.930 238.550 ;
        RECT 31.380 230.350 31.530 238.550 ;
        RECT 31.980 230.350 32.130 238.550 ;
        RECT 32.580 230.350 32.730 238.550 ;
        RECT 33.180 230.350 33.330 238.550 ;
        RECT 33.780 230.350 33.930 238.550 ;
        RECT 30.030 229.200 30.330 229.650 ;
        RECT 26.480 229.050 30.330 229.200 ;
        RECT 30.030 228.600 30.330 229.050 ;
        RECT 26.480 228.450 30.330 228.600 ;
        RECT 30.030 228.000 30.330 228.450 ;
        RECT 26.480 227.850 30.330 228.000 ;
        RECT 30.030 227.400 30.330 227.850 ;
        RECT 26.480 227.250 30.330 227.400 ;
        RECT 30.030 226.800 30.330 227.250 ;
        RECT 19.130 226.650 22.980 226.800 ;
        RECT 26.480 226.650 30.330 226.800 ;
        RECT 19.130 226.200 19.430 226.650 ;
        RECT 30.030 226.200 30.330 226.650 ;
        RECT 19.130 226.050 22.980 226.200 ;
        RECT 26.480 226.050 30.330 226.200 ;
        RECT 19.130 225.600 19.430 226.050 ;
        RECT 30.030 225.600 30.330 226.050 ;
        RECT 19.130 225.450 22.980 225.600 ;
        RECT 26.480 225.450 30.330 225.600 ;
        RECT 19.130 225.000 19.430 225.450 ;
        RECT 30.030 225.000 30.330 225.450 ;
        RECT 19.130 224.850 22.980 225.000 ;
        RECT 26.480 224.850 30.330 225.000 ;
        RECT 19.130 224.400 19.430 224.850 ;
        RECT 30.030 224.400 30.330 224.850 ;
        RECT 19.130 224.250 22.980 224.400 ;
        RECT 26.480 224.250 30.330 224.400 ;
        RECT 19.130 223.800 19.430 224.250 ;
        RECT 30.030 223.800 30.330 224.250 ;
        RECT 19.130 223.650 22.980 223.800 ;
        RECT 26.480 223.650 30.330 223.800 ;
        RECT 19.130 223.200 19.430 223.650 ;
        RECT 30.030 223.200 30.330 223.650 ;
        RECT 19.130 223.050 22.980 223.200 ;
        RECT 26.480 223.050 30.330 223.200 ;
        RECT 19.130 222.600 19.430 223.050 ;
        RECT 30.030 222.600 30.330 223.050 ;
        RECT 19.130 222.450 22.980 222.600 ;
        RECT 26.480 222.450 30.330 222.600 ;
        RECT 19.130 222.000 19.430 222.450 ;
        RECT 30.030 222.000 30.330 222.450 ;
        RECT 19.130 221.450 22.930 222.000 ;
        RECT 6.530 221.400 22.930 221.450 ;
        RECT 26.530 221.450 30.330 222.000 ;
        RECT 30.780 221.450 30.930 229.650 ;
        RECT 31.380 221.450 31.530 229.650 ;
        RECT 31.980 221.450 32.130 229.650 ;
        RECT 32.580 221.450 32.730 229.650 ;
        RECT 33.180 221.450 33.330 229.650 ;
        RECT 33.780 221.450 33.930 229.650 ;
        RECT 34.380 221.450 35.080 238.550 ;
        RECT 35.530 230.350 35.680 238.550 ;
        RECT 36.130 230.350 36.280 238.550 ;
        RECT 36.730 230.350 36.880 238.550 ;
        RECT 37.330 230.350 37.480 238.550 ;
        RECT 37.930 230.350 38.080 238.550 ;
        RECT 38.530 230.350 38.680 238.550 ;
        RECT 39.130 238.000 42.930 238.550 ;
        RECT 46.530 238.550 62.930 238.600 ;
        RECT 46.530 238.000 50.330 238.550 ;
        RECT 39.130 237.550 39.430 238.000 ;
        RECT 50.030 237.550 50.330 238.000 ;
        RECT 39.130 237.400 42.980 237.550 ;
        RECT 46.480 237.400 50.330 237.550 ;
        RECT 39.130 236.950 39.430 237.400 ;
        RECT 50.030 236.950 50.330 237.400 ;
        RECT 39.130 236.800 42.980 236.950 ;
        RECT 46.480 236.800 50.330 236.950 ;
        RECT 39.130 236.350 39.430 236.800 ;
        RECT 50.030 236.350 50.330 236.800 ;
        RECT 39.130 236.200 42.980 236.350 ;
        RECT 46.480 236.200 50.330 236.350 ;
        RECT 39.130 235.750 39.430 236.200 ;
        RECT 50.030 235.750 50.330 236.200 ;
        RECT 39.130 235.600 42.980 235.750 ;
        RECT 46.480 235.600 50.330 235.750 ;
        RECT 39.130 235.150 39.430 235.600 ;
        RECT 50.030 235.150 50.330 235.600 ;
        RECT 39.130 235.000 42.980 235.150 ;
        RECT 46.480 235.000 50.330 235.150 ;
        RECT 39.130 234.550 39.430 235.000 ;
        RECT 50.030 234.550 50.330 235.000 ;
        RECT 39.130 234.400 42.980 234.550 ;
        RECT 46.480 234.400 50.330 234.550 ;
        RECT 39.130 233.950 39.430 234.400 ;
        RECT 50.030 233.950 50.330 234.400 ;
        RECT 39.130 233.800 42.980 233.950 ;
        RECT 46.480 233.800 50.330 233.950 ;
        RECT 39.130 233.350 39.430 233.800 ;
        RECT 50.030 233.350 50.330 233.800 ;
        RECT 39.130 233.200 42.980 233.350 ;
        RECT 46.480 233.200 50.330 233.350 ;
        RECT 39.130 232.750 39.430 233.200 ;
        RECT 39.130 232.600 42.980 232.750 ;
        RECT 39.130 232.150 39.430 232.600 ;
        RECT 39.130 232.000 42.980 232.150 ;
        RECT 39.130 231.550 39.430 232.000 ;
        RECT 39.130 231.400 42.980 231.550 ;
        RECT 39.130 230.950 39.430 231.400 ;
        RECT 39.130 230.800 42.980 230.950 ;
        RECT 39.130 230.350 39.430 230.800 ;
        RECT 35.530 221.450 35.680 229.650 ;
        RECT 36.130 221.450 36.280 229.650 ;
        RECT 36.730 221.450 36.880 229.650 ;
        RECT 37.330 221.450 37.480 229.650 ;
        RECT 37.930 221.450 38.080 229.650 ;
        RECT 38.530 221.450 38.680 229.650 ;
        RECT 39.130 229.200 39.430 229.650 ;
        RECT 39.130 229.050 42.980 229.200 ;
        RECT 39.130 228.600 39.430 229.050 ;
        RECT 39.130 228.450 42.980 228.600 ;
        RECT 39.130 228.000 39.430 228.450 ;
        RECT 39.130 227.850 42.980 228.000 ;
        RECT 39.130 227.400 39.430 227.850 ;
        RECT 39.130 227.250 42.980 227.400 ;
        RECT 39.130 226.800 39.430 227.250 ;
        RECT 43.830 226.800 45.630 233.200 ;
        RECT 50.030 232.750 50.330 233.200 ;
        RECT 46.480 232.600 50.330 232.750 ;
        RECT 50.030 232.150 50.330 232.600 ;
        RECT 46.480 232.000 50.330 232.150 ;
        RECT 50.030 231.550 50.330 232.000 ;
        RECT 46.480 231.400 50.330 231.550 ;
        RECT 50.030 230.950 50.330 231.400 ;
        RECT 46.480 230.800 50.330 230.950 ;
        RECT 50.030 230.350 50.330 230.800 ;
        RECT 50.780 230.350 50.930 238.550 ;
        RECT 51.380 230.350 51.530 238.550 ;
        RECT 51.980 230.350 52.130 238.550 ;
        RECT 52.580 230.350 52.730 238.550 ;
        RECT 53.180 230.350 53.330 238.550 ;
        RECT 53.780 230.350 53.930 238.550 ;
        RECT 50.030 229.200 50.330 229.650 ;
        RECT 46.480 229.050 50.330 229.200 ;
        RECT 50.030 228.600 50.330 229.050 ;
        RECT 46.480 228.450 50.330 228.600 ;
        RECT 50.030 228.000 50.330 228.450 ;
        RECT 46.480 227.850 50.330 228.000 ;
        RECT 50.030 227.400 50.330 227.850 ;
        RECT 46.480 227.250 50.330 227.400 ;
        RECT 50.030 226.800 50.330 227.250 ;
        RECT 39.130 226.650 42.980 226.800 ;
        RECT 46.480 226.650 50.330 226.800 ;
        RECT 39.130 226.200 39.430 226.650 ;
        RECT 50.030 226.200 50.330 226.650 ;
        RECT 39.130 226.050 42.980 226.200 ;
        RECT 46.480 226.050 50.330 226.200 ;
        RECT 39.130 225.600 39.430 226.050 ;
        RECT 50.030 225.600 50.330 226.050 ;
        RECT 39.130 225.450 42.980 225.600 ;
        RECT 46.480 225.450 50.330 225.600 ;
        RECT 39.130 225.000 39.430 225.450 ;
        RECT 50.030 225.000 50.330 225.450 ;
        RECT 39.130 224.850 42.980 225.000 ;
        RECT 46.480 224.850 50.330 225.000 ;
        RECT 39.130 224.400 39.430 224.850 ;
        RECT 50.030 224.400 50.330 224.850 ;
        RECT 39.130 224.250 42.980 224.400 ;
        RECT 46.480 224.250 50.330 224.400 ;
        RECT 39.130 223.800 39.430 224.250 ;
        RECT 50.030 223.800 50.330 224.250 ;
        RECT 39.130 223.650 42.980 223.800 ;
        RECT 46.480 223.650 50.330 223.800 ;
        RECT 39.130 223.200 39.430 223.650 ;
        RECT 50.030 223.200 50.330 223.650 ;
        RECT 39.130 223.050 42.980 223.200 ;
        RECT 46.480 223.050 50.330 223.200 ;
        RECT 39.130 222.600 39.430 223.050 ;
        RECT 50.030 222.600 50.330 223.050 ;
        RECT 39.130 222.450 42.980 222.600 ;
        RECT 46.480 222.450 50.330 222.600 ;
        RECT 39.130 222.000 39.430 222.450 ;
        RECT 50.030 222.000 50.330 222.450 ;
        RECT 39.130 221.450 42.930 222.000 ;
        RECT 26.530 221.400 42.930 221.450 ;
        RECT 46.530 221.450 50.330 222.000 ;
        RECT 50.780 221.450 50.930 229.650 ;
        RECT 51.380 221.450 51.530 229.650 ;
        RECT 51.980 221.450 52.130 229.650 ;
        RECT 52.580 221.450 52.730 229.650 ;
        RECT 53.180 221.450 53.330 229.650 ;
        RECT 53.780 221.450 53.930 229.650 ;
        RECT 54.380 221.450 55.080 238.550 ;
        RECT 55.530 230.350 55.680 238.550 ;
        RECT 56.130 230.350 56.280 238.550 ;
        RECT 56.730 230.350 56.880 238.550 ;
        RECT 57.330 230.350 57.480 238.550 ;
        RECT 57.930 230.350 58.080 238.550 ;
        RECT 58.530 230.350 58.680 238.550 ;
        RECT 59.130 238.000 62.930 238.550 ;
        RECT 66.530 238.550 82.930 238.600 ;
        RECT 66.530 238.000 70.330 238.550 ;
        RECT 59.130 237.550 59.430 238.000 ;
        RECT 70.030 237.550 70.330 238.000 ;
        RECT 59.130 237.400 62.980 237.550 ;
        RECT 66.480 237.400 70.330 237.550 ;
        RECT 59.130 236.950 59.430 237.400 ;
        RECT 70.030 236.950 70.330 237.400 ;
        RECT 59.130 236.800 62.980 236.950 ;
        RECT 66.480 236.800 70.330 236.950 ;
        RECT 59.130 236.350 59.430 236.800 ;
        RECT 70.030 236.350 70.330 236.800 ;
        RECT 59.130 236.200 62.980 236.350 ;
        RECT 66.480 236.200 70.330 236.350 ;
        RECT 59.130 235.750 59.430 236.200 ;
        RECT 70.030 235.750 70.330 236.200 ;
        RECT 59.130 235.600 62.980 235.750 ;
        RECT 66.480 235.600 70.330 235.750 ;
        RECT 59.130 235.150 59.430 235.600 ;
        RECT 70.030 235.150 70.330 235.600 ;
        RECT 59.130 235.000 62.980 235.150 ;
        RECT 66.480 235.000 70.330 235.150 ;
        RECT 59.130 234.550 59.430 235.000 ;
        RECT 70.030 234.550 70.330 235.000 ;
        RECT 59.130 234.400 62.980 234.550 ;
        RECT 66.480 234.400 70.330 234.550 ;
        RECT 59.130 233.950 59.430 234.400 ;
        RECT 70.030 233.950 70.330 234.400 ;
        RECT 59.130 233.800 62.980 233.950 ;
        RECT 66.480 233.800 70.330 233.950 ;
        RECT 59.130 233.350 59.430 233.800 ;
        RECT 70.030 233.350 70.330 233.800 ;
        RECT 59.130 233.200 62.980 233.350 ;
        RECT 66.480 233.200 70.330 233.350 ;
        RECT 59.130 232.750 59.430 233.200 ;
        RECT 59.130 232.600 62.980 232.750 ;
        RECT 59.130 232.150 59.430 232.600 ;
        RECT 59.130 232.000 62.980 232.150 ;
        RECT 59.130 231.550 59.430 232.000 ;
        RECT 59.130 231.400 62.980 231.550 ;
        RECT 59.130 230.950 59.430 231.400 ;
        RECT 59.130 230.800 62.980 230.950 ;
        RECT 59.130 230.350 59.430 230.800 ;
        RECT 55.530 221.450 55.680 229.650 ;
        RECT 56.130 221.450 56.280 229.650 ;
        RECT 56.730 221.450 56.880 229.650 ;
        RECT 57.330 221.450 57.480 229.650 ;
        RECT 57.930 221.450 58.080 229.650 ;
        RECT 58.530 221.450 58.680 229.650 ;
        RECT 59.130 229.200 59.430 229.650 ;
        RECT 59.130 229.050 62.980 229.200 ;
        RECT 59.130 228.600 59.430 229.050 ;
        RECT 59.130 228.450 62.980 228.600 ;
        RECT 59.130 228.000 59.430 228.450 ;
        RECT 59.130 227.850 62.980 228.000 ;
        RECT 59.130 227.400 59.430 227.850 ;
        RECT 59.130 227.250 62.980 227.400 ;
        RECT 59.130 226.800 59.430 227.250 ;
        RECT 63.830 226.800 65.630 233.200 ;
        RECT 70.030 232.750 70.330 233.200 ;
        RECT 66.480 232.600 70.330 232.750 ;
        RECT 70.030 232.150 70.330 232.600 ;
        RECT 66.480 232.000 70.330 232.150 ;
        RECT 70.030 231.550 70.330 232.000 ;
        RECT 66.480 231.400 70.330 231.550 ;
        RECT 70.030 230.950 70.330 231.400 ;
        RECT 66.480 230.800 70.330 230.950 ;
        RECT 70.030 230.350 70.330 230.800 ;
        RECT 70.780 230.350 70.930 238.550 ;
        RECT 71.380 230.350 71.530 238.550 ;
        RECT 71.980 230.350 72.130 238.550 ;
        RECT 72.580 230.350 72.730 238.550 ;
        RECT 73.180 230.350 73.330 238.550 ;
        RECT 73.780 230.350 73.930 238.550 ;
        RECT 70.030 229.200 70.330 229.650 ;
        RECT 66.480 229.050 70.330 229.200 ;
        RECT 70.030 228.600 70.330 229.050 ;
        RECT 66.480 228.450 70.330 228.600 ;
        RECT 70.030 228.000 70.330 228.450 ;
        RECT 66.480 227.850 70.330 228.000 ;
        RECT 70.030 227.400 70.330 227.850 ;
        RECT 66.480 227.250 70.330 227.400 ;
        RECT 70.030 226.800 70.330 227.250 ;
        RECT 59.130 226.650 62.980 226.800 ;
        RECT 66.480 226.650 70.330 226.800 ;
        RECT 59.130 226.200 59.430 226.650 ;
        RECT 70.030 226.200 70.330 226.650 ;
        RECT 59.130 226.050 62.980 226.200 ;
        RECT 66.480 226.050 70.330 226.200 ;
        RECT 59.130 225.600 59.430 226.050 ;
        RECT 70.030 225.600 70.330 226.050 ;
        RECT 59.130 225.450 62.980 225.600 ;
        RECT 66.480 225.450 70.330 225.600 ;
        RECT 59.130 225.000 59.430 225.450 ;
        RECT 70.030 225.000 70.330 225.450 ;
        RECT 59.130 224.850 62.980 225.000 ;
        RECT 66.480 224.850 70.330 225.000 ;
        RECT 59.130 224.400 59.430 224.850 ;
        RECT 70.030 224.400 70.330 224.850 ;
        RECT 59.130 224.250 62.980 224.400 ;
        RECT 66.480 224.250 70.330 224.400 ;
        RECT 59.130 223.800 59.430 224.250 ;
        RECT 70.030 223.800 70.330 224.250 ;
        RECT 59.130 223.650 62.980 223.800 ;
        RECT 66.480 223.650 70.330 223.800 ;
        RECT 59.130 223.200 59.430 223.650 ;
        RECT 70.030 223.200 70.330 223.650 ;
        RECT 59.130 223.050 62.980 223.200 ;
        RECT 66.480 223.050 70.330 223.200 ;
        RECT 59.130 222.600 59.430 223.050 ;
        RECT 70.030 222.600 70.330 223.050 ;
        RECT 59.130 222.450 62.980 222.600 ;
        RECT 66.480 222.450 70.330 222.600 ;
        RECT 59.130 222.000 59.430 222.450 ;
        RECT 70.030 222.000 70.330 222.450 ;
        RECT 59.130 221.450 62.930 222.000 ;
        RECT 46.530 221.400 62.930 221.450 ;
        RECT 66.530 221.450 70.330 222.000 ;
        RECT 70.780 221.450 70.930 229.650 ;
        RECT 71.380 221.450 71.530 229.650 ;
        RECT 71.980 221.450 72.130 229.650 ;
        RECT 72.580 221.450 72.730 229.650 ;
        RECT 73.180 221.450 73.330 229.650 ;
        RECT 73.780 221.450 73.930 229.650 ;
        RECT 74.380 221.450 75.080 238.550 ;
        RECT 75.530 230.350 75.680 238.550 ;
        RECT 76.130 230.350 76.280 238.550 ;
        RECT 76.730 230.350 76.880 238.550 ;
        RECT 77.330 230.350 77.480 238.550 ;
        RECT 77.930 230.350 78.080 238.550 ;
        RECT 78.530 230.350 78.680 238.550 ;
        RECT 79.130 238.000 82.930 238.550 ;
        RECT 86.530 238.550 102.930 238.600 ;
        RECT 86.530 238.000 90.330 238.550 ;
        RECT 79.130 237.550 79.430 238.000 ;
        RECT 90.030 237.550 90.330 238.000 ;
        RECT 79.130 237.400 82.980 237.550 ;
        RECT 86.480 237.400 90.330 237.550 ;
        RECT 79.130 236.950 79.430 237.400 ;
        RECT 90.030 236.950 90.330 237.400 ;
        RECT 79.130 236.800 82.980 236.950 ;
        RECT 86.480 236.800 90.330 236.950 ;
        RECT 79.130 236.350 79.430 236.800 ;
        RECT 90.030 236.350 90.330 236.800 ;
        RECT 79.130 236.200 82.980 236.350 ;
        RECT 86.480 236.200 90.330 236.350 ;
        RECT 79.130 235.750 79.430 236.200 ;
        RECT 90.030 235.750 90.330 236.200 ;
        RECT 79.130 235.600 82.980 235.750 ;
        RECT 86.480 235.600 90.330 235.750 ;
        RECT 79.130 235.150 79.430 235.600 ;
        RECT 90.030 235.150 90.330 235.600 ;
        RECT 79.130 235.000 82.980 235.150 ;
        RECT 86.480 235.000 90.330 235.150 ;
        RECT 79.130 234.550 79.430 235.000 ;
        RECT 90.030 234.550 90.330 235.000 ;
        RECT 79.130 234.400 82.980 234.550 ;
        RECT 86.480 234.400 90.330 234.550 ;
        RECT 79.130 233.950 79.430 234.400 ;
        RECT 90.030 233.950 90.330 234.400 ;
        RECT 79.130 233.800 82.980 233.950 ;
        RECT 86.480 233.800 90.330 233.950 ;
        RECT 79.130 233.350 79.430 233.800 ;
        RECT 90.030 233.350 90.330 233.800 ;
        RECT 79.130 233.200 82.980 233.350 ;
        RECT 86.480 233.200 90.330 233.350 ;
        RECT 79.130 232.750 79.430 233.200 ;
        RECT 79.130 232.600 82.980 232.750 ;
        RECT 79.130 232.150 79.430 232.600 ;
        RECT 79.130 232.000 82.980 232.150 ;
        RECT 79.130 231.550 79.430 232.000 ;
        RECT 79.130 231.400 82.980 231.550 ;
        RECT 79.130 230.950 79.430 231.400 ;
        RECT 79.130 230.800 82.980 230.950 ;
        RECT 79.130 230.350 79.430 230.800 ;
        RECT 75.530 221.450 75.680 229.650 ;
        RECT 76.130 221.450 76.280 229.650 ;
        RECT 76.730 221.450 76.880 229.650 ;
        RECT 77.330 221.450 77.480 229.650 ;
        RECT 77.930 221.450 78.080 229.650 ;
        RECT 78.530 221.450 78.680 229.650 ;
        RECT 79.130 229.200 79.430 229.650 ;
        RECT 79.130 229.050 82.980 229.200 ;
        RECT 79.130 228.600 79.430 229.050 ;
        RECT 79.130 228.450 82.980 228.600 ;
        RECT 79.130 228.000 79.430 228.450 ;
        RECT 79.130 227.850 82.980 228.000 ;
        RECT 79.130 227.400 79.430 227.850 ;
        RECT 79.130 227.250 82.980 227.400 ;
        RECT 79.130 226.800 79.430 227.250 ;
        RECT 83.830 226.800 85.630 233.200 ;
        RECT 90.030 232.750 90.330 233.200 ;
        RECT 86.480 232.600 90.330 232.750 ;
        RECT 90.030 232.150 90.330 232.600 ;
        RECT 86.480 232.000 90.330 232.150 ;
        RECT 90.030 231.550 90.330 232.000 ;
        RECT 86.480 231.400 90.330 231.550 ;
        RECT 90.030 230.950 90.330 231.400 ;
        RECT 86.480 230.800 90.330 230.950 ;
        RECT 90.030 230.350 90.330 230.800 ;
        RECT 90.780 230.350 90.930 238.550 ;
        RECT 91.380 230.350 91.530 238.550 ;
        RECT 91.980 230.350 92.130 238.550 ;
        RECT 92.580 230.350 92.730 238.550 ;
        RECT 93.180 230.350 93.330 238.550 ;
        RECT 93.780 230.350 93.930 238.550 ;
        RECT 90.030 229.200 90.330 229.650 ;
        RECT 86.480 229.050 90.330 229.200 ;
        RECT 90.030 228.600 90.330 229.050 ;
        RECT 86.480 228.450 90.330 228.600 ;
        RECT 90.030 228.000 90.330 228.450 ;
        RECT 86.480 227.850 90.330 228.000 ;
        RECT 90.030 227.400 90.330 227.850 ;
        RECT 86.480 227.250 90.330 227.400 ;
        RECT 90.030 226.800 90.330 227.250 ;
        RECT 79.130 226.650 82.980 226.800 ;
        RECT 86.480 226.650 90.330 226.800 ;
        RECT 79.130 226.200 79.430 226.650 ;
        RECT 90.030 226.200 90.330 226.650 ;
        RECT 79.130 226.050 82.980 226.200 ;
        RECT 86.480 226.050 90.330 226.200 ;
        RECT 79.130 225.600 79.430 226.050 ;
        RECT 90.030 225.600 90.330 226.050 ;
        RECT 79.130 225.450 82.980 225.600 ;
        RECT 86.480 225.450 90.330 225.600 ;
        RECT 79.130 225.000 79.430 225.450 ;
        RECT 90.030 225.000 90.330 225.450 ;
        RECT 79.130 224.850 82.980 225.000 ;
        RECT 86.480 224.850 90.330 225.000 ;
        RECT 79.130 224.400 79.430 224.850 ;
        RECT 90.030 224.400 90.330 224.850 ;
        RECT 79.130 224.250 82.980 224.400 ;
        RECT 86.480 224.250 90.330 224.400 ;
        RECT 79.130 223.800 79.430 224.250 ;
        RECT 90.030 223.800 90.330 224.250 ;
        RECT 79.130 223.650 82.980 223.800 ;
        RECT 86.480 223.650 90.330 223.800 ;
        RECT 79.130 223.200 79.430 223.650 ;
        RECT 90.030 223.200 90.330 223.650 ;
        RECT 79.130 223.050 82.980 223.200 ;
        RECT 86.480 223.050 90.330 223.200 ;
        RECT 79.130 222.600 79.430 223.050 ;
        RECT 90.030 222.600 90.330 223.050 ;
        RECT 79.130 222.450 82.980 222.600 ;
        RECT 86.480 222.450 90.330 222.600 ;
        RECT 79.130 222.000 79.430 222.450 ;
        RECT 90.030 222.000 90.330 222.450 ;
        RECT 79.130 221.450 82.930 222.000 ;
        RECT 66.530 221.400 82.930 221.450 ;
        RECT 86.530 221.450 90.330 222.000 ;
        RECT 90.780 221.450 90.930 229.650 ;
        RECT 91.380 221.450 91.530 229.650 ;
        RECT 91.980 221.450 92.130 229.650 ;
        RECT 92.580 221.450 92.730 229.650 ;
        RECT 93.180 221.450 93.330 229.650 ;
        RECT 93.780 221.450 93.930 229.650 ;
        RECT 94.380 221.450 95.080 238.550 ;
        RECT 95.530 230.350 95.680 238.550 ;
        RECT 96.130 230.350 96.280 238.550 ;
        RECT 96.730 230.350 96.880 238.550 ;
        RECT 97.330 230.350 97.480 238.550 ;
        RECT 97.930 230.350 98.080 238.550 ;
        RECT 98.530 230.350 98.680 238.550 ;
        RECT 99.130 238.000 102.930 238.550 ;
        RECT 106.530 238.550 122.930 238.600 ;
        RECT 106.530 238.000 110.330 238.550 ;
        RECT 99.130 237.550 99.430 238.000 ;
        RECT 110.030 237.550 110.330 238.000 ;
        RECT 99.130 237.400 102.980 237.550 ;
        RECT 106.480 237.400 110.330 237.550 ;
        RECT 99.130 236.950 99.430 237.400 ;
        RECT 110.030 236.950 110.330 237.400 ;
        RECT 99.130 236.800 102.980 236.950 ;
        RECT 106.480 236.800 110.330 236.950 ;
        RECT 99.130 236.350 99.430 236.800 ;
        RECT 110.030 236.350 110.330 236.800 ;
        RECT 99.130 236.200 102.980 236.350 ;
        RECT 106.480 236.200 110.330 236.350 ;
        RECT 99.130 235.750 99.430 236.200 ;
        RECT 110.030 235.750 110.330 236.200 ;
        RECT 99.130 235.600 102.980 235.750 ;
        RECT 106.480 235.600 110.330 235.750 ;
        RECT 99.130 235.150 99.430 235.600 ;
        RECT 110.030 235.150 110.330 235.600 ;
        RECT 99.130 235.000 102.980 235.150 ;
        RECT 106.480 235.000 110.330 235.150 ;
        RECT 99.130 234.550 99.430 235.000 ;
        RECT 110.030 234.550 110.330 235.000 ;
        RECT 99.130 234.400 102.980 234.550 ;
        RECT 106.480 234.400 110.330 234.550 ;
        RECT 99.130 233.950 99.430 234.400 ;
        RECT 110.030 233.950 110.330 234.400 ;
        RECT 99.130 233.800 102.980 233.950 ;
        RECT 106.480 233.800 110.330 233.950 ;
        RECT 99.130 233.350 99.430 233.800 ;
        RECT 110.030 233.350 110.330 233.800 ;
        RECT 99.130 233.200 102.980 233.350 ;
        RECT 106.480 233.200 110.330 233.350 ;
        RECT 99.130 232.750 99.430 233.200 ;
        RECT 99.130 232.600 102.980 232.750 ;
        RECT 99.130 232.150 99.430 232.600 ;
        RECT 99.130 232.000 102.980 232.150 ;
        RECT 99.130 231.550 99.430 232.000 ;
        RECT 99.130 231.400 102.980 231.550 ;
        RECT 99.130 230.950 99.430 231.400 ;
        RECT 99.130 230.800 102.980 230.950 ;
        RECT 99.130 230.350 99.430 230.800 ;
        RECT 95.530 221.450 95.680 229.650 ;
        RECT 96.130 221.450 96.280 229.650 ;
        RECT 96.730 221.450 96.880 229.650 ;
        RECT 97.330 221.450 97.480 229.650 ;
        RECT 97.930 221.450 98.080 229.650 ;
        RECT 98.530 221.450 98.680 229.650 ;
        RECT 99.130 229.200 99.430 229.650 ;
        RECT 99.130 229.050 102.980 229.200 ;
        RECT 99.130 228.600 99.430 229.050 ;
        RECT 99.130 228.450 102.980 228.600 ;
        RECT 99.130 228.000 99.430 228.450 ;
        RECT 99.130 227.850 102.980 228.000 ;
        RECT 99.130 227.400 99.430 227.850 ;
        RECT 99.130 227.250 102.980 227.400 ;
        RECT 99.130 226.800 99.430 227.250 ;
        RECT 103.830 226.800 105.630 233.200 ;
        RECT 110.030 232.750 110.330 233.200 ;
        RECT 106.480 232.600 110.330 232.750 ;
        RECT 110.030 232.150 110.330 232.600 ;
        RECT 106.480 232.000 110.330 232.150 ;
        RECT 110.030 231.550 110.330 232.000 ;
        RECT 106.480 231.400 110.330 231.550 ;
        RECT 110.030 230.950 110.330 231.400 ;
        RECT 106.480 230.800 110.330 230.950 ;
        RECT 110.030 230.350 110.330 230.800 ;
        RECT 110.780 230.350 110.930 238.550 ;
        RECT 111.380 230.350 111.530 238.550 ;
        RECT 111.980 230.350 112.130 238.550 ;
        RECT 112.580 230.350 112.730 238.550 ;
        RECT 113.180 230.350 113.330 238.550 ;
        RECT 113.780 230.350 113.930 238.550 ;
        RECT 110.030 229.200 110.330 229.650 ;
        RECT 106.480 229.050 110.330 229.200 ;
        RECT 110.030 228.600 110.330 229.050 ;
        RECT 106.480 228.450 110.330 228.600 ;
        RECT 110.030 228.000 110.330 228.450 ;
        RECT 106.480 227.850 110.330 228.000 ;
        RECT 110.030 227.400 110.330 227.850 ;
        RECT 106.480 227.250 110.330 227.400 ;
        RECT 110.030 226.800 110.330 227.250 ;
        RECT 99.130 226.650 102.980 226.800 ;
        RECT 106.480 226.650 110.330 226.800 ;
        RECT 99.130 226.200 99.430 226.650 ;
        RECT 110.030 226.200 110.330 226.650 ;
        RECT 99.130 226.050 102.980 226.200 ;
        RECT 106.480 226.050 110.330 226.200 ;
        RECT 99.130 225.600 99.430 226.050 ;
        RECT 110.030 225.600 110.330 226.050 ;
        RECT 99.130 225.450 102.980 225.600 ;
        RECT 106.480 225.450 110.330 225.600 ;
        RECT 99.130 225.000 99.430 225.450 ;
        RECT 110.030 225.000 110.330 225.450 ;
        RECT 99.130 224.850 102.980 225.000 ;
        RECT 106.480 224.850 110.330 225.000 ;
        RECT 99.130 224.400 99.430 224.850 ;
        RECT 110.030 224.400 110.330 224.850 ;
        RECT 99.130 224.250 102.980 224.400 ;
        RECT 106.480 224.250 110.330 224.400 ;
        RECT 99.130 223.800 99.430 224.250 ;
        RECT 110.030 223.800 110.330 224.250 ;
        RECT 99.130 223.650 102.980 223.800 ;
        RECT 106.480 223.650 110.330 223.800 ;
        RECT 99.130 223.200 99.430 223.650 ;
        RECT 110.030 223.200 110.330 223.650 ;
        RECT 99.130 223.050 102.980 223.200 ;
        RECT 106.480 223.050 110.330 223.200 ;
        RECT 99.130 222.600 99.430 223.050 ;
        RECT 110.030 222.600 110.330 223.050 ;
        RECT 99.130 222.450 102.980 222.600 ;
        RECT 106.480 222.450 110.330 222.600 ;
        RECT 99.130 222.000 99.430 222.450 ;
        RECT 110.030 222.000 110.330 222.450 ;
        RECT 99.130 221.450 102.930 222.000 ;
        RECT 86.530 221.400 102.930 221.450 ;
        RECT 106.530 221.450 110.330 222.000 ;
        RECT 110.780 221.450 110.930 229.650 ;
        RECT 111.380 221.450 111.530 229.650 ;
        RECT 111.980 221.450 112.130 229.650 ;
        RECT 112.580 221.450 112.730 229.650 ;
        RECT 113.180 221.450 113.330 229.650 ;
        RECT 113.780 221.450 113.930 229.650 ;
        RECT 114.380 221.450 115.080 238.550 ;
        RECT 115.530 230.350 115.680 238.550 ;
        RECT 116.130 230.350 116.280 238.550 ;
        RECT 116.730 230.350 116.880 238.550 ;
        RECT 117.330 230.350 117.480 238.550 ;
        RECT 117.930 230.350 118.080 238.550 ;
        RECT 118.530 230.350 118.680 238.550 ;
        RECT 119.130 238.000 122.930 238.550 ;
        RECT 119.130 237.550 119.430 238.000 ;
        RECT 119.130 237.400 122.980 237.550 ;
        RECT 119.130 236.950 119.430 237.400 ;
        RECT 119.130 236.800 122.980 236.950 ;
        RECT 119.130 236.350 119.430 236.800 ;
        RECT 119.130 236.200 122.980 236.350 ;
        RECT 119.130 235.750 119.430 236.200 ;
        RECT 119.130 235.600 122.980 235.750 ;
        RECT 119.130 235.150 119.430 235.600 ;
        RECT 119.130 235.000 122.980 235.150 ;
        RECT 119.130 234.550 119.430 235.000 ;
        RECT 119.130 234.400 122.980 234.550 ;
        RECT 119.130 233.950 119.430 234.400 ;
        RECT 119.130 233.800 122.980 233.950 ;
        RECT 119.130 233.350 119.430 233.800 ;
        RECT 119.130 233.200 122.980 233.350 ;
        RECT 119.130 232.750 119.430 233.200 ;
        RECT 119.130 232.600 122.980 232.750 ;
        RECT 119.130 232.150 119.430 232.600 ;
        RECT 119.130 232.000 122.980 232.150 ;
        RECT 119.130 231.550 119.430 232.000 ;
        RECT 119.130 231.400 122.980 231.550 ;
        RECT 119.130 230.950 119.430 231.400 ;
        RECT 119.130 230.800 122.980 230.950 ;
        RECT 119.130 230.350 119.430 230.800 ;
        RECT 115.530 221.450 115.680 229.650 ;
        RECT 116.130 221.450 116.280 229.650 ;
        RECT 116.730 221.450 116.880 229.650 ;
        RECT 117.330 221.450 117.480 229.650 ;
        RECT 117.930 221.450 118.080 229.650 ;
        RECT 118.530 221.450 118.680 229.650 ;
        RECT 119.130 229.200 119.430 229.650 ;
        RECT 119.130 229.050 122.980 229.200 ;
        RECT 119.130 228.600 119.430 229.050 ;
        RECT 119.130 228.450 122.980 228.600 ;
        RECT 119.130 228.000 119.430 228.450 ;
        RECT 119.130 227.850 122.980 228.000 ;
        RECT 119.130 227.400 119.430 227.850 ;
        RECT 119.130 227.250 122.980 227.400 ;
        RECT 119.130 226.800 119.430 227.250 ;
        RECT 123.830 226.800 124.730 233.200 ;
        RECT 129.850 229.640 131.850 230.915 ;
        RECT 119.130 226.650 122.980 226.800 ;
        RECT 119.130 226.200 119.430 226.650 ;
        RECT 119.130 226.050 122.980 226.200 ;
        RECT 119.130 225.600 119.430 226.050 ;
        RECT 119.130 225.450 122.980 225.600 ;
        RECT 119.130 225.000 119.430 225.450 ;
        RECT 119.130 224.850 122.980 225.000 ;
        RECT 119.130 224.400 119.430 224.850 ;
        RECT 119.130 224.250 122.980 224.400 ;
        RECT 119.130 223.800 119.430 224.250 ;
        RECT 119.130 223.650 122.980 223.800 ;
        RECT 119.130 223.200 119.430 223.650 ;
        RECT 119.130 223.050 122.980 223.200 ;
        RECT 119.130 222.600 119.430 223.050 ;
        RECT 119.130 222.450 122.980 222.600 ;
        RECT 119.130 222.000 119.430 222.450 ;
        RECT 119.130 221.450 122.930 222.000 ;
        RECT 106.530 221.400 122.930 221.450 ;
        RECT 9.630 220.900 19.830 221.400 ;
        RECT 29.630 220.900 39.830 221.400 ;
        RECT 49.630 220.900 59.830 221.400 ;
        RECT 69.630 220.900 79.830 221.400 ;
        RECT 89.630 220.900 99.830 221.400 ;
        RECT 109.630 220.900 119.830 221.400 ;
        RECT 11.530 219.100 17.930 220.900 ;
        RECT 31.530 219.100 37.930 220.900 ;
        RECT 51.530 219.100 57.930 220.900 ;
        RECT 71.530 219.100 77.930 220.900 ;
        RECT 91.530 219.100 97.930 220.900 ;
        RECT 111.530 219.100 117.930 220.900 ;
        RECT 9.630 218.600 19.830 219.100 ;
        RECT 29.630 218.600 39.830 219.100 ;
        RECT 49.630 218.600 59.830 219.100 ;
        RECT 69.630 218.600 79.830 219.100 ;
        RECT 89.630 218.600 99.830 219.100 ;
        RECT 109.630 218.600 119.830 219.100 ;
        RECT 6.530 218.550 22.930 218.600 ;
        RECT 6.530 218.000 10.330 218.550 ;
        RECT 10.030 217.550 10.330 218.000 ;
        RECT 6.480 217.400 10.330 217.550 ;
        RECT 10.030 216.950 10.330 217.400 ;
        RECT 6.480 216.800 10.330 216.950 ;
        RECT 10.030 216.350 10.330 216.800 ;
        RECT 6.480 216.200 10.330 216.350 ;
        RECT 10.030 215.750 10.330 216.200 ;
        RECT 6.480 215.600 10.330 215.750 ;
        RECT 10.030 215.150 10.330 215.600 ;
        RECT 6.480 215.000 10.330 215.150 ;
        RECT 10.030 214.550 10.330 215.000 ;
        RECT 6.480 214.400 10.330 214.550 ;
        RECT 10.030 213.950 10.330 214.400 ;
        RECT 6.480 213.800 10.330 213.950 ;
        RECT 10.030 213.350 10.330 213.800 ;
        RECT 6.480 213.200 10.330 213.350 ;
        RECT 4.730 206.800 5.630 213.200 ;
        RECT 10.030 212.750 10.330 213.200 ;
        RECT 6.480 212.600 10.330 212.750 ;
        RECT 10.030 212.150 10.330 212.600 ;
        RECT 6.480 212.000 10.330 212.150 ;
        RECT 10.030 211.550 10.330 212.000 ;
        RECT 6.480 211.400 10.330 211.550 ;
        RECT 10.030 210.950 10.330 211.400 ;
        RECT 6.480 210.800 10.330 210.950 ;
        RECT 10.030 210.350 10.330 210.800 ;
        RECT 10.780 210.350 10.930 218.550 ;
        RECT 11.380 210.350 11.530 218.550 ;
        RECT 11.980 210.350 12.130 218.550 ;
        RECT 12.580 210.350 12.730 218.550 ;
        RECT 13.180 210.350 13.330 218.550 ;
        RECT 13.780 210.350 13.930 218.550 ;
        RECT 10.030 209.200 10.330 209.650 ;
        RECT 6.480 209.050 10.330 209.200 ;
        RECT 10.030 208.600 10.330 209.050 ;
        RECT 6.480 208.450 10.330 208.600 ;
        RECT 10.030 208.000 10.330 208.450 ;
        RECT 6.480 207.850 10.330 208.000 ;
        RECT 10.030 207.400 10.330 207.850 ;
        RECT 6.480 207.250 10.330 207.400 ;
        RECT 10.030 206.800 10.330 207.250 ;
        RECT 6.480 206.650 10.330 206.800 ;
        RECT 10.030 206.200 10.330 206.650 ;
        RECT 6.480 206.050 10.330 206.200 ;
        RECT 10.030 205.600 10.330 206.050 ;
        RECT 6.480 205.450 10.330 205.600 ;
        RECT 10.030 205.000 10.330 205.450 ;
        RECT 6.480 204.850 10.330 205.000 ;
        RECT 10.030 204.400 10.330 204.850 ;
        RECT 6.480 204.250 10.330 204.400 ;
        RECT 10.030 203.800 10.330 204.250 ;
        RECT 6.480 203.650 10.330 203.800 ;
        RECT 10.030 203.200 10.330 203.650 ;
        RECT 6.480 203.050 10.330 203.200 ;
        RECT 10.030 202.600 10.330 203.050 ;
        RECT 6.480 202.450 10.330 202.600 ;
        RECT 10.030 202.000 10.330 202.450 ;
        RECT 6.530 201.450 10.330 202.000 ;
        RECT 10.780 201.450 10.930 209.650 ;
        RECT 11.380 201.450 11.530 209.650 ;
        RECT 11.980 201.450 12.130 209.650 ;
        RECT 12.580 201.450 12.730 209.650 ;
        RECT 13.180 201.450 13.330 209.650 ;
        RECT 13.780 201.450 13.930 209.650 ;
        RECT 14.380 201.450 15.080 218.550 ;
        RECT 15.530 210.350 15.680 218.550 ;
        RECT 16.130 210.350 16.280 218.550 ;
        RECT 16.730 210.350 16.880 218.550 ;
        RECT 17.330 210.350 17.480 218.550 ;
        RECT 17.930 210.350 18.080 218.550 ;
        RECT 18.530 210.350 18.680 218.550 ;
        RECT 19.130 218.000 22.930 218.550 ;
        RECT 26.530 218.550 42.930 218.600 ;
        RECT 26.530 218.000 30.330 218.550 ;
        RECT 19.130 217.550 19.430 218.000 ;
        RECT 30.030 217.550 30.330 218.000 ;
        RECT 19.130 217.400 22.980 217.550 ;
        RECT 26.480 217.400 30.330 217.550 ;
        RECT 19.130 216.950 19.430 217.400 ;
        RECT 30.030 216.950 30.330 217.400 ;
        RECT 19.130 216.800 22.980 216.950 ;
        RECT 26.480 216.800 30.330 216.950 ;
        RECT 19.130 216.350 19.430 216.800 ;
        RECT 30.030 216.350 30.330 216.800 ;
        RECT 19.130 216.200 22.980 216.350 ;
        RECT 26.480 216.200 30.330 216.350 ;
        RECT 19.130 215.750 19.430 216.200 ;
        RECT 30.030 215.750 30.330 216.200 ;
        RECT 19.130 215.600 22.980 215.750 ;
        RECT 26.480 215.600 30.330 215.750 ;
        RECT 19.130 215.150 19.430 215.600 ;
        RECT 30.030 215.150 30.330 215.600 ;
        RECT 19.130 215.000 22.980 215.150 ;
        RECT 26.480 215.000 30.330 215.150 ;
        RECT 19.130 214.550 19.430 215.000 ;
        RECT 30.030 214.550 30.330 215.000 ;
        RECT 19.130 214.400 22.980 214.550 ;
        RECT 26.480 214.400 30.330 214.550 ;
        RECT 19.130 213.950 19.430 214.400 ;
        RECT 30.030 213.950 30.330 214.400 ;
        RECT 19.130 213.800 22.980 213.950 ;
        RECT 26.480 213.800 30.330 213.950 ;
        RECT 19.130 213.350 19.430 213.800 ;
        RECT 30.030 213.350 30.330 213.800 ;
        RECT 19.130 213.200 22.980 213.350 ;
        RECT 26.480 213.200 30.330 213.350 ;
        RECT 19.130 212.750 19.430 213.200 ;
        RECT 19.130 212.600 22.980 212.750 ;
        RECT 19.130 212.150 19.430 212.600 ;
        RECT 19.130 212.000 22.980 212.150 ;
        RECT 19.130 211.550 19.430 212.000 ;
        RECT 19.130 211.400 22.980 211.550 ;
        RECT 19.130 210.950 19.430 211.400 ;
        RECT 19.130 210.800 22.980 210.950 ;
        RECT 19.130 210.350 19.430 210.800 ;
        RECT 15.530 201.450 15.680 209.650 ;
        RECT 16.130 201.450 16.280 209.650 ;
        RECT 16.730 201.450 16.880 209.650 ;
        RECT 17.330 201.450 17.480 209.650 ;
        RECT 17.930 201.450 18.080 209.650 ;
        RECT 18.530 201.450 18.680 209.650 ;
        RECT 19.130 209.200 19.430 209.650 ;
        RECT 19.130 209.050 22.980 209.200 ;
        RECT 19.130 208.600 19.430 209.050 ;
        RECT 19.130 208.450 22.980 208.600 ;
        RECT 19.130 208.000 19.430 208.450 ;
        RECT 19.130 207.850 22.980 208.000 ;
        RECT 19.130 207.400 19.430 207.850 ;
        RECT 19.130 207.250 22.980 207.400 ;
        RECT 19.130 206.800 19.430 207.250 ;
        RECT 23.830 206.800 25.630 213.200 ;
        RECT 30.030 212.750 30.330 213.200 ;
        RECT 26.480 212.600 30.330 212.750 ;
        RECT 30.030 212.150 30.330 212.600 ;
        RECT 26.480 212.000 30.330 212.150 ;
        RECT 30.030 211.550 30.330 212.000 ;
        RECT 26.480 211.400 30.330 211.550 ;
        RECT 30.030 210.950 30.330 211.400 ;
        RECT 26.480 210.800 30.330 210.950 ;
        RECT 30.030 210.350 30.330 210.800 ;
        RECT 30.780 210.350 30.930 218.550 ;
        RECT 31.380 210.350 31.530 218.550 ;
        RECT 31.980 210.350 32.130 218.550 ;
        RECT 32.580 210.350 32.730 218.550 ;
        RECT 33.180 210.350 33.330 218.550 ;
        RECT 33.780 210.350 33.930 218.550 ;
        RECT 30.030 209.200 30.330 209.650 ;
        RECT 26.480 209.050 30.330 209.200 ;
        RECT 30.030 208.600 30.330 209.050 ;
        RECT 26.480 208.450 30.330 208.600 ;
        RECT 30.030 208.000 30.330 208.450 ;
        RECT 26.480 207.850 30.330 208.000 ;
        RECT 30.030 207.400 30.330 207.850 ;
        RECT 26.480 207.250 30.330 207.400 ;
        RECT 30.030 206.800 30.330 207.250 ;
        RECT 19.130 206.650 22.980 206.800 ;
        RECT 26.480 206.650 30.330 206.800 ;
        RECT 19.130 206.200 19.430 206.650 ;
        RECT 30.030 206.200 30.330 206.650 ;
        RECT 19.130 206.050 22.980 206.200 ;
        RECT 26.480 206.050 30.330 206.200 ;
        RECT 19.130 205.600 19.430 206.050 ;
        RECT 30.030 205.600 30.330 206.050 ;
        RECT 19.130 205.450 22.980 205.600 ;
        RECT 26.480 205.450 30.330 205.600 ;
        RECT 19.130 205.000 19.430 205.450 ;
        RECT 30.030 205.000 30.330 205.450 ;
        RECT 19.130 204.850 22.980 205.000 ;
        RECT 26.480 204.850 30.330 205.000 ;
        RECT 19.130 204.400 19.430 204.850 ;
        RECT 30.030 204.400 30.330 204.850 ;
        RECT 19.130 204.250 22.980 204.400 ;
        RECT 26.480 204.250 30.330 204.400 ;
        RECT 19.130 203.800 19.430 204.250 ;
        RECT 30.030 203.800 30.330 204.250 ;
        RECT 19.130 203.650 22.980 203.800 ;
        RECT 26.480 203.650 30.330 203.800 ;
        RECT 19.130 203.200 19.430 203.650 ;
        RECT 30.030 203.200 30.330 203.650 ;
        RECT 19.130 203.050 22.980 203.200 ;
        RECT 26.480 203.050 30.330 203.200 ;
        RECT 19.130 202.600 19.430 203.050 ;
        RECT 30.030 202.600 30.330 203.050 ;
        RECT 19.130 202.450 22.980 202.600 ;
        RECT 26.480 202.450 30.330 202.600 ;
        RECT 19.130 202.000 19.430 202.450 ;
        RECT 30.030 202.000 30.330 202.450 ;
        RECT 19.130 201.450 22.930 202.000 ;
        RECT 6.530 201.400 22.930 201.450 ;
        RECT 26.530 201.450 30.330 202.000 ;
        RECT 30.780 201.450 30.930 209.650 ;
        RECT 31.380 201.450 31.530 209.650 ;
        RECT 31.980 201.450 32.130 209.650 ;
        RECT 32.580 201.450 32.730 209.650 ;
        RECT 33.180 201.450 33.330 209.650 ;
        RECT 33.780 201.450 33.930 209.650 ;
        RECT 34.380 201.450 35.080 218.550 ;
        RECT 35.530 210.350 35.680 218.550 ;
        RECT 36.130 210.350 36.280 218.550 ;
        RECT 36.730 210.350 36.880 218.550 ;
        RECT 37.330 210.350 37.480 218.550 ;
        RECT 37.930 210.350 38.080 218.550 ;
        RECT 38.530 210.350 38.680 218.550 ;
        RECT 39.130 218.000 42.930 218.550 ;
        RECT 46.530 218.550 62.930 218.600 ;
        RECT 46.530 218.000 50.330 218.550 ;
        RECT 39.130 217.550 39.430 218.000 ;
        RECT 50.030 217.550 50.330 218.000 ;
        RECT 39.130 217.400 42.980 217.550 ;
        RECT 46.480 217.400 50.330 217.550 ;
        RECT 39.130 216.950 39.430 217.400 ;
        RECT 50.030 216.950 50.330 217.400 ;
        RECT 39.130 216.800 42.980 216.950 ;
        RECT 46.480 216.800 50.330 216.950 ;
        RECT 39.130 216.350 39.430 216.800 ;
        RECT 50.030 216.350 50.330 216.800 ;
        RECT 39.130 216.200 42.980 216.350 ;
        RECT 46.480 216.200 50.330 216.350 ;
        RECT 39.130 215.750 39.430 216.200 ;
        RECT 50.030 215.750 50.330 216.200 ;
        RECT 39.130 215.600 42.980 215.750 ;
        RECT 46.480 215.600 50.330 215.750 ;
        RECT 39.130 215.150 39.430 215.600 ;
        RECT 50.030 215.150 50.330 215.600 ;
        RECT 39.130 215.000 42.980 215.150 ;
        RECT 46.480 215.000 50.330 215.150 ;
        RECT 39.130 214.550 39.430 215.000 ;
        RECT 50.030 214.550 50.330 215.000 ;
        RECT 39.130 214.400 42.980 214.550 ;
        RECT 46.480 214.400 50.330 214.550 ;
        RECT 39.130 213.950 39.430 214.400 ;
        RECT 50.030 213.950 50.330 214.400 ;
        RECT 39.130 213.800 42.980 213.950 ;
        RECT 46.480 213.800 50.330 213.950 ;
        RECT 39.130 213.350 39.430 213.800 ;
        RECT 50.030 213.350 50.330 213.800 ;
        RECT 39.130 213.200 42.980 213.350 ;
        RECT 46.480 213.200 50.330 213.350 ;
        RECT 39.130 212.750 39.430 213.200 ;
        RECT 39.130 212.600 42.980 212.750 ;
        RECT 39.130 212.150 39.430 212.600 ;
        RECT 39.130 212.000 42.980 212.150 ;
        RECT 39.130 211.550 39.430 212.000 ;
        RECT 39.130 211.400 42.980 211.550 ;
        RECT 39.130 210.950 39.430 211.400 ;
        RECT 39.130 210.800 42.980 210.950 ;
        RECT 39.130 210.350 39.430 210.800 ;
        RECT 35.530 201.450 35.680 209.650 ;
        RECT 36.130 201.450 36.280 209.650 ;
        RECT 36.730 201.450 36.880 209.650 ;
        RECT 37.330 201.450 37.480 209.650 ;
        RECT 37.930 201.450 38.080 209.650 ;
        RECT 38.530 201.450 38.680 209.650 ;
        RECT 39.130 209.200 39.430 209.650 ;
        RECT 39.130 209.050 42.980 209.200 ;
        RECT 39.130 208.600 39.430 209.050 ;
        RECT 39.130 208.450 42.980 208.600 ;
        RECT 39.130 208.000 39.430 208.450 ;
        RECT 39.130 207.850 42.980 208.000 ;
        RECT 39.130 207.400 39.430 207.850 ;
        RECT 39.130 207.250 42.980 207.400 ;
        RECT 39.130 206.800 39.430 207.250 ;
        RECT 43.830 206.800 45.630 213.200 ;
        RECT 50.030 212.750 50.330 213.200 ;
        RECT 46.480 212.600 50.330 212.750 ;
        RECT 50.030 212.150 50.330 212.600 ;
        RECT 46.480 212.000 50.330 212.150 ;
        RECT 50.030 211.550 50.330 212.000 ;
        RECT 46.480 211.400 50.330 211.550 ;
        RECT 50.030 210.950 50.330 211.400 ;
        RECT 46.480 210.800 50.330 210.950 ;
        RECT 50.030 210.350 50.330 210.800 ;
        RECT 50.780 210.350 50.930 218.550 ;
        RECT 51.380 210.350 51.530 218.550 ;
        RECT 51.980 210.350 52.130 218.550 ;
        RECT 52.580 210.350 52.730 218.550 ;
        RECT 53.180 210.350 53.330 218.550 ;
        RECT 53.780 210.350 53.930 218.550 ;
        RECT 50.030 209.200 50.330 209.650 ;
        RECT 46.480 209.050 50.330 209.200 ;
        RECT 50.030 208.600 50.330 209.050 ;
        RECT 46.480 208.450 50.330 208.600 ;
        RECT 50.030 208.000 50.330 208.450 ;
        RECT 46.480 207.850 50.330 208.000 ;
        RECT 50.030 207.400 50.330 207.850 ;
        RECT 46.480 207.250 50.330 207.400 ;
        RECT 50.030 206.800 50.330 207.250 ;
        RECT 39.130 206.650 42.980 206.800 ;
        RECT 46.480 206.650 50.330 206.800 ;
        RECT 39.130 206.200 39.430 206.650 ;
        RECT 50.030 206.200 50.330 206.650 ;
        RECT 39.130 206.050 42.980 206.200 ;
        RECT 46.480 206.050 50.330 206.200 ;
        RECT 39.130 205.600 39.430 206.050 ;
        RECT 50.030 205.600 50.330 206.050 ;
        RECT 39.130 205.450 42.980 205.600 ;
        RECT 46.480 205.450 50.330 205.600 ;
        RECT 39.130 205.000 39.430 205.450 ;
        RECT 50.030 205.000 50.330 205.450 ;
        RECT 39.130 204.850 42.980 205.000 ;
        RECT 46.480 204.850 50.330 205.000 ;
        RECT 39.130 204.400 39.430 204.850 ;
        RECT 50.030 204.400 50.330 204.850 ;
        RECT 39.130 204.250 42.980 204.400 ;
        RECT 46.480 204.250 50.330 204.400 ;
        RECT 39.130 203.800 39.430 204.250 ;
        RECT 50.030 203.800 50.330 204.250 ;
        RECT 39.130 203.650 42.980 203.800 ;
        RECT 46.480 203.650 50.330 203.800 ;
        RECT 39.130 203.200 39.430 203.650 ;
        RECT 50.030 203.200 50.330 203.650 ;
        RECT 39.130 203.050 42.980 203.200 ;
        RECT 46.480 203.050 50.330 203.200 ;
        RECT 39.130 202.600 39.430 203.050 ;
        RECT 50.030 202.600 50.330 203.050 ;
        RECT 39.130 202.450 42.980 202.600 ;
        RECT 46.480 202.450 50.330 202.600 ;
        RECT 39.130 202.000 39.430 202.450 ;
        RECT 50.030 202.000 50.330 202.450 ;
        RECT 39.130 201.450 42.930 202.000 ;
        RECT 26.530 201.400 42.930 201.450 ;
        RECT 46.530 201.450 50.330 202.000 ;
        RECT 50.780 201.450 50.930 209.650 ;
        RECT 51.380 201.450 51.530 209.650 ;
        RECT 51.980 201.450 52.130 209.650 ;
        RECT 52.580 201.450 52.730 209.650 ;
        RECT 53.180 201.450 53.330 209.650 ;
        RECT 53.780 201.450 53.930 209.650 ;
        RECT 54.380 201.450 55.080 218.550 ;
        RECT 55.530 210.350 55.680 218.550 ;
        RECT 56.130 210.350 56.280 218.550 ;
        RECT 56.730 210.350 56.880 218.550 ;
        RECT 57.330 210.350 57.480 218.550 ;
        RECT 57.930 210.350 58.080 218.550 ;
        RECT 58.530 210.350 58.680 218.550 ;
        RECT 59.130 218.000 62.930 218.550 ;
        RECT 66.530 218.550 82.930 218.600 ;
        RECT 66.530 218.000 70.330 218.550 ;
        RECT 59.130 217.550 59.430 218.000 ;
        RECT 70.030 217.550 70.330 218.000 ;
        RECT 59.130 217.400 62.980 217.550 ;
        RECT 66.480 217.400 70.330 217.550 ;
        RECT 59.130 216.950 59.430 217.400 ;
        RECT 70.030 216.950 70.330 217.400 ;
        RECT 59.130 216.800 62.980 216.950 ;
        RECT 66.480 216.800 70.330 216.950 ;
        RECT 59.130 216.350 59.430 216.800 ;
        RECT 70.030 216.350 70.330 216.800 ;
        RECT 59.130 216.200 62.980 216.350 ;
        RECT 66.480 216.200 70.330 216.350 ;
        RECT 59.130 215.750 59.430 216.200 ;
        RECT 70.030 215.750 70.330 216.200 ;
        RECT 59.130 215.600 62.980 215.750 ;
        RECT 66.480 215.600 70.330 215.750 ;
        RECT 59.130 215.150 59.430 215.600 ;
        RECT 70.030 215.150 70.330 215.600 ;
        RECT 59.130 215.000 62.980 215.150 ;
        RECT 66.480 215.000 70.330 215.150 ;
        RECT 59.130 214.550 59.430 215.000 ;
        RECT 70.030 214.550 70.330 215.000 ;
        RECT 59.130 214.400 62.980 214.550 ;
        RECT 66.480 214.400 70.330 214.550 ;
        RECT 59.130 213.950 59.430 214.400 ;
        RECT 70.030 213.950 70.330 214.400 ;
        RECT 59.130 213.800 62.980 213.950 ;
        RECT 66.480 213.800 70.330 213.950 ;
        RECT 59.130 213.350 59.430 213.800 ;
        RECT 70.030 213.350 70.330 213.800 ;
        RECT 59.130 213.200 62.980 213.350 ;
        RECT 66.480 213.200 70.330 213.350 ;
        RECT 59.130 212.750 59.430 213.200 ;
        RECT 59.130 212.600 62.980 212.750 ;
        RECT 59.130 212.150 59.430 212.600 ;
        RECT 59.130 212.000 62.980 212.150 ;
        RECT 59.130 211.550 59.430 212.000 ;
        RECT 59.130 211.400 62.980 211.550 ;
        RECT 59.130 210.950 59.430 211.400 ;
        RECT 59.130 210.800 62.980 210.950 ;
        RECT 59.130 210.350 59.430 210.800 ;
        RECT 55.530 201.450 55.680 209.650 ;
        RECT 56.130 201.450 56.280 209.650 ;
        RECT 56.730 201.450 56.880 209.650 ;
        RECT 57.330 201.450 57.480 209.650 ;
        RECT 57.930 201.450 58.080 209.650 ;
        RECT 58.530 201.450 58.680 209.650 ;
        RECT 59.130 209.200 59.430 209.650 ;
        RECT 59.130 209.050 62.980 209.200 ;
        RECT 59.130 208.600 59.430 209.050 ;
        RECT 59.130 208.450 62.980 208.600 ;
        RECT 59.130 208.000 59.430 208.450 ;
        RECT 59.130 207.850 62.980 208.000 ;
        RECT 59.130 207.400 59.430 207.850 ;
        RECT 59.130 207.250 62.980 207.400 ;
        RECT 59.130 206.800 59.430 207.250 ;
        RECT 63.830 206.800 65.630 213.200 ;
        RECT 70.030 212.750 70.330 213.200 ;
        RECT 66.480 212.600 70.330 212.750 ;
        RECT 70.030 212.150 70.330 212.600 ;
        RECT 66.480 212.000 70.330 212.150 ;
        RECT 70.030 211.550 70.330 212.000 ;
        RECT 66.480 211.400 70.330 211.550 ;
        RECT 70.030 210.950 70.330 211.400 ;
        RECT 66.480 210.800 70.330 210.950 ;
        RECT 70.030 210.350 70.330 210.800 ;
        RECT 70.780 210.350 70.930 218.550 ;
        RECT 71.380 210.350 71.530 218.550 ;
        RECT 71.980 210.350 72.130 218.550 ;
        RECT 72.580 210.350 72.730 218.550 ;
        RECT 73.180 210.350 73.330 218.550 ;
        RECT 73.780 210.350 73.930 218.550 ;
        RECT 70.030 209.200 70.330 209.650 ;
        RECT 66.480 209.050 70.330 209.200 ;
        RECT 70.030 208.600 70.330 209.050 ;
        RECT 66.480 208.450 70.330 208.600 ;
        RECT 70.030 208.000 70.330 208.450 ;
        RECT 66.480 207.850 70.330 208.000 ;
        RECT 70.030 207.400 70.330 207.850 ;
        RECT 66.480 207.250 70.330 207.400 ;
        RECT 70.030 206.800 70.330 207.250 ;
        RECT 59.130 206.650 62.980 206.800 ;
        RECT 66.480 206.650 70.330 206.800 ;
        RECT 59.130 206.200 59.430 206.650 ;
        RECT 70.030 206.200 70.330 206.650 ;
        RECT 59.130 206.050 62.980 206.200 ;
        RECT 66.480 206.050 70.330 206.200 ;
        RECT 59.130 205.600 59.430 206.050 ;
        RECT 70.030 205.600 70.330 206.050 ;
        RECT 59.130 205.450 62.980 205.600 ;
        RECT 66.480 205.450 70.330 205.600 ;
        RECT 59.130 205.000 59.430 205.450 ;
        RECT 70.030 205.000 70.330 205.450 ;
        RECT 59.130 204.850 62.980 205.000 ;
        RECT 66.480 204.850 70.330 205.000 ;
        RECT 59.130 204.400 59.430 204.850 ;
        RECT 70.030 204.400 70.330 204.850 ;
        RECT 59.130 204.250 62.980 204.400 ;
        RECT 66.480 204.250 70.330 204.400 ;
        RECT 59.130 203.800 59.430 204.250 ;
        RECT 70.030 203.800 70.330 204.250 ;
        RECT 59.130 203.650 62.980 203.800 ;
        RECT 66.480 203.650 70.330 203.800 ;
        RECT 59.130 203.200 59.430 203.650 ;
        RECT 70.030 203.200 70.330 203.650 ;
        RECT 59.130 203.050 62.980 203.200 ;
        RECT 66.480 203.050 70.330 203.200 ;
        RECT 59.130 202.600 59.430 203.050 ;
        RECT 70.030 202.600 70.330 203.050 ;
        RECT 59.130 202.450 62.980 202.600 ;
        RECT 66.480 202.450 70.330 202.600 ;
        RECT 59.130 202.000 59.430 202.450 ;
        RECT 70.030 202.000 70.330 202.450 ;
        RECT 59.130 201.450 62.930 202.000 ;
        RECT 46.530 201.400 62.930 201.450 ;
        RECT 66.530 201.450 70.330 202.000 ;
        RECT 70.780 201.450 70.930 209.650 ;
        RECT 71.380 201.450 71.530 209.650 ;
        RECT 71.980 201.450 72.130 209.650 ;
        RECT 72.580 201.450 72.730 209.650 ;
        RECT 73.180 201.450 73.330 209.650 ;
        RECT 73.780 201.450 73.930 209.650 ;
        RECT 74.380 201.450 75.080 218.550 ;
        RECT 75.530 210.350 75.680 218.550 ;
        RECT 76.130 210.350 76.280 218.550 ;
        RECT 76.730 210.350 76.880 218.550 ;
        RECT 77.330 210.350 77.480 218.550 ;
        RECT 77.930 210.350 78.080 218.550 ;
        RECT 78.530 210.350 78.680 218.550 ;
        RECT 79.130 218.000 82.930 218.550 ;
        RECT 86.530 218.550 102.930 218.600 ;
        RECT 86.530 218.000 90.330 218.550 ;
        RECT 79.130 217.550 79.430 218.000 ;
        RECT 90.030 217.550 90.330 218.000 ;
        RECT 79.130 217.400 82.980 217.550 ;
        RECT 86.480 217.400 90.330 217.550 ;
        RECT 79.130 216.950 79.430 217.400 ;
        RECT 90.030 216.950 90.330 217.400 ;
        RECT 79.130 216.800 82.980 216.950 ;
        RECT 86.480 216.800 90.330 216.950 ;
        RECT 79.130 216.350 79.430 216.800 ;
        RECT 90.030 216.350 90.330 216.800 ;
        RECT 79.130 216.200 82.980 216.350 ;
        RECT 86.480 216.200 90.330 216.350 ;
        RECT 79.130 215.750 79.430 216.200 ;
        RECT 90.030 215.750 90.330 216.200 ;
        RECT 79.130 215.600 82.980 215.750 ;
        RECT 86.480 215.600 90.330 215.750 ;
        RECT 79.130 215.150 79.430 215.600 ;
        RECT 90.030 215.150 90.330 215.600 ;
        RECT 79.130 215.000 82.980 215.150 ;
        RECT 86.480 215.000 90.330 215.150 ;
        RECT 79.130 214.550 79.430 215.000 ;
        RECT 90.030 214.550 90.330 215.000 ;
        RECT 79.130 214.400 82.980 214.550 ;
        RECT 86.480 214.400 90.330 214.550 ;
        RECT 79.130 213.950 79.430 214.400 ;
        RECT 90.030 213.950 90.330 214.400 ;
        RECT 79.130 213.800 82.980 213.950 ;
        RECT 86.480 213.800 90.330 213.950 ;
        RECT 79.130 213.350 79.430 213.800 ;
        RECT 90.030 213.350 90.330 213.800 ;
        RECT 79.130 213.200 82.980 213.350 ;
        RECT 86.480 213.200 90.330 213.350 ;
        RECT 79.130 212.750 79.430 213.200 ;
        RECT 79.130 212.600 82.980 212.750 ;
        RECT 79.130 212.150 79.430 212.600 ;
        RECT 79.130 212.000 82.980 212.150 ;
        RECT 79.130 211.550 79.430 212.000 ;
        RECT 79.130 211.400 82.980 211.550 ;
        RECT 79.130 210.950 79.430 211.400 ;
        RECT 79.130 210.800 82.980 210.950 ;
        RECT 79.130 210.350 79.430 210.800 ;
        RECT 75.530 201.450 75.680 209.650 ;
        RECT 76.130 201.450 76.280 209.650 ;
        RECT 76.730 201.450 76.880 209.650 ;
        RECT 77.330 201.450 77.480 209.650 ;
        RECT 77.930 201.450 78.080 209.650 ;
        RECT 78.530 201.450 78.680 209.650 ;
        RECT 79.130 209.200 79.430 209.650 ;
        RECT 79.130 209.050 82.980 209.200 ;
        RECT 79.130 208.600 79.430 209.050 ;
        RECT 79.130 208.450 82.980 208.600 ;
        RECT 79.130 208.000 79.430 208.450 ;
        RECT 79.130 207.850 82.980 208.000 ;
        RECT 79.130 207.400 79.430 207.850 ;
        RECT 79.130 207.250 82.980 207.400 ;
        RECT 79.130 206.800 79.430 207.250 ;
        RECT 83.830 206.800 85.630 213.200 ;
        RECT 90.030 212.750 90.330 213.200 ;
        RECT 86.480 212.600 90.330 212.750 ;
        RECT 90.030 212.150 90.330 212.600 ;
        RECT 86.480 212.000 90.330 212.150 ;
        RECT 90.030 211.550 90.330 212.000 ;
        RECT 86.480 211.400 90.330 211.550 ;
        RECT 90.030 210.950 90.330 211.400 ;
        RECT 86.480 210.800 90.330 210.950 ;
        RECT 90.030 210.350 90.330 210.800 ;
        RECT 90.780 210.350 90.930 218.550 ;
        RECT 91.380 210.350 91.530 218.550 ;
        RECT 91.980 210.350 92.130 218.550 ;
        RECT 92.580 210.350 92.730 218.550 ;
        RECT 93.180 210.350 93.330 218.550 ;
        RECT 93.780 210.350 93.930 218.550 ;
        RECT 90.030 209.200 90.330 209.650 ;
        RECT 86.480 209.050 90.330 209.200 ;
        RECT 90.030 208.600 90.330 209.050 ;
        RECT 86.480 208.450 90.330 208.600 ;
        RECT 90.030 208.000 90.330 208.450 ;
        RECT 86.480 207.850 90.330 208.000 ;
        RECT 90.030 207.400 90.330 207.850 ;
        RECT 86.480 207.250 90.330 207.400 ;
        RECT 90.030 206.800 90.330 207.250 ;
        RECT 79.130 206.650 82.980 206.800 ;
        RECT 86.480 206.650 90.330 206.800 ;
        RECT 79.130 206.200 79.430 206.650 ;
        RECT 90.030 206.200 90.330 206.650 ;
        RECT 79.130 206.050 82.980 206.200 ;
        RECT 86.480 206.050 90.330 206.200 ;
        RECT 79.130 205.600 79.430 206.050 ;
        RECT 90.030 205.600 90.330 206.050 ;
        RECT 79.130 205.450 82.980 205.600 ;
        RECT 86.480 205.450 90.330 205.600 ;
        RECT 79.130 205.000 79.430 205.450 ;
        RECT 90.030 205.000 90.330 205.450 ;
        RECT 79.130 204.850 82.980 205.000 ;
        RECT 86.480 204.850 90.330 205.000 ;
        RECT 79.130 204.400 79.430 204.850 ;
        RECT 90.030 204.400 90.330 204.850 ;
        RECT 79.130 204.250 82.980 204.400 ;
        RECT 86.480 204.250 90.330 204.400 ;
        RECT 79.130 203.800 79.430 204.250 ;
        RECT 90.030 203.800 90.330 204.250 ;
        RECT 79.130 203.650 82.980 203.800 ;
        RECT 86.480 203.650 90.330 203.800 ;
        RECT 79.130 203.200 79.430 203.650 ;
        RECT 90.030 203.200 90.330 203.650 ;
        RECT 79.130 203.050 82.980 203.200 ;
        RECT 86.480 203.050 90.330 203.200 ;
        RECT 79.130 202.600 79.430 203.050 ;
        RECT 90.030 202.600 90.330 203.050 ;
        RECT 79.130 202.450 82.980 202.600 ;
        RECT 86.480 202.450 90.330 202.600 ;
        RECT 79.130 202.000 79.430 202.450 ;
        RECT 90.030 202.000 90.330 202.450 ;
        RECT 79.130 201.450 82.930 202.000 ;
        RECT 66.530 201.400 82.930 201.450 ;
        RECT 86.530 201.450 90.330 202.000 ;
        RECT 90.780 201.450 90.930 209.650 ;
        RECT 91.380 201.450 91.530 209.650 ;
        RECT 91.980 201.450 92.130 209.650 ;
        RECT 92.580 201.450 92.730 209.650 ;
        RECT 93.180 201.450 93.330 209.650 ;
        RECT 93.780 201.450 93.930 209.650 ;
        RECT 94.380 201.450 95.080 218.550 ;
        RECT 95.530 210.350 95.680 218.550 ;
        RECT 96.130 210.350 96.280 218.550 ;
        RECT 96.730 210.350 96.880 218.550 ;
        RECT 97.330 210.350 97.480 218.550 ;
        RECT 97.930 210.350 98.080 218.550 ;
        RECT 98.530 210.350 98.680 218.550 ;
        RECT 99.130 218.000 102.930 218.550 ;
        RECT 106.530 218.550 122.930 218.600 ;
        RECT 106.530 218.000 110.330 218.550 ;
        RECT 99.130 217.550 99.430 218.000 ;
        RECT 110.030 217.550 110.330 218.000 ;
        RECT 99.130 217.400 102.980 217.550 ;
        RECT 106.480 217.400 110.330 217.550 ;
        RECT 99.130 216.950 99.430 217.400 ;
        RECT 110.030 216.950 110.330 217.400 ;
        RECT 99.130 216.800 102.980 216.950 ;
        RECT 106.480 216.800 110.330 216.950 ;
        RECT 99.130 216.350 99.430 216.800 ;
        RECT 110.030 216.350 110.330 216.800 ;
        RECT 99.130 216.200 102.980 216.350 ;
        RECT 106.480 216.200 110.330 216.350 ;
        RECT 99.130 215.750 99.430 216.200 ;
        RECT 110.030 215.750 110.330 216.200 ;
        RECT 99.130 215.600 102.980 215.750 ;
        RECT 106.480 215.600 110.330 215.750 ;
        RECT 99.130 215.150 99.430 215.600 ;
        RECT 110.030 215.150 110.330 215.600 ;
        RECT 99.130 215.000 102.980 215.150 ;
        RECT 106.480 215.000 110.330 215.150 ;
        RECT 99.130 214.550 99.430 215.000 ;
        RECT 110.030 214.550 110.330 215.000 ;
        RECT 99.130 214.400 102.980 214.550 ;
        RECT 106.480 214.400 110.330 214.550 ;
        RECT 99.130 213.950 99.430 214.400 ;
        RECT 110.030 213.950 110.330 214.400 ;
        RECT 99.130 213.800 102.980 213.950 ;
        RECT 106.480 213.800 110.330 213.950 ;
        RECT 99.130 213.350 99.430 213.800 ;
        RECT 110.030 213.350 110.330 213.800 ;
        RECT 99.130 213.200 102.980 213.350 ;
        RECT 106.480 213.200 110.330 213.350 ;
        RECT 99.130 212.750 99.430 213.200 ;
        RECT 99.130 212.600 102.980 212.750 ;
        RECT 99.130 212.150 99.430 212.600 ;
        RECT 99.130 212.000 102.980 212.150 ;
        RECT 99.130 211.550 99.430 212.000 ;
        RECT 99.130 211.400 102.980 211.550 ;
        RECT 99.130 210.950 99.430 211.400 ;
        RECT 99.130 210.800 102.980 210.950 ;
        RECT 99.130 210.350 99.430 210.800 ;
        RECT 95.530 201.450 95.680 209.650 ;
        RECT 96.130 201.450 96.280 209.650 ;
        RECT 96.730 201.450 96.880 209.650 ;
        RECT 97.330 201.450 97.480 209.650 ;
        RECT 97.930 201.450 98.080 209.650 ;
        RECT 98.530 201.450 98.680 209.650 ;
        RECT 99.130 209.200 99.430 209.650 ;
        RECT 99.130 209.050 102.980 209.200 ;
        RECT 99.130 208.600 99.430 209.050 ;
        RECT 99.130 208.450 102.980 208.600 ;
        RECT 99.130 208.000 99.430 208.450 ;
        RECT 99.130 207.850 102.980 208.000 ;
        RECT 99.130 207.400 99.430 207.850 ;
        RECT 99.130 207.250 102.980 207.400 ;
        RECT 99.130 206.800 99.430 207.250 ;
        RECT 103.830 206.800 105.630 213.200 ;
        RECT 110.030 212.750 110.330 213.200 ;
        RECT 106.480 212.600 110.330 212.750 ;
        RECT 110.030 212.150 110.330 212.600 ;
        RECT 106.480 212.000 110.330 212.150 ;
        RECT 110.030 211.550 110.330 212.000 ;
        RECT 106.480 211.400 110.330 211.550 ;
        RECT 110.030 210.950 110.330 211.400 ;
        RECT 106.480 210.800 110.330 210.950 ;
        RECT 110.030 210.350 110.330 210.800 ;
        RECT 110.780 210.350 110.930 218.550 ;
        RECT 111.380 210.350 111.530 218.550 ;
        RECT 111.980 210.350 112.130 218.550 ;
        RECT 112.580 210.350 112.730 218.550 ;
        RECT 113.180 210.350 113.330 218.550 ;
        RECT 113.780 210.350 113.930 218.550 ;
        RECT 110.030 209.200 110.330 209.650 ;
        RECT 106.480 209.050 110.330 209.200 ;
        RECT 110.030 208.600 110.330 209.050 ;
        RECT 106.480 208.450 110.330 208.600 ;
        RECT 110.030 208.000 110.330 208.450 ;
        RECT 106.480 207.850 110.330 208.000 ;
        RECT 110.030 207.400 110.330 207.850 ;
        RECT 106.480 207.250 110.330 207.400 ;
        RECT 110.030 206.800 110.330 207.250 ;
        RECT 99.130 206.650 102.980 206.800 ;
        RECT 106.480 206.650 110.330 206.800 ;
        RECT 99.130 206.200 99.430 206.650 ;
        RECT 110.030 206.200 110.330 206.650 ;
        RECT 99.130 206.050 102.980 206.200 ;
        RECT 106.480 206.050 110.330 206.200 ;
        RECT 99.130 205.600 99.430 206.050 ;
        RECT 110.030 205.600 110.330 206.050 ;
        RECT 99.130 205.450 102.980 205.600 ;
        RECT 106.480 205.450 110.330 205.600 ;
        RECT 99.130 205.000 99.430 205.450 ;
        RECT 110.030 205.000 110.330 205.450 ;
        RECT 99.130 204.850 102.980 205.000 ;
        RECT 106.480 204.850 110.330 205.000 ;
        RECT 99.130 204.400 99.430 204.850 ;
        RECT 110.030 204.400 110.330 204.850 ;
        RECT 99.130 204.250 102.980 204.400 ;
        RECT 106.480 204.250 110.330 204.400 ;
        RECT 99.130 203.800 99.430 204.250 ;
        RECT 110.030 203.800 110.330 204.250 ;
        RECT 99.130 203.650 102.980 203.800 ;
        RECT 106.480 203.650 110.330 203.800 ;
        RECT 99.130 203.200 99.430 203.650 ;
        RECT 110.030 203.200 110.330 203.650 ;
        RECT 99.130 203.050 102.980 203.200 ;
        RECT 106.480 203.050 110.330 203.200 ;
        RECT 99.130 202.600 99.430 203.050 ;
        RECT 110.030 202.600 110.330 203.050 ;
        RECT 99.130 202.450 102.980 202.600 ;
        RECT 106.480 202.450 110.330 202.600 ;
        RECT 99.130 202.000 99.430 202.450 ;
        RECT 110.030 202.000 110.330 202.450 ;
        RECT 99.130 201.450 102.930 202.000 ;
        RECT 86.530 201.400 102.930 201.450 ;
        RECT 106.530 201.450 110.330 202.000 ;
        RECT 110.780 201.450 110.930 209.650 ;
        RECT 111.380 201.450 111.530 209.650 ;
        RECT 111.980 201.450 112.130 209.650 ;
        RECT 112.580 201.450 112.730 209.650 ;
        RECT 113.180 201.450 113.330 209.650 ;
        RECT 113.780 201.450 113.930 209.650 ;
        RECT 114.380 201.450 115.080 218.550 ;
        RECT 115.530 210.350 115.680 218.550 ;
        RECT 116.130 210.350 116.280 218.550 ;
        RECT 116.730 210.350 116.880 218.550 ;
        RECT 117.330 210.350 117.480 218.550 ;
        RECT 117.930 210.350 118.080 218.550 ;
        RECT 118.530 210.350 118.680 218.550 ;
        RECT 119.130 218.000 122.930 218.550 ;
        RECT 119.130 217.550 119.430 218.000 ;
        RECT 119.130 217.400 122.980 217.550 ;
        RECT 119.130 216.950 119.430 217.400 ;
        RECT 119.130 216.800 122.980 216.950 ;
        RECT 119.130 216.350 119.430 216.800 ;
        RECT 119.130 216.200 122.980 216.350 ;
        RECT 119.130 215.750 119.430 216.200 ;
        RECT 119.130 215.600 122.980 215.750 ;
        RECT 119.130 215.150 119.430 215.600 ;
        RECT 119.130 215.000 122.980 215.150 ;
        RECT 119.130 214.550 119.430 215.000 ;
        RECT 119.130 214.400 122.980 214.550 ;
        RECT 119.130 213.950 119.430 214.400 ;
        RECT 119.130 213.800 122.980 213.950 ;
        RECT 119.130 213.350 119.430 213.800 ;
        RECT 119.130 213.200 122.980 213.350 ;
        RECT 119.130 212.750 119.430 213.200 ;
        RECT 119.130 212.600 122.980 212.750 ;
        RECT 119.130 212.150 119.430 212.600 ;
        RECT 119.130 212.000 122.980 212.150 ;
        RECT 119.130 211.550 119.430 212.000 ;
        RECT 119.130 211.400 122.980 211.550 ;
        RECT 119.130 210.950 119.430 211.400 ;
        RECT 119.130 210.800 122.980 210.950 ;
        RECT 119.130 210.350 119.430 210.800 ;
        RECT 115.530 201.450 115.680 209.650 ;
        RECT 116.130 201.450 116.280 209.650 ;
        RECT 116.730 201.450 116.880 209.650 ;
        RECT 117.330 201.450 117.480 209.650 ;
        RECT 117.930 201.450 118.080 209.650 ;
        RECT 118.530 201.450 118.680 209.650 ;
        RECT 119.130 209.200 119.430 209.650 ;
        RECT 119.130 209.050 122.980 209.200 ;
        RECT 119.130 208.600 119.430 209.050 ;
        RECT 119.130 208.450 122.980 208.600 ;
        RECT 119.130 208.000 119.430 208.450 ;
        RECT 119.130 207.850 122.980 208.000 ;
        RECT 119.130 207.400 119.430 207.850 ;
        RECT 119.130 207.250 122.980 207.400 ;
        RECT 119.130 206.800 119.430 207.250 ;
        RECT 123.830 206.800 124.730 213.200 ;
        RECT 129.850 208.350 131.850 209.625 ;
        RECT 119.130 206.650 122.980 206.800 ;
        RECT 119.130 206.200 119.430 206.650 ;
        RECT 119.130 206.050 122.980 206.200 ;
        RECT 119.130 205.600 119.430 206.050 ;
        RECT 119.130 205.450 122.980 205.600 ;
        RECT 119.130 205.000 119.430 205.450 ;
        RECT 119.130 204.850 122.980 205.000 ;
        RECT 119.130 204.400 119.430 204.850 ;
        RECT 119.130 204.250 122.980 204.400 ;
        RECT 119.130 203.800 119.430 204.250 ;
        RECT 119.130 203.650 122.980 203.800 ;
        RECT 119.130 203.200 119.430 203.650 ;
        RECT 119.130 203.050 122.980 203.200 ;
        RECT 119.130 202.600 119.430 203.050 ;
        RECT 119.130 202.450 122.980 202.600 ;
        RECT 119.130 202.000 119.430 202.450 ;
        RECT 119.130 201.450 122.930 202.000 ;
        RECT 106.530 201.400 122.930 201.450 ;
        RECT 9.630 200.900 19.830 201.400 ;
        RECT 29.630 200.900 39.830 201.400 ;
        RECT 49.630 200.900 59.830 201.400 ;
        RECT 69.630 200.900 79.830 201.400 ;
        RECT 89.630 200.900 99.830 201.400 ;
        RECT 109.630 200.900 119.830 201.400 ;
        RECT 11.530 200.000 17.930 200.900 ;
        RECT 31.530 200.000 37.930 200.900 ;
        RECT 51.530 200.000 57.930 200.900 ;
        RECT 71.530 200.000 77.930 200.900 ;
        RECT 91.530 200.000 97.930 200.900 ;
        RECT 111.530 200.000 117.930 200.900 ;
        RECT 12.340 178.555 14.335 200.000 ;
        RECT 9.335 177.190 14.340 178.555 ;
        RECT 9.340 177.050 11.335 177.190 ;
        RECT 9.340 176.350 11.675 177.050 ;
        RECT 9.340 144.680 11.335 176.350 ;
        RECT 9.340 143.550 13.710 144.680 ;
        RECT 9.330 142.425 13.710 143.550 ;
        RECT 11.530 140.000 13.710 142.425 ;
        RECT 11.530 139.100 17.930 140.000 ;
        RECT 31.530 139.100 37.930 140.000 ;
        RECT 51.530 139.100 57.930 140.000 ;
        RECT 71.530 139.100 77.930 140.000 ;
        RECT 91.530 139.100 97.930 140.000 ;
        RECT 111.530 139.100 117.930 140.000 ;
        RECT 9.630 138.600 19.830 139.100 ;
        RECT 29.630 138.600 39.830 139.100 ;
        RECT 49.630 138.600 59.830 139.100 ;
        RECT 69.630 138.600 79.830 139.100 ;
        RECT 89.630 138.600 99.830 139.100 ;
        RECT 109.630 138.600 119.830 139.100 ;
        RECT 6.530 138.550 22.930 138.600 ;
        RECT 6.530 138.000 10.330 138.550 ;
        RECT 10.030 137.550 10.330 138.000 ;
        RECT 6.480 137.400 10.330 137.550 ;
        RECT 10.030 136.950 10.330 137.400 ;
        RECT 6.480 136.800 10.330 136.950 ;
        RECT 10.030 136.350 10.330 136.800 ;
        RECT 6.480 136.200 10.330 136.350 ;
        RECT 10.030 135.750 10.330 136.200 ;
        RECT 6.480 135.600 10.330 135.750 ;
        RECT 10.030 135.150 10.330 135.600 ;
        RECT 6.480 135.000 10.330 135.150 ;
        RECT 10.030 134.550 10.330 135.000 ;
        RECT 6.480 134.400 10.330 134.550 ;
        RECT 10.030 133.950 10.330 134.400 ;
        RECT 6.480 133.800 10.330 133.950 ;
        RECT 10.030 133.350 10.330 133.800 ;
        RECT 6.480 133.200 10.330 133.350 ;
        RECT 4.730 126.800 5.630 133.200 ;
        RECT 10.030 132.750 10.330 133.200 ;
        RECT 6.480 132.600 10.330 132.750 ;
        RECT 10.030 132.150 10.330 132.600 ;
        RECT 6.480 132.000 10.330 132.150 ;
        RECT 10.030 131.550 10.330 132.000 ;
        RECT 6.480 131.400 10.330 131.550 ;
        RECT 10.030 130.950 10.330 131.400 ;
        RECT 6.480 130.800 10.330 130.950 ;
        RECT 10.030 130.350 10.330 130.800 ;
        RECT 10.780 130.350 10.930 138.550 ;
        RECT 11.380 130.350 11.530 138.550 ;
        RECT 11.980 130.350 12.130 138.550 ;
        RECT 12.580 130.350 12.730 138.550 ;
        RECT 13.180 130.350 13.330 138.550 ;
        RECT 13.780 130.350 13.930 138.550 ;
        RECT 10.030 129.200 10.330 129.650 ;
        RECT 6.480 129.050 10.330 129.200 ;
        RECT 10.030 128.600 10.330 129.050 ;
        RECT 6.480 128.450 10.330 128.600 ;
        RECT 10.030 128.000 10.330 128.450 ;
        RECT 6.480 127.850 10.330 128.000 ;
        RECT 10.030 127.400 10.330 127.850 ;
        RECT 6.480 127.250 10.330 127.400 ;
        RECT 10.030 126.800 10.330 127.250 ;
        RECT 6.480 126.650 10.330 126.800 ;
        RECT 10.030 126.200 10.330 126.650 ;
        RECT 6.480 126.050 10.330 126.200 ;
        RECT 10.030 125.600 10.330 126.050 ;
        RECT 6.480 125.450 10.330 125.600 ;
        RECT 10.030 125.000 10.330 125.450 ;
        RECT 6.480 124.850 10.330 125.000 ;
        RECT 10.030 124.400 10.330 124.850 ;
        RECT 6.480 124.250 10.330 124.400 ;
        RECT 10.030 123.800 10.330 124.250 ;
        RECT 6.480 123.650 10.330 123.800 ;
        RECT 10.030 123.200 10.330 123.650 ;
        RECT 6.480 123.050 10.330 123.200 ;
        RECT 10.030 122.600 10.330 123.050 ;
        RECT 6.480 122.450 10.330 122.600 ;
        RECT 10.030 122.000 10.330 122.450 ;
        RECT 6.530 121.450 10.330 122.000 ;
        RECT 10.780 121.450 10.930 129.650 ;
        RECT 11.380 121.450 11.530 129.650 ;
        RECT 11.980 121.450 12.130 129.650 ;
        RECT 12.580 121.450 12.730 129.650 ;
        RECT 13.180 121.450 13.330 129.650 ;
        RECT 13.780 121.450 13.930 129.650 ;
        RECT 14.380 121.450 15.080 138.550 ;
        RECT 15.530 130.350 15.680 138.550 ;
        RECT 16.130 130.350 16.280 138.550 ;
        RECT 16.730 130.350 16.880 138.550 ;
        RECT 17.330 130.350 17.480 138.550 ;
        RECT 17.930 130.350 18.080 138.550 ;
        RECT 18.530 130.350 18.680 138.550 ;
        RECT 19.130 138.000 22.930 138.550 ;
        RECT 26.530 138.550 42.930 138.600 ;
        RECT 26.530 138.000 30.330 138.550 ;
        RECT 19.130 137.550 19.430 138.000 ;
        RECT 30.030 137.550 30.330 138.000 ;
        RECT 19.130 137.400 22.980 137.550 ;
        RECT 26.480 137.400 30.330 137.550 ;
        RECT 19.130 136.950 19.430 137.400 ;
        RECT 30.030 136.950 30.330 137.400 ;
        RECT 19.130 136.800 22.980 136.950 ;
        RECT 26.480 136.800 30.330 136.950 ;
        RECT 19.130 136.350 19.430 136.800 ;
        RECT 30.030 136.350 30.330 136.800 ;
        RECT 19.130 136.200 22.980 136.350 ;
        RECT 26.480 136.200 30.330 136.350 ;
        RECT 19.130 135.750 19.430 136.200 ;
        RECT 30.030 135.750 30.330 136.200 ;
        RECT 19.130 135.600 22.980 135.750 ;
        RECT 26.480 135.600 30.330 135.750 ;
        RECT 19.130 135.150 19.430 135.600 ;
        RECT 30.030 135.150 30.330 135.600 ;
        RECT 19.130 135.000 22.980 135.150 ;
        RECT 26.480 135.000 30.330 135.150 ;
        RECT 19.130 134.550 19.430 135.000 ;
        RECT 30.030 134.550 30.330 135.000 ;
        RECT 19.130 134.400 22.980 134.550 ;
        RECT 26.480 134.400 30.330 134.550 ;
        RECT 19.130 133.950 19.430 134.400 ;
        RECT 30.030 133.950 30.330 134.400 ;
        RECT 19.130 133.800 22.980 133.950 ;
        RECT 26.480 133.800 30.330 133.950 ;
        RECT 19.130 133.350 19.430 133.800 ;
        RECT 30.030 133.350 30.330 133.800 ;
        RECT 19.130 133.200 22.980 133.350 ;
        RECT 26.480 133.200 30.330 133.350 ;
        RECT 19.130 132.750 19.430 133.200 ;
        RECT 19.130 132.600 22.980 132.750 ;
        RECT 19.130 132.150 19.430 132.600 ;
        RECT 19.130 132.000 22.980 132.150 ;
        RECT 19.130 131.550 19.430 132.000 ;
        RECT 19.130 131.400 22.980 131.550 ;
        RECT 19.130 130.950 19.430 131.400 ;
        RECT 19.130 130.800 22.980 130.950 ;
        RECT 19.130 130.350 19.430 130.800 ;
        RECT 15.530 121.450 15.680 129.650 ;
        RECT 16.130 121.450 16.280 129.650 ;
        RECT 16.730 121.450 16.880 129.650 ;
        RECT 17.330 121.450 17.480 129.650 ;
        RECT 17.930 121.450 18.080 129.650 ;
        RECT 18.530 121.450 18.680 129.650 ;
        RECT 19.130 129.200 19.430 129.650 ;
        RECT 19.130 129.050 22.980 129.200 ;
        RECT 19.130 128.600 19.430 129.050 ;
        RECT 19.130 128.450 22.980 128.600 ;
        RECT 19.130 128.000 19.430 128.450 ;
        RECT 19.130 127.850 22.980 128.000 ;
        RECT 19.130 127.400 19.430 127.850 ;
        RECT 19.130 127.250 22.980 127.400 ;
        RECT 19.130 126.800 19.430 127.250 ;
        RECT 23.830 126.800 25.630 133.200 ;
        RECT 30.030 132.750 30.330 133.200 ;
        RECT 26.480 132.600 30.330 132.750 ;
        RECT 30.030 132.150 30.330 132.600 ;
        RECT 26.480 132.000 30.330 132.150 ;
        RECT 30.030 131.550 30.330 132.000 ;
        RECT 26.480 131.400 30.330 131.550 ;
        RECT 30.030 130.950 30.330 131.400 ;
        RECT 26.480 130.800 30.330 130.950 ;
        RECT 30.030 130.350 30.330 130.800 ;
        RECT 30.780 130.350 30.930 138.550 ;
        RECT 31.380 130.350 31.530 138.550 ;
        RECT 31.980 130.350 32.130 138.550 ;
        RECT 32.580 130.350 32.730 138.550 ;
        RECT 33.180 130.350 33.330 138.550 ;
        RECT 33.780 130.350 33.930 138.550 ;
        RECT 30.030 129.200 30.330 129.650 ;
        RECT 26.480 129.050 30.330 129.200 ;
        RECT 30.030 128.600 30.330 129.050 ;
        RECT 26.480 128.450 30.330 128.600 ;
        RECT 30.030 128.000 30.330 128.450 ;
        RECT 26.480 127.850 30.330 128.000 ;
        RECT 30.030 127.400 30.330 127.850 ;
        RECT 26.480 127.250 30.330 127.400 ;
        RECT 30.030 126.800 30.330 127.250 ;
        RECT 19.130 126.650 22.980 126.800 ;
        RECT 26.480 126.650 30.330 126.800 ;
        RECT 19.130 126.200 19.430 126.650 ;
        RECT 30.030 126.200 30.330 126.650 ;
        RECT 19.130 126.050 22.980 126.200 ;
        RECT 26.480 126.050 30.330 126.200 ;
        RECT 19.130 125.600 19.430 126.050 ;
        RECT 30.030 125.600 30.330 126.050 ;
        RECT 19.130 125.450 22.980 125.600 ;
        RECT 26.480 125.450 30.330 125.600 ;
        RECT 19.130 125.000 19.430 125.450 ;
        RECT 30.030 125.000 30.330 125.450 ;
        RECT 19.130 124.850 22.980 125.000 ;
        RECT 26.480 124.850 30.330 125.000 ;
        RECT 19.130 124.400 19.430 124.850 ;
        RECT 30.030 124.400 30.330 124.850 ;
        RECT 19.130 124.250 22.980 124.400 ;
        RECT 26.480 124.250 30.330 124.400 ;
        RECT 19.130 123.800 19.430 124.250 ;
        RECT 30.030 123.800 30.330 124.250 ;
        RECT 19.130 123.650 22.980 123.800 ;
        RECT 26.480 123.650 30.330 123.800 ;
        RECT 19.130 123.200 19.430 123.650 ;
        RECT 30.030 123.200 30.330 123.650 ;
        RECT 19.130 123.050 22.980 123.200 ;
        RECT 26.480 123.050 30.330 123.200 ;
        RECT 19.130 122.600 19.430 123.050 ;
        RECT 30.030 122.600 30.330 123.050 ;
        RECT 19.130 122.450 22.980 122.600 ;
        RECT 26.480 122.450 30.330 122.600 ;
        RECT 19.130 122.000 19.430 122.450 ;
        RECT 30.030 122.000 30.330 122.450 ;
        RECT 19.130 121.450 22.930 122.000 ;
        RECT 6.530 121.400 22.930 121.450 ;
        RECT 26.530 121.450 30.330 122.000 ;
        RECT 30.780 121.450 30.930 129.650 ;
        RECT 31.380 121.450 31.530 129.650 ;
        RECT 31.980 121.450 32.130 129.650 ;
        RECT 32.580 121.450 32.730 129.650 ;
        RECT 33.180 121.450 33.330 129.650 ;
        RECT 33.780 121.450 33.930 129.650 ;
        RECT 34.380 121.450 35.080 138.550 ;
        RECT 35.530 130.350 35.680 138.550 ;
        RECT 36.130 130.350 36.280 138.550 ;
        RECT 36.730 130.350 36.880 138.550 ;
        RECT 37.330 130.350 37.480 138.550 ;
        RECT 37.930 130.350 38.080 138.550 ;
        RECT 38.530 130.350 38.680 138.550 ;
        RECT 39.130 138.000 42.930 138.550 ;
        RECT 46.530 138.550 62.930 138.600 ;
        RECT 46.530 138.000 50.330 138.550 ;
        RECT 39.130 137.550 39.430 138.000 ;
        RECT 50.030 137.550 50.330 138.000 ;
        RECT 39.130 137.400 42.980 137.550 ;
        RECT 46.480 137.400 50.330 137.550 ;
        RECT 39.130 136.950 39.430 137.400 ;
        RECT 50.030 136.950 50.330 137.400 ;
        RECT 39.130 136.800 42.980 136.950 ;
        RECT 46.480 136.800 50.330 136.950 ;
        RECT 39.130 136.350 39.430 136.800 ;
        RECT 50.030 136.350 50.330 136.800 ;
        RECT 39.130 136.200 42.980 136.350 ;
        RECT 46.480 136.200 50.330 136.350 ;
        RECT 39.130 135.750 39.430 136.200 ;
        RECT 50.030 135.750 50.330 136.200 ;
        RECT 39.130 135.600 42.980 135.750 ;
        RECT 46.480 135.600 50.330 135.750 ;
        RECT 39.130 135.150 39.430 135.600 ;
        RECT 50.030 135.150 50.330 135.600 ;
        RECT 39.130 135.000 42.980 135.150 ;
        RECT 46.480 135.000 50.330 135.150 ;
        RECT 39.130 134.550 39.430 135.000 ;
        RECT 50.030 134.550 50.330 135.000 ;
        RECT 39.130 134.400 42.980 134.550 ;
        RECT 46.480 134.400 50.330 134.550 ;
        RECT 39.130 133.950 39.430 134.400 ;
        RECT 50.030 133.950 50.330 134.400 ;
        RECT 39.130 133.800 42.980 133.950 ;
        RECT 46.480 133.800 50.330 133.950 ;
        RECT 39.130 133.350 39.430 133.800 ;
        RECT 50.030 133.350 50.330 133.800 ;
        RECT 39.130 133.200 42.980 133.350 ;
        RECT 46.480 133.200 50.330 133.350 ;
        RECT 39.130 132.750 39.430 133.200 ;
        RECT 39.130 132.600 42.980 132.750 ;
        RECT 39.130 132.150 39.430 132.600 ;
        RECT 39.130 132.000 42.980 132.150 ;
        RECT 39.130 131.550 39.430 132.000 ;
        RECT 39.130 131.400 42.980 131.550 ;
        RECT 39.130 130.950 39.430 131.400 ;
        RECT 39.130 130.800 42.980 130.950 ;
        RECT 39.130 130.350 39.430 130.800 ;
        RECT 35.530 121.450 35.680 129.650 ;
        RECT 36.130 121.450 36.280 129.650 ;
        RECT 36.730 121.450 36.880 129.650 ;
        RECT 37.330 121.450 37.480 129.650 ;
        RECT 37.930 121.450 38.080 129.650 ;
        RECT 38.530 121.450 38.680 129.650 ;
        RECT 39.130 129.200 39.430 129.650 ;
        RECT 39.130 129.050 42.980 129.200 ;
        RECT 39.130 128.600 39.430 129.050 ;
        RECT 39.130 128.450 42.980 128.600 ;
        RECT 39.130 128.000 39.430 128.450 ;
        RECT 39.130 127.850 42.980 128.000 ;
        RECT 39.130 127.400 39.430 127.850 ;
        RECT 39.130 127.250 42.980 127.400 ;
        RECT 39.130 126.800 39.430 127.250 ;
        RECT 43.830 126.800 45.630 133.200 ;
        RECT 50.030 132.750 50.330 133.200 ;
        RECT 46.480 132.600 50.330 132.750 ;
        RECT 50.030 132.150 50.330 132.600 ;
        RECT 46.480 132.000 50.330 132.150 ;
        RECT 50.030 131.550 50.330 132.000 ;
        RECT 46.480 131.400 50.330 131.550 ;
        RECT 50.030 130.950 50.330 131.400 ;
        RECT 46.480 130.800 50.330 130.950 ;
        RECT 50.030 130.350 50.330 130.800 ;
        RECT 50.780 130.350 50.930 138.550 ;
        RECT 51.380 130.350 51.530 138.550 ;
        RECT 51.980 130.350 52.130 138.550 ;
        RECT 52.580 130.350 52.730 138.550 ;
        RECT 53.180 130.350 53.330 138.550 ;
        RECT 53.780 130.350 53.930 138.550 ;
        RECT 50.030 129.200 50.330 129.650 ;
        RECT 46.480 129.050 50.330 129.200 ;
        RECT 50.030 128.600 50.330 129.050 ;
        RECT 46.480 128.450 50.330 128.600 ;
        RECT 50.030 128.000 50.330 128.450 ;
        RECT 46.480 127.850 50.330 128.000 ;
        RECT 50.030 127.400 50.330 127.850 ;
        RECT 46.480 127.250 50.330 127.400 ;
        RECT 50.030 126.800 50.330 127.250 ;
        RECT 39.130 126.650 42.980 126.800 ;
        RECT 46.480 126.650 50.330 126.800 ;
        RECT 39.130 126.200 39.430 126.650 ;
        RECT 50.030 126.200 50.330 126.650 ;
        RECT 39.130 126.050 42.980 126.200 ;
        RECT 46.480 126.050 50.330 126.200 ;
        RECT 39.130 125.600 39.430 126.050 ;
        RECT 50.030 125.600 50.330 126.050 ;
        RECT 39.130 125.450 42.980 125.600 ;
        RECT 46.480 125.450 50.330 125.600 ;
        RECT 39.130 125.000 39.430 125.450 ;
        RECT 50.030 125.000 50.330 125.450 ;
        RECT 39.130 124.850 42.980 125.000 ;
        RECT 46.480 124.850 50.330 125.000 ;
        RECT 39.130 124.400 39.430 124.850 ;
        RECT 50.030 124.400 50.330 124.850 ;
        RECT 39.130 124.250 42.980 124.400 ;
        RECT 46.480 124.250 50.330 124.400 ;
        RECT 39.130 123.800 39.430 124.250 ;
        RECT 50.030 123.800 50.330 124.250 ;
        RECT 39.130 123.650 42.980 123.800 ;
        RECT 46.480 123.650 50.330 123.800 ;
        RECT 39.130 123.200 39.430 123.650 ;
        RECT 50.030 123.200 50.330 123.650 ;
        RECT 39.130 123.050 42.980 123.200 ;
        RECT 46.480 123.050 50.330 123.200 ;
        RECT 39.130 122.600 39.430 123.050 ;
        RECT 50.030 122.600 50.330 123.050 ;
        RECT 39.130 122.450 42.980 122.600 ;
        RECT 46.480 122.450 50.330 122.600 ;
        RECT 39.130 122.000 39.430 122.450 ;
        RECT 50.030 122.000 50.330 122.450 ;
        RECT 39.130 121.450 42.930 122.000 ;
        RECT 26.530 121.400 42.930 121.450 ;
        RECT 46.530 121.450 50.330 122.000 ;
        RECT 50.780 121.450 50.930 129.650 ;
        RECT 51.380 121.450 51.530 129.650 ;
        RECT 51.980 121.450 52.130 129.650 ;
        RECT 52.580 121.450 52.730 129.650 ;
        RECT 53.180 121.450 53.330 129.650 ;
        RECT 53.780 121.450 53.930 129.650 ;
        RECT 54.380 121.450 55.080 138.550 ;
        RECT 55.530 130.350 55.680 138.550 ;
        RECT 56.130 130.350 56.280 138.550 ;
        RECT 56.730 130.350 56.880 138.550 ;
        RECT 57.330 130.350 57.480 138.550 ;
        RECT 57.930 130.350 58.080 138.550 ;
        RECT 58.530 130.350 58.680 138.550 ;
        RECT 59.130 138.000 62.930 138.550 ;
        RECT 66.530 138.550 82.930 138.600 ;
        RECT 66.530 138.000 70.330 138.550 ;
        RECT 59.130 137.550 59.430 138.000 ;
        RECT 70.030 137.550 70.330 138.000 ;
        RECT 59.130 137.400 62.980 137.550 ;
        RECT 66.480 137.400 70.330 137.550 ;
        RECT 59.130 136.950 59.430 137.400 ;
        RECT 70.030 136.950 70.330 137.400 ;
        RECT 59.130 136.800 62.980 136.950 ;
        RECT 66.480 136.800 70.330 136.950 ;
        RECT 59.130 136.350 59.430 136.800 ;
        RECT 70.030 136.350 70.330 136.800 ;
        RECT 59.130 136.200 62.980 136.350 ;
        RECT 66.480 136.200 70.330 136.350 ;
        RECT 59.130 135.750 59.430 136.200 ;
        RECT 70.030 135.750 70.330 136.200 ;
        RECT 59.130 135.600 62.980 135.750 ;
        RECT 66.480 135.600 70.330 135.750 ;
        RECT 59.130 135.150 59.430 135.600 ;
        RECT 70.030 135.150 70.330 135.600 ;
        RECT 59.130 135.000 62.980 135.150 ;
        RECT 66.480 135.000 70.330 135.150 ;
        RECT 59.130 134.550 59.430 135.000 ;
        RECT 70.030 134.550 70.330 135.000 ;
        RECT 59.130 134.400 62.980 134.550 ;
        RECT 66.480 134.400 70.330 134.550 ;
        RECT 59.130 133.950 59.430 134.400 ;
        RECT 70.030 133.950 70.330 134.400 ;
        RECT 59.130 133.800 62.980 133.950 ;
        RECT 66.480 133.800 70.330 133.950 ;
        RECT 59.130 133.350 59.430 133.800 ;
        RECT 70.030 133.350 70.330 133.800 ;
        RECT 59.130 133.200 62.980 133.350 ;
        RECT 66.480 133.200 70.330 133.350 ;
        RECT 59.130 132.750 59.430 133.200 ;
        RECT 59.130 132.600 62.980 132.750 ;
        RECT 59.130 132.150 59.430 132.600 ;
        RECT 59.130 132.000 62.980 132.150 ;
        RECT 59.130 131.550 59.430 132.000 ;
        RECT 59.130 131.400 62.980 131.550 ;
        RECT 59.130 130.950 59.430 131.400 ;
        RECT 59.130 130.800 62.980 130.950 ;
        RECT 59.130 130.350 59.430 130.800 ;
        RECT 55.530 121.450 55.680 129.650 ;
        RECT 56.130 121.450 56.280 129.650 ;
        RECT 56.730 121.450 56.880 129.650 ;
        RECT 57.330 121.450 57.480 129.650 ;
        RECT 57.930 121.450 58.080 129.650 ;
        RECT 58.530 121.450 58.680 129.650 ;
        RECT 59.130 129.200 59.430 129.650 ;
        RECT 59.130 129.050 62.980 129.200 ;
        RECT 59.130 128.600 59.430 129.050 ;
        RECT 59.130 128.450 62.980 128.600 ;
        RECT 59.130 128.000 59.430 128.450 ;
        RECT 59.130 127.850 62.980 128.000 ;
        RECT 59.130 127.400 59.430 127.850 ;
        RECT 59.130 127.250 62.980 127.400 ;
        RECT 59.130 126.800 59.430 127.250 ;
        RECT 63.830 126.800 65.630 133.200 ;
        RECT 70.030 132.750 70.330 133.200 ;
        RECT 66.480 132.600 70.330 132.750 ;
        RECT 70.030 132.150 70.330 132.600 ;
        RECT 66.480 132.000 70.330 132.150 ;
        RECT 70.030 131.550 70.330 132.000 ;
        RECT 66.480 131.400 70.330 131.550 ;
        RECT 70.030 130.950 70.330 131.400 ;
        RECT 66.480 130.800 70.330 130.950 ;
        RECT 70.030 130.350 70.330 130.800 ;
        RECT 70.780 130.350 70.930 138.550 ;
        RECT 71.380 130.350 71.530 138.550 ;
        RECT 71.980 130.350 72.130 138.550 ;
        RECT 72.580 130.350 72.730 138.550 ;
        RECT 73.180 130.350 73.330 138.550 ;
        RECT 73.780 130.350 73.930 138.550 ;
        RECT 70.030 129.200 70.330 129.650 ;
        RECT 66.480 129.050 70.330 129.200 ;
        RECT 70.030 128.600 70.330 129.050 ;
        RECT 66.480 128.450 70.330 128.600 ;
        RECT 70.030 128.000 70.330 128.450 ;
        RECT 66.480 127.850 70.330 128.000 ;
        RECT 70.030 127.400 70.330 127.850 ;
        RECT 66.480 127.250 70.330 127.400 ;
        RECT 70.030 126.800 70.330 127.250 ;
        RECT 59.130 126.650 62.980 126.800 ;
        RECT 66.480 126.650 70.330 126.800 ;
        RECT 59.130 126.200 59.430 126.650 ;
        RECT 70.030 126.200 70.330 126.650 ;
        RECT 59.130 126.050 62.980 126.200 ;
        RECT 66.480 126.050 70.330 126.200 ;
        RECT 59.130 125.600 59.430 126.050 ;
        RECT 70.030 125.600 70.330 126.050 ;
        RECT 59.130 125.450 62.980 125.600 ;
        RECT 66.480 125.450 70.330 125.600 ;
        RECT 59.130 125.000 59.430 125.450 ;
        RECT 70.030 125.000 70.330 125.450 ;
        RECT 59.130 124.850 62.980 125.000 ;
        RECT 66.480 124.850 70.330 125.000 ;
        RECT 59.130 124.400 59.430 124.850 ;
        RECT 70.030 124.400 70.330 124.850 ;
        RECT 59.130 124.250 62.980 124.400 ;
        RECT 66.480 124.250 70.330 124.400 ;
        RECT 59.130 123.800 59.430 124.250 ;
        RECT 70.030 123.800 70.330 124.250 ;
        RECT 59.130 123.650 62.980 123.800 ;
        RECT 66.480 123.650 70.330 123.800 ;
        RECT 59.130 123.200 59.430 123.650 ;
        RECT 70.030 123.200 70.330 123.650 ;
        RECT 59.130 123.050 62.980 123.200 ;
        RECT 66.480 123.050 70.330 123.200 ;
        RECT 59.130 122.600 59.430 123.050 ;
        RECT 70.030 122.600 70.330 123.050 ;
        RECT 59.130 122.450 62.980 122.600 ;
        RECT 66.480 122.450 70.330 122.600 ;
        RECT 59.130 122.000 59.430 122.450 ;
        RECT 70.030 122.000 70.330 122.450 ;
        RECT 59.130 121.450 62.930 122.000 ;
        RECT 46.530 121.400 62.930 121.450 ;
        RECT 66.530 121.450 70.330 122.000 ;
        RECT 70.780 121.450 70.930 129.650 ;
        RECT 71.380 121.450 71.530 129.650 ;
        RECT 71.980 121.450 72.130 129.650 ;
        RECT 72.580 121.450 72.730 129.650 ;
        RECT 73.180 121.450 73.330 129.650 ;
        RECT 73.780 121.450 73.930 129.650 ;
        RECT 74.380 121.450 75.080 138.550 ;
        RECT 75.530 130.350 75.680 138.550 ;
        RECT 76.130 130.350 76.280 138.550 ;
        RECT 76.730 130.350 76.880 138.550 ;
        RECT 77.330 130.350 77.480 138.550 ;
        RECT 77.930 130.350 78.080 138.550 ;
        RECT 78.530 130.350 78.680 138.550 ;
        RECT 79.130 138.000 82.930 138.550 ;
        RECT 86.530 138.550 102.930 138.600 ;
        RECT 86.530 138.000 90.330 138.550 ;
        RECT 79.130 137.550 79.430 138.000 ;
        RECT 90.030 137.550 90.330 138.000 ;
        RECT 79.130 137.400 82.980 137.550 ;
        RECT 86.480 137.400 90.330 137.550 ;
        RECT 79.130 136.950 79.430 137.400 ;
        RECT 90.030 136.950 90.330 137.400 ;
        RECT 79.130 136.800 82.980 136.950 ;
        RECT 86.480 136.800 90.330 136.950 ;
        RECT 79.130 136.350 79.430 136.800 ;
        RECT 90.030 136.350 90.330 136.800 ;
        RECT 79.130 136.200 82.980 136.350 ;
        RECT 86.480 136.200 90.330 136.350 ;
        RECT 79.130 135.750 79.430 136.200 ;
        RECT 90.030 135.750 90.330 136.200 ;
        RECT 79.130 135.600 82.980 135.750 ;
        RECT 86.480 135.600 90.330 135.750 ;
        RECT 79.130 135.150 79.430 135.600 ;
        RECT 90.030 135.150 90.330 135.600 ;
        RECT 79.130 135.000 82.980 135.150 ;
        RECT 86.480 135.000 90.330 135.150 ;
        RECT 79.130 134.550 79.430 135.000 ;
        RECT 90.030 134.550 90.330 135.000 ;
        RECT 79.130 134.400 82.980 134.550 ;
        RECT 86.480 134.400 90.330 134.550 ;
        RECT 79.130 133.950 79.430 134.400 ;
        RECT 90.030 133.950 90.330 134.400 ;
        RECT 79.130 133.800 82.980 133.950 ;
        RECT 86.480 133.800 90.330 133.950 ;
        RECT 79.130 133.350 79.430 133.800 ;
        RECT 90.030 133.350 90.330 133.800 ;
        RECT 79.130 133.200 82.980 133.350 ;
        RECT 86.480 133.200 90.330 133.350 ;
        RECT 79.130 132.750 79.430 133.200 ;
        RECT 79.130 132.600 82.980 132.750 ;
        RECT 79.130 132.150 79.430 132.600 ;
        RECT 79.130 132.000 82.980 132.150 ;
        RECT 79.130 131.550 79.430 132.000 ;
        RECT 79.130 131.400 82.980 131.550 ;
        RECT 79.130 130.950 79.430 131.400 ;
        RECT 79.130 130.800 82.980 130.950 ;
        RECT 79.130 130.350 79.430 130.800 ;
        RECT 75.530 121.450 75.680 129.650 ;
        RECT 76.130 121.450 76.280 129.650 ;
        RECT 76.730 121.450 76.880 129.650 ;
        RECT 77.330 121.450 77.480 129.650 ;
        RECT 77.930 121.450 78.080 129.650 ;
        RECT 78.530 121.450 78.680 129.650 ;
        RECT 79.130 129.200 79.430 129.650 ;
        RECT 79.130 129.050 82.980 129.200 ;
        RECT 79.130 128.600 79.430 129.050 ;
        RECT 79.130 128.450 82.980 128.600 ;
        RECT 79.130 128.000 79.430 128.450 ;
        RECT 79.130 127.850 82.980 128.000 ;
        RECT 79.130 127.400 79.430 127.850 ;
        RECT 79.130 127.250 82.980 127.400 ;
        RECT 79.130 126.800 79.430 127.250 ;
        RECT 83.830 126.800 85.630 133.200 ;
        RECT 90.030 132.750 90.330 133.200 ;
        RECT 86.480 132.600 90.330 132.750 ;
        RECT 90.030 132.150 90.330 132.600 ;
        RECT 86.480 132.000 90.330 132.150 ;
        RECT 90.030 131.550 90.330 132.000 ;
        RECT 86.480 131.400 90.330 131.550 ;
        RECT 90.030 130.950 90.330 131.400 ;
        RECT 86.480 130.800 90.330 130.950 ;
        RECT 90.030 130.350 90.330 130.800 ;
        RECT 90.780 130.350 90.930 138.550 ;
        RECT 91.380 130.350 91.530 138.550 ;
        RECT 91.980 130.350 92.130 138.550 ;
        RECT 92.580 130.350 92.730 138.550 ;
        RECT 93.180 130.350 93.330 138.550 ;
        RECT 93.780 130.350 93.930 138.550 ;
        RECT 90.030 129.200 90.330 129.650 ;
        RECT 86.480 129.050 90.330 129.200 ;
        RECT 90.030 128.600 90.330 129.050 ;
        RECT 86.480 128.450 90.330 128.600 ;
        RECT 90.030 128.000 90.330 128.450 ;
        RECT 86.480 127.850 90.330 128.000 ;
        RECT 90.030 127.400 90.330 127.850 ;
        RECT 86.480 127.250 90.330 127.400 ;
        RECT 90.030 126.800 90.330 127.250 ;
        RECT 79.130 126.650 82.980 126.800 ;
        RECT 86.480 126.650 90.330 126.800 ;
        RECT 79.130 126.200 79.430 126.650 ;
        RECT 90.030 126.200 90.330 126.650 ;
        RECT 79.130 126.050 82.980 126.200 ;
        RECT 86.480 126.050 90.330 126.200 ;
        RECT 79.130 125.600 79.430 126.050 ;
        RECT 90.030 125.600 90.330 126.050 ;
        RECT 79.130 125.450 82.980 125.600 ;
        RECT 86.480 125.450 90.330 125.600 ;
        RECT 79.130 125.000 79.430 125.450 ;
        RECT 90.030 125.000 90.330 125.450 ;
        RECT 79.130 124.850 82.980 125.000 ;
        RECT 86.480 124.850 90.330 125.000 ;
        RECT 79.130 124.400 79.430 124.850 ;
        RECT 90.030 124.400 90.330 124.850 ;
        RECT 79.130 124.250 82.980 124.400 ;
        RECT 86.480 124.250 90.330 124.400 ;
        RECT 79.130 123.800 79.430 124.250 ;
        RECT 90.030 123.800 90.330 124.250 ;
        RECT 79.130 123.650 82.980 123.800 ;
        RECT 86.480 123.650 90.330 123.800 ;
        RECT 79.130 123.200 79.430 123.650 ;
        RECT 90.030 123.200 90.330 123.650 ;
        RECT 79.130 123.050 82.980 123.200 ;
        RECT 86.480 123.050 90.330 123.200 ;
        RECT 79.130 122.600 79.430 123.050 ;
        RECT 90.030 122.600 90.330 123.050 ;
        RECT 79.130 122.450 82.980 122.600 ;
        RECT 86.480 122.450 90.330 122.600 ;
        RECT 79.130 122.000 79.430 122.450 ;
        RECT 90.030 122.000 90.330 122.450 ;
        RECT 79.130 121.450 82.930 122.000 ;
        RECT 66.530 121.400 82.930 121.450 ;
        RECT 86.530 121.450 90.330 122.000 ;
        RECT 90.780 121.450 90.930 129.650 ;
        RECT 91.380 121.450 91.530 129.650 ;
        RECT 91.980 121.450 92.130 129.650 ;
        RECT 92.580 121.450 92.730 129.650 ;
        RECT 93.180 121.450 93.330 129.650 ;
        RECT 93.780 121.450 93.930 129.650 ;
        RECT 94.380 121.450 95.080 138.550 ;
        RECT 95.530 130.350 95.680 138.550 ;
        RECT 96.130 130.350 96.280 138.550 ;
        RECT 96.730 130.350 96.880 138.550 ;
        RECT 97.330 130.350 97.480 138.550 ;
        RECT 97.930 130.350 98.080 138.550 ;
        RECT 98.530 130.350 98.680 138.550 ;
        RECT 99.130 138.000 102.930 138.550 ;
        RECT 106.530 138.550 122.930 138.600 ;
        RECT 106.530 138.000 110.330 138.550 ;
        RECT 99.130 137.550 99.430 138.000 ;
        RECT 110.030 137.550 110.330 138.000 ;
        RECT 99.130 137.400 102.980 137.550 ;
        RECT 106.480 137.400 110.330 137.550 ;
        RECT 99.130 136.950 99.430 137.400 ;
        RECT 110.030 136.950 110.330 137.400 ;
        RECT 99.130 136.800 102.980 136.950 ;
        RECT 106.480 136.800 110.330 136.950 ;
        RECT 99.130 136.350 99.430 136.800 ;
        RECT 110.030 136.350 110.330 136.800 ;
        RECT 99.130 136.200 102.980 136.350 ;
        RECT 106.480 136.200 110.330 136.350 ;
        RECT 99.130 135.750 99.430 136.200 ;
        RECT 110.030 135.750 110.330 136.200 ;
        RECT 99.130 135.600 102.980 135.750 ;
        RECT 106.480 135.600 110.330 135.750 ;
        RECT 99.130 135.150 99.430 135.600 ;
        RECT 110.030 135.150 110.330 135.600 ;
        RECT 99.130 135.000 102.980 135.150 ;
        RECT 106.480 135.000 110.330 135.150 ;
        RECT 99.130 134.550 99.430 135.000 ;
        RECT 110.030 134.550 110.330 135.000 ;
        RECT 99.130 134.400 102.980 134.550 ;
        RECT 106.480 134.400 110.330 134.550 ;
        RECT 99.130 133.950 99.430 134.400 ;
        RECT 110.030 133.950 110.330 134.400 ;
        RECT 99.130 133.800 102.980 133.950 ;
        RECT 106.480 133.800 110.330 133.950 ;
        RECT 99.130 133.350 99.430 133.800 ;
        RECT 110.030 133.350 110.330 133.800 ;
        RECT 99.130 133.200 102.980 133.350 ;
        RECT 106.480 133.200 110.330 133.350 ;
        RECT 99.130 132.750 99.430 133.200 ;
        RECT 99.130 132.600 102.980 132.750 ;
        RECT 99.130 132.150 99.430 132.600 ;
        RECT 99.130 132.000 102.980 132.150 ;
        RECT 99.130 131.550 99.430 132.000 ;
        RECT 99.130 131.400 102.980 131.550 ;
        RECT 99.130 130.950 99.430 131.400 ;
        RECT 99.130 130.800 102.980 130.950 ;
        RECT 99.130 130.350 99.430 130.800 ;
        RECT 95.530 121.450 95.680 129.650 ;
        RECT 96.130 121.450 96.280 129.650 ;
        RECT 96.730 121.450 96.880 129.650 ;
        RECT 97.330 121.450 97.480 129.650 ;
        RECT 97.930 121.450 98.080 129.650 ;
        RECT 98.530 121.450 98.680 129.650 ;
        RECT 99.130 129.200 99.430 129.650 ;
        RECT 99.130 129.050 102.980 129.200 ;
        RECT 99.130 128.600 99.430 129.050 ;
        RECT 99.130 128.450 102.980 128.600 ;
        RECT 99.130 128.000 99.430 128.450 ;
        RECT 99.130 127.850 102.980 128.000 ;
        RECT 99.130 127.400 99.430 127.850 ;
        RECT 99.130 127.250 102.980 127.400 ;
        RECT 99.130 126.800 99.430 127.250 ;
        RECT 103.830 126.800 105.630 133.200 ;
        RECT 110.030 132.750 110.330 133.200 ;
        RECT 106.480 132.600 110.330 132.750 ;
        RECT 110.030 132.150 110.330 132.600 ;
        RECT 106.480 132.000 110.330 132.150 ;
        RECT 110.030 131.550 110.330 132.000 ;
        RECT 106.480 131.400 110.330 131.550 ;
        RECT 110.030 130.950 110.330 131.400 ;
        RECT 106.480 130.800 110.330 130.950 ;
        RECT 110.030 130.350 110.330 130.800 ;
        RECT 110.780 130.350 110.930 138.550 ;
        RECT 111.380 130.350 111.530 138.550 ;
        RECT 111.980 130.350 112.130 138.550 ;
        RECT 112.580 130.350 112.730 138.550 ;
        RECT 113.180 130.350 113.330 138.550 ;
        RECT 113.780 130.350 113.930 138.550 ;
        RECT 110.030 129.200 110.330 129.650 ;
        RECT 106.480 129.050 110.330 129.200 ;
        RECT 110.030 128.600 110.330 129.050 ;
        RECT 106.480 128.450 110.330 128.600 ;
        RECT 110.030 128.000 110.330 128.450 ;
        RECT 106.480 127.850 110.330 128.000 ;
        RECT 110.030 127.400 110.330 127.850 ;
        RECT 106.480 127.250 110.330 127.400 ;
        RECT 110.030 126.800 110.330 127.250 ;
        RECT 99.130 126.650 102.980 126.800 ;
        RECT 106.480 126.650 110.330 126.800 ;
        RECT 99.130 126.200 99.430 126.650 ;
        RECT 110.030 126.200 110.330 126.650 ;
        RECT 99.130 126.050 102.980 126.200 ;
        RECT 106.480 126.050 110.330 126.200 ;
        RECT 99.130 125.600 99.430 126.050 ;
        RECT 110.030 125.600 110.330 126.050 ;
        RECT 99.130 125.450 102.980 125.600 ;
        RECT 106.480 125.450 110.330 125.600 ;
        RECT 99.130 125.000 99.430 125.450 ;
        RECT 110.030 125.000 110.330 125.450 ;
        RECT 99.130 124.850 102.980 125.000 ;
        RECT 106.480 124.850 110.330 125.000 ;
        RECT 99.130 124.400 99.430 124.850 ;
        RECT 110.030 124.400 110.330 124.850 ;
        RECT 99.130 124.250 102.980 124.400 ;
        RECT 106.480 124.250 110.330 124.400 ;
        RECT 99.130 123.800 99.430 124.250 ;
        RECT 110.030 123.800 110.330 124.250 ;
        RECT 99.130 123.650 102.980 123.800 ;
        RECT 106.480 123.650 110.330 123.800 ;
        RECT 99.130 123.200 99.430 123.650 ;
        RECT 110.030 123.200 110.330 123.650 ;
        RECT 99.130 123.050 102.980 123.200 ;
        RECT 106.480 123.050 110.330 123.200 ;
        RECT 99.130 122.600 99.430 123.050 ;
        RECT 110.030 122.600 110.330 123.050 ;
        RECT 99.130 122.450 102.980 122.600 ;
        RECT 106.480 122.450 110.330 122.600 ;
        RECT 99.130 122.000 99.430 122.450 ;
        RECT 110.030 122.000 110.330 122.450 ;
        RECT 99.130 121.450 102.930 122.000 ;
        RECT 86.530 121.400 102.930 121.450 ;
        RECT 106.530 121.450 110.330 122.000 ;
        RECT 110.780 121.450 110.930 129.650 ;
        RECT 111.380 121.450 111.530 129.650 ;
        RECT 111.980 121.450 112.130 129.650 ;
        RECT 112.580 121.450 112.730 129.650 ;
        RECT 113.180 121.450 113.330 129.650 ;
        RECT 113.780 121.450 113.930 129.650 ;
        RECT 114.380 121.450 115.080 138.550 ;
        RECT 115.530 130.350 115.680 138.550 ;
        RECT 116.130 130.350 116.280 138.550 ;
        RECT 116.730 130.350 116.880 138.550 ;
        RECT 117.330 130.350 117.480 138.550 ;
        RECT 117.930 130.350 118.080 138.550 ;
        RECT 118.530 130.350 118.680 138.550 ;
        RECT 119.130 138.000 122.930 138.550 ;
        RECT 119.130 137.550 119.430 138.000 ;
        RECT 119.130 137.400 122.980 137.550 ;
        RECT 119.130 136.950 119.430 137.400 ;
        RECT 119.130 136.800 122.980 136.950 ;
        RECT 119.130 136.350 119.430 136.800 ;
        RECT 119.130 136.200 122.980 136.350 ;
        RECT 119.130 135.750 119.430 136.200 ;
        RECT 119.130 135.600 122.980 135.750 ;
        RECT 119.130 135.150 119.430 135.600 ;
        RECT 119.130 135.000 122.980 135.150 ;
        RECT 119.130 134.550 119.430 135.000 ;
        RECT 119.130 134.400 122.980 134.550 ;
        RECT 119.130 133.950 119.430 134.400 ;
        RECT 119.130 133.800 122.980 133.950 ;
        RECT 119.130 133.350 119.430 133.800 ;
        RECT 119.130 133.200 122.980 133.350 ;
        RECT 119.130 132.750 119.430 133.200 ;
        RECT 119.130 132.600 122.980 132.750 ;
        RECT 119.130 132.150 119.430 132.600 ;
        RECT 119.130 132.000 122.980 132.150 ;
        RECT 119.130 131.550 119.430 132.000 ;
        RECT 119.130 131.400 122.980 131.550 ;
        RECT 119.130 130.950 119.430 131.400 ;
        RECT 119.130 130.800 122.980 130.950 ;
        RECT 119.130 130.350 119.430 130.800 ;
        RECT 115.530 121.450 115.680 129.650 ;
        RECT 116.130 121.450 116.280 129.650 ;
        RECT 116.730 121.450 116.880 129.650 ;
        RECT 117.330 121.450 117.480 129.650 ;
        RECT 117.930 121.450 118.080 129.650 ;
        RECT 118.530 121.450 118.680 129.650 ;
        RECT 119.130 129.200 119.430 129.650 ;
        RECT 119.130 129.050 122.980 129.200 ;
        RECT 119.130 128.600 119.430 129.050 ;
        RECT 119.130 128.450 122.980 128.600 ;
        RECT 119.130 128.000 119.430 128.450 ;
        RECT 119.130 127.850 122.980 128.000 ;
        RECT 119.130 127.400 119.430 127.850 ;
        RECT 119.130 127.250 122.980 127.400 ;
        RECT 119.130 126.800 119.430 127.250 ;
        RECT 123.830 126.800 124.730 133.200 ;
        RECT 129.850 129.500 131.850 130.775 ;
        RECT 119.130 126.650 122.980 126.800 ;
        RECT 119.130 126.200 119.430 126.650 ;
        RECT 119.130 126.050 122.980 126.200 ;
        RECT 119.130 125.600 119.430 126.050 ;
        RECT 119.130 125.450 122.980 125.600 ;
        RECT 119.130 125.000 119.430 125.450 ;
        RECT 119.130 124.850 122.980 125.000 ;
        RECT 119.130 124.400 119.430 124.850 ;
        RECT 119.130 124.250 122.980 124.400 ;
        RECT 119.130 123.800 119.430 124.250 ;
        RECT 119.130 123.650 122.980 123.800 ;
        RECT 119.130 123.200 119.430 123.650 ;
        RECT 119.130 123.050 122.980 123.200 ;
        RECT 119.130 122.600 119.430 123.050 ;
        RECT 119.130 122.450 122.980 122.600 ;
        RECT 119.130 122.000 119.430 122.450 ;
        RECT 119.130 121.450 122.930 122.000 ;
        RECT 106.530 121.400 122.930 121.450 ;
        RECT 9.630 120.900 19.830 121.400 ;
        RECT 29.630 120.900 39.830 121.400 ;
        RECT 49.630 120.900 59.830 121.400 ;
        RECT 69.630 120.900 79.830 121.400 ;
        RECT 89.630 120.900 99.830 121.400 ;
        RECT 109.630 120.900 119.830 121.400 ;
        RECT 11.530 119.100 17.930 120.900 ;
        RECT 31.530 119.100 37.930 120.900 ;
        RECT 51.530 119.100 57.930 120.900 ;
        RECT 71.530 119.100 77.930 120.900 ;
        RECT 91.530 119.100 97.930 120.900 ;
        RECT 111.530 119.100 117.930 120.900 ;
        RECT 9.630 118.600 19.830 119.100 ;
        RECT 29.630 118.600 39.830 119.100 ;
        RECT 49.630 118.600 59.830 119.100 ;
        RECT 69.630 118.600 79.830 119.100 ;
        RECT 89.630 118.600 99.830 119.100 ;
        RECT 109.630 118.600 119.830 119.100 ;
        RECT 6.530 118.550 22.930 118.600 ;
        RECT 6.530 118.000 10.330 118.550 ;
        RECT 10.030 117.550 10.330 118.000 ;
        RECT 6.480 117.400 10.330 117.550 ;
        RECT 10.030 116.950 10.330 117.400 ;
        RECT 6.480 116.800 10.330 116.950 ;
        RECT 10.030 116.350 10.330 116.800 ;
        RECT 6.480 116.200 10.330 116.350 ;
        RECT 10.030 115.750 10.330 116.200 ;
        RECT 6.480 115.600 10.330 115.750 ;
        RECT 10.030 115.150 10.330 115.600 ;
        RECT 6.480 115.000 10.330 115.150 ;
        RECT 10.030 114.550 10.330 115.000 ;
        RECT 6.480 114.400 10.330 114.550 ;
        RECT 10.030 113.950 10.330 114.400 ;
        RECT 6.480 113.800 10.330 113.950 ;
        RECT 10.030 113.350 10.330 113.800 ;
        RECT 6.480 113.200 10.330 113.350 ;
        RECT 4.730 106.800 5.630 113.200 ;
        RECT 10.030 112.750 10.330 113.200 ;
        RECT 6.480 112.600 10.330 112.750 ;
        RECT 10.030 112.150 10.330 112.600 ;
        RECT 6.480 112.000 10.330 112.150 ;
        RECT 10.030 111.550 10.330 112.000 ;
        RECT 6.480 111.400 10.330 111.550 ;
        RECT 10.030 110.950 10.330 111.400 ;
        RECT 6.480 110.800 10.330 110.950 ;
        RECT 10.030 110.350 10.330 110.800 ;
        RECT 10.780 110.350 10.930 118.550 ;
        RECT 11.380 110.350 11.530 118.550 ;
        RECT 11.980 110.350 12.130 118.550 ;
        RECT 12.580 110.350 12.730 118.550 ;
        RECT 13.180 110.350 13.330 118.550 ;
        RECT 13.780 110.350 13.930 118.550 ;
        RECT 10.030 109.200 10.330 109.650 ;
        RECT 6.480 109.050 10.330 109.200 ;
        RECT 10.030 108.600 10.330 109.050 ;
        RECT 6.480 108.450 10.330 108.600 ;
        RECT 10.030 108.000 10.330 108.450 ;
        RECT 6.480 107.850 10.330 108.000 ;
        RECT 10.030 107.400 10.330 107.850 ;
        RECT 6.480 107.250 10.330 107.400 ;
        RECT 10.030 106.800 10.330 107.250 ;
        RECT 6.480 106.650 10.330 106.800 ;
        RECT 10.030 106.200 10.330 106.650 ;
        RECT 6.480 106.050 10.330 106.200 ;
        RECT 10.030 105.600 10.330 106.050 ;
        RECT 6.480 105.450 10.330 105.600 ;
        RECT 10.030 105.000 10.330 105.450 ;
        RECT 6.480 104.850 10.330 105.000 ;
        RECT 10.030 104.400 10.330 104.850 ;
        RECT 6.480 104.250 10.330 104.400 ;
        RECT 10.030 103.800 10.330 104.250 ;
        RECT 6.480 103.650 10.330 103.800 ;
        RECT 10.030 103.200 10.330 103.650 ;
        RECT 6.480 103.050 10.330 103.200 ;
        RECT 10.030 102.600 10.330 103.050 ;
        RECT 6.480 102.450 10.330 102.600 ;
        RECT 10.030 102.000 10.330 102.450 ;
        RECT 6.530 101.450 10.330 102.000 ;
        RECT 10.780 101.450 10.930 109.650 ;
        RECT 11.380 101.450 11.530 109.650 ;
        RECT 11.980 101.450 12.130 109.650 ;
        RECT 12.580 101.450 12.730 109.650 ;
        RECT 13.180 101.450 13.330 109.650 ;
        RECT 13.780 101.450 13.930 109.650 ;
        RECT 14.380 101.450 15.080 118.550 ;
        RECT 15.530 110.350 15.680 118.550 ;
        RECT 16.130 110.350 16.280 118.550 ;
        RECT 16.730 110.350 16.880 118.550 ;
        RECT 17.330 110.350 17.480 118.550 ;
        RECT 17.930 110.350 18.080 118.550 ;
        RECT 18.530 110.350 18.680 118.550 ;
        RECT 19.130 118.000 22.930 118.550 ;
        RECT 26.530 118.550 42.930 118.600 ;
        RECT 26.530 118.000 30.330 118.550 ;
        RECT 19.130 117.550 19.430 118.000 ;
        RECT 30.030 117.550 30.330 118.000 ;
        RECT 19.130 117.400 22.980 117.550 ;
        RECT 26.480 117.400 30.330 117.550 ;
        RECT 19.130 116.950 19.430 117.400 ;
        RECT 30.030 116.950 30.330 117.400 ;
        RECT 19.130 116.800 22.980 116.950 ;
        RECT 26.480 116.800 30.330 116.950 ;
        RECT 19.130 116.350 19.430 116.800 ;
        RECT 30.030 116.350 30.330 116.800 ;
        RECT 19.130 116.200 22.980 116.350 ;
        RECT 26.480 116.200 30.330 116.350 ;
        RECT 19.130 115.750 19.430 116.200 ;
        RECT 30.030 115.750 30.330 116.200 ;
        RECT 19.130 115.600 22.980 115.750 ;
        RECT 26.480 115.600 30.330 115.750 ;
        RECT 19.130 115.150 19.430 115.600 ;
        RECT 30.030 115.150 30.330 115.600 ;
        RECT 19.130 115.000 22.980 115.150 ;
        RECT 26.480 115.000 30.330 115.150 ;
        RECT 19.130 114.550 19.430 115.000 ;
        RECT 30.030 114.550 30.330 115.000 ;
        RECT 19.130 114.400 22.980 114.550 ;
        RECT 26.480 114.400 30.330 114.550 ;
        RECT 19.130 113.950 19.430 114.400 ;
        RECT 30.030 113.950 30.330 114.400 ;
        RECT 19.130 113.800 22.980 113.950 ;
        RECT 26.480 113.800 30.330 113.950 ;
        RECT 19.130 113.350 19.430 113.800 ;
        RECT 30.030 113.350 30.330 113.800 ;
        RECT 19.130 113.200 22.980 113.350 ;
        RECT 26.480 113.200 30.330 113.350 ;
        RECT 19.130 112.750 19.430 113.200 ;
        RECT 19.130 112.600 22.980 112.750 ;
        RECT 19.130 112.150 19.430 112.600 ;
        RECT 19.130 112.000 22.980 112.150 ;
        RECT 19.130 111.550 19.430 112.000 ;
        RECT 19.130 111.400 22.980 111.550 ;
        RECT 19.130 110.950 19.430 111.400 ;
        RECT 19.130 110.800 22.980 110.950 ;
        RECT 19.130 110.350 19.430 110.800 ;
        RECT 15.530 101.450 15.680 109.650 ;
        RECT 16.130 101.450 16.280 109.650 ;
        RECT 16.730 101.450 16.880 109.650 ;
        RECT 17.330 101.450 17.480 109.650 ;
        RECT 17.930 101.450 18.080 109.650 ;
        RECT 18.530 101.450 18.680 109.650 ;
        RECT 19.130 109.200 19.430 109.650 ;
        RECT 19.130 109.050 22.980 109.200 ;
        RECT 19.130 108.600 19.430 109.050 ;
        RECT 19.130 108.450 22.980 108.600 ;
        RECT 19.130 108.000 19.430 108.450 ;
        RECT 19.130 107.850 22.980 108.000 ;
        RECT 19.130 107.400 19.430 107.850 ;
        RECT 19.130 107.250 22.980 107.400 ;
        RECT 19.130 106.800 19.430 107.250 ;
        RECT 23.830 106.800 25.630 113.200 ;
        RECT 30.030 112.750 30.330 113.200 ;
        RECT 26.480 112.600 30.330 112.750 ;
        RECT 30.030 112.150 30.330 112.600 ;
        RECT 26.480 112.000 30.330 112.150 ;
        RECT 30.030 111.550 30.330 112.000 ;
        RECT 26.480 111.400 30.330 111.550 ;
        RECT 30.030 110.950 30.330 111.400 ;
        RECT 26.480 110.800 30.330 110.950 ;
        RECT 30.030 110.350 30.330 110.800 ;
        RECT 30.780 110.350 30.930 118.550 ;
        RECT 31.380 110.350 31.530 118.550 ;
        RECT 31.980 110.350 32.130 118.550 ;
        RECT 32.580 110.350 32.730 118.550 ;
        RECT 33.180 110.350 33.330 118.550 ;
        RECT 33.780 110.350 33.930 118.550 ;
        RECT 30.030 109.200 30.330 109.650 ;
        RECT 26.480 109.050 30.330 109.200 ;
        RECT 30.030 108.600 30.330 109.050 ;
        RECT 26.480 108.450 30.330 108.600 ;
        RECT 30.030 108.000 30.330 108.450 ;
        RECT 26.480 107.850 30.330 108.000 ;
        RECT 30.030 107.400 30.330 107.850 ;
        RECT 26.480 107.250 30.330 107.400 ;
        RECT 30.030 106.800 30.330 107.250 ;
        RECT 19.130 106.650 22.980 106.800 ;
        RECT 26.480 106.650 30.330 106.800 ;
        RECT 19.130 106.200 19.430 106.650 ;
        RECT 30.030 106.200 30.330 106.650 ;
        RECT 19.130 106.050 22.980 106.200 ;
        RECT 26.480 106.050 30.330 106.200 ;
        RECT 19.130 105.600 19.430 106.050 ;
        RECT 30.030 105.600 30.330 106.050 ;
        RECT 19.130 105.450 22.980 105.600 ;
        RECT 26.480 105.450 30.330 105.600 ;
        RECT 19.130 105.000 19.430 105.450 ;
        RECT 30.030 105.000 30.330 105.450 ;
        RECT 19.130 104.850 22.980 105.000 ;
        RECT 26.480 104.850 30.330 105.000 ;
        RECT 19.130 104.400 19.430 104.850 ;
        RECT 30.030 104.400 30.330 104.850 ;
        RECT 19.130 104.250 22.980 104.400 ;
        RECT 26.480 104.250 30.330 104.400 ;
        RECT 19.130 103.800 19.430 104.250 ;
        RECT 30.030 103.800 30.330 104.250 ;
        RECT 19.130 103.650 22.980 103.800 ;
        RECT 26.480 103.650 30.330 103.800 ;
        RECT 19.130 103.200 19.430 103.650 ;
        RECT 30.030 103.200 30.330 103.650 ;
        RECT 19.130 103.050 22.980 103.200 ;
        RECT 26.480 103.050 30.330 103.200 ;
        RECT 19.130 102.600 19.430 103.050 ;
        RECT 30.030 102.600 30.330 103.050 ;
        RECT 19.130 102.450 22.980 102.600 ;
        RECT 26.480 102.450 30.330 102.600 ;
        RECT 19.130 102.000 19.430 102.450 ;
        RECT 30.030 102.000 30.330 102.450 ;
        RECT 19.130 101.450 22.930 102.000 ;
        RECT 6.530 101.400 22.930 101.450 ;
        RECT 26.530 101.450 30.330 102.000 ;
        RECT 30.780 101.450 30.930 109.650 ;
        RECT 31.380 101.450 31.530 109.650 ;
        RECT 31.980 101.450 32.130 109.650 ;
        RECT 32.580 101.450 32.730 109.650 ;
        RECT 33.180 101.450 33.330 109.650 ;
        RECT 33.780 101.450 33.930 109.650 ;
        RECT 34.380 101.450 35.080 118.550 ;
        RECT 35.530 110.350 35.680 118.550 ;
        RECT 36.130 110.350 36.280 118.550 ;
        RECT 36.730 110.350 36.880 118.550 ;
        RECT 37.330 110.350 37.480 118.550 ;
        RECT 37.930 110.350 38.080 118.550 ;
        RECT 38.530 110.350 38.680 118.550 ;
        RECT 39.130 118.000 42.930 118.550 ;
        RECT 46.530 118.550 62.930 118.600 ;
        RECT 46.530 118.000 50.330 118.550 ;
        RECT 39.130 117.550 39.430 118.000 ;
        RECT 50.030 117.550 50.330 118.000 ;
        RECT 39.130 117.400 42.980 117.550 ;
        RECT 46.480 117.400 50.330 117.550 ;
        RECT 39.130 116.950 39.430 117.400 ;
        RECT 50.030 116.950 50.330 117.400 ;
        RECT 39.130 116.800 42.980 116.950 ;
        RECT 46.480 116.800 50.330 116.950 ;
        RECT 39.130 116.350 39.430 116.800 ;
        RECT 50.030 116.350 50.330 116.800 ;
        RECT 39.130 116.200 42.980 116.350 ;
        RECT 46.480 116.200 50.330 116.350 ;
        RECT 39.130 115.750 39.430 116.200 ;
        RECT 50.030 115.750 50.330 116.200 ;
        RECT 39.130 115.600 42.980 115.750 ;
        RECT 46.480 115.600 50.330 115.750 ;
        RECT 39.130 115.150 39.430 115.600 ;
        RECT 50.030 115.150 50.330 115.600 ;
        RECT 39.130 115.000 42.980 115.150 ;
        RECT 46.480 115.000 50.330 115.150 ;
        RECT 39.130 114.550 39.430 115.000 ;
        RECT 50.030 114.550 50.330 115.000 ;
        RECT 39.130 114.400 42.980 114.550 ;
        RECT 46.480 114.400 50.330 114.550 ;
        RECT 39.130 113.950 39.430 114.400 ;
        RECT 50.030 113.950 50.330 114.400 ;
        RECT 39.130 113.800 42.980 113.950 ;
        RECT 46.480 113.800 50.330 113.950 ;
        RECT 39.130 113.350 39.430 113.800 ;
        RECT 50.030 113.350 50.330 113.800 ;
        RECT 39.130 113.200 42.980 113.350 ;
        RECT 46.480 113.200 50.330 113.350 ;
        RECT 39.130 112.750 39.430 113.200 ;
        RECT 39.130 112.600 42.980 112.750 ;
        RECT 39.130 112.150 39.430 112.600 ;
        RECT 39.130 112.000 42.980 112.150 ;
        RECT 39.130 111.550 39.430 112.000 ;
        RECT 39.130 111.400 42.980 111.550 ;
        RECT 39.130 110.950 39.430 111.400 ;
        RECT 39.130 110.800 42.980 110.950 ;
        RECT 39.130 110.350 39.430 110.800 ;
        RECT 35.530 101.450 35.680 109.650 ;
        RECT 36.130 101.450 36.280 109.650 ;
        RECT 36.730 101.450 36.880 109.650 ;
        RECT 37.330 101.450 37.480 109.650 ;
        RECT 37.930 101.450 38.080 109.650 ;
        RECT 38.530 101.450 38.680 109.650 ;
        RECT 39.130 109.200 39.430 109.650 ;
        RECT 39.130 109.050 42.980 109.200 ;
        RECT 39.130 108.600 39.430 109.050 ;
        RECT 39.130 108.450 42.980 108.600 ;
        RECT 39.130 108.000 39.430 108.450 ;
        RECT 39.130 107.850 42.980 108.000 ;
        RECT 39.130 107.400 39.430 107.850 ;
        RECT 39.130 107.250 42.980 107.400 ;
        RECT 39.130 106.800 39.430 107.250 ;
        RECT 43.830 106.800 45.630 113.200 ;
        RECT 50.030 112.750 50.330 113.200 ;
        RECT 46.480 112.600 50.330 112.750 ;
        RECT 50.030 112.150 50.330 112.600 ;
        RECT 46.480 112.000 50.330 112.150 ;
        RECT 50.030 111.550 50.330 112.000 ;
        RECT 46.480 111.400 50.330 111.550 ;
        RECT 50.030 110.950 50.330 111.400 ;
        RECT 46.480 110.800 50.330 110.950 ;
        RECT 50.030 110.350 50.330 110.800 ;
        RECT 50.780 110.350 50.930 118.550 ;
        RECT 51.380 110.350 51.530 118.550 ;
        RECT 51.980 110.350 52.130 118.550 ;
        RECT 52.580 110.350 52.730 118.550 ;
        RECT 53.180 110.350 53.330 118.550 ;
        RECT 53.780 110.350 53.930 118.550 ;
        RECT 50.030 109.200 50.330 109.650 ;
        RECT 46.480 109.050 50.330 109.200 ;
        RECT 50.030 108.600 50.330 109.050 ;
        RECT 46.480 108.450 50.330 108.600 ;
        RECT 50.030 108.000 50.330 108.450 ;
        RECT 46.480 107.850 50.330 108.000 ;
        RECT 50.030 107.400 50.330 107.850 ;
        RECT 46.480 107.250 50.330 107.400 ;
        RECT 50.030 106.800 50.330 107.250 ;
        RECT 39.130 106.650 42.980 106.800 ;
        RECT 46.480 106.650 50.330 106.800 ;
        RECT 39.130 106.200 39.430 106.650 ;
        RECT 50.030 106.200 50.330 106.650 ;
        RECT 39.130 106.050 42.980 106.200 ;
        RECT 46.480 106.050 50.330 106.200 ;
        RECT 39.130 105.600 39.430 106.050 ;
        RECT 50.030 105.600 50.330 106.050 ;
        RECT 39.130 105.450 42.980 105.600 ;
        RECT 46.480 105.450 50.330 105.600 ;
        RECT 39.130 105.000 39.430 105.450 ;
        RECT 50.030 105.000 50.330 105.450 ;
        RECT 39.130 104.850 42.980 105.000 ;
        RECT 46.480 104.850 50.330 105.000 ;
        RECT 39.130 104.400 39.430 104.850 ;
        RECT 50.030 104.400 50.330 104.850 ;
        RECT 39.130 104.250 42.980 104.400 ;
        RECT 46.480 104.250 50.330 104.400 ;
        RECT 39.130 103.800 39.430 104.250 ;
        RECT 50.030 103.800 50.330 104.250 ;
        RECT 39.130 103.650 42.980 103.800 ;
        RECT 46.480 103.650 50.330 103.800 ;
        RECT 39.130 103.200 39.430 103.650 ;
        RECT 50.030 103.200 50.330 103.650 ;
        RECT 39.130 103.050 42.980 103.200 ;
        RECT 46.480 103.050 50.330 103.200 ;
        RECT 39.130 102.600 39.430 103.050 ;
        RECT 50.030 102.600 50.330 103.050 ;
        RECT 39.130 102.450 42.980 102.600 ;
        RECT 46.480 102.450 50.330 102.600 ;
        RECT 39.130 102.000 39.430 102.450 ;
        RECT 50.030 102.000 50.330 102.450 ;
        RECT 39.130 101.450 42.930 102.000 ;
        RECT 26.530 101.400 42.930 101.450 ;
        RECT 46.530 101.450 50.330 102.000 ;
        RECT 50.780 101.450 50.930 109.650 ;
        RECT 51.380 101.450 51.530 109.650 ;
        RECT 51.980 101.450 52.130 109.650 ;
        RECT 52.580 101.450 52.730 109.650 ;
        RECT 53.180 101.450 53.330 109.650 ;
        RECT 53.780 101.450 53.930 109.650 ;
        RECT 54.380 101.450 55.080 118.550 ;
        RECT 55.530 110.350 55.680 118.550 ;
        RECT 56.130 110.350 56.280 118.550 ;
        RECT 56.730 110.350 56.880 118.550 ;
        RECT 57.330 110.350 57.480 118.550 ;
        RECT 57.930 110.350 58.080 118.550 ;
        RECT 58.530 110.350 58.680 118.550 ;
        RECT 59.130 118.000 62.930 118.550 ;
        RECT 66.530 118.550 82.930 118.600 ;
        RECT 66.530 118.000 70.330 118.550 ;
        RECT 59.130 117.550 59.430 118.000 ;
        RECT 70.030 117.550 70.330 118.000 ;
        RECT 59.130 117.400 62.980 117.550 ;
        RECT 66.480 117.400 70.330 117.550 ;
        RECT 59.130 116.950 59.430 117.400 ;
        RECT 70.030 116.950 70.330 117.400 ;
        RECT 59.130 116.800 62.980 116.950 ;
        RECT 66.480 116.800 70.330 116.950 ;
        RECT 59.130 116.350 59.430 116.800 ;
        RECT 70.030 116.350 70.330 116.800 ;
        RECT 59.130 116.200 62.980 116.350 ;
        RECT 66.480 116.200 70.330 116.350 ;
        RECT 59.130 115.750 59.430 116.200 ;
        RECT 70.030 115.750 70.330 116.200 ;
        RECT 59.130 115.600 62.980 115.750 ;
        RECT 66.480 115.600 70.330 115.750 ;
        RECT 59.130 115.150 59.430 115.600 ;
        RECT 70.030 115.150 70.330 115.600 ;
        RECT 59.130 115.000 62.980 115.150 ;
        RECT 66.480 115.000 70.330 115.150 ;
        RECT 59.130 114.550 59.430 115.000 ;
        RECT 70.030 114.550 70.330 115.000 ;
        RECT 59.130 114.400 62.980 114.550 ;
        RECT 66.480 114.400 70.330 114.550 ;
        RECT 59.130 113.950 59.430 114.400 ;
        RECT 70.030 113.950 70.330 114.400 ;
        RECT 59.130 113.800 62.980 113.950 ;
        RECT 66.480 113.800 70.330 113.950 ;
        RECT 59.130 113.350 59.430 113.800 ;
        RECT 70.030 113.350 70.330 113.800 ;
        RECT 59.130 113.200 62.980 113.350 ;
        RECT 66.480 113.200 70.330 113.350 ;
        RECT 59.130 112.750 59.430 113.200 ;
        RECT 59.130 112.600 62.980 112.750 ;
        RECT 59.130 112.150 59.430 112.600 ;
        RECT 59.130 112.000 62.980 112.150 ;
        RECT 59.130 111.550 59.430 112.000 ;
        RECT 59.130 111.400 62.980 111.550 ;
        RECT 59.130 110.950 59.430 111.400 ;
        RECT 59.130 110.800 62.980 110.950 ;
        RECT 59.130 110.350 59.430 110.800 ;
        RECT 55.530 101.450 55.680 109.650 ;
        RECT 56.130 101.450 56.280 109.650 ;
        RECT 56.730 101.450 56.880 109.650 ;
        RECT 57.330 101.450 57.480 109.650 ;
        RECT 57.930 101.450 58.080 109.650 ;
        RECT 58.530 101.450 58.680 109.650 ;
        RECT 59.130 109.200 59.430 109.650 ;
        RECT 59.130 109.050 62.980 109.200 ;
        RECT 59.130 108.600 59.430 109.050 ;
        RECT 59.130 108.450 62.980 108.600 ;
        RECT 59.130 108.000 59.430 108.450 ;
        RECT 59.130 107.850 62.980 108.000 ;
        RECT 59.130 107.400 59.430 107.850 ;
        RECT 59.130 107.250 62.980 107.400 ;
        RECT 59.130 106.800 59.430 107.250 ;
        RECT 63.830 106.800 65.630 113.200 ;
        RECT 70.030 112.750 70.330 113.200 ;
        RECT 66.480 112.600 70.330 112.750 ;
        RECT 70.030 112.150 70.330 112.600 ;
        RECT 66.480 112.000 70.330 112.150 ;
        RECT 70.030 111.550 70.330 112.000 ;
        RECT 66.480 111.400 70.330 111.550 ;
        RECT 70.030 110.950 70.330 111.400 ;
        RECT 66.480 110.800 70.330 110.950 ;
        RECT 70.030 110.350 70.330 110.800 ;
        RECT 70.780 110.350 70.930 118.550 ;
        RECT 71.380 110.350 71.530 118.550 ;
        RECT 71.980 110.350 72.130 118.550 ;
        RECT 72.580 110.350 72.730 118.550 ;
        RECT 73.180 110.350 73.330 118.550 ;
        RECT 73.780 110.350 73.930 118.550 ;
        RECT 70.030 109.200 70.330 109.650 ;
        RECT 66.480 109.050 70.330 109.200 ;
        RECT 70.030 108.600 70.330 109.050 ;
        RECT 66.480 108.450 70.330 108.600 ;
        RECT 70.030 108.000 70.330 108.450 ;
        RECT 66.480 107.850 70.330 108.000 ;
        RECT 70.030 107.400 70.330 107.850 ;
        RECT 66.480 107.250 70.330 107.400 ;
        RECT 70.030 106.800 70.330 107.250 ;
        RECT 59.130 106.650 62.980 106.800 ;
        RECT 66.480 106.650 70.330 106.800 ;
        RECT 59.130 106.200 59.430 106.650 ;
        RECT 70.030 106.200 70.330 106.650 ;
        RECT 59.130 106.050 62.980 106.200 ;
        RECT 66.480 106.050 70.330 106.200 ;
        RECT 59.130 105.600 59.430 106.050 ;
        RECT 70.030 105.600 70.330 106.050 ;
        RECT 59.130 105.450 62.980 105.600 ;
        RECT 66.480 105.450 70.330 105.600 ;
        RECT 59.130 105.000 59.430 105.450 ;
        RECT 70.030 105.000 70.330 105.450 ;
        RECT 59.130 104.850 62.980 105.000 ;
        RECT 66.480 104.850 70.330 105.000 ;
        RECT 59.130 104.400 59.430 104.850 ;
        RECT 70.030 104.400 70.330 104.850 ;
        RECT 59.130 104.250 62.980 104.400 ;
        RECT 66.480 104.250 70.330 104.400 ;
        RECT 59.130 103.800 59.430 104.250 ;
        RECT 70.030 103.800 70.330 104.250 ;
        RECT 59.130 103.650 62.980 103.800 ;
        RECT 66.480 103.650 70.330 103.800 ;
        RECT 59.130 103.200 59.430 103.650 ;
        RECT 70.030 103.200 70.330 103.650 ;
        RECT 59.130 103.050 62.980 103.200 ;
        RECT 66.480 103.050 70.330 103.200 ;
        RECT 59.130 102.600 59.430 103.050 ;
        RECT 70.030 102.600 70.330 103.050 ;
        RECT 59.130 102.450 62.980 102.600 ;
        RECT 66.480 102.450 70.330 102.600 ;
        RECT 59.130 102.000 59.430 102.450 ;
        RECT 70.030 102.000 70.330 102.450 ;
        RECT 59.130 101.450 62.930 102.000 ;
        RECT 46.530 101.400 62.930 101.450 ;
        RECT 66.530 101.450 70.330 102.000 ;
        RECT 70.780 101.450 70.930 109.650 ;
        RECT 71.380 101.450 71.530 109.650 ;
        RECT 71.980 101.450 72.130 109.650 ;
        RECT 72.580 101.450 72.730 109.650 ;
        RECT 73.180 101.450 73.330 109.650 ;
        RECT 73.780 101.450 73.930 109.650 ;
        RECT 74.380 101.450 75.080 118.550 ;
        RECT 75.530 110.350 75.680 118.550 ;
        RECT 76.130 110.350 76.280 118.550 ;
        RECT 76.730 110.350 76.880 118.550 ;
        RECT 77.330 110.350 77.480 118.550 ;
        RECT 77.930 110.350 78.080 118.550 ;
        RECT 78.530 110.350 78.680 118.550 ;
        RECT 79.130 118.000 82.930 118.550 ;
        RECT 86.530 118.550 102.930 118.600 ;
        RECT 86.530 118.000 90.330 118.550 ;
        RECT 79.130 117.550 79.430 118.000 ;
        RECT 90.030 117.550 90.330 118.000 ;
        RECT 79.130 117.400 82.980 117.550 ;
        RECT 86.480 117.400 90.330 117.550 ;
        RECT 79.130 116.950 79.430 117.400 ;
        RECT 90.030 116.950 90.330 117.400 ;
        RECT 79.130 116.800 82.980 116.950 ;
        RECT 86.480 116.800 90.330 116.950 ;
        RECT 79.130 116.350 79.430 116.800 ;
        RECT 90.030 116.350 90.330 116.800 ;
        RECT 79.130 116.200 82.980 116.350 ;
        RECT 86.480 116.200 90.330 116.350 ;
        RECT 79.130 115.750 79.430 116.200 ;
        RECT 90.030 115.750 90.330 116.200 ;
        RECT 79.130 115.600 82.980 115.750 ;
        RECT 86.480 115.600 90.330 115.750 ;
        RECT 79.130 115.150 79.430 115.600 ;
        RECT 90.030 115.150 90.330 115.600 ;
        RECT 79.130 115.000 82.980 115.150 ;
        RECT 86.480 115.000 90.330 115.150 ;
        RECT 79.130 114.550 79.430 115.000 ;
        RECT 90.030 114.550 90.330 115.000 ;
        RECT 79.130 114.400 82.980 114.550 ;
        RECT 86.480 114.400 90.330 114.550 ;
        RECT 79.130 113.950 79.430 114.400 ;
        RECT 90.030 113.950 90.330 114.400 ;
        RECT 79.130 113.800 82.980 113.950 ;
        RECT 86.480 113.800 90.330 113.950 ;
        RECT 79.130 113.350 79.430 113.800 ;
        RECT 90.030 113.350 90.330 113.800 ;
        RECT 79.130 113.200 82.980 113.350 ;
        RECT 86.480 113.200 90.330 113.350 ;
        RECT 79.130 112.750 79.430 113.200 ;
        RECT 79.130 112.600 82.980 112.750 ;
        RECT 79.130 112.150 79.430 112.600 ;
        RECT 79.130 112.000 82.980 112.150 ;
        RECT 79.130 111.550 79.430 112.000 ;
        RECT 79.130 111.400 82.980 111.550 ;
        RECT 79.130 110.950 79.430 111.400 ;
        RECT 79.130 110.800 82.980 110.950 ;
        RECT 79.130 110.350 79.430 110.800 ;
        RECT 75.530 101.450 75.680 109.650 ;
        RECT 76.130 101.450 76.280 109.650 ;
        RECT 76.730 101.450 76.880 109.650 ;
        RECT 77.330 101.450 77.480 109.650 ;
        RECT 77.930 101.450 78.080 109.650 ;
        RECT 78.530 101.450 78.680 109.650 ;
        RECT 79.130 109.200 79.430 109.650 ;
        RECT 79.130 109.050 82.980 109.200 ;
        RECT 79.130 108.600 79.430 109.050 ;
        RECT 79.130 108.450 82.980 108.600 ;
        RECT 79.130 108.000 79.430 108.450 ;
        RECT 79.130 107.850 82.980 108.000 ;
        RECT 79.130 107.400 79.430 107.850 ;
        RECT 79.130 107.250 82.980 107.400 ;
        RECT 79.130 106.800 79.430 107.250 ;
        RECT 83.830 106.800 85.630 113.200 ;
        RECT 90.030 112.750 90.330 113.200 ;
        RECT 86.480 112.600 90.330 112.750 ;
        RECT 90.030 112.150 90.330 112.600 ;
        RECT 86.480 112.000 90.330 112.150 ;
        RECT 90.030 111.550 90.330 112.000 ;
        RECT 86.480 111.400 90.330 111.550 ;
        RECT 90.030 110.950 90.330 111.400 ;
        RECT 86.480 110.800 90.330 110.950 ;
        RECT 90.030 110.350 90.330 110.800 ;
        RECT 90.780 110.350 90.930 118.550 ;
        RECT 91.380 110.350 91.530 118.550 ;
        RECT 91.980 110.350 92.130 118.550 ;
        RECT 92.580 110.350 92.730 118.550 ;
        RECT 93.180 110.350 93.330 118.550 ;
        RECT 93.780 110.350 93.930 118.550 ;
        RECT 90.030 109.200 90.330 109.650 ;
        RECT 86.480 109.050 90.330 109.200 ;
        RECT 90.030 108.600 90.330 109.050 ;
        RECT 86.480 108.450 90.330 108.600 ;
        RECT 90.030 108.000 90.330 108.450 ;
        RECT 86.480 107.850 90.330 108.000 ;
        RECT 90.030 107.400 90.330 107.850 ;
        RECT 86.480 107.250 90.330 107.400 ;
        RECT 90.030 106.800 90.330 107.250 ;
        RECT 79.130 106.650 82.980 106.800 ;
        RECT 86.480 106.650 90.330 106.800 ;
        RECT 79.130 106.200 79.430 106.650 ;
        RECT 90.030 106.200 90.330 106.650 ;
        RECT 79.130 106.050 82.980 106.200 ;
        RECT 86.480 106.050 90.330 106.200 ;
        RECT 79.130 105.600 79.430 106.050 ;
        RECT 90.030 105.600 90.330 106.050 ;
        RECT 79.130 105.450 82.980 105.600 ;
        RECT 86.480 105.450 90.330 105.600 ;
        RECT 79.130 105.000 79.430 105.450 ;
        RECT 90.030 105.000 90.330 105.450 ;
        RECT 79.130 104.850 82.980 105.000 ;
        RECT 86.480 104.850 90.330 105.000 ;
        RECT 79.130 104.400 79.430 104.850 ;
        RECT 90.030 104.400 90.330 104.850 ;
        RECT 79.130 104.250 82.980 104.400 ;
        RECT 86.480 104.250 90.330 104.400 ;
        RECT 79.130 103.800 79.430 104.250 ;
        RECT 90.030 103.800 90.330 104.250 ;
        RECT 79.130 103.650 82.980 103.800 ;
        RECT 86.480 103.650 90.330 103.800 ;
        RECT 79.130 103.200 79.430 103.650 ;
        RECT 90.030 103.200 90.330 103.650 ;
        RECT 79.130 103.050 82.980 103.200 ;
        RECT 86.480 103.050 90.330 103.200 ;
        RECT 79.130 102.600 79.430 103.050 ;
        RECT 90.030 102.600 90.330 103.050 ;
        RECT 79.130 102.450 82.980 102.600 ;
        RECT 86.480 102.450 90.330 102.600 ;
        RECT 79.130 102.000 79.430 102.450 ;
        RECT 90.030 102.000 90.330 102.450 ;
        RECT 79.130 101.450 82.930 102.000 ;
        RECT 66.530 101.400 82.930 101.450 ;
        RECT 86.530 101.450 90.330 102.000 ;
        RECT 90.780 101.450 90.930 109.650 ;
        RECT 91.380 101.450 91.530 109.650 ;
        RECT 91.980 101.450 92.130 109.650 ;
        RECT 92.580 101.450 92.730 109.650 ;
        RECT 93.180 101.450 93.330 109.650 ;
        RECT 93.780 101.450 93.930 109.650 ;
        RECT 94.380 101.450 95.080 118.550 ;
        RECT 95.530 110.350 95.680 118.550 ;
        RECT 96.130 110.350 96.280 118.550 ;
        RECT 96.730 110.350 96.880 118.550 ;
        RECT 97.330 110.350 97.480 118.550 ;
        RECT 97.930 110.350 98.080 118.550 ;
        RECT 98.530 110.350 98.680 118.550 ;
        RECT 99.130 118.000 102.930 118.550 ;
        RECT 106.530 118.550 122.930 118.600 ;
        RECT 106.530 118.000 110.330 118.550 ;
        RECT 99.130 117.550 99.430 118.000 ;
        RECT 110.030 117.550 110.330 118.000 ;
        RECT 99.130 117.400 102.980 117.550 ;
        RECT 106.480 117.400 110.330 117.550 ;
        RECT 99.130 116.950 99.430 117.400 ;
        RECT 110.030 116.950 110.330 117.400 ;
        RECT 99.130 116.800 102.980 116.950 ;
        RECT 106.480 116.800 110.330 116.950 ;
        RECT 99.130 116.350 99.430 116.800 ;
        RECT 110.030 116.350 110.330 116.800 ;
        RECT 99.130 116.200 102.980 116.350 ;
        RECT 106.480 116.200 110.330 116.350 ;
        RECT 99.130 115.750 99.430 116.200 ;
        RECT 110.030 115.750 110.330 116.200 ;
        RECT 99.130 115.600 102.980 115.750 ;
        RECT 106.480 115.600 110.330 115.750 ;
        RECT 99.130 115.150 99.430 115.600 ;
        RECT 110.030 115.150 110.330 115.600 ;
        RECT 99.130 115.000 102.980 115.150 ;
        RECT 106.480 115.000 110.330 115.150 ;
        RECT 99.130 114.550 99.430 115.000 ;
        RECT 110.030 114.550 110.330 115.000 ;
        RECT 99.130 114.400 102.980 114.550 ;
        RECT 106.480 114.400 110.330 114.550 ;
        RECT 99.130 113.950 99.430 114.400 ;
        RECT 110.030 113.950 110.330 114.400 ;
        RECT 99.130 113.800 102.980 113.950 ;
        RECT 106.480 113.800 110.330 113.950 ;
        RECT 99.130 113.350 99.430 113.800 ;
        RECT 110.030 113.350 110.330 113.800 ;
        RECT 99.130 113.200 102.980 113.350 ;
        RECT 106.480 113.200 110.330 113.350 ;
        RECT 99.130 112.750 99.430 113.200 ;
        RECT 99.130 112.600 102.980 112.750 ;
        RECT 99.130 112.150 99.430 112.600 ;
        RECT 99.130 112.000 102.980 112.150 ;
        RECT 99.130 111.550 99.430 112.000 ;
        RECT 99.130 111.400 102.980 111.550 ;
        RECT 99.130 110.950 99.430 111.400 ;
        RECT 99.130 110.800 102.980 110.950 ;
        RECT 99.130 110.350 99.430 110.800 ;
        RECT 95.530 101.450 95.680 109.650 ;
        RECT 96.130 101.450 96.280 109.650 ;
        RECT 96.730 101.450 96.880 109.650 ;
        RECT 97.330 101.450 97.480 109.650 ;
        RECT 97.930 101.450 98.080 109.650 ;
        RECT 98.530 101.450 98.680 109.650 ;
        RECT 99.130 109.200 99.430 109.650 ;
        RECT 99.130 109.050 102.980 109.200 ;
        RECT 99.130 108.600 99.430 109.050 ;
        RECT 99.130 108.450 102.980 108.600 ;
        RECT 99.130 108.000 99.430 108.450 ;
        RECT 99.130 107.850 102.980 108.000 ;
        RECT 99.130 107.400 99.430 107.850 ;
        RECT 99.130 107.250 102.980 107.400 ;
        RECT 99.130 106.800 99.430 107.250 ;
        RECT 103.830 106.800 105.630 113.200 ;
        RECT 110.030 112.750 110.330 113.200 ;
        RECT 106.480 112.600 110.330 112.750 ;
        RECT 110.030 112.150 110.330 112.600 ;
        RECT 106.480 112.000 110.330 112.150 ;
        RECT 110.030 111.550 110.330 112.000 ;
        RECT 106.480 111.400 110.330 111.550 ;
        RECT 110.030 110.950 110.330 111.400 ;
        RECT 106.480 110.800 110.330 110.950 ;
        RECT 110.030 110.350 110.330 110.800 ;
        RECT 110.780 110.350 110.930 118.550 ;
        RECT 111.380 110.350 111.530 118.550 ;
        RECT 111.980 110.350 112.130 118.550 ;
        RECT 112.580 110.350 112.730 118.550 ;
        RECT 113.180 110.350 113.330 118.550 ;
        RECT 113.780 110.350 113.930 118.550 ;
        RECT 110.030 109.200 110.330 109.650 ;
        RECT 106.480 109.050 110.330 109.200 ;
        RECT 110.030 108.600 110.330 109.050 ;
        RECT 106.480 108.450 110.330 108.600 ;
        RECT 110.030 108.000 110.330 108.450 ;
        RECT 106.480 107.850 110.330 108.000 ;
        RECT 110.030 107.400 110.330 107.850 ;
        RECT 106.480 107.250 110.330 107.400 ;
        RECT 110.030 106.800 110.330 107.250 ;
        RECT 99.130 106.650 102.980 106.800 ;
        RECT 106.480 106.650 110.330 106.800 ;
        RECT 99.130 106.200 99.430 106.650 ;
        RECT 110.030 106.200 110.330 106.650 ;
        RECT 99.130 106.050 102.980 106.200 ;
        RECT 106.480 106.050 110.330 106.200 ;
        RECT 99.130 105.600 99.430 106.050 ;
        RECT 110.030 105.600 110.330 106.050 ;
        RECT 99.130 105.450 102.980 105.600 ;
        RECT 106.480 105.450 110.330 105.600 ;
        RECT 99.130 105.000 99.430 105.450 ;
        RECT 110.030 105.000 110.330 105.450 ;
        RECT 99.130 104.850 102.980 105.000 ;
        RECT 106.480 104.850 110.330 105.000 ;
        RECT 99.130 104.400 99.430 104.850 ;
        RECT 110.030 104.400 110.330 104.850 ;
        RECT 99.130 104.250 102.980 104.400 ;
        RECT 106.480 104.250 110.330 104.400 ;
        RECT 99.130 103.800 99.430 104.250 ;
        RECT 110.030 103.800 110.330 104.250 ;
        RECT 99.130 103.650 102.980 103.800 ;
        RECT 106.480 103.650 110.330 103.800 ;
        RECT 99.130 103.200 99.430 103.650 ;
        RECT 110.030 103.200 110.330 103.650 ;
        RECT 99.130 103.050 102.980 103.200 ;
        RECT 106.480 103.050 110.330 103.200 ;
        RECT 99.130 102.600 99.430 103.050 ;
        RECT 110.030 102.600 110.330 103.050 ;
        RECT 99.130 102.450 102.980 102.600 ;
        RECT 106.480 102.450 110.330 102.600 ;
        RECT 99.130 102.000 99.430 102.450 ;
        RECT 110.030 102.000 110.330 102.450 ;
        RECT 99.130 101.450 102.930 102.000 ;
        RECT 86.530 101.400 102.930 101.450 ;
        RECT 106.530 101.450 110.330 102.000 ;
        RECT 110.780 101.450 110.930 109.650 ;
        RECT 111.380 101.450 111.530 109.650 ;
        RECT 111.980 101.450 112.130 109.650 ;
        RECT 112.580 101.450 112.730 109.650 ;
        RECT 113.180 101.450 113.330 109.650 ;
        RECT 113.780 101.450 113.930 109.650 ;
        RECT 114.380 101.450 115.080 118.550 ;
        RECT 115.530 110.350 115.680 118.550 ;
        RECT 116.130 110.350 116.280 118.550 ;
        RECT 116.730 110.350 116.880 118.550 ;
        RECT 117.330 110.350 117.480 118.550 ;
        RECT 117.930 110.350 118.080 118.550 ;
        RECT 118.530 110.350 118.680 118.550 ;
        RECT 119.130 118.000 122.930 118.550 ;
        RECT 119.130 117.550 119.430 118.000 ;
        RECT 119.130 117.400 122.980 117.550 ;
        RECT 119.130 116.950 119.430 117.400 ;
        RECT 119.130 116.800 122.980 116.950 ;
        RECT 119.130 116.350 119.430 116.800 ;
        RECT 119.130 116.200 122.980 116.350 ;
        RECT 119.130 115.750 119.430 116.200 ;
        RECT 119.130 115.600 122.980 115.750 ;
        RECT 119.130 115.150 119.430 115.600 ;
        RECT 119.130 115.000 122.980 115.150 ;
        RECT 119.130 114.550 119.430 115.000 ;
        RECT 119.130 114.400 122.980 114.550 ;
        RECT 119.130 113.950 119.430 114.400 ;
        RECT 119.130 113.800 122.980 113.950 ;
        RECT 119.130 113.350 119.430 113.800 ;
        RECT 119.130 113.200 122.980 113.350 ;
        RECT 119.130 112.750 119.430 113.200 ;
        RECT 119.130 112.600 122.980 112.750 ;
        RECT 119.130 112.150 119.430 112.600 ;
        RECT 119.130 112.000 122.980 112.150 ;
        RECT 119.130 111.550 119.430 112.000 ;
        RECT 119.130 111.400 122.980 111.550 ;
        RECT 119.130 110.950 119.430 111.400 ;
        RECT 119.130 110.800 122.980 110.950 ;
        RECT 119.130 110.350 119.430 110.800 ;
        RECT 115.530 101.450 115.680 109.650 ;
        RECT 116.130 101.450 116.280 109.650 ;
        RECT 116.730 101.450 116.880 109.650 ;
        RECT 117.330 101.450 117.480 109.650 ;
        RECT 117.930 101.450 118.080 109.650 ;
        RECT 118.530 101.450 118.680 109.650 ;
        RECT 119.130 109.200 119.430 109.650 ;
        RECT 119.130 109.050 122.980 109.200 ;
        RECT 119.130 108.600 119.430 109.050 ;
        RECT 119.130 108.450 122.980 108.600 ;
        RECT 119.130 108.000 119.430 108.450 ;
        RECT 119.130 107.850 122.980 108.000 ;
        RECT 119.130 107.400 119.430 107.850 ;
        RECT 119.130 107.250 122.980 107.400 ;
        RECT 119.130 106.800 119.430 107.250 ;
        RECT 123.830 106.800 124.730 113.200 ;
        RECT 129.850 108.705 131.850 109.980 ;
        RECT 119.130 106.650 122.980 106.800 ;
        RECT 119.130 106.200 119.430 106.650 ;
        RECT 119.130 106.050 122.980 106.200 ;
        RECT 119.130 105.600 119.430 106.050 ;
        RECT 119.130 105.450 122.980 105.600 ;
        RECT 119.130 105.000 119.430 105.450 ;
        RECT 119.130 104.850 122.980 105.000 ;
        RECT 119.130 104.400 119.430 104.850 ;
        RECT 119.130 104.250 122.980 104.400 ;
        RECT 119.130 103.800 119.430 104.250 ;
        RECT 119.130 103.650 122.980 103.800 ;
        RECT 119.130 103.200 119.430 103.650 ;
        RECT 119.130 103.050 122.980 103.200 ;
        RECT 119.130 102.600 119.430 103.050 ;
        RECT 119.130 102.450 122.980 102.600 ;
        RECT 119.130 102.000 119.430 102.450 ;
        RECT 119.130 101.450 122.930 102.000 ;
        RECT 106.530 101.400 122.930 101.450 ;
        RECT 9.630 100.900 19.830 101.400 ;
        RECT 29.630 100.900 39.830 101.400 ;
        RECT 49.630 100.900 59.830 101.400 ;
        RECT 69.630 100.900 79.830 101.400 ;
        RECT 89.630 100.900 99.830 101.400 ;
        RECT 109.630 100.900 119.830 101.400 ;
        RECT 11.530 99.100 17.930 100.900 ;
        RECT 31.530 99.100 37.930 100.900 ;
        RECT 51.530 99.100 57.930 100.900 ;
        RECT 71.530 99.100 77.930 100.900 ;
        RECT 91.530 99.100 97.930 100.900 ;
        RECT 111.530 99.100 117.930 100.900 ;
        RECT 9.630 98.600 19.830 99.100 ;
        RECT 29.630 98.600 39.830 99.100 ;
        RECT 49.630 98.600 59.830 99.100 ;
        RECT 69.630 98.600 79.830 99.100 ;
        RECT 89.630 98.600 99.830 99.100 ;
        RECT 109.630 98.600 119.830 99.100 ;
        RECT 6.530 98.550 22.930 98.600 ;
        RECT 6.530 98.000 10.330 98.550 ;
        RECT 10.030 97.550 10.330 98.000 ;
        RECT 6.480 97.400 10.330 97.550 ;
        RECT 10.030 96.950 10.330 97.400 ;
        RECT 6.480 96.800 10.330 96.950 ;
        RECT 10.030 96.350 10.330 96.800 ;
        RECT 6.480 96.200 10.330 96.350 ;
        RECT 10.030 95.750 10.330 96.200 ;
        RECT 6.480 95.600 10.330 95.750 ;
        RECT 10.030 95.150 10.330 95.600 ;
        RECT 6.480 95.000 10.330 95.150 ;
        RECT 10.030 94.550 10.330 95.000 ;
        RECT 6.480 94.400 10.330 94.550 ;
        RECT 10.030 93.950 10.330 94.400 ;
        RECT 6.480 93.800 10.330 93.950 ;
        RECT 10.030 93.350 10.330 93.800 ;
        RECT 6.480 93.200 10.330 93.350 ;
        RECT 4.730 86.800 5.630 93.200 ;
        RECT 10.030 92.750 10.330 93.200 ;
        RECT 6.480 92.600 10.330 92.750 ;
        RECT 10.030 92.150 10.330 92.600 ;
        RECT 6.480 92.000 10.330 92.150 ;
        RECT 10.030 91.550 10.330 92.000 ;
        RECT 6.480 91.400 10.330 91.550 ;
        RECT 10.030 90.950 10.330 91.400 ;
        RECT 6.480 90.800 10.330 90.950 ;
        RECT 10.030 90.350 10.330 90.800 ;
        RECT 10.780 90.350 10.930 98.550 ;
        RECT 11.380 90.350 11.530 98.550 ;
        RECT 11.980 90.350 12.130 98.550 ;
        RECT 12.580 90.350 12.730 98.550 ;
        RECT 13.180 90.350 13.330 98.550 ;
        RECT 13.780 90.350 13.930 98.550 ;
        RECT 10.030 89.200 10.330 89.650 ;
        RECT 6.480 89.050 10.330 89.200 ;
        RECT 10.030 88.600 10.330 89.050 ;
        RECT 6.480 88.450 10.330 88.600 ;
        RECT 10.030 88.000 10.330 88.450 ;
        RECT 6.480 87.850 10.330 88.000 ;
        RECT 10.030 87.400 10.330 87.850 ;
        RECT 6.480 87.250 10.330 87.400 ;
        RECT 10.030 86.800 10.330 87.250 ;
        RECT 6.480 86.650 10.330 86.800 ;
        RECT 10.030 86.200 10.330 86.650 ;
        RECT 6.480 86.050 10.330 86.200 ;
        RECT 10.030 85.600 10.330 86.050 ;
        RECT 6.480 85.450 10.330 85.600 ;
        RECT 10.030 85.000 10.330 85.450 ;
        RECT 6.480 84.850 10.330 85.000 ;
        RECT 10.030 84.400 10.330 84.850 ;
        RECT 6.480 84.250 10.330 84.400 ;
        RECT 10.030 83.800 10.330 84.250 ;
        RECT 6.480 83.650 10.330 83.800 ;
        RECT 10.030 83.200 10.330 83.650 ;
        RECT 6.480 83.050 10.330 83.200 ;
        RECT 10.030 82.600 10.330 83.050 ;
        RECT 6.480 82.450 10.330 82.600 ;
        RECT 10.030 82.000 10.330 82.450 ;
        RECT 6.530 81.450 10.330 82.000 ;
        RECT 10.780 81.450 10.930 89.650 ;
        RECT 11.380 81.450 11.530 89.650 ;
        RECT 11.980 81.450 12.130 89.650 ;
        RECT 12.580 81.450 12.730 89.650 ;
        RECT 13.180 81.450 13.330 89.650 ;
        RECT 13.780 81.450 13.930 89.650 ;
        RECT 14.380 81.450 15.080 98.550 ;
        RECT 15.530 90.350 15.680 98.550 ;
        RECT 16.130 90.350 16.280 98.550 ;
        RECT 16.730 90.350 16.880 98.550 ;
        RECT 17.330 90.350 17.480 98.550 ;
        RECT 17.930 90.350 18.080 98.550 ;
        RECT 18.530 90.350 18.680 98.550 ;
        RECT 19.130 98.000 22.930 98.550 ;
        RECT 26.530 98.550 42.930 98.600 ;
        RECT 26.530 98.000 30.330 98.550 ;
        RECT 19.130 97.550 19.430 98.000 ;
        RECT 30.030 97.550 30.330 98.000 ;
        RECT 19.130 97.400 22.980 97.550 ;
        RECT 26.480 97.400 30.330 97.550 ;
        RECT 19.130 96.950 19.430 97.400 ;
        RECT 30.030 96.950 30.330 97.400 ;
        RECT 19.130 96.800 22.980 96.950 ;
        RECT 26.480 96.800 30.330 96.950 ;
        RECT 19.130 96.350 19.430 96.800 ;
        RECT 30.030 96.350 30.330 96.800 ;
        RECT 19.130 96.200 22.980 96.350 ;
        RECT 26.480 96.200 30.330 96.350 ;
        RECT 19.130 95.750 19.430 96.200 ;
        RECT 30.030 95.750 30.330 96.200 ;
        RECT 19.130 95.600 22.980 95.750 ;
        RECT 26.480 95.600 30.330 95.750 ;
        RECT 19.130 95.150 19.430 95.600 ;
        RECT 30.030 95.150 30.330 95.600 ;
        RECT 19.130 95.000 22.980 95.150 ;
        RECT 26.480 95.000 30.330 95.150 ;
        RECT 19.130 94.550 19.430 95.000 ;
        RECT 30.030 94.550 30.330 95.000 ;
        RECT 19.130 94.400 22.980 94.550 ;
        RECT 26.480 94.400 30.330 94.550 ;
        RECT 19.130 93.950 19.430 94.400 ;
        RECT 30.030 93.950 30.330 94.400 ;
        RECT 19.130 93.800 22.980 93.950 ;
        RECT 26.480 93.800 30.330 93.950 ;
        RECT 19.130 93.350 19.430 93.800 ;
        RECT 30.030 93.350 30.330 93.800 ;
        RECT 19.130 93.200 22.980 93.350 ;
        RECT 26.480 93.200 30.330 93.350 ;
        RECT 19.130 92.750 19.430 93.200 ;
        RECT 19.130 92.600 22.980 92.750 ;
        RECT 19.130 92.150 19.430 92.600 ;
        RECT 19.130 92.000 22.980 92.150 ;
        RECT 19.130 91.550 19.430 92.000 ;
        RECT 19.130 91.400 22.980 91.550 ;
        RECT 19.130 90.950 19.430 91.400 ;
        RECT 19.130 90.800 22.980 90.950 ;
        RECT 19.130 90.350 19.430 90.800 ;
        RECT 15.530 81.450 15.680 89.650 ;
        RECT 16.130 81.450 16.280 89.650 ;
        RECT 16.730 81.450 16.880 89.650 ;
        RECT 17.330 81.450 17.480 89.650 ;
        RECT 17.930 81.450 18.080 89.650 ;
        RECT 18.530 81.450 18.680 89.650 ;
        RECT 19.130 89.200 19.430 89.650 ;
        RECT 19.130 89.050 22.980 89.200 ;
        RECT 19.130 88.600 19.430 89.050 ;
        RECT 19.130 88.450 22.980 88.600 ;
        RECT 19.130 88.000 19.430 88.450 ;
        RECT 19.130 87.850 22.980 88.000 ;
        RECT 19.130 87.400 19.430 87.850 ;
        RECT 19.130 87.250 22.980 87.400 ;
        RECT 19.130 86.800 19.430 87.250 ;
        RECT 23.830 86.800 25.630 93.200 ;
        RECT 30.030 92.750 30.330 93.200 ;
        RECT 26.480 92.600 30.330 92.750 ;
        RECT 30.030 92.150 30.330 92.600 ;
        RECT 26.480 92.000 30.330 92.150 ;
        RECT 30.030 91.550 30.330 92.000 ;
        RECT 26.480 91.400 30.330 91.550 ;
        RECT 30.030 90.950 30.330 91.400 ;
        RECT 26.480 90.800 30.330 90.950 ;
        RECT 30.030 90.350 30.330 90.800 ;
        RECT 30.780 90.350 30.930 98.550 ;
        RECT 31.380 90.350 31.530 98.550 ;
        RECT 31.980 90.350 32.130 98.550 ;
        RECT 32.580 90.350 32.730 98.550 ;
        RECT 33.180 90.350 33.330 98.550 ;
        RECT 33.780 90.350 33.930 98.550 ;
        RECT 30.030 89.200 30.330 89.650 ;
        RECT 26.480 89.050 30.330 89.200 ;
        RECT 30.030 88.600 30.330 89.050 ;
        RECT 26.480 88.450 30.330 88.600 ;
        RECT 30.030 88.000 30.330 88.450 ;
        RECT 26.480 87.850 30.330 88.000 ;
        RECT 30.030 87.400 30.330 87.850 ;
        RECT 26.480 87.250 30.330 87.400 ;
        RECT 30.030 86.800 30.330 87.250 ;
        RECT 19.130 86.650 22.980 86.800 ;
        RECT 26.480 86.650 30.330 86.800 ;
        RECT 19.130 86.200 19.430 86.650 ;
        RECT 30.030 86.200 30.330 86.650 ;
        RECT 19.130 86.050 22.980 86.200 ;
        RECT 26.480 86.050 30.330 86.200 ;
        RECT 19.130 85.600 19.430 86.050 ;
        RECT 30.030 85.600 30.330 86.050 ;
        RECT 19.130 85.450 22.980 85.600 ;
        RECT 26.480 85.450 30.330 85.600 ;
        RECT 19.130 85.000 19.430 85.450 ;
        RECT 30.030 85.000 30.330 85.450 ;
        RECT 19.130 84.850 22.980 85.000 ;
        RECT 26.480 84.850 30.330 85.000 ;
        RECT 19.130 84.400 19.430 84.850 ;
        RECT 30.030 84.400 30.330 84.850 ;
        RECT 19.130 84.250 22.980 84.400 ;
        RECT 26.480 84.250 30.330 84.400 ;
        RECT 19.130 83.800 19.430 84.250 ;
        RECT 30.030 83.800 30.330 84.250 ;
        RECT 19.130 83.650 22.980 83.800 ;
        RECT 26.480 83.650 30.330 83.800 ;
        RECT 19.130 83.200 19.430 83.650 ;
        RECT 30.030 83.200 30.330 83.650 ;
        RECT 19.130 83.050 22.980 83.200 ;
        RECT 26.480 83.050 30.330 83.200 ;
        RECT 19.130 82.600 19.430 83.050 ;
        RECT 30.030 82.600 30.330 83.050 ;
        RECT 19.130 82.450 22.980 82.600 ;
        RECT 26.480 82.450 30.330 82.600 ;
        RECT 19.130 82.000 19.430 82.450 ;
        RECT 30.030 82.000 30.330 82.450 ;
        RECT 19.130 81.450 22.930 82.000 ;
        RECT 6.530 81.400 22.930 81.450 ;
        RECT 26.530 81.450 30.330 82.000 ;
        RECT 30.780 81.450 30.930 89.650 ;
        RECT 31.380 81.450 31.530 89.650 ;
        RECT 31.980 81.450 32.130 89.650 ;
        RECT 32.580 81.450 32.730 89.650 ;
        RECT 33.180 81.450 33.330 89.650 ;
        RECT 33.780 81.450 33.930 89.650 ;
        RECT 34.380 81.450 35.080 98.550 ;
        RECT 35.530 90.350 35.680 98.550 ;
        RECT 36.130 90.350 36.280 98.550 ;
        RECT 36.730 90.350 36.880 98.550 ;
        RECT 37.330 90.350 37.480 98.550 ;
        RECT 37.930 90.350 38.080 98.550 ;
        RECT 38.530 90.350 38.680 98.550 ;
        RECT 39.130 98.000 42.930 98.550 ;
        RECT 46.530 98.550 62.930 98.600 ;
        RECT 46.530 98.000 50.330 98.550 ;
        RECT 39.130 97.550 39.430 98.000 ;
        RECT 50.030 97.550 50.330 98.000 ;
        RECT 39.130 97.400 42.980 97.550 ;
        RECT 46.480 97.400 50.330 97.550 ;
        RECT 39.130 96.950 39.430 97.400 ;
        RECT 50.030 96.950 50.330 97.400 ;
        RECT 39.130 96.800 42.980 96.950 ;
        RECT 46.480 96.800 50.330 96.950 ;
        RECT 39.130 96.350 39.430 96.800 ;
        RECT 50.030 96.350 50.330 96.800 ;
        RECT 39.130 96.200 42.980 96.350 ;
        RECT 46.480 96.200 50.330 96.350 ;
        RECT 39.130 95.750 39.430 96.200 ;
        RECT 50.030 95.750 50.330 96.200 ;
        RECT 39.130 95.600 42.980 95.750 ;
        RECT 46.480 95.600 50.330 95.750 ;
        RECT 39.130 95.150 39.430 95.600 ;
        RECT 50.030 95.150 50.330 95.600 ;
        RECT 39.130 95.000 42.980 95.150 ;
        RECT 46.480 95.000 50.330 95.150 ;
        RECT 39.130 94.550 39.430 95.000 ;
        RECT 50.030 94.550 50.330 95.000 ;
        RECT 39.130 94.400 42.980 94.550 ;
        RECT 46.480 94.400 50.330 94.550 ;
        RECT 39.130 93.950 39.430 94.400 ;
        RECT 50.030 93.950 50.330 94.400 ;
        RECT 39.130 93.800 42.980 93.950 ;
        RECT 46.480 93.800 50.330 93.950 ;
        RECT 39.130 93.350 39.430 93.800 ;
        RECT 50.030 93.350 50.330 93.800 ;
        RECT 39.130 93.200 42.980 93.350 ;
        RECT 46.480 93.200 50.330 93.350 ;
        RECT 39.130 92.750 39.430 93.200 ;
        RECT 39.130 92.600 42.980 92.750 ;
        RECT 39.130 92.150 39.430 92.600 ;
        RECT 39.130 92.000 42.980 92.150 ;
        RECT 39.130 91.550 39.430 92.000 ;
        RECT 39.130 91.400 42.980 91.550 ;
        RECT 39.130 90.950 39.430 91.400 ;
        RECT 39.130 90.800 42.980 90.950 ;
        RECT 39.130 90.350 39.430 90.800 ;
        RECT 35.530 81.450 35.680 89.650 ;
        RECT 36.130 81.450 36.280 89.650 ;
        RECT 36.730 81.450 36.880 89.650 ;
        RECT 37.330 81.450 37.480 89.650 ;
        RECT 37.930 81.450 38.080 89.650 ;
        RECT 38.530 81.450 38.680 89.650 ;
        RECT 39.130 89.200 39.430 89.650 ;
        RECT 39.130 89.050 42.980 89.200 ;
        RECT 39.130 88.600 39.430 89.050 ;
        RECT 39.130 88.450 42.980 88.600 ;
        RECT 39.130 88.000 39.430 88.450 ;
        RECT 39.130 87.850 42.980 88.000 ;
        RECT 39.130 87.400 39.430 87.850 ;
        RECT 39.130 87.250 42.980 87.400 ;
        RECT 39.130 86.800 39.430 87.250 ;
        RECT 43.830 86.800 45.630 93.200 ;
        RECT 50.030 92.750 50.330 93.200 ;
        RECT 46.480 92.600 50.330 92.750 ;
        RECT 50.030 92.150 50.330 92.600 ;
        RECT 46.480 92.000 50.330 92.150 ;
        RECT 50.030 91.550 50.330 92.000 ;
        RECT 46.480 91.400 50.330 91.550 ;
        RECT 50.030 90.950 50.330 91.400 ;
        RECT 46.480 90.800 50.330 90.950 ;
        RECT 50.030 90.350 50.330 90.800 ;
        RECT 50.780 90.350 50.930 98.550 ;
        RECT 51.380 90.350 51.530 98.550 ;
        RECT 51.980 90.350 52.130 98.550 ;
        RECT 52.580 90.350 52.730 98.550 ;
        RECT 53.180 90.350 53.330 98.550 ;
        RECT 53.780 90.350 53.930 98.550 ;
        RECT 50.030 89.200 50.330 89.650 ;
        RECT 46.480 89.050 50.330 89.200 ;
        RECT 50.030 88.600 50.330 89.050 ;
        RECT 46.480 88.450 50.330 88.600 ;
        RECT 50.030 88.000 50.330 88.450 ;
        RECT 46.480 87.850 50.330 88.000 ;
        RECT 50.030 87.400 50.330 87.850 ;
        RECT 46.480 87.250 50.330 87.400 ;
        RECT 50.030 86.800 50.330 87.250 ;
        RECT 39.130 86.650 42.980 86.800 ;
        RECT 46.480 86.650 50.330 86.800 ;
        RECT 39.130 86.200 39.430 86.650 ;
        RECT 50.030 86.200 50.330 86.650 ;
        RECT 39.130 86.050 42.980 86.200 ;
        RECT 46.480 86.050 50.330 86.200 ;
        RECT 39.130 85.600 39.430 86.050 ;
        RECT 50.030 85.600 50.330 86.050 ;
        RECT 39.130 85.450 42.980 85.600 ;
        RECT 46.480 85.450 50.330 85.600 ;
        RECT 39.130 85.000 39.430 85.450 ;
        RECT 50.030 85.000 50.330 85.450 ;
        RECT 39.130 84.850 42.980 85.000 ;
        RECT 46.480 84.850 50.330 85.000 ;
        RECT 39.130 84.400 39.430 84.850 ;
        RECT 50.030 84.400 50.330 84.850 ;
        RECT 39.130 84.250 42.980 84.400 ;
        RECT 46.480 84.250 50.330 84.400 ;
        RECT 39.130 83.800 39.430 84.250 ;
        RECT 50.030 83.800 50.330 84.250 ;
        RECT 39.130 83.650 42.980 83.800 ;
        RECT 46.480 83.650 50.330 83.800 ;
        RECT 39.130 83.200 39.430 83.650 ;
        RECT 50.030 83.200 50.330 83.650 ;
        RECT 39.130 83.050 42.980 83.200 ;
        RECT 46.480 83.050 50.330 83.200 ;
        RECT 39.130 82.600 39.430 83.050 ;
        RECT 50.030 82.600 50.330 83.050 ;
        RECT 39.130 82.450 42.980 82.600 ;
        RECT 46.480 82.450 50.330 82.600 ;
        RECT 39.130 82.000 39.430 82.450 ;
        RECT 50.030 82.000 50.330 82.450 ;
        RECT 39.130 81.450 42.930 82.000 ;
        RECT 26.530 81.400 42.930 81.450 ;
        RECT 46.530 81.450 50.330 82.000 ;
        RECT 50.780 81.450 50.930 89.650 ;
        RECT 51.380 81.450 51.530 89.650 ;
        RECT 51.980 81.450 52.130 89.650 ;
        RECT 52.580 81.450 52.730 89.650 ;
        RECT 53.180 81.450 53.330 89.650 ;
        RECT 53.780 81.450 53.930 89.650 ;
        RECT 54.380 81.450 55.080 98.550 ;
        RECT 55.530 90.350 55.680 98.550 ;
        RECT 56.130 90.350 56.280 98.550 ;
        RECT 56.730 90.350 56.880 98.550 ;
        RECT 57.330 90.350 57.480 98.550 ;
        RECT 57.930 90.350 58.080 98.550 ;
        RECT 58.530 90.350 58.680 98.550 ;
        RECT 59.130 98.000 62.930 98.550 ;
        RECT 66.530 98.550 82.930 98.600 ;
        RECT 66.530 98.000 70.330 98.550 ;
        RECT 59.130 97.550 59.430 98.000 ;
        RECT 70.030 97.550 70.330 98.000 ;
        RECT 59.130 97.400 62.980 97.550 ;
        RECT 66.480 97.400 70.330 97.550 ;
        RECT 59.130 96.950 59.430 97.400 ;
        RECT 70.030 96.950 70.330 97.400 ;
        RECT 59.130 96.800 62.980 96.950 ;
        RECT 66.480 96.800 70.330 96.950 ;
        RECT 59.130 96.350 59.430 96.800 ;
        RECT 70.030 96.350 70.330 96.800 ;
        RECT 59.130 96.200 62.980 96.350 ;
        RECT 66.480 96.200 70.330 96.350 ;
        RECT 59.130 95.750 59.430 96.200 ;
        RECT 70.030 95.750 70.330 96.200 ;
        RECT 59.130 95.600 62.980 95.750 ;
        RECT 66.480 95.600 70.330 95.750 ;
        RECT 59.130 95.150 59.430 95.600 ;
        RECT 70.030 95.150 70.330 95.600 ;
        RECT 59.130 95.000 62.980 95.150 ;
        RECT 66.480 95.000 70.330 95.150 ;
        RECT 59.130 94.550 59.430 95.000 ;
        RECT 70.030 94.550 70.330 95.000 ;
        RECT 59.130 94.400 62.980 94.550 ;
        RECT 66.480 94.400 70.330 94.550 ;
        RECT 59.130 93.950 59.430 94.400 ;
        RECT 70.030 93.950 70.330 94.400 ;
        RECT 59.130 93.800 62.980 93.950 ;
        RECT 66.480 93.800 70.330 93.950 ;
        RECT 59.130 93.350 59.430 93.800 ;
        RECT 70.030 93.350 70.330 93.800 ;
        RECT 59.130 93.200 62.980 93.350 ;
        RECT 66.480 93.200 70.330 93.350 ;
        RECT 59.130 92.750 59.430 93.200 ;
        RECT 59.130 92.600 62.980 92.750 ;
        RECT 59.130 92.150 59.430 92.600 ;
        RECT 59.130 92.000 62.980 92.150 ;
        RECT 59.130 91.550 59.430 92.000 ;
        RECT 59.130 91.400 62.980 91.550 ;
        RECT 59.130 90.950 59.430 91.400 ;
        RECT 59.130 90.800 62.980 90.950 ;
        RECT 59.130 90.350 59.430 90.800 ;
        RECT 55.530 81.450 55.680 89.650 ;
        RECT 56.130 81.450 56.280 89.650 ;
        RECT 56.730 81.450 56.880 89.650 ;
        RECT 57.330 81.450 57.480 89.650 ;
        RECT 57.930 81.450 58.080 89.650 ;
        RECT 58.530 81.450 58.680 89.650 ;
        RECT 59.130 89.200 59.430 89.650 ;
        RECT 59.130 89.050 62.980 89.200 ;
        RECT 59.130 88.600 59.430 89.050 ;
        RECT 59.130 88.450 62.980 88.600 ;
        RECT 59.130 88.000 59.430 88.450 ;
        RECT 59.130 87.850 62.980 88.000 ;
        RECT 59.130 87.400 59.430 87.850 ;
        RECT 59.130 87.250 62.980 87.400 ;
        RECT 59.130 86.800 59.430 87.250 ;
        RECT 63.830 86.800 65.630 93.200 ;
        RECT 70.030 92.750 70.330 93.200 ;
        RECT 66.480 92.600 70.330 92.750 ;
        RECT 70.030 92.150 70.330 92.600 ;
        RECT 66.480 92.000 70.330 92.150 ;
        RECT 70.030 91.550 70.330 92.000 ;
        RECT 66.480 91.400 70.330 91.550 ;
        RECT 70.030 90.950 70.330 91.400 ;
        RECT 66.480 90.800 70.330 90.950 ;
        RECT 70.030 90.350 70.330 90.800 ;
        RECT 70.780 90.350 70.930 98.550 ;
        RECT 71.380 90.350 71.530 98.550 ;
        RECT 71.980 90.350 72.130 98.550 ;
        RECT 72.580 90.350 72.730 98.550 ;
        RECT 73.180 90.350 73.330 98.550 ;
        RECT 73.780 90.350 73.930 98.550 ;
        RECT 70.030 89.200 70.330 89.650 ;
        RECT 66.480 89.050 70.330 89.200 ;
        RECT 70.030 88.600 70.330 89.050 ;
        RECT 66.480 88.450 70.330 88.600 ;
        RECT 70.030 88.000 70.330 88.450 ;
        RECT 66.480 87.850 70.330 88.000 ;
        RECT 70.030 87.400 70.330 87.850 ;
        RECT 66.480 87.250 70.330 87.400 ;
        RECT 70.030 86.800 70.330 87.250 ;
        RECT 59.130 86.650 62.980 86.800 ;
        RECT 66.480 86.650 70.330 86.800 ;
        RECT 59.130 86.200 59.430 86.650 ;
        RECT 70.030 86.200 70.330 86.650 ;
        RECT 59.130 86.050 62.980 86.200 ;
        RECT 66.480 86.050 70.330 86.200 ;
        RECT 59.130 85.600 59.430 86.050 ;
        RECT 70.030 85.600 70.330 86.050 ;
        RECT 59.130 85.450 62.980 85.600 ;
        RECT 66.480 85.450 70.330 85.600 ;
        RECT 59.130 85.000 59.430 85.450 ;
        RECT 70.030 85.000 70.330 85.450 ;
        RECT 59.130 84.850 62.980 85.000 ;
        RECT 66.480 84.850 70.330 85.000 ;
        RECT 59.130 84.400 59.430 84.850 ;
        RECT 70.030 84.400 70.330 84.850 ;
        RECT 59.130 84.250 62.980 84.400 ;
        RECT 66.480 84.250 70.330 84.400 ;
        RECT 59.130 83.800 59.430 84.250 ;
        RECT 70.030 83.800 70.330 84.250 ;
        RECT 59.130 83.650 62.980 83.800 ;
        RECT 66.480 83.650 70.330 83.800 ;
        RECT 59.130 83.200 59.430 83.650 ;
        RECT 70.030 83.200 70.330 83.650 ;
        RECT 59.130 83.050 62.980 83.200 ;
        RECT 66.480 83.050 70.330 83.200 ;
        RECT 59.130 82.600 59.430 83.050 ;
        RECT 70.030 82.600 70.330 83.050 ;
        RECT 59.130 82.450 62.980 82.600 ;
        RECT 66.480 82.450 70.330 82.600 ;
        RECT 59.130 82.000 59.430 82.450 ;
        RECT 70.030 82.000 70.330 82.450 ;
        RECT 59.130 81.450 62.930 82.000 ;
        RECT 46.530 81.400 62.930 81.450 ;
        RECT 66.530 81.450 70.330 82.000 ;
        RECT 70.780 81.450 70.930 89.650 ;
        RECT 71.380 81.450 71.530 89.650 ;
        RECT 71.980 81.450 72.130 89.650 ;
        RECT 72.580 81.450 72.730 89.650 ;
        RECT 73.180 81.450 73.330 89.650 ;
        RECT 73.780 81.450 73.930 89.650 ;
        RECT 74.380 81.450 75.080 98.550 ;
        RECT 75.530 90.350 75.680 98.550 ;
        RECT 76.130 90.350 76.280 98.550 ;
        RECT 76.730 90.350 76.880 98.550 ;
        RECT 77.330 90.350 77.480 98.550 ;
        RECT 77.930 90.350 78.080 98.550 ;
        RECT 78.530 90.350 78.680 98.550 ;
        RECT 79.130 98.000 82.930 98.550 ;
        RECT 86.530 98.550 102.930 98.600 ;
        RECT 86.530 98.000 90.330 98.550 ;
        RECT 79.130 97.550 79.430 98.000 ;
        RECT 90.030 97.550 90.330 98.000 ;
        RECT 79.130 97.400 82.980 97.550 ;
        RECT 86.480 97.400 90.330 97.550 ;
        RECT 79.130 96.950 79.430 97.400 ;
        RECT 90.030 96.950 90.330 97.400 ;
        RECT 79.130 96.800 82.980 96.950 ;
        RECT 86.480 96.800 90.330 96.950 ;
        RECT 79.130 96.350 79.430 96.800 ;
        RECT 90.030 96.350 90.330 96.800 ;
        RECT 79.130 96.200 82.980 96.350 ;
        RECT 86.480 96.200 90.330 96.350 ;
        RECT 79.130 95.750 79.430 96.200 ;
        RECT 90.030 95.750 90.330 96.200 ;
        RECT 79.130 95.600 82.980 95.750 ;
        RECT 86.480 95.600 90.330 95.750 ;
        RECT 79.130 95.150 79.430 95.600 ;
        RECT 90.030 95.150 90.330 95.600 ;
        RECT 79.130 95.000 82.980 95.150 ;
        RECT 86.480 95.000 90.330 95.150 ;
        RECT 79.130 94.550 79.430 95.000 ;
        RECT 90.030 94.550 90.330 95.000 ;
        RECT 79.130 94.400 82.980 94.550 ;
        RECT 86.480 94.400 90.330 94.550 ;
        RECT 79.130 93.950 79.430 94.400 ;
        RECT 90.030 93.950 90.330 94.400 ;
        RECT 79.130 93.800 82.980 93.950 ;
        RECT 86.480 93.800 90.330 93.950 ;
        RECT 79.130 93.350 79.430 93.800 ;
        RECT 90.030 93.350 90.330 93.800 ;
        RECT 79.130 93.200 82.980 93.350 ;
        RECT 86.480 93.200 90.330 93.350 ;
        RECT 79.130 92.750 79.430 93.200 ;
        RECT 79.130 92.600 82.980 92.750 ;
        RECT 79.130 92.150 79.430 92.600 ;
        RECT 79.130 92.000 82.980 92.150 ;
        RECT 79.130 91.550 79.430 92.000 ;
        RECT 79.130 91.400 82.980 91.550 ;
        RECT 79.130 90.950 79.430 91.400 ;
        RECT 79.130 90.800 82.980 90.950 ;
        RECT 79.130 90.350 79.430 90.800 ;
        RECT 75.530 81.450 75.680 89.650 ;
        RECT 76.130 81.450 76.280 89.650 ;
        RECT 76.730 81.450 76.880 89.650 ;
        RECT 77.330 81.450 77.480 89.650 ;
        RECT 77.930 81.450 78.080 89.650 ;
        RECT 78.530 81.450 78.680 89.650 ;
        RECT 79.130 89.200 79.430 89.650 ;
        RECT 79.130 89.050 82.980 89.200 ;
        RECT 79.130 88.600 79.430 89.050 ;
        RECT 79.130 88.450 82.980 88.600 ;
        RECT 79.130 88.000 79.430 88.450 ;
        RECT 79.130 87.850 82.980 88.000 ;
        RECT 79.130 87.400 79.430 87.850 ;
        RECT 79.130 87.250 82.980 87.400 ;
        RECT 79.130 86.800 79.430 87.250 ;
        RECT 83.830 86.800 85.630 93.200 ;
        RECT 90.030 92.750 90.330 93.200 ;
        RECT 86.480 92.600 90.330 92.750 ;
        RECT 90.030 92.150 90.330 92.600 ;
        RECT 86.480 92.000 90.330 92.150 ;
        RECT 90.030 91.550 90.330 92.000 ;
        RECT 86.480 91.400 90.330 91.550 ;
        RECT 90.030 90.950 90.330 91.400 ;
        RECT 86.480 90.800 90.330 90.950 ;
        RECT 90.030 90.350 90.330 90.800 ;
        RECT 90.780 90.350 90.930 98.550 ;
        RECT 91.380 90.350 91.530 98.550 ;
        RECT 91.980 90.350 92.130 98.550 ;
        RECT 92.580 90.350 92.730 98.550 ;
        RECT 93.180 90.350 93.330 98.550 ;
        RECT 93.780 90.350 93.930 98.550 ;
        RECT 90.030 89.200 90.330 89.650 ;
        RECT 86.480 89.050 90.330 89.200 ;
        RECT 90.030 88.600 90.330 89.050 ;
        RECT 86.480 88.450 90.330 88.600 ;
        RECT 90.030 88.000 90.330 88.450 ;
        RECT 86.480 87.850 90.330 88.000 ;
        RECT 90.030 87.400 90.330 87.850 ;
        RECT 86.480 87.250 90.330 87.400 ;
        RECT 90.030 86.800 90.330 87.250 ;
        RECT 79.130 86.650 82.980 86.800 ;
        RECT 86.480 86.650 90.330 86.800 ;
        RECT 79.130 86.200 79.430 86.650 ;
        RECT 90.030 86.200 90.330 86.650 ;
        RECT 79.130 86.050 82.980 86.200 ;
        RECT 86.480 86.050 90.330 86.200 ;
        RECT 79.130 85.600 79.430 86.050 ;
        RECT 90.030 85.600 90.330 86.050 ;
        RECT 79.130 85.450 82.980 85.600 ;
        RECT 86.480 85.450 90.330 85.600 ;
        RECT 79.130 85.000 79.430 85.450 ;
        RECT 90.030 85.000 90.330 85.450 ;
        RECT 79.130 84.850 82.980 85.000 ;
        RECT 86.480 84.850 90.330 85.000 ;
        RECT 79.130 84.400 79.430 84.850 ;
        RECT 90.030 84.400 90.330 84.850 ;
        RECT 79.130 84.250 82.980 84.400 ;
        RECT 86.480 84.250 90.330 84.400 ;
        RECT 79.130 83.800 79.430 84.250 ;
        RECT 90.030 83.800 90.330 84.250 ;
        RECT 79.130 83.650 82.980 83.800 ;
        RECT 86.480 83.650 90.330 83.800 ;
        RECT 79.130 83.200 79.430 83.650 ;
        RECT 90.030 83.200 90.330 83.650 ;
        RECT 79.130 83.050 82.980 83.200 ;
        RECT 86.480 83.050 90.330 83.200 ;
        RECT 79.130 82.600 79.430 83.050 ;
        RECT 90.030 82.600 90.330 83.050 ;
        RECT 79.130 82.450 82.980 82.600 ;
        RECT 86.480 82.450 90.330 82.600 ;
        RECT 79.130 82.000 79.430 82.450 ;
        RECT 90.030 82.000 90.330 82.450 ;
        RECT 79.130 81.450 82.930 82.000 ;
        RECT 66.530 81.400 82.930 81.450 ;
        RECT 86.530 81.450 90.330 82.000 ;
        RECT 90.780 81.450 90.930 89.650 ;
        RECT 91.380 81.450 91.530 89.650 ;
        RECT 91.980 81.450 92.130 89.650 ;
        RECT 92.580 81.450 92.730 89.650 ;
        RECT 93.180 81.450 93.330 89.650 ;
        RECT 93.780 81.450 93.930 89.650 ;
        RECT 94.380 81.450 95.080 98.550 ;
        RECT 95.530 90.350 95.680 98.550 ;
        RECT 96.130 90.350 96.280 98.550 ;
        RECT 96.730 90.350 96.880 98.550 ;
        RECT 97.330 90.350 97.480 98.550 ;
        RECT 97.930 90.350 98.080 98.550 ;
        RECT 98.530 90.350 98.680 98.550 ;
        RECT 99.130 98.000 102.930 98.550 ;
        RECT 106.530 98.550 122.930 98.600 ;
        RECT 106.530 98.000 110.330 98.550 ;
        RECT 99.130 97.550 99.430 98.000 ;
        RECT 110.030 97.550 110.330 98.000 ;
        RECT 99.130 97.400 102.980 97.550 ;
        RECT 106.480 97.400 110.330 97.550 ;
        RECT 99.130 96.950 99.430 97.400 ;
        RECT 110.030 96.950 110.330 97.400 ;
        RECT 99.130 96.800 102.980 96.950 ;
        RECT 106.480 96.800 110.330 96.950 ;
        RECT 99.130 96.350 99.430 96.800 ;
        RECT 110.030 96.350 110.330 96.800 ;
        RECT 99.130 96.200 102.980 96.350 ;
        RECT 106.480 96.200 110.330 96.350 ;
        RECT 99.130 95.750 99.430 96.200 ;
        RECT 110.030 95.750 110.330 96.200 ;
        RECT 99.130 95.600 102.980 95.750 ;
        RECT 106.480 95.600 110.330 95.750 ;
        RECT 99.130 95.150 99.430 95.600 ;
        RECT 110.030 95.150 110.330 95.600 ;
        RECT 99.130 95.000 102.980 95.150 ;
        RECT 106.480 95.000 110.330 95.150 ;
        RECT 99.130 94.550 99.430 95.000 ;
        RECT 110.030 94.550 110.330 95.000 ;
        RECT 99.130 94.400 102.980 94.550 ;
        RECT 106.480 94.400 110.330 94.550 ;
        RECT 99.130 93.950 99.430 94.400 ;
        RECT 110.030 93.950 110.330 94.400 ;
        RECT 99.130 93.800 102.980 93.950 ;
        RECT 106.480 93.800 110.330 93.950 ;
        RECT 99.130 93.350 99.430 93.800 ;
        RECT 110.030 93.350 110.330 93.800 ;
        RECT 99.130 93.200 102.980 93.350 ;
        RECT 106.480 93.200 110.330 93.350 ;
        RECT 99.130 92.750 99.430 93.200 ;
        RECT 99.130 92.600 102.980 92.750 ;
        RECT 99.130 92.150 99.430 92.600 ;
        RECT 99.130 92.000 102.980 92.150 ;
        RECT 99.130 91.550 99.430 92.000 ;
        RECT 99.130 91.400 102.980 91.550 ;
        RECT 99.130 90.950 99.430 91.400 ;
        RECT 99.130 90.800 102.980 90.950 ;
        RECT 99.130 90.350 99.430 90.800 ;
        RECT 95.530 81.450 95.680 89.650 ;
        RECT 96.130 81.450 96.280 89.650 ;
        RECT 96.730 81.450 96.880 89.650 ;
        RECT 97.330 81.450 97.480 89.650 ;
        RECT 97.930 81.450 98.080 89.650 ;
        RECT 98.530 81.450 98.680 89.650 ;
        RECT 99.130 89.200 99.430 89.650 ;
        RECT 99.130 89.050 102.980 89.200 ;
        RECT 99.130 88.600 99.430 89.050 ;
        RECT 99.130 88.450 102.980 88.600 ;
        RECT 99.130 88.000 99.430 88.450 ;
        RECT 99.130 87.850 102.980 88.000 ;
        RECT 99.130 87.400 99.430 87.850 ;
        RECT 99.130 87.250 102.980 87.400 ;
        RECT 99.130 86.800 99.430 87.250 ;
        RECT 103.830 86.800 105.630 93.200 ;
        RECT 110.030 92.750 110.330 93.200 ;
        RECT 106.480 92.600 110.330 92.750 ;
        RECT 110.030 92.150 110.330 92.600 ;
        RECT 106.480 92.000 110.330 92.150 ;
        RECT 110.030 91.550 110.330 92.000 ;
        RECT 106.480 91.400 110.330 91.550 ;
        RECT 110.030 90.950 110.330 91.400 ;
        RECT 106.480 90.800 110.330 90.950 ;
        RECT 110.030 90.350 110.330 90.800 ;
        RECT 110.780 90.350 110.930 98.550 ;
        RECT 111.380 90.350 111.530 98.550 ;
        RECT 111.980 90.350 112.130 98.550 ;
        RECT 112.580 90.350 112.730 98.550 ;
        RECT 113.180 90.350 113.330 98.550 ;
        RECT 113.780 90.350 113.930 98.550 ;
        RECT 110.030 89.200 110.330 89.650 ;
        RECT 106.480 89.050 110.330 89.200 ;
        RECT 110.030 88.600 110.330 89.050 ;
        RECT 106.480 88.450 110.330 88.600 ;
        RECT 110.030 88.000 110.330 88.450 ;
        RECT 106.480 87.850 110.330 88.000 ;
        RECT 110.030 87.400 110.330 87.850 ;
        RECT 106.480 87.250 110.330 87.400 ;
        RECT 110.030 86.800 110.330 87.250 ;
        RECT 99.130 86.650 102.980 86.800 ;
        RECT 106.480 86.650 110.330 86.800 ;
        RECT 99.130 86.200 99.430 86.650 ;
        RECT 110.030 86.200 110.330 86.650 ;
        RECT 99.130 86.050 102.980 86.200 ;
        RECT 106.480 86.050 110.330 86.200 ;
        RECT 99.130 85.600 99.430 86.050 ;
        RECT 110.030 85.600 110.330 86.050 ;
        RECT 99.130 85.450 102.980 85.600 ;
        RECT 106.480 85.450 110.330 85.600 ;
        RECT 99.130 85.000 99.430 85.450 ;
        RECT 110.030 85.000 110.330 85.450 ;
        RECT 99.130 84.850 102.980 85.000 ;
        RECT 106.480 84.850 110.330 85.000 ;
        RECT 99.130 84.400 99.430 84.850 ;
        RECT 110.030 84.400 110.330 84.850 ;
        RECT 99.130 84.250 102.980 84.400 ;
        RECT 106.480 84.250 110.330 84.400 ;
        RECT 99.130 83.800 99.430 84.250 ;
        RECT 110.030 83.800 110.330 84.250 ;
        RECT 99.130 83.650 102.980 83.800 ;
        RECT 106.480 83.650 110.330 83.800 ;
        RECT 99.130 83.200 99.430 83.650 ;
        RECT 110.030 83.200 110.330 83.650 ;
        RECT 99.130 83.050 102.980 83.200 ;
        RECT 106.480 83.050 110.330 83.200 ;
        RECT 99.130 82.600 99.430 83.050 ;
        RECT 110.030 82.600 110.330 83.050 ;
        RECT 99.130 82.450 102.980 82.600 ;
        RECT 106.480 82.450 110.330 82.600 ;
        RECT 99.130 82.000 99.430 82.450 ;
        RECT 110.030 82.000 110.330 82.450 ;
        RECT 99.130 81.450 102.930 82.000 ;
        RECT 86.530 81.400 102.930 81.450 ;
        RECT 106.530 81.450 110.330 82.000 ;
        RECT 110.780 81.450 110.930 89.650 ;
        RECT 111.380 81.450 111.530 89.650 ;
        RECT 111.980 81.450 112.130 89.650 ;
        RECT 112.580 81.450 112.730 89.650 ;
        RECT 113.180 81.450 113.330 89.650 ;
        RECT 113.780 81.450 113.930 89.650 ;
        RECT 114.380 81.450 115.080 98.550 ;
        RECT 115.530 90.350 115.680 98.550 ;
        RECT 116.130 90.350 116.280 98.550 ;
        RECT 116.730 90.350 116.880 98.550 ;
        RECT 117.330 90.350 117.480 98.550 ;
        RECT 117.930 90.350 118.080 98.550 ;
        RECT 118.530 90.350 118.680 98.550 ;
        RECT 119.130 98.000 122.930 98.550 ;
        RECT 119.130 97.550 119.430 98.000 ;
        RECT 119.130 97.400 122.980 97.550 ;
        RECT 119.130 96.950 119.430 97.400 ;
        RECT 119.130 96.800 122.980 96.950 ;
        RECT 119.130 96.350 119.430 96.800 ;
        RECT 119.130 96.200 122.980 96.350 ;
        RECT 119.130 95.750 119.430 96.200 ;
        RECT 119.130 95.600 122.980 95.750 ;
        RECT 119.130 95.150 119.430 95.600 ;
        RECT 119.130 95.000 122.980 95.150 ;
        RECT 119.130 94.550 119.430 95.000 ;
        RECT 119.130 94.400 122.980 94.550 ;
        RECT 119.130 93.950 119.430 94.400 ;
        RECT 119.130 93.800 122.980 93.950 ;
        RECT 119.130 93.350 119.430 93.800 ;
        RECT 119.130 93.200 122.980 93.350 ;
        RECT 119.130 92.750 119.430 93.200 ;
        RECT 119.130 92.600 122.980 92.750 ;
        RECT 119.130 92.150 119.430 92.600 ;
        RECT 119.130 92.000 122.980 92.150 ;
        RECT 119.130 91.550 119.430 92.000 ;
        RECT 119.130 91.400 122.980 91.550 ;
        RECT 119.130 90.950 119.430 91.400 ;
        RECT 119.130 90.800 122.980 90.950 ;
        RECT 119.130 90.350 119.430 90.800 ;
        RECT 115.530 81.450 115.680 89.650 ;
        RECT 116.130 81.450 116.280 89.650 ;
        RECT 116.730 81.450 116.880 89.650 ;
        RECT 117.330 81.450 117.480 89.650 ;
        RECT 117.930 81.450 118.080 89.650 ;
        RECT 118.530 81.450 118.680 89.650 ;
        RECT 119.130 89.200 119.430 89.650 ;
        RECT 119.130 89.050 122.980 89.200 ;
        RECT 119.130 88.600 119.430 89.050 ;
        RECT 119.130 88.450 122.980 88.600 ;
        RECT 119.130 88.000 119.430 88.450 ;
        RECT 119.130 87.850 122.980 88.000 ;
        RECT 119.130 87.400 119.430 87.850 ;
        RECT 119.130 87.250 122.980 87.400 ;
        RECT 119.130 86.800 119.430 87.250 ;
        RECT 123.830 86.800 124.730 93.200 ;
        RECT 129.850 89.755 131.850 91.030 ;
        RECT 119.130 86.650 122.980 86.800 ;
        RECT 119.130 86.200 119.430 86.650 ;
        RECT 119.130 86.050 122.980 86.200 ;
        RECT 119.130 85.600 119.430 86.050 ;
        RECT 119.130 85.450 122.980 85.600 ;
        RECT 119.130 85.000 119.430 85.450 ;
        RECT 119.130 84.850 122.980 85.000 ;
        RECT 119.130 84.400 119.430 84.850 ;
        RECT 119.130 84.250 122.980 84.400 ;
        RECT 119.130 83.800 119.430 84.250 ;
        RECT 119.130 83.650 122.980 83.800 ;
        RECT 119.130 83.200 119.430 83.650 ;
        RECT 119.130 83.050 122.980 83.200 ;
        RECT 119.130 82.600 119.430 83.050 ;
        RECT 119.130 82.450 122.980 82.600 ;
        RECT 119.130 82.000 119.430 82.450 ;
        RECT 119.130 81.450 122.930 82.000 ;
        RECT 106.530 81.400 122.930 81.450 ;
        RECT 9.630 80.900 19.830 81.400 ;
        RECT 29.630 80.900 39.830 81.400 ;
        RECT 49.630 80.900 59.830 81.400 ;
        RECT 69.630 80.900 79.830 81.400 ;
        RECT 89.630 80.900 99.830 81.400 ;
        RECT 109.630 80.900 119.830 81.400 ;
        RECT 11.530 79.100 17.930 80.900 ;
        RECT 31.530 79.100 37.930 80.900 ;
        RECT 51.530 79.100 57.930 80.900 ;
        RECT 71.530 79.100 77.930 80.900 ;
        RECT 91.530 79.100 97.930 80.900 ;
        RECT 111.530 79.100 117.930 80.900 ;
        RECT 9.630 78.600 19.830 79.100 ;
        RECT 29.630 78.600 39.830 79.100 ;
        RECT 49.630 78.600 59.830 79.100 ;
        RECT 69.630 78.600 79.830 79.100 ;
        RECT 89.630 78.600 99.830 79.100 ;
        RECT 109.630 78.600 119.830 79.100 ;
        RECT 6.530 78.550 22.930 78.600 ;
        RECT 6.530 78.000 10.330 78.550 ;
        RECT 10.030 77.550 10.330 78.000 ;
        RECT 6.480 77.400 10.330 77.550 ;
        RECT 10.030 76.950 10.330 77.400 ;
        RECT 6.480 76.800 10.330 76.950 ;
        RECT 10.030 76.350 10.330 76.800 ;
        RECT 6.480 76.200 10.330 76.350 ;
        RECT 10.030 75.750 10.330 76.200 ;
        RECT 6.480 75.600 10.330 75.750 ;
        RECT 10.030 75.150 10.330 75.600 ;
        RECT 6.480 75.000 10.330 75.150 ;
        RECT 10.030 74.550 10.330 75.000 ;
        RECT 6.480 74.400 10.330 74.550 ;
        RECT 10.030 73.950 10.330 74.400 ;
        RECT 6.480 73.800 10.330 73.950 ;
        RECT 10.030 73.350 10.330 73.800 ;
        RECT 6.480 73.200 10.330 73.350 ;
        RECT 4.730 66.800 5.630 73.200 ;
        RECT 10.030 72.750 10.330 73.200 ;
        RECT 6.480 72.600 10.330 72.750 ;
        RECT 10.030 72.150 10.330 72.600 ;
        RECT 6.480 72.000 10.330 72.150 ;
        RECT 10.030 71.550 10.330 72.000 ;
        RECT 6.480 71.400 10.330 71.550 ;
        RECT 10.030 70.950 10.330 71.400 ;
        RECT 6.480 70.800 10.330 70.950 ;
        RECT 10.030 70.350 10.330 70.800 ;
        RECT 10.780 70.350 10.930 78.550 ;
        RECT 11.380 70.350 11.530 78.550 ;
        RECT 11.980 70.350 12.130 78.550 ;
        RECT 12.580 70.350 12.730 78.550 ;
        RECT 13.180 70.350 13.330 78.550 ;
        RECT 13.780 70.350 13.930 78.550 ;
        RECT 10.030 69.200 10.330 69.650 ;
        RECT 6.480 69.050 10.330 69.200 ;
        RECT 10.030 68.600 10.330 69.050 ;
        RECT 6.480 68.450 10.330 68.600 ;
        RECT 10.030 68.000 10.330 68.450 ;
        RECT 6.480 67.850 10.330 68.000 ;
        RECT 10.030 67.400 10.330 67.850 ;
        RECT 6.480 67.250 10.330 67.400 ;
        RECT 10.030 66.800 10.330 67.250 ;
        RECT 6.480 66.650 10.330 66.800 ;
        RECT 10.030 66.200 10.330 66.650 ;
        RECT 6.480 66.050 10.330 66.200 ;
        RECT 10.030 65.600 10.330 66.050 ;
        RECT 6.480 65.450 10.330 65.600 ;
        RECT 10.030 65.000 10.330 65.450 ;
        RECT 6.480 64.850 10.330 65.000 ;
        RECT 10.030 64.400 10.330 64.850 ;
        RECT 6.480 64.250 10.330 64.400 ;
        RECT 10.030 63.800 10.330 64.250 ;
        RECT 6.480 63.650 10.330 63.800 ;
        RECT 10.030 63.200 10.330 63.650 ;
        RECT 6.480 63.050 10.330 63.200 ;
        RECT 10.030 62.600 10.330 63.050 ;
        RECT 6.480 62.450 10.330 62.600 ;
        RECT 10.030 62.000 10.330 62.450 ;
        RECT 6.530 61.450 10.330 62.000 ;
        RECT 10.780 61.450 10.930 69.650 ;
        RECT 11.380 61.450 11.530 69.650 ;
        RECT 11.980 61.450 12.130 69.650 ;
        RECT 12.580 61.450 12.730 69.650 ;
        RECT 13.180 61.450 13.330 69.650 ;
        RECT 13.780 61.450 13.930 69.650 ;
        RECT 14.380 61.450 15.080 78.550 ;
        RECT 15.530 70.350 15.680 78.550 ;
        RECT 16.130 70.350 16.280 78.550 ;
        RECT 16.730 70.350 16.880 78.550 ;
        RECT 17.330 70.350 17.480 78.550 ;
        RECT 17.930 70.350 18.080 78.550 ;
        RECT 18.530 70.350 18.680 78.550 ;
        RECT 19.130 78.000 22.930 78.550 ;
        RECT 26.530 78.550 42.930 78.600 ;
        RECT 26.530 78.000 30.330 78.550 ;
        RECT 19.130 77.550 19.430 78.000 ;
        RECT 30.030 77.550 30.330 78.000 ;
        RECT 19.130 77.400 22.980 77.550 ;
        RECT 26.480 77.400 30.330 77.550 ;
        RECT 19.130 76.950 19.430 77.400 ;
        RECT 30.030 76.950 30.330 77.400 ;
        RECT 19.130 76.800 22.980 76.950 ;
        RECT 26.480 76.800 30.330 76.950 ;
        RECT 19.130 76.350 19.430 76.800 ;
        RECT 30.030 76.350 30.330 76.800 ;
        RECT 19.130 76.200 22.980 76.350 ;
        RECT 26.480 76.200 30.330 76.350 ;
        RECT 19.130 75.750 19.430 76.200 ;
        RECT 30.030 75.750 30.330 76.200 ;
        RECT 19.130 75.600 22.980 75.750 ;
        RECT 26.480 75.600 30.330 75.750 ;
        RECT 19.130 75.150 19.430 75.600 ;
        RECT 30.030 75.150 30.330 75.600 ;
        RECT 19.130 75.000 22.980 75.150 ;
        RECT 26.480 75.000 30.330 75.150 ;
        RECT 19.130 74.550 19.430 75.000 ;
        RECT 30.030 74.550 30.330 75.000 ;
        RECT 19.130 74.400 22.980 74.550 ;
        RECT 26.480 74.400 30.330 74.550 ;
        RECT 19.130 73.950 19.430 74.400 ;
        RECT 30.030 73.950 30.330 74.400 ;
        RECT 19.130 73.800 22.980 73.950 ;
        RECT 26.480 73.800 30.330 73.950 ;
        RECT 19.130 73.350 19.430 73.800 ;
        RECT 30.030 73.350 30.330 73.800 ;
        RECT 19.130 73.200 22.980 73.350 ;
        RECT 26.480 73.200 30.330 73.350 ;
        RECT 19.130 72.750 19.430 73.200 ;
        RECT 19.130 72.600 22.980 72.750 ;
        RECT 19.130 72.150 19.430 72.600 ;
        RECT 19.130 72.000 22.980 72.150 ;
        RECT 19.130 71.550 19.430 72.000 ;
        RECT 19.130 71.400 22.980 71.550 ;
        RECT 19.130 70.950 19.430 71.400 ;
        RECT 19.130 70.800 22.980 70.950 ;
        RECT 19.130 70.350 19.430 70.800 ;
        RECT 15.530 61.450 15.680 69.650 ;
        RECT 16.130 61.450 16.280 69.650 ;
        RECT 16.730 61.450 16.880 69.650 ;
        RECT 17.330 61.450 17.480 69.650 ;
        RECT 17.930 61.450 18.080 69.650 ;
        RECT 18.530 61.450 18.680 69.650 ;
        RECT 19.130 69.200 19.430 69.650 ;
        RECT 19.130 69.050 22.980 69.200 ;
        RECT 19.130 68.600 19.430 69.050 ;
        RECT 19.130 68.450 22.980 68.600 ;
        RECT 19.130 68.000 19.430 68.450 ;
        RECT 19.130 67.850 22.980 68.000 ;
        RECT 19.130 67.400 19.430 67.850 ;
        RECT 19.130 67.250 22.980 67.400 ;
        RECT 19.130 66.800 19.430 67.250 ;
        RECT 23.830 66.800 25.630 73.200 ;
        RECT 30.030 72.750 30.330 73.200 ;
        RECT 26.480 72.600 30.330 72.750 ;
        RECT 30.030 72.150 30.330 72.600 ;
        RECT 26.480 72.000 30.330 72.150 ;
        RECT 30.030 71.550 30.330 72.000 ;
        RECT 26.480 71.400 30.330 71.550 ;
        RECT 30.030 70.950 30.330 71.400 ;
        RECT 26.480 70.800 30.330 70.950 ;
        RECT 30.030 70.350 30.330 70.800 ;
        RECT 30.780 70.350 30.930 78.550 ;
        RECT 31.380 70.350 31.530 78.550 ;
        RECT 31.980 70.350 32.130 78.550 ;
        RECT 32.580 70.350 32.730 78.550 ;
        RECT 33.180 70.350 33.330 78.550 ;
        RECT 33.780 70.350 33.930 78.550 ;
        RECT 30.030 69.200 30.330 69.650 ;
        RECT 26.480 69.050 30.330 69.200 ;
        RECT 30.030 68.600 30.330 69.050 ;
        RECT 26.480 68.450 30.330 68.600 ;
        RECT 30.030 68.000 30.330 68.450 ;
        RECT 26.480 67.850 30.330 68.000 ;
        RECT 30.030 67.400 30.330 67.850 ;
        RECT 26.480 67.250 30.330 67.400 ;
        RECT 30.030 66.800 30.330 67.250 ;
        RECT 19.130 66.650 22.980 66.800 ;
        RECT 26.480 66.650 30.330 66.800 ;
        RECT 19.130 66.200 19.430 66.650 ;
        RECT 30.030 66.200 30.330 66.650 ;
        RECT 19.130 66.050 22.980 66.200 ;
        RECT 26.480 66.050 30.330 66.200 ;
        RECT 19.130 65.600 19.430 66.050 ;
        RECT 30.030 65.600 30.330 66.050 ;
        RECT 19.130 65.450 22.980 65.600 ;
        RECT 26.480 65.450 30.330 65.600 ;
        RECT 19.130 65.000 19.430 65.450 ;
        RECT 30.030 65.000 30.330 65.450 ;
        RECT 19.130 64.850 22.980 65.000 ;
        RECT 26.480 64.850 30.330 65.000 ;
        RECT 19.130 64.400 19.430 64.850 ;
        RECT 30.030 64.400 30.330 64.850 ;
        RECT 19.130 64.250 22.980 64.400 ;
        RECT 26.480 64.250 30.330 64.400 ;
        RECT 19.130 63.800 19.430 64.250 ;
        RECT 30.030 63.800 30.330 64.250 ;
        RECT 19.130 63.650 22.980 63.800 ;
        RECT 26.480 63.650 30.330 63.800 ;
        RECT 19.130 63.200 19.430 63.650 ;
        RECT 30.030 63.200 30.330 63.650 ;
        RECT 19.130 63.050 22.980 63.200 ;
        RECT 26.480 63.050 30.330 63.200 ;
        RECT 19.130 62.600 19.430 63.050 ;
        RECT 30.030 62.600 30.330 63.050 ;
        RECT 19.130 62.450 22.980 62.600 ;
        RECT 26.480 62.450 30.330 62.600 ;
        RECT 19.130 62.000 19.430 62.450 ;
        RECT 30.030 62.000 30.330 62.450 ;
        RECT 19.130 61.450 22.930 62.000 ;
        RECT 6.530 61.400 22.930 61.450 ;
        RECT 26.530 61.450 30.330 62.000 ;
        RECT 30.780 61.450 30.930 69.650 ;
        RECT 31.380 61.450 31.530 69.650 ;
        RECT 31.980 61.450 32.130 69.650 ;
        RECT 32.580 61.450 32.730 69.650 ;
        RECT 33.180 61.450 33.330 69.650 ;
        RECT 33.780 61.450 33.930 69.650 ;
        RECT 34.380 61.450 35.080 78.550 ;
        RECT 35.530 70.350 35.680 78.550 ;
        RECT 36.130 70.350 36.280 78.550 ;
        RECT 36.730 70.350 36.880 78.550 ;
        RECT 37.330 70.350 37.480 78.550 ;
        RECT 37.930 70.350 38.080 78.550 ;
        RECT 38.530 70.350 38.680 78.550 ;
        RECT 39.130 78.000 42.930 78.550 ;
        RECT 46.530 78.550 62.930 78.600 ;
        RECT 46.530 78.000 50.330 78.550 ;
        RECT 39.130 77.550 39.430 78.000 ;
        RECT 50.030 77.550 50.330 78.000 ;
        RECT 39.130 77.400 42.980 77.550 ;
        RECT 46.480 77.400 50.330 77.550 ;
        RECT 39.130 76.950 39.430 77.400 ;
        RECT 50.030 76.950 50.330 77.400 ;
        RECT 39.130 76.800 42.980 76.950 ;
        RECT 46.480 76.800 50.330 76.950 ;
        RECT 39.130 76.350 39.430 76.800 ;
        RECT 50.030 76.350 50.330 76.800 ;
        RECT 39.130 76.200 42.980 76.350 ;
        RECT 46.480 76.200 50.330 76.350 ;
        RECT 39.130 75.750 39.430 76.200 ;
        RECT 50.030 75.750 50.330 76.200 ;
        RECT 39.130 75.600 42.980 75.750 ;
        RECT 46.480 75.600 50.330 75.750 ;
        RECT 39.130 75.150 39.430 75.600 ;
        RECT 50.030 75.150 50.330 75.600 ;
        RECT 39.130 75.000 42.980 75.150 ;
        RECT 46.480 75.000 50.330 75.150 ;
        RECT 39.130 74.550 39.430 75.000 ;
        RECT 50.030 74.550 50.330 75.000 ;
        RECT 39.130 74.400 42.980 74.550 ;
        RECT 46.480 74.400 50.330 74.550 ;
        RECT 39.130 73.950 39.430 74.400 ;
        RECT 50.030 73.950 50.330 74.400 ;
        RECT 39.130 73.800 42.980 73.950 ;
        RECT 46.480 73.800 50.330 73.950 ;
        RECT 39.130 73.350 39.430 73.800 ;
        RECT 50.030 73.350 50.330 73.800 ;
        RECT 39.130 73.200 42.980 73.350 ;
        RECT 46.480 73.200 50.330 73.350 ;
        RECT 39.130 72.750 39.430 73.200 ;
        RECT 39.130 72.600 42.980 72.750 ;
        RECT 39.130 72.150 39.430 72.600 ;
        RECT 39.130 72.000 42.980 72.150 ;
        RECT 39.130 71.550 39.430 72.000 ;
        RECT 39.130 71.400 42.980 71.550 ;
        RECT 39.130 70.950 39.430 71.400 ;
        RECT 39.130 70.800 42.980 70.950 ;
        RECT 39.130 70.350 39.430 70.800 ;
        RECT 35.530 61.450 35.680 69.650 ;
        RECT 36.130 61.450 36.280 69.650 ;
        RECT 36.730 61.450 36.880 69.650 ;
        RECT 37.330 61.450 37.480 69.650 ;
        RECT 37.930 61.450 38.080 69.650 ;
        RECT 38.530 61.450 38.680 69.650 ;
        RECT 39.130 69.200 39.430 69.650 ;
        RECT 39.130 69.050 42.980 69.200 ;
        RECT 39.130 68.600 39.430 69.050 ;
        RECT 39.130 68.450 42.980 68.600 ;
        RECT 39.130 68.000 39.430 68.450 ;
        RECT 39.130 67.850 42.980 68.000 ;
        RECT 39.130 67.400 39.430 67.850 ;
        RECT 39.130 67.250 42.980 67.400 ;
        RECT 39.130 66.800 39.430 67.250 ;
        RECT 43.830 66.800 45.630 73.200 ;
        RECT 50.030 72.750 50.330 73.200 ;
        RECT 46.480 72.600 50.330 72.750 ;
        RECT 50.030 72.150 50.330 72.600 ;
        RECT 46.480 72.000 50.330 72.150 ;
        RECT 50.030 71.550 50.330 72.000 ;
        RECT 46.480 71.400 50.330 71.550 ;
        RECT 50.030 70.950 50.330 71.400 ;
        RECT 46.480 70.800 50.330 70.950 ;
        RECT 50.030 70.350 50.330 70.800 ;
        RECT 50.780 70.350 50.930 78.550 ;
        RECT 51.380 70.350 51.530 78.550 ;
        RECT 51.980 70.350 52.130 78.550 ;
        RECT 52.580 70.350 52.730 78.550 ;
        RECT 53.180 70.350 53.330 78.550 ;
        RECT 53.780 70.350 53.930 78.550 ;
        RECT 50.030 69.200 50.330 69.650 ;
        RECT 46.480 69.050 50.330 69.200 ;
        RECT 50.030 68.600 50.330 69.050 ;
        RECT 46.480 68.450 50.330 68.600 ;
        RECT 50.030 68.000 50.330 68.450 ;
        RECT 46.480 67.850 50.330 68.000 ;
        RECT 50.030 67.400 50.330 67.850 ;
        RECT 46.480 67.250 50.330 67.400 ;
        RECT 50.030 66.800 50.330 67.250 ;
        RECT 39.130 66.650 42.980 66.800 ;
        RECT 46.480 66.650 50.330 66.800 ;
        RECT 39.130 66.200 39.430 66.650 ;
        RECT 50.030 66.200 50.330 66.650 ;
        RECT 39.130 66.050 42.980 66.200 ;
        RECT 46.480 66.050 50.330 66.200 ;
        RECT 39.130 65.600 39.430 66.050 ;
        RECT 50.030 65.600 50.330 66.050 ;
        RECT 39.130 65.450 42.980 65.600 ;
        RECT 46.480 65.450 50.330 65.600 ;
        RECT 39.130 65.000 39.430 65.450 ;
        RECT 50.030 65.000 50.330 65.450 ;
        RECT 39.130 64.850 42.980 65.000 ;
        RECT 46.480 64.850 50.330 65.000 ;
        RECT 39.130 64.400 39.430 64.850 ;
        RECT 50.030 64.400 50.330 64.850 ;
        RECT 39.130 64.250 42.980 64.400 ;
        RECT 46.480 64.250 50.330 64.400 ;
        RECT 39.130 63.800 39.430 64.250 ;
        RECT 50.030 63.800 50.330 64.250 ;
        RECT 39.130 63.650 42.980 63.800 ;
        RECT 46.480 63.650 50.330 63.800 ;
        RECT 39.130 63.200 39.430 63.650 ;
        RECT 50.030 63.200 50.330 63.650 ;
        RECT 39.130 63.050 42.980 63.200 ;
        RECT 46.480 63.050 50.330 63.200 ;
        RECT 39.130 62.600 39.430 63.050 ;
        RECT 50.030 62.600 50.330 63.050 ;
        RECT 39.130 62.450 42.980 62.600 ;
        RECT 46.480 62.450 50.330 62.600 ;
        RECT 39.130 62.000 39.430 62.450 ;
        RECT 50.030 62.000 50.330 62.450 ;
        RECT 39.130 61.450 42.930 62.000 ;
        RECT 26.530 61.400 42.930 61.450 ;
        RECT 46.530 61.450 50.330 62.000 ;
        RECT 50.780 61.450 50.930 69.650 ;
        RECT 51.380 61.450 51.530 69.650 ;
        RECT 51.980 61.450 52.130 69.650 ;
        RECT 52.580 61.450 52.730 69.650 ;
        RECT 53.180 61.450 53.330 69.650 ;
        RECT 53.780 61.450 53.930 69.650 ;
        RECT 54.380 61.450 55.080 78.550 ;
        RECT 55.530 70.350 55.680 78.550 ;
        RECT 56.130 70.350 56.280 78.550 ;
        RECT 56.730 70.350 56.880 78.550 ;
        RECT 57.330 70.350 57.480 78.550 ;
        RECT 57.930 70.350 58.080 78.550 ;
        RECT 58.530 70.350 58.680 78.550 ;
        RECT 59.130 78.000 62.930 78.550 ;
        RECT 66.530 78.550 82.930 78.600 ;
        RECT 66.530 78.000 70.330 78.550 ;
        RECT 59.130 77.550 59.430 78.000 ;
        RECT 70.030 77.550 70.330 78.000 ;
        RECT 59.130 77.400 62.980 77.550 ;
        RECT 66.480 77.400 70.330 77.550 ;
        RECT 59.130 76.950 59.430 77.400 ;
        RECT 70.030 76.950 70.330 77.400 ;
        RECT 59.130 76.800 62.980 76.950 ;
        RECT 66.480 76.800 70.330 76.950 ;
        RECT 59.130 76.350 59.430 76.800 ;
        RECT 70.030 76.350 70.330 76.800 ;
        RECT 59.130 76.200 62.980 76.350 ;
        RECT 66.480 76.200 70.330 76.350 ;
        RECT 59.130 75.750 59.430 76.200 ;
        RECT 70.030 75.750 70.330 76.200 ;
        RECT 59.130 75.600 62.980 75.750 ;
        RECT 66.480 75.600 70.330 75.750 ;
        RECT 59.130 75.150 59.430 75.600 ;
        RECT 70.030 75.150 70.330 75.600 ;
        RECT 59.130 75.000 62.980 75.150 ;
        RECT 66.480 75.000 70.330 75.150 ;
        RECT 59.130 74.550 59.430 75.000 ;
        RECT 70.030 74.550 70.330 75.000 ;
        RECT 59.130 74.400 62.980 74.550 ;
        RECT 66.480 74.400 70.330 74.550 ;
        RECT 59.130 73.950 59.430 74.400 ;
        RECT 70.030 73.950 70.330 74.400 ;
        RECT 59.130 73.800 62.980 73.950 ;
        RECT 66.480 73.800 70.330 73.950 ;
        RECT 59.130 73.350 59.430 73.800 ;
        RECT 70.030 73.350 70.330 73.800 ;
        RECT 59.130 73.200 62.980 73.350 ;
        RECT 66.480 73.200 70.330 73.350 ;
        RECT 59.130 72.750 59.430 73.200 ;
        RECT 59.130 72.600 62.980 72.750 ;
        RECT 59.130 72.150 59.430 72.600 ;
        RECT 59.130 72.000 62.980 72.150 ;
        RECT 59.130 71.550 59.430 72.000 ;
        RECT 59.130 71.400 62.980 71.550 ;
        RECT 59.130 70.950 59.430 71.400 ;
        RECT 59.130 70.800 62.980 70.950 ;
        RECT 59.130 70.350 59.430 70.800 ;
        RECT 55.530 61.450 55.680 69.650 ;
        RECT 56.130 61.450 56.280 69.650 ;
        RECT 56.730 61.450 56.880 69.650 ;
        RECT 57.330 61.450 57.480 69.650 ;
        RECT 57.930 61.450 58.080 69.650 ;
        RECT 58.530 61.450 58.680 69.650 ;
        RECT 59.130 69.200 59.430 69.650 ;
        RECT 59.130 69.050 62.980 69.200 ;
        RECT 59.130 68.600 59.430 69.050 ;
        RECT 59.130 68.450 62.980 68.600 ;
        RECT 59.130 68.000 59.430 68.450 ;
        RECT 59.130 67.850 62.980 68.000 ;
        RECT 59.130 67.400 59.430 67.850 ;
        RECT 59.130 67.250 62.980 67.400 ;
        RECT 59.130 66.800 59.430 67.250 ;
        RECT 63.830 66.800 65.630 73.200 ;
        RECT 70.030 72.750 70.330 73.200 ;
        RECT 66.480 72.600 70.330 72.750 ;
        RECT 70.030 72.150 70.330 72.600 ;
        RECT 66.480 72.000 70.330 72.150 ;
        RECT 70.030 71.550 70.330 72.000 ;
        RECT 66.480 71.400 70.330 71.550 ;
        RECT 70.030 70.950 70.330 71.400 ;
        RECT 66.480 70.800 70.330 70.950 ;
        RECT 70.030 70.350 70.330 70.800 ;
        RECT 70.780 70.350 70.930 78.550 ;
        RECT 71.380 70.350 71.530 78.550 ;
        RECT 71.980 70.350 72.130 78.550 ;
        RECT 72.580 70.350 72.730 78.550 ;
        RECT 73.180 70.350 73.330 78.550 ;
        RECT 73.780 70.350 73.930 78.550 ;
        RECT 70.030 69.200 70.330 69.650 ;
        RECT 66.480 69.050 70.330 69.200 ;
        RECT 70.030 68.600 70.330 69.050 ;
        RECT 66.480 68.450 70.330 68.600 ;
        RECT 70.030 68.000 70.330 68.450 ;
        RECT 66.480 67.850 70.330 68.000 ;
        RECT 70.030 67.400 70.330 67.850 ;
        RECT 66.480 67.250 70.330 67.400 ;
        RECT 70.030 66.800 70.330 67.250 ;
        RECT 59.130 66.650 62.980 66.800 ;
        RECT 66.480 66.650 70.330 66.800 ;
        RECT 59.130 66.200 59.430 66.650 ;
        RECT 70.030 66.200 70.330 66.650 ;
        RECT 59.130 66.050 62.980 66.200 ;
        RECT 66.480 66.050 70.330 66.200 ;
        RECT 59.130 65.600 59.430 66.050 ;
        RECT 70.030 65.600 70.330 66.050 ;
        RECT 59.130 65.450 62.980 65.600 ;
        RECT 66.480 65.450 70.330 65.600 ;
        RECT 59.130 65.000 59.430 65.450 ;
        RECT 70.030 65.000 70.330 65.450 ;
        RECT 59.130 64.850 62.980 65.000 ;
        RECT 66.480 64.850 70.330 65.000 ;
        RECT 59.130 64.400 59.430 64.850 ;
        RECT 70.030 64.400 70.330 64.850 ;
        RECT 59.130 64.250 62.980 64.400 ;
        RECT 66.480 64.250 70.330 64.400 ;
        RECT 59.130 63.800 59.430 64.250 ;
        RECT 70.030 63.800 70.330 64.250 ;
        RECT 59.130 63.650 62.980 63.800 ;
        RECT 66.480 63.650 70.330 63.800 ;
        RECT 59.130 63.200 59.430 63.650 ;
        RECT 70.030 63.200 70.330 63.650 ;
        RECT 59.130 63.050 62.980 63.200 ;
        RECT 66.480 63.050 70.330 63.200 ;
        RECT 59.130 62.600 59.430 63.050 ;
        RECT 70.030 62.600 70.330 63.050 ;
        RECT 59.130 62.450 62.980 62.600 ;
        RECT 66.480 62.450 70.330 62.600 ;
        RECT 59.130 62.000 59.430 62.450 ;
        RECT 70.030 62.000 70.330 62.450 ;
        RECT 59.130 61.450 62.930 62.000 ;
        RECT 46.530 61.400 62.930 61.450 ;
        RECT 66.530 61.450 70.330 62.000 ;
        RECT 70.780 61.450 70.930 69.650 ;
        RECT 71.380 61.450 71.530 69.650 ;
        RECT 71.980 61.450 72.130 69.650 ;
        RECT 72.580 61.450 72.730 69.650 ;
        RECT 73.180 61.450 73.330 69.650 ;
        RECT 73.780 61.450 73.930 69.650 ;
        RECT 74.380 61.450 75.080 78.550 ;
        RECT 75.530 70.350 75.680 78.550 ;
        RECT 76.130 70.350 76.280 78.550 ;
        RECT 76.730 70.350 76.880 78.550 ;
        RECT 77.330 70.350 77.480 78.550 ;
        RECT 77.930 70.350 78.080 78.550 ;
        RECT 78.530 70.350 78.680 78.550 ;
        RECT 79.130 78.000 82.930 78.550 ;
        RECT 86.530 78.550 102.930 78.600 ;
        RECT 86.530 78.000 90.330 78.550 ;
        RECT 79.130 77.550 79.430 78.000 ;
        RECT 90.030 77.550 90.330 78.000 ;
        RECT 79.130 77.400 82.980 77.550 ;
        RECT 86.480 77.400 90.330 77.550 ;
        RECT 79.130 76.950 79.430 77.400 ;
        RECT 90.030 76.950 90.330 77.400 ;
        RECT 79.130 76.800 82.980 76.950 ;
        RECT 86.480 76.800 90.330 76.950 ;
        RECT 79.130 76.350 79.430 76.800 ;
        RECT 90.030 76.350 90.330 76.800 ;
        RECT 79.130 76.200 82.980 76.350 ;
        RECT 86.480 76.200 90.330 76.350 ;
        RECT 79.130 75.750 79.430 76.200 ;
        RECT 90.030 75.750 90.330 76.200 ;
        RECT 79.130 75.600 82.980 75.750 ;
        RECT 86.480 75.600 90.330 75.750 ;
        RECT 79.130 75.150 79.430 75.600 ;
        RECT 90.030 75.150 90.330 75.600 ;
        RECT 79.130 75.000 82.980 75.150 ;
        RECT 86.480 75.000 90.330 75.150 ;
        RECT 79.130 74.550 79.430 75.000 ;
        RECT 90.030 74.550 90.330 75.000 ;
        RECT 79.130 74.400 82.980 74.550 ;
        RECT 86.480 74.400 90.330 74.550 ;
        RECT 79.130 73.950 79.430 74.400 ;
        RECT 90.030 73.950 90.330 74.400 ;
        RECT 79.130 73.800 82.980 73.950 ;
        RECT 86.480 73.800 90.330 73.950 ;
        RECT 79.130 73.350 79.430 73.800 ;
        RECT 90.030 73.350 90.330 73.800 ;
        RECT 79.130 73.200 82.980 73.350 ;
        RECT 86.480 73.200 90.330 73.350 ;
        RECT 79.130 72.750 79.430 73.200 ;
        RECT 79.130 72.600 82.980 72.750 ;
        RECT 79.130 72.150 79.430 72.600 ;
        RECT 79.130 72.000 82.980 72.150 ;
        RECT 79.130 71.550 79.430 72.000 ;
        RECT 79.130 71.400 82.980 71.550 ;
        RECT 79.130 70.950 79.430 71.400 ;
        RECT 79.130 70.800 82.980 70.950 ;
        RECT 79.130 70.350 79.430 70.800 ;
        RECT 75.530 61.450 75.680 69.650 ;
        RECT 76.130 61.450 76.280 69.650 ;
        RECT 76.730 61.450 76.880 69.650 ;
        RECT 77.330 61.450 77.480 69.650 ;
        RECT 77.930 61.450 78.080 69.650 ;
        RECT 78.530 61.450 78.680 69.650 ;
        RECT 79.130 69.200 79.430 69.650 ;
        RECT 79.130 69.050 82.980 69.200 ;
        RECT 79.130 68.600 79.430 69.050 ;
        RECT 79.130 68.450 82.980 68.600 ;
        RECT 79.130 68.000 79.430 68.450 ;
        RECT 79.130 67.850 82.980 68.000 ;
        RECT 79.130 67.400 79.430 67.850 ;
        RECT 79.130 67.250 82.980 67.400 ;
        RECT 79.130 66.800 79.430 67.250 ;
        RECT 83.830 66.800 85.630 73.200 ;
        RECT 90.030 72.750 90.330 73.200 ;
        RECT 86.480 72.600 90.330 72.750 ;
        RECT 90.030 72.150 90.330 72.600 ;
        RECT 86.480 72.000 90.330 72.150 ;
        RECT 90.030 71.550 90.330 72.000 ;
        RECT 86.480 71.400 90.330 71.550 ;
        RECT 90.030 70.950 90.330 71.400 ;
        RECT 86.480 70.800 90.330 70.950 ;
        RECT 90.030 70.350 90.330 70.800 ;
        RECT 90.780 70.350 90.930 78.550 ;
        RECT 91.380 70.350 91.530 78.550 ;
        RECT 91.980 70.350 92.130 78.550 ;
        RECT 92.580 70.350 92.730 78.550 ;
        RECT 93.180 70.350 93.330 78.550 ;
        RECT 93.780 70.350 93.930 78.550 ;
        RECT 90.030 69.200 90.330 69.650 ;
        RECT 86.480 69.050 90.330 69.200 ;
        RECT 90.030 68.600 90.330 69.050 ;
        RECT 86.480 68.450 90.330 68.600 ;
        RECT 90.030 68.000 90.330 68.450 ;
        RECT 86.480 67.850 90.330 68.000 ;
        RECT 90.030 67.400 90.330 67.850 ;
        RECT 86.480 67.250 90.330 67.400 ;
        RECT 90.030 66.800 90.330 67.250 ;
        RECT 79.130 66.650 82.980 66.800 ;
        RECT 86.480 66.650 90.330 66.800 ;
        RECT 79.130 66.200 79.430 66.650 ;
        RECT 90.030 66.200 90.330 66.650 ;
        RECT 79.130 66.050 82.980 66.200 ;
        RECT 86.480 66.050 90.330 66.200 ;
        RECT 79.130 65.600 79.430 66.050 ;
        RECT 90.030 65.600 90.330 66.050 ;
        RECT 79.130 65.450 82.980 65.600 ;
        RECT 86.480 65.450 90.330 65.600 ;
        RECT 79.130 65.000 79.430 65.450 ;
        RECT 90.030 65.000 90.330 65.450 ;
        RECT 79.130 64.850 82.980 65.000 ;
        RECT 86.480 64.850 90.330 65.000 ;
        RECT 79.130 64.400 79.430 64.850 ;
        RECT 90.030 64.400 90.330 64.850 ;
        RECT 79.130 64.250 82.980 64.400 ;
        RECT 86.480 64.250 90.330 64.400 ;
        RECT 79.130 63.800 79.430 64.250 ;
        RECT 90.030 63.800 90.330 64.250 ;
        RECT 79.130 63.650 82.980 63.800 ;
        RECT 86.480 63.650 90.330 63.800 ;
        RECT 79.130 63.200 79.430 63.650 ;
        RECT 90.030 63.200 90.330 63.650 ;
        RECT 79.130 63.050 82.980 63.200 ;
        RECT 86.480 63.050 90.330 63.200 ;
        RECT 79.130 62.600 79.430 63.050 ;
        RECT 90.030 62.600 90.330 63.050 ;
        RECT 79.130 62.450 82.980 62.600 ;
        RECT 86.480 62.450 90.330 62.600 ;
        RECT 79.130 62.000 79.430 62.450 ;
        RECT 90.030 62.000 90.330 62.450 ;
        RECT 79.130 61.450 82.930 62.000 ;
        RECT 66.530 61.400 82.930 61.450 ;
        RECT 86.530 61.450 90.330 62.000 ;
        RECT 90.780 61.450 90.930 69.650 ;
        RECT 91.380 61.450 91.530 69.650 ;
        RECT 91.980 61.450 92.130 69.650 ;
        RECT 92.580 61.450 92.730 69.650 ;
        RECT 93.180 61.450 93.330 69.650 ;
        RECT 93.780 61.450 93.930 69.650 ;
        RECT 94.380 61.450 95.080 78.550 ;
        RECT 95.530 70.350 95.680 78.550 ;
        RECT 96.130 70.350 96.280 78.550 ;
        RECT 96.730 70.350 96.880 78.550 ;
        RECT 97.330 70.350 97.480 78.550 ;
        RECT 97.930 70.350 98.080 78.550 ;
        RECT 98.530 70.350 98.680 78.550 ;
        RECT 99.130 78.000 102.930 78.550 ;
        RECT 106.530 78.550 122.930 78.600 ;
        RECT 106.530 78.000 110.330 78.550 ;
        RECT 99.130 77.550 99.430 78.000 ;
        RECT 110.030 77.550 110.330 78.000 ;
        RECT 99.130 77.400 102.980 77.550 ;
        RECT 106.480 77.400 110.330 77.550 ;
        RECT 99.130 76.950 99.430 77.400 ;
        RECT 110.030 76.950 110.330 77.400 ;
        RECT 99.130 76.800 102.980 76.950 ;
        RECT 106.480 76.800 110.330 76.950 ;
        RECT 99.130 76.350 99.430 76.800 ;
        RECT 110.030 76.350 110.330 76.800 ;
        RECT 99.130 76.200 102.980 76.350 ;
        RECT 106.480 76.200 110.330 76.350 ;
        RECT 99.130 75.750 99.430 76.200 ;
        RECT 110.030 75.750 110.330 76.200 ;
        RECT 99.130 75.600 102.980 75.750 ;
        RECT 106.480 75.600 110.330 75.750 ;
        RECT 99.130 75.150 99.430 75.600 ;
        RECT 110.030 75.150 110.330 75.600 ;
        RECT 99.130 75.000 102.980 75.150 ;
        RECT 106.480 75.000 110.330 75.150 ;
        RECT 99.130 74.550 99.430 75.000 ;
        RECT 110.030 74.550 110.330 75.000 ;
        RECT 99.130 74.400 102.980 74.550 ;
        RECT 106.480 74.400 110.330 74.550 ;
        RECT 99.130 73.950 99.430 74.400 ;
        RECT 110.030 73.950 110.330 74.400 ;
        RECT 99.130 73.800 102.980 73.950 ;
        RECT 106.480 73.800 110.330 73.950 ;
        RECT 99.130 73.350 99.430 73.800 ;
        RECT 110.030 73.350 110.330 73.800 ;
        RECT 99.130 73.200 102.980 73.350 ;
        RECT 106.480 73.200 110.330 73.350 ;
        RECT 99.130 72.750 99.430 73.200 ;
        RECT 99.130 72.600 102.980 72.750 ;
        RECT 99.130 72.150 99.430 72.600 ;
        RECT 99.130 72.000 102.980 72.150 ;
        RECT 99.130 71.550 99.430 72.000 ;
        RECT 99.130 71.400 102.980 71.550 ;
        RECT 99.130 70.950 99.430 71.400 ;
        RECT 99.130 70.800 102.980 70.950 ;
        RECT 99.130 70.350 99.430 70.800 ;
        RECT 95.530 61.450 95.680 69.650 ;
        RECT 96.130 61.450 96.280 69.650 ;
        RECT 96.730 61.450 96.880 69.650 ;
        RECT 97.330 61.450 97.480 69.650 ;
        RECT 97.930 61.450 98.080 69.650 ;
        RECT 98.530 61.450 98.680 69.650 ;
        RECT 99.130 69.200 99.430 69.650 ;
        RECT 99.130 69.050 102.980 69.200 ;
        RECT 99.130 68.600 99.430 69.050 ;
        RECT 99.130 68.450 102.980 68.600 ;
        RECT 99.130 68.000 99.430 68.450 ;
        RECT 99.130 67.850 102.980 68.000 ;
        RECT 99.130 67.400 99.430 67.850 ;
        RECT 99.130 67.250 102.980 67.400 ;
        RECT 99.130 66.800 99.430 67.250 ;
        RECT 103.830 66.800 105.630 73.200 ;
        RECT 110.030 72.750 110.330 73.200 ;
        RECT 106.480 72.600 110.330 72.750 ;
        RECT 110.030 72.150 110.330 72.600 ;
        RECT 106.480 72.000 110.330 72.150 ;
        RECT 110.030 71.550 110.330 72.000 ;
        RECT 106.480 71.400 110.330 71.550 ;
        RECT 110.030 70.950 110.330 71.400 ;
        RECT 106.480 70.800 110.330 70.950 ;
        RECT 110.030 70.350 110.330 70.800 ;
        RECT 110.780 70.350 110.930 78.550 ;
        RECT 111.380 70.350 111.530 78.550 ;
        RECT 111.980 70.350 112.130 78.550 ;
        RECT 112.580 70.350 112.730 78.550 ;
        RECT 113.180 70.350 113.330 78.550 ;
        RECT 113.780 70.350 113.930 78.550 ;
        RECT 110.030 69.200 110.330 69.650 ;
        RECT 106.480 69.050 110.330 69.200 ;
        RECT 110.030 68.600 110.330 69.050 ;
        RECT 106.480 68.450 110.330 68.600 ;
        RECT 110.030 68.000 110.330 68.450 ;
        RECT 106.480 67.850 110.330 68.000 ;
        RECT 110.030 67.400 110.330 67.850 ;
        RECT 106.480 67.250 110.330 67.400 ;
        RECT 110.030 66.800 110.330 67.250 ;
        RECT 99.130 66.650 102.980 66.800 ;
        RECT 106.480 66.650 110.330 66.800 ;
        RECT 99.130 66.200 99.430 66.650 ;
        RECT 110.030 66.200 110.330 66.650 ;
        RECT 99.130 66.050 102.980 66.200 ;
        RECT 106.480 66.050 110.330 66.200 ;
        RECT 99.130 65.600 99.430 66.050 ;
        RECT 110.030 65.600 110.330 66.050 ;
        RECT 99.130 65.450 102.980 65.600 ;
        RECT 106.480 65.450 110.330 65.600 ;
        RECT 99.130 65.000 99.430 65.450 ;
        RECT 110.030 65.000 110.330 65.450 ;
        RECT 99.130 64.850 102.980 65.000 ;
        RECT 106.480 64.850 110.330 65.000 ;
        RECT 99.130 64.400 99.430 64.850 ;
        RECT 110.030 64.400 110.330 64.850 ;
        RECT 99.130 64.250 102.980 64.400 ;
        RECT 106.480 64.250 110.330 64.400 ;
        RECT 99.130 63.800 99.430 64.250 ;
        RECT 110.030 63.800 110.330 64.250 ;
        RECT 99.130 63.650 102.980 63.800 ;
        RECT 106.480 63.650 110.330 63.800 ;
        RECT 99.130 63.200 99.430 63.650 ;
        RECT 110.030 63.200 110.330 63.650 ;
        RECT 99.130 63.050 102.980 63.200 ;
        RECT 106.480 63.050 110.330 63.200 ;
        RECT 99.130 62.600 99.430 63.050 ;
        RECT 110.030 62.600 110.330 63.050 ;
        RECT 99.130 62.450 102.980 62.600 ;
        RECT 106.480 62.450 110.330 62.600 ;
        RECT 99.130 62.000 99.430 62.450 ;
        RECT 110.030 62.000 110.330 62.450 ;
        RECT 99.130 61.450 102.930 62.000 ;
        RECT 86.530 61.400 102.930 61.450 ;
        RECT 106.530 61.450 110.330 62.000 ;
        RECT 110.780 61.450 110.930 69.650 ;
        RECT 111.380 61.450 111.530 69.650 ;
        RECT 111.980 61.450 112.130 69.650 ;
        RECT 112.580 61.450 112.730 69.650 ;
        RECT 113.180 61.450 113.330 69.650 ;
        RECT 113.780 61.450 113.930 69.650 ;
        RECT 114.380 61.450 115.080 78.550 ;
        RECT 115.530 70.350 115.680 78.550 ;
        RECT 116.130 70.350 116.280 78.550 ;
        RECT 116.730 70.350 116.880 78.550 ;
        RECT 117.330 70.350 117.480 78.550 ;
        RECT 117.930 70.350 118.080 78.550 ;
        RECT 118.530 70.350 118.680 78.550 ;
        RECT 119.130 78.000 122.930 78.550 ;
        RECT 119.130 77.550 119.430 78.000 ;
        RECT 119.130 77.400 122.980 77.550 ;
        RECT 119.130 76.950 119.430 77.400 ;
        RECT 119.130 76.800 122.980 76.950 ;
        RECT 119.130 76.350 119.430 76.800 ;
        RECT 119.130 76.200 122.980 76.350 ;
        RECT 119.130 75.750 119.430 76.200 ;
        RECT 119.130 75.600 122.980 75.750 ;
        RECT 119.130 75.150 119.430 75.600 ;
        RECT 119.130 75.000 122.980 75.150 ;
        RECT 119.130 74.550 119.430 75.000 ;
        RECT 119.130 74.400 122.980 74.550 ;
        RECT 119.130 73.950 119.430 74.400 ;
        RECT 119.130 73.800 122.980 73.950 ;
        RECT 119.130 73.350 119.430 73.800 ;
        RECT 119.130 73.200 122.980 73.350 ;
        RECT 119.130 72.750 119.430 73.200 ;
        RECT 119.130 72.600 122.980 72.750 ;
        RECT 119.130 72.150 119.430 72.600 ;
        RECT 119.130 72.000 122.980 72.150 ;
        RECT 119.130 71.550 119.430 72.000 ;
        RECT 119.130 71.400 122.980 71.550 ;
        RECT 119.130 70.950 119.430 71.400 ;
        RECT 119.130 70.800 122.980 70.950 ;
        RECT 119.130 70.350 119.430 70.800 ;
        RECT 115.530 61.450 115.680 69.650 ;
        RECT 116.130 61.450 116.280 69.650 ;
        RECT 116.730 61.450 116.880 69.650 ;
        RECT 117.330 61.450 117.480 69.650 ;
        RECT 117.930 61.450 118.080 69.650 ;
        RECT 118.530 61.450 118.680 69.650 ;
        RECT 119.130 69.200 119.430 69.650 ;
        RECT 119.130 69.050 122.980 69.200 ;
        RECT 119.130 68.600 119.430 69.050 ;
        RECT 119.130 68.450 122.980 68.600 ;
        RECT 119.130 68.000 119.430 68.450 ;
        RECT 119.130 67.850 122.980 68.000 ;
        RECT 119.130 67.400 119.430 67.850 ;
        RECT 119.130 67.250 122.980 67.400 ;
        RECT 119.130 66.800 119.430 67.250 ;
        RECT 123.830 66.800 124.730 73.200 ;
        RECT 129.850 69.220 131.850 70.495 ;
        RECT 119.130 66.650 122.980 66.800 ;
        RECT 119.130 66.200 119.430 66.650 ;
        RECT 119.130 66.050 122.980 66.200 ;
        RECT 119.130 65.600 119.430 66.050 ;
        RECT 119.130 65.450 122.980 65.600 ;
        RECT 119.130 65.000 119.430 65.450 ;
        RECT 119.130 64.850 122.980 65.000 ;
        RECT 119.130 64.400 119.430 64.850 ;
        RECT 119.130 64.250 122.980 64.400 ;
        RECT 119.130 63.800 119.430 64.250 ;
        RECT 119.130 63.650 122.980 63.800 ;
        RECT 119.130 63.200 119.430 63.650 ;
        RECT 119.130 63.050 122.980 63.200 ;
        RECT 119.130 62.600 119.430 63.050 ;
        RECT 119.130 62.450 122.980 62.600 ;
        RECT 119.130 62.000 119.430 62.450 ;
        RECT 119.130 61.450 122.930 62.000 ;
        RECT 106.530 61.400 122.930 61.450 ;
        RECT 9.630 60.900 19.830 61.400 ;
        RECT 29.630 60.900 39.830 61.400 ;
        RECT 49.630 60.900 59.830 61.400 ;
        RECT 69.630 60.900 79.830 61.400 ;
        RECT 89.630 60.900 99.830 61.400 ;
        RECT 109.630 60.900 119.830 61.400 ;
        RECT 11.530 59.100 17.930 60.900 ;
        RECT 31.530 59.100 37.930 60.900 ;
        RECT 51.530 59.100 57.930 60.900 ;
        RECT 71.530 59.100 77.930 60.900 ;
        RECT 91.530 59.100 97.930 60.900 ;
        RECT 111.530 59.100 117.930 60.900 ;
        RECT 9.630 58.600 19.830 59.100 ;
        RECT 29.630 58.600 39.830 59.100 ;
        RECT 49.630 58.600 59.830 59.100 ;
        RECT 69.630 58.600 79.830 59.100 ;
        RECT 89.630 58.600 99.830 59.100 ;
        RECT 109.630 58.600 119.830 59.100 ;
        RECT 6.530 58.550 22.930 58.600 ;
        RECT 6.530 58.000 10.330 58.550 ;
        RECT 10.030 57.550 10.330 58.000 ;
        RECT 6.480 57.400 10.330 57.550 ;
        RECT 10.030 56.950 10.330 57.400 ;
        RECT 6.480 56.800 10.330 56.950 ;
        RECT 10.030 56.350 10.330 56.800 ;
        RECT 6.480 56.200 10.330 56.350 ;
        RECT 10.030 55.750 10.330 56.200 ;
        RECT 6.480 55.600 10.330 55.750 ;
        RECT 10.030 55.150 10.330 55.600 ;
        RECT 6.480 55.000 10.330 55.150 ;
        RECT 10.030 54.550 10.330 55.000 ;
        RECT 6.480 54.400 10.330 54.550 ;
        RECT 10.030 53.950 10.330 54.400 ;
        RECT 6.480 53.800 10.330 53.950 ;
        RECT 10.030 53.350 10.330 53.800 ;
        RECT 6.480 53.200 10.330 53.350 ;
        RECT 4.730 46.800 5.630 53.200 ;
        RECT 10.030 52.750 10.330 53.200 ;
        RECT 6.480 52.600 10.330 52.750 ;
        RECT 10.030 52.150 10.330 52.600 ;
        RECT 6.480 52.000 10.330 52.150 ;
        RECT 10.030 51.550 10.330 52.000 ;
        RECT 6.480 51.400 10.330 51.550 ;
        RECT 10.030 50.950 10.330 51.400 ;
        RECT 6.480 50.800 10.330 50.950 ;
        RECT 10.030 50.350 10.330 50.800 ;
        RECT 10.780 50.350 10.930 58.550 ;
        RECT 11.380 50.350 11.530 58.550 ;
        RECT 11.980 50.350 12.130 58.550 ;
        RECT 12.580 50.350 12.730 58.550 ;
        RECT 13.180 50.350 13.330 58.550 ;
        RECT 13.780 50.350 13.930 58.550 ;
        RECT 10.030 49.200 10.330 49.650 ;
        RECT 6.480 49.050 10.330 49.200 ;
        RECT 10.030 48.600 10.330 49.050 ;
        RECT 6.480 48.450 10.330 48.600 ;
        RECT 10.030 48.000 10.330 48.450 ;
        RECT 6.480 47.850 10.330 48.000 ;
        RECT 10.030 47.400 10.330 47.850 ;
        RECT 6.480 47.250 10.330 47.400 ;
        RECT 10.030 46.800 10.330 47.250 ;
        RECT 6.480 46.650 10.330 46.800 ;
        RECT 10.030 46.200 10.330 46.650 ;
        RECT 6.480 46.050 10.330 46.200 ;
        RECT 10.030 45.600 10.330 46.050 ;
        RECT 6.480 45.450 10.330 45.600 ;
        RECT 10.030 45.000 10.330 45.450 ;
        RECT 6.480 44.850 10.330 45.000 ;
        RECT 10.030 44.400 10.330 44.850 ;
        RECT 6.480 44.250 10.330 44.400 ;
        RECT 10.030 43.800 10.330 44.250 ;
        RECT 6.480 43.650 10.330 43.800 ;
        RECT 10.030 43.200 10.330 43.650 ;
        RECT 6.480 43.050 10.330 43.200 ;
        RECT 10.030 42.600 10.330 43.050 ;
        RECT 6.480 42.450 10.330 42.600 ;
        RECT 10.030 42.000 10.330 42.450 ;
        RECT 6.530 41.450 10.330 42.000 ;
        RECT 10.780 41.450 10.930 49.650 ;
        RECT 11.380 41.450 11.530 49.650 ;
        RECT 11.980 41.450 12.130 49.650 ;
        RECT 12.580 41.450 12.730 49.650 ;
        RECT 13.180 41.450 13.330 49.650 ;
        RECT 13.780 41.450 13.930 49.650 ;
        RECT 14.380 41.450 15.080 58.550 ;
        RECT 15.530 50.350 15.680 58.550 ;
        RECT 16.130 50.350 16.280 58.550 ;
        RECT 16.730 50.350 16.880 58.550 ;
        RECT 17.330 50.350 17.480 58.550 ;
        RECT 17.930 50.350 18.080 58.550 ;
        RECT 18.530 50.350 18.680 58.550 ;
        RECT 19.130 58.000 22.930 58.550 ;
        RECT 26.530 58.550 42.930 58.600 ;
        RECT 26.530 58.000 30.330 58.550 ;
        RECT 19.130 57.550 19.430 58.000 ;
        RECT 30.030 57.550 30.330 58.000 ;
        RECT 19.130 57.400 22.980 57.550 ;
        RECT 26.480 57.400 30.330 57.550 ;
        RECT 19.130 56.950 19.430 57.400 ;
        RECT 30.030 56.950 30.330 57.400 ;
        RECT 19.130 56.800 22.980 56.950 ;
        RECT 26.480 56.800 30.330 56.950 ;
        RECT 19.130 56.350 19.430 56.800 ;
        RECT 30.030 56.350 30.330 56.800 ;
        RECT 19.130 56.200 22.980 56.350 ;
        RECT 26.480 56.200 30.330 56.350 ;
        RECT 19.130 55.750 19.430 56.200 ;
        RECT 30.030 55.750 30.330 56.200 ;
        RECT 19.130 55.600 22.980 55.750 ;
        RECT 26.480 55.600 30.330 55.750 ;
        RECT 19.130 55.150 19.430 55.600 ;
        RECT 30.030 55.150 30.330 55.600 ;
        RECT 19.130 55.000 22.980 55.150 ;
        RECT 26.480 55.000 30.330 55.150 ;
        RECT 19.130 54.550 19.430 55.000 ;
        RECT 30.030 54.550 30.330 55.000 ;
        RECT 19.130 54.400 22.980 54.550 ;
        RECT 26.480 54.400 30.330 54.550 ;
        RECT 19.130 53.950 19.430 54.400 ;
        RECT 30.030 53.950 30.330 54.400 ;
        RECT 19.130 53.800 22.980 53.950 ;
        RECT 26.480 53.800 30.330 53.950 ;
        RECT 19.130 53.350 19.430 53.800 ;
        RECT 30.030 53.350 30.330 53.800 ;
        RECT 19.130 53.200 22.980 53.350 ;
        RECT 26.480 53.200 30.330 53.350 ;
        RECT 19.130 52.750 19.430 53.200 ;
        RECT 19.130 52.600 22.980 52.750 ;
        RECT 19.130 52.150 19.430 52.600 ;
        RECT 19.130 52.000 22.980 52.150 ;
        RECT 19.130 51.550 19.430 52.000 ;
        RECT 19.130 51.400 22.980 51.550 ;
        RECT 19.130 50.950 19.430 51.400 ;
        RECT 19.130 50.800 22.980 50.950 ;
        RECT 19.130 50.350 19.430 50.800 ;
        RECT 15.530 41.450 15.680 49.650 ;
        RECT 16.130 41.450 16.280 49.650 ;
        RECT 16.730 41.450 16.880 49.650 ;
        RECT 17.330 41.450 17.480 49.650 ;
        RECT 17.930 41.450 18.080 49.650 ;
        RECT 18.530 41.450 18.680 49.650 ;
        RECT 19.130 49.200 19.430 49.650 ;
        RECT 19.130 49.050 22.980 49.200 ;
        RECT 19.130 48.600 19.430 49.050 ;
        RECT 19.130 48.450 22.980 48.600 ;
        RECT 19.130 48.000 19.430 48.450 ;
        RECT 19.130 47.850 22.980 48.000 ;
        RECT 19.130 47.400 19.430 47.850 ;
        RECT 19.130 47.250 22.980 47.400 ;
        RECT 19.130 46.800 19.430 47.250 ;
        RECT 23.830 46.800 25.630 53.200 ;
        RECT 30.030 52.750 30.330 53.200 ;
        RECT 26.480 52.600 30.330 52.750 ;
        RECT 30.030 52.150 30.330 52.600 ;
        RECT 26.480 52.000 30.330 52.150 ;
        RECT 30.030 51.550 30.330 52.000 ;
        RECT 26.480 51.400 30.330 51.550 ;
        RECT 30.030 50.950 30.330 51.400 ;
        RECT 26.480 50.800 30.330 50.950 ;
        RECT 30.030 50.350 30.330 50.800 ;
        RECT 30.780 50.350 30.930 58.550 ;
        RECT 31.380 50.350 31.530 58.550 ;
        RECT 31.980 50.350 32.130 58.550 ;
        RECT 32.580 50.350 32.730 58.550 ;
        RECT 33.180 50.350 33.330 58.550 ;
        RECT 33.780 50.350 33.930 58.550 ;
        RECT 30.030 49.200 30.330 49.650 ;
        RECT 26.480 49.050 30.330 49.200 ;
        RECT 30.030 48.600 30.330 49.050 ;
        RECT 26.480 48.450 30.330 48.600 ;
        RECT 30.030 48.000 30.330 48.450 ;
        RECT 26.480 47.850 30.330 48.000 ;
        RECT 30.030 47.400 30.330 47.850 ;
        RECT 26.480 47.250 30.330 47.400 ;
        RECT 30.030 46.800 30.330 47.250 ;
        RECT 19.130 46.650 22.980 46.800 ;
        RECT 26.480 46.650 30.330 46.800 ;
        RECT 19.130 46.200 19.430 46.650 ;
        RECT 30.030 46.200 30.330 46.650 ;
        RECT 19.130 46.050 22.980 46.200 ;
        RECT 26.480 46.050 30.330 46.200 ;
        RECT 19.130 45.600 19.430 46.050 ;
        RECT 30.030 45.600 30.330 46.050 ;
        RECT 19.130 45.450 22.980 45.600 ;
        RECT 26.480 45.450 30.330 45.600 ;
        RECT 19.130 45.000 19.430 45.450 ;
        RECT 30.030 45.000 30.330 45.450 ;
        RECT 19.130 44.850 22.980 45.000 ;
        RECT 26.480 44.850 30.330 45.000 ;
        RECT 19.130 44.400 19.430 44.850 ;
        RECT 30.030 44.400 30.330 44.850 ;
        RECT 19.130 44.250 22.980 44.400 ;
        RECT 26.480 44.250 30.330 44.400 ;
        RECT 19.130 43.800 19.430 44.250 ;
        RECT 30.030 43.800 30.330 44.250 ;
        RECT 19.130 43.650 22.980 43.800 ;
        RECT 26.480 43.650 30.330 43.800 ;
        RECT 19.130 43.200 19.430 43.650 ;
        RECT 30.030 43.200 30.330 43.650 ;
        RECT 19.130 43.050 22.980 43.200 ;
        RECT 26.480 43.050 30.330 43.200 ;
        RECT 19.130 42.600 19.430 43.050 ;
        RECT 30.030 42.600 30.330 43.050 ;
        RECT 19.130 42.450 22.980 42.600 ;
        RECT 26.480 42.450 30.330 42.600 ;
        RECT 19.130 42.000 19.430 42.450 ;
        RECT 30.030 42.000 30.330 42.450 ;
        RECT 19.130 41.450 22.930 42.000 ;
        RECT 6.530 41.400 22.930 41.450 ;
        RECT 26.530 41.450 30.330 42.000 ;
        RECT 30.780 41.450 30.930 49.650 ;
        RECT 31.380 41.450 31.530 49.650 ;
        RECT 31.980 41.450 32.130 49.650 ;
        RECT 32.580 41.450 32.730 49.650 ;
        RECT 33.180 41.450 33.330 49.650 ;
        RECT 33.780 41.450 33.930 49.650 ;
        RECT 34.380 41.450 35.080 58.550 ;
        RECT 35.530 50.350 35.680 58.550 ;
        RECT 36.130 50.350 36.280 58.550 ;
        RECT 36.730 50.350 36.880 58.550 ;
        RECT 37.330 50.350 37.480 58.550 ;
        RECT 37.930 50.350 38.080 58.550 ;
        RECT 38.530 50.350 38.680 58.550 ;
        RECT 39.130 58.000 42.930 58.550 ;
        RECT 46.530 58.550 62.930 58.600 ;
        RECT 46.530 58.000 50.330 58.550 ;
        RECT 39.130 57.550 39.430 58.000 ;
        RECT 50.030 57.550 50.330 58.000 ;
        RECT 39.130 57.400 42.980 57.550 ;
        RECT 46.480 57.400 50.330 57.550 ;
        RECT 39.130 56.950 39.430 57.400 ;
        RECT 50.030 56.950 50.330 57.400 ;
        RECT 39.130 56.800 42.980 56.950 ;
        RECT 46.480 56.800 50.330 56.950 ;
        RECT 39.130 56.350 39.430 56.800 ;
        RECT 50.030 56.350 50.330 56.800 ;
        RECT 39.130 56.200 42.980 56.350 ;
        RECT 46.480 56.200 50.330 56.350 ;
        RECT 39.130 55.750 39.430 56.200 ;
        RECT 50.030 55.750 50.330 56.200 ;
        RECT 39.130 55.600 42.980 55.750 ;
        RECT 46.480 55.600 50.330 55.750 ;
        RECT 39.130 55.150 39.430 55.600 ;
        RECT 50.030 55.150 50.330 55.600 ;
        RECT 39.130 55.000 42.980 55.150 ;
        RECT 46.480 55.000 50.330 55.150 ;
        RECT 39.130 54.550 39.430 55.000 ;
        RECT 50.030 54.550 50.330 55.000 ;
        RECT 39.130 54.400 42.980 54.550 ;
        RECT 46.480 54.400 50.330 54.550 ;
        RECT 39.130 53.950 39.430 54.400 ;
        RECT 50.030 53.950 50.330 54.400 ;
        RECT 39.130 53.800 42.980 53.950 ;
        RECT 46.480 53.800 50.330 53.950 ;
        RECT 39.130 53.350 39.430 53.800 ;
        RECT 50.030 53.350 50.330 53.800 ;
        RECT 39.130 53.200 42.980 53.350 ;
        RECT 46.480 53.200 50.330 53.350 ;
        RECT 39.130 52.750 39.430 53.200 ;
        RECT 39.130 52.600 42.980 52.750 ;
        RECT 39.130 52.150 39.430 52.600 ;
        RECT 39.130 52.000 42.980 52.150 ;
        RECT 39.130 51.550 39.430 52.000 ;
        RECT 39.130 51.400 42.980 51.550 ;
        RECT 39.130 50.950 39.430 51.400 ;
        RECT 39.130 50.800 42.980 50.950 ;
        RECT 39.130 50.350 39.430 50.800 ;
        RECT 35.530 41.450 35.680 49.650 ;
        RECT 36.130 41.450 36.280 49.650 ;
        RECT 36.730 41.450 36.880 49.650 ;
        RECT 37.330 41.450 37.480 49.650 ;
        RECT 37.930 41.450 38.080 49.650 ;
        RECT 38.530 41.450 38.680 49.650 ;
        RECT 39.130 49.200 39.430 49.650 ;
        RECT 39.130 49.050 42.980 49.200 ;
        RECT 39.130 48.600 39.430 49.050 ;
        RECT 39.130 48.450 42.980 48.600 ;
        RECT 39.130 48.000 39.430 48.450 ;
        RECT 39.130 47.850 42.980 48.000 ;
        RECT 39.130 47.400 39.430 47.850 ;
        RECT 39.130 47.250 42.980 47.400 ;
        RECT 39.130 46.800 39.430 47.250 ;
        RECT 43.830 46.800 45.630 53.200 ;
        RECT 50.030 52.750 50.330 53.200 ;
        RECT 46.480 52.600 50.330 52.750 ;
        RECT 50.030 52.150 50.330 52.600 ;
        RECT 46.480 52.000 50.330 52.150 ;
        RECT 50.030 51.550 50.330 52.000 ;
        RECT 46.480 51.400 50.330 51.550 ;
        RECT 50.030 50.950 50.330 51.400 ;
        RECT 46.480 50.800 50.330 50.950 ;
        RECT 50.030 50.350 50.330 50.800 ;
        RECT 50.780 50.350 50.930 58.550 ;
        RECT 51.380 50.350 51.530 58.550 ;
        RECT 51.980 50.350 52.130 58.550 ;
        RECT 52.580 50.350 52.730 58.550 ;
        RECT 53.180 50.350 53.330 58.550 ;
        RECT 53.780 50.350 53.930 58.550 ;
        RECT 50.030 49.200 50.330 49.650 ;
        RECT 46.480 49.050 50.330 49.200 ;
        RECT 50.030 48.600 50.330 49.050 ;
        RECT 46.480 48.450 50.330 48.600 ;
        RECT 50.030 48.000 50.330 48.450 ;
        RECT 46.480 47.850 50.330 48.000 ;
        RECT 50.030 47.400 50.330 47.850 ;
        RECT 46.480 47.250 50.330 47.400 ;
        RECT 50.030 46.800 50.330 47.250 ;
        RECT 39.130 46.650 42.980 46.800 ;
        RECT 46.480 46.650 50.330 46.800 ;
        RECT 39.130 46.200 39.430 46.650 ;
        RECT 50.030 46.200 50.330 46.650 ;
        RECT 39.130 46.050 42.980 46.200 ;
        RECT 46.480 46.050 50.330 46.200 ;
        RECT 39.130 45.600 39.430 46.050 ;
        RECT 50.030 45.600 50.330 46.050 ;
        RECT 39.130 45.450 42.980 45.600 ;
        RECT 46.480 45.450 50.330 45.600 ;
        RECT 39.130 45.000 39.430 45.450 ;
        RECT 50.030 45.000 50.330 45.450 ;
        RECT 39.130 44.850 42.980 45.000 ;
        RECT 46.480 44.850 50.330 45.000 ;
        RECT 39.130 44.400 39.430 44.850 ;
        RECT 50.030 44.400 50.330 44.850 ;
        RECT 39.130 44.250 42.980 44.400 ;
        RECT 46.480 44.250 50.330 44.400 ;
        RECT 39.130 43.800 39.430 44.250 ;
        RECT 50.030 43.800 50.330 44.250 ;
        RECT 39.130 43.650 42.980 43.800 ;
        RECT 46.480 43.650 50.330 43.800 ;
        RECT 39.130 43.200 39.430 43.650 ;
        RECT 50.030 43.200 50.330 43.650 ;
        RECT 39.130 43.050 42.980 43.200 ;
        RECT 46.480 43.050 50.330 43.200 ;
        RECT 39.130 42.600 39.430 43.050 ;
        RECT 50.030 42.600 50.330 43.050 ;
        RECT 39.130 42.450 42.980 42.600 ;
        RECT 46.480 42.450 50.330 42.600 ;
        RECT 39.130 42.000 39.430 42.450 ;
        RECT 50.030 42.000 50.330 42.450 ;
        RECT 39.130 41.450 42.930 42.000 ;
        RECT 26.530 41.400 42.930 41.450 ;
        RECT 46.530 41.450 50.330 42.000 ;
        RECT 50.780 41.450 50.930 49.650 ;
        RECT 51.380 41.450 51.530 49.650 ;
        RECT 51.980 41.450 52.130 49.650 ;
        RECT 52.580 41.450 52.730 49.650 ;
        RECT 53.180 41.450 53.330 49.650 ;
        RECT 53.780 41.450 53.930 49.650 ;
        RECT 54.380 41.450 55.080 58.550 ;
        RECT 55.530 50.350 55.680 58.550 ;
        RECT 56.130 50.350 56.280 58.550 ;
        RECT 56.730 50.350 56.880 58.550 ;
        RECT 57.330 50.350 57.480 58.550 ;
        RECT 57.930 50.350 58.080 58.550 ;
        RECT 58.530 50.350 58.680 58.550 ;
        RECT 59.130 58.000 62.930 58.550 ;
        RECT 66.530 58.550 82.930 58.600 ;
        RECT 66.530 58.000 70.330 58.550 ;
        RECT 59.130 57.550 59.430 58.000 ;
        RECT 70.030 57.550 70.330 58.000 ;
        RECT 59.130 57.400 62.980 57.550 ;
        RECT 66.480 57.400 70.330 57.550 ;
        RECT 59.130 56.950 59.430 57.400 ;
        RECT 70.030 56.950 70.330 57.400 ;
        RECT 59.130 56.800 62.980 56.950 ;
        RECT 66.480 56.800 70.330 56.950 ;
        RECT 59.130 56.350 59.430 56.800 ;
        RECT 70.030 56.350 70.330 56.800 ;
        RECT 59.130 56.200 62.980 56.350 ;
        RECT 66.480 56.200 70.330 56.350 ;
        RECT 59.130 55.750 59.430 56.200 ;
        RECT 70.030 55.750 70.330 56.200 ;
        RECT 59.130 55.600 62.980 55.750 ;
        RECT 66.480 55.600 70.330 55.750 ;
        RECT 59.130 55.150 59.430 55.600 ;
        RECT 70.030 55.150 70.330 55.600 ;
        RECT 59.130 55.000 62.980 55.150 ;
        RECT 66.480 55.000 70.330 55.150 ;
        RECT 59.130 54.550 59.430 55.000 ;
        RECT 70.030 54.550 70.330 55.000 ;
        RECT 59.130 54.400 62.980 54.550 ;
        RECT 66.480 54.400 70.330 54.550 ;
        RECT 59.130 53.950 59.430 54.400 ;
        RECT 70.030 53.950 70.330 54.400 ;
        RECT 59.130 53.800 62.980 53.950 ;
        RECT 66.480 53.800 70.330 53.950 ;
        RECT 59.130 53.350 59.430 53.800 ;
        RECT 70.030 53.350 70.330 53.800 ;
        RECT 59.130 53.200 62.980 53.350 ;
        RECT 66.480 53.200 70.330 53.350 ;
        RECT 59.130 52.750 59.430 53.200 ;
        RECT 59.130 52.600 62.980 52.750 ;
        RECT 59.130 52.150 59.430 52.600 ;
        RECT 59.130 52.000 62.980 52.150 ;
        RECT 59.130 51.550 59.430 52.000 ;
        RECT 59.130 51.400 62.980 51.550 ;
        RECT 59.130 50.950 59.430 51.400 ;
        RECT 59.130 50.800 62.980 50.950 ;
        RECT 59.130 50.350 59.430 50.800 ;
        RECT 55.530 41.450 55.680 49.650 ;
        RECT 56.130 41.450 56.280 49.650 ;
        RECT 56.730 41.450 56.880 49.650 ;
        RECT 57.330 41.450 57.480 49.650 ;
        RECT 57.930 41.450 58.080 49.650 ;
        RECT 58.530 41.450 58.680 49.650 ;
        RECT 59.130 49.200 59.430 49.650 ;
        RECT 59.130 49.050 62.980 49.200 ;
        RECT 59.130 48.600 59.430 49.050 ;
        RECT 59.130 48.450 62.980 48.600 ;
        RECT 59.130 48.000 59.430 48.450 ;
        RECT 59.130 47.850 62.980 48.000 ;
        RECT 59.130 47.400 59.430 47.850 ;
        RECT 59.130 47.250 62.980 47.400 ;
        RECT 59.130 46.800 59.430 47.250 ;
        RECT 63.830 46.800 65.630 53.200 ;
        RECT 70.030 52.750 70.330 53.200 ;
        RECT 66.480 52.600 70.330 52.750 ;
        RECT 70.030 52.150 70.330 52.600 ;
        RECT 66.480 52.000 70.330 52.150 ;
        RECT 70.030 51.550 70.330 52.000 ;
        RECT 66.480 51.400 70.330 51.550 ;
        RECT 70.030 50.950 70.330 51.400 ;
        RECT 66.480 50.800 70.330 50.950 ;
        RECT 70.030 50.350 70.330 50.800 ;
        RECT 70.780 50.350 70.930 58.550 ;
        RECT 71.380 50.350 71.530 58.550 ;
        RECT 71.980 50.350 72.130 58.550 ;
        RECT 72.580 50.350 72.730 58.550 ;
        RECT 73.180 50.350 73.330 58.550 ;
        RECT 73.780 50.350 73.930 58.550 ;
        RECT 70.030 49.200 70.330 49.650 ;
        RECT 66.480 49.050 70.330 49.200 ;
        RECT 70.030 48.600 70.330 49.050 ;
        RECT 66.480 48.450 70.330 48.600 ;
        RECT 70.030 48.000 70.330 48.450 ;
        RECT 66.480 47.850 70.330 48.000 ;
        RECT 70.030 47.400 70.330 47.850 ;
        RECT 66.480 47.250 70.330 47.400 ;
        RECT 70.030 46.800 70.330 47.250 ;
        RECT 59.130 46.650 62.980 46.800 ;
        RECT 66.480 46.650 70.330 46.800 ;
        RECT 59.130 46.200 59.430 46.650 ;
        RECT 70.030 46.200 70.330 46.650 ;
        RECT 59.130 46.050 62.980 46.200 ;
        RECT 66.480 46.050 70.330 46.200 ;
        RECT 59.130 45.600 59.430 46.050 ;
        RECT 70.030 45.600 70.330 46.050 ;
        RECT 59.130 45.450 62.980 45.600 ;
        RECT 66.480 45.450 70.330 45.600 ;
        RECT 59.130 45.000 59.430 45.450 ;
        RECT 70.030 45.000 70.330 45.450 ;
        RECT 59.130 44.850 62.980 45.000 ;
        RECT 66.480 44.850 70.330 45.000 ;
        RECT 59.130 44.400 59.430 44.850 ;
        RECT 70.030 44.400 70.330 44.850 ;
        RECT 59.130 44.250 62.980 44.400 ;
        RECT 66.480 44.250 70.330 44.400 ;
        RECT 59.130 43.800 59.430 44.250 ;
        RECT 70.030 43.800 70.330 44.250 ;
        RECT 59.130 43.650 62.980 43.800 ;
        RECT 66.480 43.650 70.330 43.800 ;
        RECT 59.130 43.200 59.430 43.650 ;
        RECT 70.030 43.200 70.330 43.650 ;
        RECT 59.130 43.050 62.980 43.200 ;
        RECT 66.480 43.050 70.330 43.200 ;
        RECT 59.130 42.600 59.430 43.050 ;
        RECT 70.030 42.600 70.330 43.050 ;
        RECT 59.130 42.450 62.980 42.600 ;
        RECT 66.480 42.450 70.330 42.600 ;
        RECT 59.130 42.000 59.430 42.450 ;
        RECT 70.030 42.000 70.330 42.450 ;
        RECT 59.130 41.450 62.930 42.000 ;
        RECT 46.530 41.400 62.930 41.450 ;
        RECT 66.530 41.450 70.330 42.000 ;
        RECT 70.780 41.450 70.930 49.650 ;
        RECT 71.380 41.450 71.530 49.650 ;
        RECT 71.980 41.450 72.130 49.650 ;
        RECT 72.580 41.450 72.730 49.650 ;
        RECT 73.180 41.450 73.330 49.650 ;
        RECT 73.780 41.450 73.930 49.650 ;
        RECT 74.380 41.450 75.080 58.550 ;
        RECT 75.530 50.350 75.680 58.550 ;
        RECT 76.130 50.350 76.280 58.550 ;
        RECT 76.730 50.350 76.880 58.550 ;
        RECT 77.330 50.350 77.480 58.550 ;
        RECT 77.930 50.350 78.080 58.550 ;
        RECT 78.530 50.350 78.680 58.550 ;
        RECT 79.130 58.000 82.930 58.550 ;
        RECT 86.530 58.550 102.930 58.600 ;
        RECT 86.530 58.000 90.330 58.550 ;
        RECT 79.130 57.550 79.430 58.000 ;
        RECT 90.030 57.550 90.330 58.000 ;
        RECT 79.130 57.400 82.980 57.550 ;
        RECT 86.480 57.400 90.330 57.550 ;
        RECT 79.130 56.950 79.430 57.400 ;
        RECT 90.030 56.950 90.330 57.400 ;
        RECT 79.130 56.800 82.980 56.950 ;
        RECT 86.480 56.800 90.330 56.950 ;
        RECT 79.130 56.350 79.430 56.800 ;
        RECT 90.030 56.350 90.330 56.800 ;
        RECT 79.130 56.200 82.980 56.350 ;
        RECT 86.480 56.200 90.330 56.350 ;
        RECT 79.130 55.750 79.430 56.200 ;
        RECT 90.030 55.750 90.330 56.200 ;
        RECT 79.130 55.600 82.980 55.750 ;
        RECT 86.480 55.600 90.330 55.750 ;
        RECT 79.130 55.150 79.430 55.600 ;
        RECT 90.030 55.150 90.330 55.600 ;
        RECT 79.130 55.000 82.980 55.150 ;
        RECT 86.480 55.000 90.330 55.150 ;
        RECT 79.130 54.550 79.430 55.000 ;
        RECT 90.030 54.550 90.330 55.000 ;
        RECT 79.130 54.400 82.980 54.550 ;
        RECT 86.480 54.400 90.330 54.550 ;
        RECT 79.130 53.950 79.430 54.400 ;
        RECT 90.030 53.950 90.330 54.400 ;
        RECT 79.130 53.800 82.980 53.950 ;
        RECT 86.480 53.800 90.330 53.950 ;
        RECT 79.130 53.350 79.430 53.800 ;
        RECT 90.030 53.350 90.330 53.800 ;
        RECT 79.130 53.200 82.980 53.350 ;
        RECT 86.480 53.200 90.330 53.350 ;
        RECT 79.130 52.750 79.430 53.200 ;
        RECT 79.130 52.600 82.980 52.750 ;
        RECT 79.130 52.150 79.430 52.600 ;
        RECT 79.130 52.000 82.980 52.150 ;
        RECT 79.130 51.550 79.430 52.000 ;
        RECT 79.130 51.400 82.980 51.550 ;
        RECT 79.130 50.950 79.430 51.400 ;
        RECT 79.130 50.800 82.980 50.950 ;
        RECT 79.130 50.350 79.430 50.800 ;
        RECT 75.530 41.450 75.680 49.650 ;
        RECT 76.130 41.450 76.280 49.650 ;
        RECT 76.730 41.450 76.880 49.650 ;
        RECT 77.330 41.450 77.480 49.650 ;
        RECT 77.930 41.450 78.080 49.650 ;
        RECT 78.530 41.450 78.680 49.650 ;
        RECT 79.130 49.200 79.430 49.650 ;
        RECT 79.130 49.050 82.980 49.200 ;
        RECT 79.130 48.600 79.430 49.050 ;
        RECT 79.130 48.450 82.980 48.600 ;
        RECT 79.130 48.000 79.430 48.450 ;
        RECT 79.130 47.850 82.980 48.000 ;
        RECT 79.130 47.400 79.430 47.850 ;
        RECT 79.130 47.250 82.980 47.400 ;
        RECT 79.130 46.800 79.430 47.250 ;
        RECT 83.830 46.800 85.630 53.200 ;
        RECT 90.030 52.750 90.330 53.200 ;
        RECT 86.480 52.600 90.330 52.750 ;
        RECT 90.030 52.150 90.330 52.600 ;
        RECT 86.480 52.000 90.330 52.150 ;
        RECT 90.030 51.550 90.330 52.000 ;
        RECT 86.480 51.400 90.330 51.550 ;
        RECT 90.030 50.950 90.330 51.400 ;
        RECT 86.480 50.800 90.330 50.950 ;
        RECT 90.030 50.350 90.330 50.800 ;
        RECT 90.780 50.350 90.930 58.550 ;
        RECT 91.380 50.350 91.530 58.550 ;
        RECT 91.980 50.350 92.130 58.550 ;
        RECT 92.580 50.350 92.730 58.550 ;
        RECT 93.180 50.350 93.330 58.550 ;
        RECT 93.780 50.350 93.930 58.550 ;
        RECT 90.030 49.200 90.330 49.650 ;
        RECT 86.480 49.050 90.330 49.200 ;
        RECT 90.030 48.600 90.330 49.050 ;
        RECT 86.480 48.450 90.330 48.600 ;
        RECT 90.030 48.000 90.330 48.450 ;
        RECT 86.480 47.850 90.330 48.000 ;
        RECT 90.030 47.400 90.330 47.850 ;
        RECT 86.480 47.250 90.330 47.400 ;
        RECT 90.030 46.800 90.330 47.250 ;
        RECT 79.130 46.650 82.980 46.800 ;
        RECT 86.480 46.650 90.330 46.800 ;
        RECT 79.130 46.200 79.430 46.650 ;
        RECT 90.030 46.200 90.330 46.650 ;
        RECT 79.130 46.050 82.980 46.200 ;
        RECT 86.480 46.050 90.330 46.200 ;
        RECT 79.130 45.600 79.430 46.050 ;
        RECT 90.030 45.600 90.330 46.050 ;
        RECT 79.130 45.450 82.980 45.600 ;
        RECT 86.480 45.450 90.330 45.600 ;
        RECT 79.130 45.000 79.430 45.450 ;
        RECT 90.030 45.000 90.330 45.450 ;
        RECT 79.130 44.850 82.980 45.000 ;
        RECT 86.480 44.850 90.330 45.000 ;
        RECT 79.130 44.400 79.430 44.850 ;
        RECT 90.030 44.400 90.330 44.850 ;
        RECT 79.130 44.250 82.980 44.400 ;
        RECT 86.480 44.250 90.330 44.400 ;
        RECT 79.130 43.800 79.430 44.250 ;
        RECT 90.030 43.800 90.330 44.250 ;
        RECT 79.130 43.650 82.980 43.800 ;
        RECT 86.480 43.650 90.330 43.800 ;
        RECT 79.130 43.200 79.430 43.650 ;
        RECT 90.030 43.200 90.330 43.650 ;
        RECT 79.130 43.050 82.980 43.200 ;
        RECT 86.480 43.050 90.330 43.200 ;
        RECT 79.130 42.600 79.430 43.050 ;
        RECT 90.030 42.600 90.330 43.050 ;
        RECT 79.130 42.450 82.980 42.600 ;
        RECT 86.480 42.450 90.330 42.600 ;
        RECT 79.130 42.000 79.430 42.450 ;
        RECT 90.030 42.000 90.330 42.450 ;
        RECT 79.130 41.450 82.930 42.000 ;
        RECT 66.530 41.400 82.930 41.450 ;
        RECT 86.530 41.450 90.330 42.000 ;
        RECT 90.780 41.450 90.930 49.650 ;
        RECT 91.380 41.450 91.530 49.650 ;
        RECT 91.980 41.450 92.130 49.650 ;
        RECT 92.580 41.450 92.730 49.650 ;
        RECT 93.180 41.450 93.330 49.650 ;
        RECT 93.780 41.450 93.930 49.650 ;
        RECT 94.380 41.450 95.080 58.550 ;
        RECT 95.530 50.350 95.680 58.550 ;
        RECT 96.130 50.350 96.280 58.550 ;
        RECT 96.730 50.350 96.880 58.550 ;
        RECT 97.330 50.350 97.480 58.550 ;
        RECT 97.930 50.350 98.080 58.550 ;
        RECT 98.530 50.350 98.680 58.550 ;
        RECT 99.130 58.000 102.930 58.550 ;
        RECT 106.530 58.550 122.930 58.600 ;
        RECT 106.530 58.000 110.330 58.550 ;
        RECT 99.130 57.550 99.430 58.000 ;
        RECT 110.030 57.550 110.330 58.000 ;
        RECT 99.130 57.400 102.980 57.550 ;
        RECT 106.480 57.400 110.330 57.550 ;
        RECT 99.130 56.950 99.430 57.400 ;
        RECT 110.030 56.950 110.330 57.400 ;
        RECT 99.130 56.800 102.980 56.950 ;
        RECT 106.480 56.800 110.330 56.950 ;
        RECT 99.130 56.350 99.430 56.800 ;
        RECT 110.030 56.350 110.330 56.800 ;
        RECT 99.130 56.200 102.980 56.350 ;
        RECT 106.480 56.200 110.330 56.350 ;
        RECT 99.130 55.750 99.430 56.200 ;
        RECT 110.030 55.750 110.330 56.200 ;
        RECT 99.130 55.600 102.980 55.750 ;
        RECT 106.480 55.600 110.330 55.750 ;
        RECT 99.130 55.150 99.430 55.600 ;
        RECT 110.030 55.150 110.330 55.600 ;
        RECT 99.130 55.000 102.980 55.150 ;
        RECT 106.480 55.000 110.330 55.150 ;
        RECT 99.130 54.550 99.430 55.000 ;
        RECT 110.030 54.550 110.330 55.000 ;
        RECT 99.130 54.400 102.980 54.550 ;
        RECT 106.480 54.400 110.330 54.550 ;
        RECT 99.130 53.950 99.430 54.400 ;
        RECT 110.030 53.950 110.330 54.400 ;
        RECT 99.130 53.800 102.980 53.950 ;
        RECT 106.480 53.800 110.330 53.950 ;
        RECT 99.130 53.350 99.430 53.800 ;
        RECT 110.030 53.350 110.330 53.800 ;
        RECT 99.130 53.200 102.980 53.350 ;
        RECT 106.480 53.200 110.330 53.350 ;
        RECT 99.130 52.750 99.430 53.200 ;
        RECT 99.130 52.600 102.980 52.750 ;
        RECT 99.130 52.150 99.430 52.600 ;
        RECT 99.130 52.000 102.980 52.150 ;
        RECT 99.130 51.550 99.430 52.000 ;
        RECT 99.130 51.400 102.980 51.550 ;
        RECT 99.130 50.950 99.430 51.400 ;
        RECT 99.130 50.800 102.980 50.950 ;
        RECT 99.130 50.350 99.430 50.800 ;
        RECT 95.530 41.450 95.680 49.650 ;
        RECT 96.130 41.450 96.280 49.650 ;
        RECT 96.730 41.450 96.880 49.650 ;
        RECT 97.330 41.450 97.480 49.650 ;
        RECT 97.930 41.450 98.080 49.650 ;
        RECT 98.530 41.450 98.680 49.650 ;
        RECT 99.130 49.200 99.430 49.650 ;
        RECT 99.130 49.050 102.980 49.200 ;
        RECT 99.130 48.600 99.430 49.050 ;
        RECT 99.130 48.450 102.980 48.600 ;
        RECT 99.130 48.000 99.430 48.450 ;
        RECT 99.130 47.850 102.980 48.000 ;
        RECT 99.130 47.400 99.430 47.850 ;
        RECT 99.130 47.250 102.980 47.400 ;
        RECT 99.130 46.800 99.430 47.250 ;
        RECT 103.830 46.800 105.630 53.200 ;
        RECT 110.030 52.750 110.330 53.200 ;
        RECT 106.480 52.600 110.330 52.750 ;
        RECT 110.030 52.150 110.330 52.600 ;
        RECT 106.480 52.000 110.330 52.150 ;
        RECT 110.030 51.550 110.330 52.000 ;
        RECT 106.480 51.400 110.330 51.550 ;
        RECT 110.030 50.950 110.330 51.400 ;
        RECT 106.480 50.800 110.330 50.950 ;
        RECT 110.030 50.350 110.330 50.800 ;
        RECT 110.780 50.350 110.930 58.550 ;
        RECT 111.380 50.350 111.530 58.550 ;
        RECT 111.980 50.350 112.130 58.550 ;
        RECT 112.580 50.350 112.730 58.550 ;
        RECT 113.180 50.350 113.330 58.550 ;
        RECT 113.780 50.350 113.930 58.550 ;
        RECT 110.030 49.200 110.330 49.650 ;
        RECT 106.480 49.050 110.330 49.200 ;
        RECT 110.030 48.600 110.330 49.050 ;
        RECT 106.480 48.450 110.330 48.600 ;
        RECT 110.030 48.000 110.330 48.450 ;
        RECT 106.480 47.850 110.330 48.000 ;
        RECT 110.030 47.400 110.330 47.850 ;
        RECT 106.480 47.250 110.330 47.400 ;
        RECT 110.030 46.800 110.330 47.250 ;
        RECT 99.130 46.650 102.980 46.800 ;
        RECT 106.480 46.650 110.330 46.800 ;
        RECT 99.130 46.200 99.430 46.650 ;
        RECT 110.030 46.200 110.330 46.650 ;
        RECT 99.130 46.050 102.980 46.200 ;
        RECT 106.480 46.050 110.330 46.200 ;
        RECT 99.130 45.600 99.430 46.050 ;
        RECT 110.030 45.600 110.330 46.050 ;
        RECT 99.130 45.450 102.980 45.600 ;
        RECT 106.480 45.450 110.330 45.600 ;
        RECT 99.130 45.000 99.430 45.450 ;
        RECT 110.030 45.000 110.330 45.450 ;
        RECT 99.130 44.850 102.980 45.000 ;
        RECT 106.480 44.850 110.330 45.000 ;
        RECT 99.130 44.400 99.430 44.850 ;
        RECT 110.030 44.400 110.330 44.850 ;
        RECT 99.130 44.250 102.980 44.400 ;
        RECT 106.480 44.250 110.330 44.400 ;
        RECT 99.130 43.800 99.430 44.250 ;
        RECT 110.030 43.800 110.330 44.250 ;
        RECT 99.130 43.650 102.980 43.800 ;
        RECT 106.480 43.650 110.330 43.800 ;
        RECT 99.130 43.200 99.430 43.650 ;
        RECT 110.030 43.200 110.330 43.650 ;
        RECT 99.130 43.050 102.980 43.200 ;
        RECT 106.480 43.050 110.330 43.200 ;
        RECT 99.130 42.600 99.430 43.050 ;
        RECT 110.030 42.600 110.330 43.050 ;
        RECT 99.130 42.450 102.980 42.600 ;
        RECT 106.480 42.450 110.330 42.600 ;
        RECT 99.130 42.000 99.430 42.450 ;
        RECT 110.030 42.000 110.330 42.450 ;
        RECT 99.130 41.450 102.930 42.000 ;
        RECT 86.530 41.400 102.930 41.450 ;
        RECT 106.530 41.450 110.330 42.000 ;
        RECT 110.780 41.450 110.930 49.650 ;
        RECT 111.380 41.450 111.530 49.650 ;
        RECT 111.980 41.450 112.130 49.650 ;
        RECT 112.580 41.450 112.730 49.650 ;
        RECT 113.180 41.450 113.330 49.650 ;
        RECT 113.780 41.450 113.930 49.650 ;
        RECT 114.380 41.450 115.080 58.550 ;
        RECT 115.530 50.350 115.680 58.550 ;
        RECT 116.130 50.350 116.280 58.550 ;
        RECT 116.730 50.350 116.880 58.550 ;
        RECT 117.330 50.350 117.480 58.550 ;
        RECT 117.930 50.350 118.080 58.550 ;
        RECT 118.530 50.350 118.680 58.550 ;
        RECT 119.130 58.000 122.930 58.550 ;
        RECT 119.130 57.550 119.430 58.000 ;
        RECT 119.130 57.400 122.980 57.550 ;
        RECT 119.130 56.950 119.430 57.400 ;
        RECT 119.130 56.800 122.980 56.950 ;
        RECT 119.130 56.350 119.430 56.800 ;
        RECT 119.130 56.200 122.980 56.350 ;
        RECT 119.130 55.750 119.430 56.200 ;
        RECT 119.130 55.600 122.980 55.750 ;
        RECT 119.130 55.150 119.430 55.600 ;
        RECT 119.130 55.000 122.980 55.150 ;
        RECT 119.130 54.550 119.430 55.000 ;
        RECT 119.130 54.400 122.980 54.550 ;
        RECT 119.130 53.950 119.430 54.400 ;
        RECT 119.130 53.800 122.980 53.950 ;
        RECT 119.130 53.350 119.430 53.800 ;
        RECT 119.130 53.200 122.980 53.350 ;
        RECT 119.130 52.750 119.430 53.200 ;
        RECT 119.130 52.600 122.980 52.750 ;
        RECT 119.130 52.150 119.430 52.600 ;
        RECT 119.130 52.000 122.980 52.150 ;
        RECT 119.130 51.550 119.430 52.000 ;
        RECT 119.130 51.400 122.980 51.550 ;
        RECT 119.130 50.950 119.430 51.400 ;
        RECT 119.130 50.800 122.980 50.950 ;
        RECT 119.130 50.350 119.430 50.800 ;
        RECT 115.530 41.450 115.680 49.650 ;
        RECT 116.130 41.450 116.280 49.650 ;
        RECT 116.730 41.450 116.880 49.650 ;
        RECT 117.330 41.450 117.480 49.650 ;
        RECT 117.930 41.450 118.080 49.650 ;
        RECT 118.530 41.450 118.680 49.650 ;
        RECT 119.130 49.200 119.430 49.650 ;
        RECT 119.130 49.050 122.980 49.200 ;
        RECT 119.130 48.600 119.430 49.050 ;
        RECT 119.130 48.450 122.980 48.600 ;
        RECT 119.130 48.000 119.430 48.450 ;
        RECT 119.130 47.850 122.980 48.000 ;
        RECT 119.130 47.400 119.430 47.850 ;
        RECT 119.130 47.250 122.980 47.400 ;
        RECT 119.130 46.800 119.430 47.250 ;
        RECT 123.830 46.800 124.730 53.200 ;
        RECT 129.850 50.130 131.850 51.405 ;
        RECT 119.130 46.650 122.980 46.800 ;
        RECT 119.130 46.200 119.430 46.650 ;
        RECT 119.130 46.050 122.980 46.200 ;
        RECT 119.130 45.600 119.430 46.050 ;
        RECT 119.130 45.450 122.980 45.600 ;
        RECT 119.130 45.000 119.430 45.450 ;
        RECT 119.130 44.850 122.980 45.000 ;
        RECT 119.130 44.400 119.430 44.850 ;
        RECT 119.130 44.250 122.980 44.400 ;
        RECT 119.130 43.800 119.430 44.250 ;
        RECT 119.130 43.650 122.980 43.800 ;
        RECT 119.130 43.200 119.430 43.650 ;
        RECT 119.130 43.050 122.980 43.200 ;
        RECT 119.130 42.600 119.430 43.050 ;
        RECT 119.130 42.450 122.980 42.600 ;
        RECT 119.130 42.000 119.430 42.450 ;
        RECT 119.130 41.450 122.930 42.000 ;
        RECT 106.530 41.400 122.930 41.450 ;
        RECT 9.630 40.900 19.830 41.400 ;
        RECT 29.630 40.900 39.830 41.400 ;
        RECT 49.630 40.900 59.830 41.400 ;
        RECT 69.630 40.900 79.830 41.400 ;
        RECT 89.630 40.900 99.830 41.400 ;
        RECT 109.630 40.900 119.830 41.400 ;
        RECT 11.530 39.100 17.930 40.900 ;
        RECT 31.530 39.100 37.930 40.900 ;
        RECT 51.530 39.100 57.930 40.900 ;
        RECT 71.530 39.100 77.930 40.900 ;
        RECT 91.530 39.100 97.930 40.900 ;
        RECT 111.530 39.100 117.930 40.900 ;
        RECT 9.630 38.600 19.830 39.100 ;
        RECT 29.630 38.600 39.830 39.100 ;
        RECT 49.630 38.600 59.830 39.100 ;
        RECT 69.630 38.600 79.830 39.100 ;
        RECT 89.630 38.600 99.830 39.100 ;
        RECT 109.630 38.600 119.830 39.100 ;
        RECT 6.530 38.550 22.930 38.600 ;
        RECT 6.530 38.000 10.330 38.550 ;
        RECT 10.030 37.550 10.330 38.000 ;
        RECT 6.480 37.400 10.330 37.550 ;
        RECT 10.030 36.950 10.330 37.400 ;
        RECT 6.480 36.800 10.330 36.950 ;
        RECT 10.030 36.350 10.330 36.800 ;
        RECT 6.480 36.200 10.330 36.350 ;
        RECT 10.030 35.750 10.330 36.200 ;
        RECT 6.480 35.600 10.330 35.750 ;
        RECT 10.030 35.150 10.330 35.600 ;
        RECT 6.480 35.000 10.330 35.150 ;
        RECT 10.030 34.550 10.330 35.000 ;
        RECT 6.480 34.400 10.330 34.550 ;
        RECT 10.030 33.950 10.330 34.400 ;
        RECT 6.480 33.800 10.330 33.950 ;
        RECT 10.030 33.350 10.330 33.800 ;
        RECT 6.480 33.200 10.330 33.350 ;
        RECT 4.730 26.800 5.630 33.200 ;
        RECT 10.030 32.750 10.330 33.200 ;
        RECT 6.480 32.600 10.330 32.750 ;
        RECT 10.030 32.150 10.330 32.600 ;
        RECT 6.480 32.000 10.330 32.150 ;
        RECT 10.030 31.550 10.330 32.000 ;
        RECT 6.480 31.400 10.330 31.550 ;
        RECT 10.030 30.950 10.330 31.400 ;
        RECT 6.480 30.800 10.330 30.950 ;
        RECT 10.030 30.350 10.330 30.800 ;
        RECT 10.780 30.350 10.930 38.550 ;
        RECT 11.380 30.350 11.530 38.550 ;
        RECT 11.980 30.350 12.130 38.550 ;
        RECT 12.580 30.350 12.730 38.550 ;
        RECT 13.180 30.350 13.330 38.550 ;
        RECT 13.780 30.350 13.930 38.550 ;
        RECT 10.030 29.200 10.330 29.650 ;
        RECT 6.480 29.050 10.330 29.200 ;
        RECT 10.030 28.600 10.330 29.050 ;
        RECT 6.480 28.450 10.330 28.600 ;
        RECT 10.030 28.000 10.330 28.450 ;
        RECT 6.480 27.850 10.330 28.000 ;
        RECT 10.030 27.400 10.330 27.850 ;
        RECT 6.480 27.250 10.330 27.400 ;
        RECT 10.030 26.800 10.330 27.250 ;
        RECT 6.480 26.650 10.330 26.800 ;
        RECT 10.030 26.200 10.330 26.650 ;
        RECT 6.480 26.050 10.330 26.200 ;
        RECT 10.030 25.600 10.330 26.050 ;
        RECT 6.480 25.450 10.330 25.600 ;
        RECT 10.030 25.000 10.330 25.450 ;
        RECT 6.480 24.850 10.330 25.000 ;
        RECT 10.030 24.400 10.330 24.850 ;
        RECT 6.480 24.250 10.330 24.400 ;
        RECT 10.030 23.800 10.330 24.250 ;
        RECT 6.480 23.650 10.330 23.800 ;
        RECT 10.030 23.200 10.330 23.650 ;
        RECT 6.480 23.050 10.330 23.200 ;
        RECT 10.030 22.600 10.330 23.050 ;
        RECT 6.480 22.450 10.330 22.600 ;
        RECT 10.030 22.000 10.330 22.450 ;
        RECT 6.530 21.450 10.330 22.000 ;
        RECT 10.780 21.450 10.930 29.650 ;
        RECT 11.380 21.450 11.530 29.650 ;
        RECT 11.980 21.450 12.130 29.650 ;
        RECT 12.580 21.450 12.730 29.650 ;
        RECT 13.180 21.450 13.330 29.650 ;
        RECT 13.780 21.450 13.930 29.650 ;
        RECT 14.380 21.450 15.080 38.550 ;
        RECT 15.530 30.350 15.680 38.550 ;
        RECT 16.130 30.350 16.280 38.550 ;
        RECT 16.730 30.350 16.880 38.550 ;
        RECT 17.330 30.350 17.480 38.550 ;
        RECT 17.930 30.350 18.080 38.550 ;
        RECT 18.530 30.350 18.680 38.550 ;
        RECT 19.130 38.000 22.930 38.550 ;
        RECT 26.530 38.550 42.930 38.600 ;
        RECT 26.530 38.000 30.330 38.550 ;
        RECT 19.130 37.550 19.430 38.000 ;
        RECT 30.030 37.550 30.330 38.000 ;
        RECT 19.130 37.400 22.980 37.550 ;
        RECT 26.480 37.400 30.330 37.550 ;
        RECT 19.130 36.950 19.430 37.400 ;
        RECT 30.030 36.950 30.330 37.400 ;
        RECT 19.130 36.800 22.980 36.950 ;
        RECT 26.480 36.800 30.330 36.950 ;
        RECT 19.130 36.350 19.430 36.800 ;
        RECT 30.030 36.350 30.330 36.800 ;
        RECT 19.130 36.200 22.980 36.350 ;
        RECT 26.480 36.200 30.330 36.350 ;
        RECT 19.130 35.750 19.430 36.200 ;
        RECT 30.030 35.750 30.330 36.200 ;
        RECT 19.130 35.600 22.980 35.750 ;
        RECT 26.480 35.600 30.330 35.750 ;
        RECT 19.130 35.150 19.430 35.600 ;
        RECT 30.030 35.150 30.330 35.600 ;
        RECT 19.130 35.000 22.980 35.150 ;
        RECT 26.480 35.000 30.330 35.150 ;
        RECT 19.130 34.550 19.430 35.000 ;
        RECT 30.030 34.550 30.330 35.000 ;
        RECT 19.130 34.400 22.980 34.550 ;
        RECT 26.480 34.400 30.330 34.550 ;
        RECT 19.130 33.950 19.430 34.400 ;
        RECT 30.030 33.950 30.330 34.400 ;
        RECT 19.130 33.800 22.980 33.950 ;
        RECT 26.480 33.800 30.330 33.950 ;
        RECT 19.130 33.350 19.430 33.800 ;
        RECT 30.030 33.350 30.330 33.800 ;
        RECT 19.130 33.200 22.980 33.350 ;
        RECT 26.480 33.200 30.330 33.350 ;
        RECT 19.130 32.750 19.430 33.200 ;
        RECT 19.130 32.600 22.980 32.750 ;
        RECT 19.130 32.150 19.430 32.600 ;
        RECT 19.130 32.000 22.980 32.150 ;
        RECT 19.130 31.550 19.430 32.000 ;
        RECT 19.130 31.400 22.980 31.550 ;
        RECT 19.130 30.950 19.430 31.400 ;
        RECT 19.130 30.800 22.980 30.950 ;
        RECT 19.130 30.350 19.430 30.800 ;
        RECT 15.530 21.450 15.680 29.650 ;
        RECT 16.130 21.450 16.280 29.650 ;
        RECT 16.730 21.450 16.880 29.650 ;
        RECT 17.330 21.450 17.480 29.650 ;
        RECT 17.930 21.450 18.080 29.650 ;
        RECT 18.530 21.450 18.680 29.650 ;
        RECT 19.130 29.200 19.430 29.650 ;
        RECT 19.130 29.050 22.980 29.200 ;
        RECT 19.130 28.600 19.430 29.050 ;
        RECT 19.130 28.450 22.980 28.600 ;
        RECT 19.130 28.000 19.430 28.450 ;
        RECT 19.130 27.850 22.980 28.000 ;
        RECT 19.130 27.400 19.430 27.850 ;
        RECT 19.130 27.250 22.980 27.400 ;
        RECT 19.130 26.800 19.430 27.250 ;
        RECT 23.830 26.800 25.630 33.200 ;
        RECT 30.030 32.750 30.330 33.200 ;
        RECT 26.480 32.600 30.330 32.750 ;
        RECT 30.030 32.150 30.330 32.600 ;
        RECT 26.480 32.000 30.330 32.150 ;
        RECT 30.030 31.550 30.330 32.000 ;
        RECT 26.480 31.400 30.330 31.550 ;
        RECT 30.030 30.950 30.330 31.400 ;
        RECT 26.480 30.800 30.330 30.950 ;
        RECT 30.030 30.350 30.330 30.800 ;
        RECT 30.780 30.350 30.930 38.550 ;
        RECT 31.380 30.350 31.530 38.550 ;
        RECT 31.980 30.350 32.130 38.550 ;
        RECT 32.580 30.350 32.730 38.550 ;
        RECT 33.180 30.350 33.330 38.550 ;
        RECT 33.780 30.350 33.930 38.550 ;
        RECT 30.030 29.200 30.330 29.650 ;
        RECT 26.480 29.050 30.330 29.200 ;
        RECT 30.030 28.600 30.330 29.050 ;
        RECT 26.480 28.450 30.330 28.600 ;
        RECT 30.030 28.000 30.330 28.450 ;
        RECT 26.480 27.850 30.330 28.000 ;
        RECT 30.030 27.400 30.330 27.850 ;
        RECT 26.480 27.250 30.330 27.400 ;
        RECT 30.030 26.800 30.330 27.250 ;
        RECT 19.130 26.650 22.980 26.800 ;
        RECT 26.480 26.650 30.330 26.800 ;
        RECT 19.130 26.200 19.430 26.650 ;
        RECT 30.030 26.200 30.330 26.650 ;
        RECT 19.130 26.050 22.980 26.200 ;
        RECT 26.480 26.050 30.330 26.200 ;
        RECT 19.130 25.600 19.430 26.050 ;
        RECT 30.030 25.600 30.330 26.050 ;
        RECT 19.130 25.450 22.980 25.600 ;
        RECT 26.480 25.450 30.330 25.600 ;
        RECT 19.130 25.000 19.430 25.450 ;
        RECT 30.030 25.000 30.330 25.450 ;
        RECT 19.130 24.850 22.980 25.000 ;
        RECT 26.480 24.850 30.330 25.000 ;
        RECT 19.130 24.400 19.430 24.850 ;
        RECT 30.030 24.400 30.330 24.850 ;
        RECT 19.130 24.250 22.980 24.400 ;
        RECT 26.480 24.250 30.330 24.400 ;
        RECT 19.130 23.800 19.430 24.250 ;
        RECT 30.030 23.800 30.330 24.250 ;
        RECT 19.130 23.650 22.980 23.800 ;
        RECT 26.480 23.650 30.330 23.800 ;
        RECT 19.130 23.200 19.430 23.650 ;
        RECT 30.030 23.200 30.330 23.650 ;
        RECT 19.130 23.050 22.980 23.200 ;
        RECT 26.480 23.050 30.330 23.200 ;
        RECT 19.130 22.600 19.430 23.050 ;
        RECT 30.030 22.600 30.330 23.050 ;
        RECT 19.130 22.450 22.980 22.600 ;
        RECT 26.480 22.450 30.330 22.600 ;
        RECT 19.130 22.000 19.430 22.450 ;
        RECT 30.030 22.000 30.330 22.450 ;
        RECT 19.130 21.450 22.930 22.000 ;
        RECT 6.530 21.400 22.930 21.450 ;
        RECT 26.530 21.450 30.330 22.000 ;
        RECT 30.780 21.450 30.930 29.650 ;
        RECT 31.380 21.450 31.530 29.650 ;
        RECT 31.980 21.450 32.130 29.650 ;
        RECT 32.580 21.450 32.730 29.650 ;
        RECT 33.180 21.450 33.330 29.650 ;
        RECT 33.780 21.450 33.930 29.650 ;
        RECT 34.380 21.450 35.080 38.550 ;
        RECT 35.530 30.350 35.680 38.550 ;
        RECT 36.130 30.350 36.280 38.550 ;
        RECT 36.730 30.350 36.880 38.550 ;
        RECT 37.330 30.350 37.480 38.550 ;
        RECT 37.930 30.350 38.080 38.550 ;
        RECT 38.530 30.350 38.680 38.550 ;
        RECT 39.130 38.000 42.930 38.550 ;
        RECT 46.530 38.550 62.930 38.600 ;
        RECT 46.530 38.000 50.330 38.550 ;
        RECT 39.130 37.550 39.430 38.000 ;
        RECT 50.030 37.550 50.330 38.000 ;
        RECT 39.130 37.400 42.980 37.550 ;
        RECT 46.480 37.400 50.330 37.550 ;
        RECT 39.130 36.950 39.430 37.400 ;
        RECT 50.030 36.950 50.330 37.400 ;
        RECT 39.130 36.800 42.980 36.950 ;
        RECT 46.480 36.800 50.330 36.950 ;
        RECT 39.130 36.350 39.430 36.800 ;
        RECT 50.030 36.350 50.330 36.800 ;
        RECT 39.130 36.200 42.980 36.350 ;
        RECT 46.480 36.200 50.330 36.350 ;
        RECT 39.130 35.750 39.430 36.200 ;
        RECT 50.030 35.750 50.330 36.200 ;
        RECT 39.130 35.600 42.980 35.750 ;
        RECT 46.480 35.600 50.330 35.750 ;
        RECT 39.130 35.150 39.430 35.600 ;
        RECT 50.030 35.150 50.330 35.600 ;
        RECT 39.130 35.000 42.980 35.150 ;
        RECT 46.480 35.000 50.330 35.150 ;
        RECT 39.130 34.550 39.430 35.000 ;
        RECT 50.030 34.550 50.330 35.000 ;
        RECT 39.130 34.400 42.980 34.550 ;
        RECT 46.480 34.400 50.330 34.550 ;
        RECT 39.130 33.950 39.430 34.400 ;
        RECT 50.030 33.950 50.330 34.400 ;
        RECT 39.130 33.800 42.980 33.950 ;
        RECT 46.480 33.800 50.330 33.950 ;
        RECT 39.130 33.350 39.430 33.800 ;
        RECT 50.030 33.350 50.330 33.800 ;
        RECT 39.130 33.200 42.980 33.350 ;
        RECT 46.480 33.200 50.330 33.350 ;
        RECT 39.130 32.750 39.430 33.200 ;
        RECT 39.130 32.600 42.980 32.750 ;
        RECT 39.130 32.150 39.430 32.600 ;
        RECT 39.130 32.000 42.980 32.150 ;
        RECT 39.130 31.550 39.430 32.000 ;
        RECT 39.130 31.400 42.980 31.550 ;
        RECT 39.130 30.950 39.430 31.400 ;
        RECT 39.130 30.800 42.980 30.950 ;
        RECT 39.130 30.350 39.430 30.800 ;
        RECT 35.530 21.450 35.680 29.650 ;
        RECT 36.130 21.450 36.280 29.650 ;
        RECT 36.730 21.450 36.880 29.650 ;
        RECT 37.330 21.450 37.480 29.650 ;
        RECT 37.930 21.450 38.080 29.650 ;
        RECT 38.530 21.450 38.680 29.650 ;
        RECT 39.130 29.200 39.430 29.650 ;
        RECT 39.130 29.050 42.980 29.200 ;
        RECT 39.130 28.600 39.430 29.050 ;
        RECT 39.130 28.450 42.980 28.600 ;
        RECT 39.130 28.000 39.430 28.450 ;
        RECT 39.130 27.850 42.980 28.000 ;
        RECT 39.130 27.400 39.430 27.850 ;
        RECT 39.130 27.250 42.980 27.400 ;
        RECT 39.130 26.800 39.430 27.250 ;
        RECT 43.830 26.800 45.630 33.200 ;
        RECT 50.030 32.750 50.330 33.200 ;
        RECT 46.480 32.600 50.330 32.750 ;
        RECT 50.030 32.150 50.330 32.600 ;
        RECT 46.480 32.000 50.330 32.150 ;
        RECT 50.030 31.550 50.330 32.000 ;
        RECT 46.480 31.400 50.330 31.550 ;
        RECT 50.030 30.950 50.330 31.400 ;
        RECT 46.480 30.800 50.330 30.950 ;
        RECT 50.030 30.350 50.330 30.800 ;
        RECT 50.780 30.350 50.930 38.550 ;
        RECT 51.380 30.350 51.530 38.550 ;
        RECT 51.980 30.350 52.130 38.550 ;
        RECT 52.580 30.350 52.730 38.550 ;
        RECT 53.180 30.350 53.330 38.550 ;
        RECT 53.780 30.350 53.930 38.550 ;
        RECT 50.030 29.200 50.330 29.650 ;
        RECT 46.480 29.050 50.330 29.200 ;
        RECT 50.030 28.600 50.330 29.050 ;
        RECT 46.480 28.450 50.330 28.600 ;
        RECT 50.030 28.000 50.330 28.450 ;
        RECT 46.480 27.850 50.330 28.000 ;
        RECT 50.030 27.400 50.330 27.850 ;
        RECT 46.480 27.250 50.330 27.400 ;
        RECT 50.030 26.800 50.330 27.250 ;
        RECT 39.130 26.650 42.980 26.800 ;
        RECT 46.480 26.650 50.330 26.800 ;
        RECT 39.130 26.200 39.430 26.650 ;
        RECT 50.030 26.200 50.330 26.650 ;
        RECT 39.130 26.050 42.980 26.200 ;
        RECT 46.480 26.050 50.330 26.200 ;
        RECT 39.130 25.600 39.430 26.050 ;
        RECT 50.030 25.600 50.330 26.050 ;
        RECT 39.130 25.450 42.980 25.600 ;
        RECT 46.480 25.450 50.330 25.600 ;
        RECT 39.130 25.000 39.430 25.450 ;
        RECT 50.030 25.000 50.330 25.450 ;
        RECT 39.130 24.850 42.980 25.000 ;
        RECT 46.480 24.850 50.330 25.000 ;
        RECT 39.130 24.400 39.430 24.850 ;
        RECT 50.030 24.400 50.330 24.850 ;
        RECT 39.130 24.250 42.980 24.400 ;
        RECT 46.480 24.250 50.330 24.400 ;
        RECT 39.130 23.800 39.430 24.250 ;
        RECT 50.030 23.800 50.330 24.250 ;
        RECT 39.130 23.650 42.980 23.800 ;
        RECT 46.480 23.650 50.330 23.800 ;
        RECT 39.130 23.200 39.430 23.650 ;
        RECT 50.030 23.200 50.330 23.650 ;
        RECT 39.130 23.050 42.980 23.200 ;
        RECT 46.480 23.050 50.330 23.200 ;
        RECT 39.130 22.600 39.430 23.050 ;
        RECT 50.030 22.600 50.330 23.050 ;
        RECT 39.130 22.450 42.980 22.600 ;
        RECT 46.480 22.450 50.330 22.600 ;
        RECT 39.130 22.000 39.430 22.450 ;
        RECT 50.030 22.000 50.330 22.450 ;
        RECT 39.130 21.450 42.930 22.000 ;
        RECT 26.530 21.400 42.930 21.450 ;
        RECT 46.530 21.450 50.330 22.000 ;
        RECT 50.780 21.450 50.930 29.650 ;
        RECT 51.380 21.450 51.530 29.650 ;
        RECT 51.980 21.450 52.130 29.650 ;
        RECT 52.580 21.450 52.730 29.650 ;
        RECT 53.180 21.450 53.330 29.650 ;
        RECT 53.780 21.450 53.930 29.650 ;
        RECT 54.380 21.450 55.080 38.550 ;
        RECT 55.530 30.350 55.680 38.550 ;
        RECT 56.130 30.350 56.280 38.550 ;
        RECT 56.730 30.350 56.880 38.550 ;
        RECT 57.330 30.350 57.480 38.550 ;
        RECT 57.930 30.350 58.080 38.550 ;
        RECT 58.530 30.350 58.680 38.550 ;
        RECT 59.130 38.000 62.930 38.550 ;
        RECT 66.530 38.550 82.930 38.600 ;
        RECT 66.530 38.000 70.330 38.550 ;
        RECT 59.130 37.550 59.430 38.000 ;
        RECT 70.030 37.550 70.330 38.000 ;
        RECT 59.130 37.400 62.980 37.550 ;
        RECT 66.480 37.400 70.330 37.550 ;
        RECT 59.130 36.950 59.430 37.400 ;
        RECT 70.030 36.950 70.330 37.400 ;
        RECT 59.130 36.800 62.980 36.950 ;
        RECT 66.480 36.800 70.330 36.950 ;
        RECT 59.130 36.350 59.430 36.800 ;
        RECT 70.030 36.350 70.330 36.800 ;
        RECT 59.130 36.200 62.980 36.350 ;
        RECT 66.480 36.200 70.330 36.350 ;
        RECT 59.130 35.750 59.430 36.200 ;
        RECT 70.030 35.750 70.330 36.200 ;
        RECT 59.130 35.600 62.980 35.750 ;
        RECT 66.480 35.600 70.330 35.750 ;
        RECT 59.130 35.150 59.430 35.600 ;
        RECT 70.030 35.150 70.330 35.600 ;
        RECT 59.130 35.000 62.980 35.150 ;
        RECT 66.480 35.000 70.330 35.150 ;
        RECT 59.130 34.550 59.430 35.000 ;
        RECT 70.030 34.550 70.330 35.000 ;
        RECT 59.130 34.400 62.980 34.550 ;
        RECT 66.480 34.400 70.330 34.550 ;
        RECT 59.130 33.950 59.430 34.400 ;
        RECT 70.030 33.950 70.330 34.400 ;
        RECT 59.130 33.800 62.980 33.950 ;
        RECT 66.480 33.800 70.330 33.950 ;
        RECT 59.130 33.350 59.430 33.800 ;
        RECT 70.030 33.350 70.330 33.800 ;
        RECT 59.130 33.200 62.980 33.350 ;
        RECT 66.480 33.200 70.330 33.350 ;
        RECT 59.130 32.750 59.430 33.200 ;
        RECT 59.130 32.600 62.980 32.750 ;
        RECT 59.130 32.150 59.430 32.600 ;
        RECT 59.130 32.000 62.980 32.150 ;
        RECT 59.130 31.550 59.430 32.000 ;
        RECT 59.130 31.400 62.980 31.550 ;
        RECT 59.130 30.950 59.430 31.400 ;
        RECT 59.130 30.800 62.980 30.950 ;
        RECT 59.130 30.350 59.430 30.800 ;
        RECT 55.530 21.450 55.680 29.650 ;
        RECT 56.130 21.450 56.280 29.650 ;
        RECT 56.730 21.450 56.880 29.650 ;
        RECT 57.330 21.450 57.480 29.650 ;
        RECT 57.930 21.450 58.080 29.650 ;
        RECT 58.530 21.450 58.680 29.650 ;
        RECT 59.130 29.200 59.430 29.650 ;
        RECT 59.130 29.050 62.980 29.200 ;
        RECT 59.130 28.600 59.430 29.050 ;
        RECT 59.130 28.450 62.980 28.600 ;
        RECT 59.130 28.000 59.430 28.450 ;
        RECT 59.130 27.850 62.980 28.000 ;
        RECT 59.130 27.400 59.430 27.850 ;
        RECT 59.130 27.250 62.980 27.400 ;
        RECT 59.130 26.800 59.430 27.250 ;
        RECT 63.830 26.800 65.630 33.200 ;
        RECT 70.030 32.750 70.330 33.200 ;
        RECT 66.480 32.600 70.330 32.750 ;
        RECT 70.030 32.150 70.330 32.600 ;
        RECT 66.480 32.000 70.330 32.150 ;
        RECT 70.030 31.550 70.330 32.000 ;
        RECT 66.480 31.400 70.330 31.550 ;
        RECT 70.030 30.950 70.330 31.400 ;
        RECT 66.480 30.800 70.330 30.950 ;
        RECT 70.030 30.350 70.330 30.800 ;
        RECT 70.780 30.350 70.930 38.550 ;
        RECT 71.380 30.350 71.530 38.550 ;
        RECT 71.980 30.350 72.130 38.550 ;
        RECT 72.580 30.350 72.730 38.550 ;
        RECT 73.180 30.350 73.330 38.550 ;
        RECT 73.780 30.350 73.930 38.550 ;
        RECT 70.030 29.200 70.330 29.650 ;
        RECT 66.480 29.050 70.330 29.200 ;
        RECT 70.030 28.600 70.330 29.050 ;
        RECT 66.480 28.450 70.330 28.600 ;
        RECT 70.030 28.000 70.330 28.450 ;
        RECT 66.480 27.850 70.330 28.000 ;
        RECT 70.030 27.400 70.330 27.850 ;
        RECT 66.480 27.250 70.330 27.400 ;
        RECT 70.030 26.800 70.330 27.250 ;
        RECT 59.130 26.650 62.980 26.800 ;
        RECT 66.480 26.650 70.330 26.800 ;
        RECT 59.130 26.200 59.430 26.650 ;
        RECT 70.030 26.200 70.330 26.650 ;
        RECT 59.130 26.050 62.980 26.200 ;
        RECT 66.480 26.050 70.330 26.200 ;
        RECT 59.130 25.600 59.430 26.050 ;
        RECT 70.030 25.600 70.330 26.050 ;
        RECT 59.130 25.450 62.980 25.600 ;
        RECT 66.480 25.450 70.330 25.600 ;
        RECT 59.130 25.000 59.430 25.450 ;
        RECT 70.030 25.000 70.330 25.450 ;
        RECT 59.130 24.850 62.980 25.000 ;
        RECT 66.480 24.850 70.330 25.000 ;
        RECT 59.130 24.400 59.430 24.850 ;
        RECT 70.030 24.400 70.330 24.850 ;
        RECT 59.130 24.250 62.980 24.400 ;
        RECT 66.480 24.250 70.330 24.400 ;
        RECT 59.130 23.800 59.430 24.250 ;
        RECT 70.030 23.800 70.330 24.250 ;
        RECT 59.130 23.650 62.980 23.800 ;
        RECT 66.480 23.650 70.330 23.800 ;
        RECT 59.130 23.200 59.430 23.650 ;
        RECT 70.030 23.200 70.330 23.650 ;
        RECT 59.130 23.050 62.980 23.200 ;
        RECT 66.480 23.050 70.330 23.200 ;
        RECT 59.130 22.600 59.430 23.050 ;
        RECT 70.030 22.600 70.330 23.050 ;
        RECT 59.130 22.450 62.980 22.600 ;
        RECT 66.480 22.450 70.330 22.600 ;
        RECT 59.130 22.000 59.430 22.450 ;
        RECT 70.030 22.000 70.330 22.450 ;
        RECT 59.130 21.450 62.930 22.000 ;
        RECT 46.530 21.400 62.930 21.450 ;
        RECT 66.530 21.450 70.330 22.000 ;
        RECT 70.780 21.450 70.930 29.650 ;
        RECT 71.380 21.450 71.530 29.650 ;
        RECT 71.980 21.450 72.130 29.650 ;
        RECT 72.580 21.450 72.730 29.650 ;
        RECT 73.180 21.450 73.330 29.650 ;
        RECT 73.780 21.450 73.930 29.650 ;
        RECT 74.380 21.450 75.080 38.550 ;
        RECT 75.530 30.350 75.680 38.550 ;
        RECT 76.130 30.350 76.280 38.550 ;
        RECT 76.730 30.350 76.880 38.550 ;
        RECT 77.330 30.350 77.480 38.550 ;
        RECT 77.930 30.350 78.080 38.550 ;
        RECT 78.530 30.350 78.680 38.550 ;
        RECT 79.130 38.000 82.930 38.550 ;
        RECT 86.530 38.550 102.930 38.600 ;
        RECT 86.530 38.000 90.330 38.550 ;
        RECT 79.130 37.550 79.430 38.000 ;
        RECT 90.030 37.550 90.330 38.000 ;
        RECT 79.130 37.400 82.980 37.550 ;
        RECT 86.480 37.400 90.330 37.550 ;
        RECT 79.130 36.950 79.430 37.400 ;
        RECT 90.030 36.950 90.330 37.400 ;
        RECT 79.130 36.800 82.980 36.950 ;
        RECT 86.480 36.800 90.330 36.950 ;
        RECT 79.130 36.350 79.430 36.800 ;
        RECT 90.030 36.350 90.330 36.800 ;
        RECT 79.130 36.200 82.980 36.350 ;
        RECT 86.480 36.200 90.330 36.350 ;
        RECT 79.130 35.750 79.430 36.200 ;
        RECT 90.030 35.750 90.330 36.200 ;
        RECT 79.130 35.600 82.980 35.750 ;
        RECT 86.480 35.600 90.330 35.750 ;
        RECT 79.130 35.150 79.430 35.600 ;
        RECT 90.030 35.150 90.330 35.600 ;
        RECT 79.130 35.000 82.980 35.150 ;
        RECT 86.480 35.000 90.330 35.150 ;
        RECT 79.130 34.550 79.430 35.000 ;
        RECT 90.030 34.550 90.330 35.000 ;
        RECT 79.130 34.400 82.980 34.550 ;
        RECT 86.480 34.400 90.330 34.550 ;
        RECT 79.130 33.950 79.430 34.400 ;
        RECT 90.030 33.950 90.330 34.400 ;
        RECT 79.130 33.800 82.980 33.950 ;
        RECT 86.480 33.800 90.330 33.950 ;
        RECT 79.130 33.350 79.430 33.800 ;
        RECT 90.030 33.350 90.330 33.800 ;
        RECT 79.130 33.200 82.980 33.350 ;
        RECT 86.480 33.200 90.330 33.350 ;
        RECT 79.130 32.750 79.430 33.200 ;
        RECT 79.130 32.600 82.980 32.750 ;
        RECT 79.130 32.150 79.430 32.600 ;
        RECT 79.130 32.000 82.980 32.150 ;
        RECT 79.130 31.550 79.430 32.000 ;
        RECT 79.130 31.400 82.980 31.550 ;
        RECT 79.130 30.950 79.430 31.400 ;
        RECT 79.130 30.800 82.980 30.950 ;
        RECT 79.130 30.350 79.430 30.800 ;
        RECT 75.530 21.450 75.680 29.650 ;
        RECT 76.130 21.450 76.280 29.650 ;
        RECT 76.730 21.450 76.880 29.650 ;
        RECT 77.330 21.450 77.480 29.650 ;
        RECT 77.930 21.450 78.080 29.650 ;
        RECT 78.530 21.450 78.680 29.650 ;
        RECT 79.130 29.200 79.430 29.650 ;
        RECT 79.130 29.050 82.980 29.200 ;
        RECT 79.130 28.600 79.430 29.050 ;
        RECT 79.130 28.450 82.980 28.600 ;
        RECT 79.130 28.000 79.430 28.450 ;
        RECT 79.130 27.850 82.980 28.000 ;
        RECT 79.130 27.400 79.430 27.850 ;
        RECT 79.130 27.250 82.980 27.400 ;
        RECT 79.130 26.800 79.430 27.250 ;
        RECT 83.830 26.800 85.630 33.200 ;
        RECT 90.030 32.750 90.330 33.200 ;
        RECT 86.480 32.600 90.330 32.750 ;
        RECT 90.030 32.150 90.330 32.600 ;
        RECT 86.480 32.000 90.330 32.150 ;
        RECT 90.030 31.550 90.330 32.000 ;
        RECT 86.480 31.400 90.330 31.550 ;
        RECT 90.030 30.950 90.330 31.400 ;
        RECT 86.480 30.800 90.330 30.950 ;
        RECT 90.030 30.350 90.330 30.800 ;
        RECT 90.780 30.350 90.930 38.550 ;
        RECT 91.380 30.350 91.530 38.550 ;
        RECT 91.980 30.350 92.130 38.550 ;
        RECT 92.580 30.350 92.730 38.550 ;
        RECT 93.180 30.350 93.330 38.550 ;
        RECT 93.780 30.350 93.930 38.550 ;
        RECT 90.030 29.200 90.330 29.650 ;
        RECT 86.480 29.050 90.330 29.200 ;
        RECT 90.030 28.600 90.330 29.050 ;
        RECT 86.480 28.450 90.330 28.600 ;
        RECT 90.030 28.000 90.330 28.450 ;
        RECT 86.480 27.850 90.330 28.000 ;
        RECT 90.030 27.400 90.330 27.850 ;
        RECT 86.480 27.250 90.330 27.400 ;
        RECT 90.030 26.800 90.330 27.250 ;
        RECT 79.130 26.650 82.980 26.800 ;
        RECT 86.480 26.650 90.330 26.800 ;
        RECT 79.130 26.200 79.430 26.650 ;
        RECT 90.030 26.200 90.330 26.650 ;
        RECT 79.130 26.050 82.980 26.200 ;
        RECT 86.480 26.050 90.330 26.200 ;
        RECT 79.130 25.600 79.430 26.050 ;
        RECT 90.030 25.600 90.330 26.050 ;
        RECT 79.130 25.450 82.980 25.600 ;
        RECT 86.480 25.450 90.330 25.600 ;
        RECT 79.130 25.000 79.430 25.450 ;
        RECT 90.030 25.000 90.330 25.450 ;
        RECT 79.130 24.850 82.980 25.000 ;
        RECT 86.480 24.850 90.330 25.000 ;
        RECT 79.130 24.400 79.430 24.850 ;
        RECT 90.030 24.400 90.330 24.850 ;
        RECT 79.130 24.250 82.980 24.400 ;
        RECT 86.480 24.250 90.330 24.400 ;
        RECT 79.130 23.800 79.430 24.250 ;
        RECT 90.030 23.800 90.330 24.250 ;
        RECT 79.130 23.650 82.980 23.800 ;
        RECT 86.480 23.650 90.330 23.800 ;
        RECT 79.130 23.200 79.430 23.650 ;
        RECT 90.030 23.200 90.330 23.650 ;
        RECT 79.130 23.050 82.980 23.200 ;
        RECT 86.480 23.050 90.330 23.200 ;
        RECT 79.130 22.600 79.430 23.050 ;
        RECT 90.030 22.600 90.330 23.050 ;
        RECT 79.130 22.450 82.980 22.600 ;
        RECT 86.480 22.450 90.330 22.600 ;
        RECT 79.130 22.000 79.430 22.450 ;
        RECT 90.030 22.000 90.330 22.450 ;
        RECT 79.130 21.450 82.930 22.000 ;
        RECT 66.530 21.400 82.930 21.450 ;
        RECT 86.530 21.450 90.330 22.000 ;
        RECT 90.780 21.450 90.930 29.650 ;
        RECT 91.380 21.450 91.530 29.650 ;
        RECT 91.980 21.450 92.130 29.650 ;
        RECT 92.580 21.450 92.730 29.650 ;
        RECT 93.180 21.450 93.330 29.650 ;
        RECT 93.780 21.450 93.930 29.650 ;
        RECT 94.380 21.450 95.080 38.550 ;
        RECT 95.530 30.350 95.680 38.550 ;
        RECT 96.130 30.350 96.280 38.550 ;
        RECT 96.730 30.350 96.880 38.550 ;
        RECT 97.330 30.350 97.480 38.550 ;
        RECT 97.930 30.350 98.080 38.550 ;
        RECT 98.530 30.350 98.680 38.550 ;
        RECT 99.130 38.000 102.930 38.550 ;
        RECT 106.530 38.550 122.930 38.600 ;
        RECT 106.530 38.000 110.330 38.550 ;
        RECT 99.130 37.550 99.430 38.000 ;
        RECT 110.030 37.550 110.330 38.000 ;
        RECT 99.130 37.400 102.980 37.550 ;
        RECT 106.480 37.400 110.330 37.550 ;
        RECT 99.130 36.950 99.430 37.400 ;
        RECT 110.030 36.950 110.330 37.400 ;
        RECT 99.130 36.800 102.980 36.950 ;
        RECT 106.480 36.800 110.330 36.950 ;
        RECT 99.130 36.350 99.430 36.800 ;
        RECT 110.030 36.350 110.330 36.800 ;
        RECT 99.130 36.200 102.980 36.350 ;
        RECT 106.480 36.200 110.330 36.350 ;
        RECT 99.130 35.750 99.430 36.200 ;
        RECT 110.030 35.750 110.330 36.200 ;
        RECT 99.130 35.600 102.980 35.750 ;
        RECT 106.480 35.600 110.330 35.750 ;
        RECT 99.130 35.150 99.430 35.600 ;
        RECT 110.030 35.150 110.330 35.600 ;
        RECT 99.130 35.000 102.980 35.150 ;
        RECT 106.480 35.000 110.330 35.150 ;
        RECT 99.130 34.550 99.430 35.000 ;
        RECT 110.030 34.550 110.330 35.000 ;
        RECT 99.130 34.400 102.980 34.550 ;
        RECT 106.480 34.400 110.330 34.550 ;
        RECT 99.130 33.950 99.430 34.400 ;
        RECT 110.030 33.950 110.330 34.400 ;
        RECT 99.130 33.800 102.980 33.950 ;
        RECT 106.480 33.800 110.330 33.950 ;
        RECT 99.130 33.350 99.430 33.800 ;
        RECT 110.030 33.350 110.330 33.800 ;
        RECT 99.130 33.200 102.980 33.350 ;
        RECT 106.480 33.200 110.330 33.350 ;
        RECT 99.130 32.750 99.430 33.200 ;
        RECT 99.130 32.600 102.980 32.750 ;
        RECT 99.130 32.150 99.430 32.600 ;
        RECT 99.130 32.000 102.980 32.150 ;
        RECT 99.130 31.550 99.430 32.000 ;
        RECT 99.130 31.400 102.980 31.550 ;
        RECT 99.130 30.950 99.430 31.400 ;
        RECT 99.130 30.800 102.980 30.950 ;
        RECT 99.130 30.350 99.430 30.800 ;
        RECT 95.530 21.450 95.680 29.650 ;
        RECT 96.130 21.450 96.280 29.650 ;
        RECT 96.730 21.450 96.880 29.650 ;
        RECT 97.330 21.450 97.480 29.650 ;
        RECT 97.930 21.450 98.080 29.650 ;
        RECT 98.530 21.450 98.680 29.650 ;
        RECT 99.130 29.200 99.430 29.650 ;
        RECT 99.130 29.050 102.980 29.200 ;
        RECT 99.130 28.600 99.430 29.050 ;
        RECT 99.130 28.450 102.980 28.600 ;
        RECT 99.130 28.000 99.430 28.450 ;
        RECT 99.130 27.850 102.980 28.000 ;
        RECT 99.130 27.400 99.430 27.850 ;
        RECT 99.130 27.250 102.980 27.400 ;
        RECT 99.130 26.800 99.430 27.250 ;
        RECT 103.830 26.800 105.630 33.200 ;
        RECT 110.030 32.750 110.330 33.200 ;
        RECT 106.480 32.600 110.330 32.750 ;
        RECT 110.030 32.150 110.330 32.600 ;
        RECT 106.480 32.000 110.330 32.150 ;
        RECT 110.030 31.550 110.330 32.000 ;
        RECT 106.480 31.400 110.330 31.550 ;
        RECT 110.030 30.950 110.330 31.400 ;
        RECT 106.480 30.800 110.330 30.950 ;
        RECT 110.030 30.350 110.330 30.800 ;
        RECT 110.780 30.350 110.930 38.550 ;
        RECT 111.380 30.350 111.530 38.550 ;
        RECT 111.980 30.350 112.130 38.550 ;
        RECT 112.580 30.350 112.730 38.550 ;
        RECT 113.180 30.350 113.330 38.550 ;
        RECT 113.780 30.350 113.930 38.550 ;
        RECT 110.030 29.200 110.330 29.650 ;
        RECT 106.480 29.050 110.330 29.200 ;
        RECT 110.030 28.600 110.330 29.050 ;
        RECT 106.480 28.450 110.330 28.600 ;
        RECT 110.030 28.000 110.330 28.450 ;
        RECT 106.480 27.850 110.330 28.000 ;
        RECT 110.030 27.400 110.330 27.850 ;
        RECT 106.480 27.250 110.330 27.400 ;
        RECT 110.030 26.800 110.330 27.250 ;
        RECT 99.130 26.650 102.980 26.800 ;
        RECT 106.480 26.650 110.330 26.800 ;
        RECT 99.130 26.200 99.430 26.650 ;
        RECT 110.030 26.200 110.330 26.650 ;
        RECT 99.130 26.050 102.980 26.200 ;
        RECT 106.480 26.050 110.330 26.200 ;
        RECT 99.130 25.600 99.430 26.050 ;
        RECT 110.030 25.600 110.330 26.050 ;
        RECT 99.130 25.450 102.980 25.600 ;
        RECT 106.480 25.450 110.330 25.600 ;
        RECT 99.130 25.000 99.430 25.450 ;
        RECT 110.030 25.000 110.330 25.450 ;
        RECT 99.130 24.850 102.980 25.000 ;
        RECT 106.480 24.850 110.330 25.000 ;
        RECT 99.130 24.400 99.430 24.850 ;
        RECT 110.030 24.400 110.330 24.850 ;
        RECT 99.130 24.250 102.980 24.400 ;
        RECT 106.480 24.250 110.330 24.400 ;
        RECT 99.130 23.800 99.430 24.250 ;
        RECT 110.030 23.800 110.330 24.250 ;
        RECT 99.130 23.650 102.980 23.800 ;
        RECT 106.480 23.650 110.330 23.800 ;
        RECT 99.130 23.200 99.430 23.650 ;
        RECT 110.030 23.200 110.330 23.650 ;
        RECT 99.130 23.050 102.980 23.200 ;
        RECT 106.480 23.050 110.330 23.200 ;
        RECT 99.130 22.600 99.430 23.050 ;
        RECT 110.030 22.600 110.330 23.050 ;
        RECT 99.130 22.450 102.980 22.600 ;
        RECT 106.480 22.450 110.330 22.600 ;
        RECT 99.130 22.000 99.430 22.450 ;
        RECT 110.030 22.000 110.330 22.450 ;
        RECT 99.130 21.450 102.930 22.000 ;
        RECT 86.530 21.400 102.930 21.450 ;
        RECT 106.530 21.450 110.330 22.000 ;
        RECT 110.780 21.450 110.930 29.650 ;
        RECT 111.380 21.450 111.530 29.650 ;
        RECT 111.980 21.450 112.130 29.650 ;
        RECT 112.580 21.450 112.730 29.650 ;
        RECT 113.180 21.450 113.330 29.650 ;
        RECT 113.780 21.450 113.930 29.650 ;
        RECT 114.380 21.450 115.080 38.550 ;
        RECT 115.530 30.350 115.680 38.550 ;
        RECT 116.130 30.350 116.280 38.550 ;
        RECT 116.730 30.350 116.880 38.550 ;
        RECT 117.330 30.350 117.480 38.550 ;
        RECT 117.930 30.350 118.080 38.550 ;
        RECT 118.530 30.350 118.680 38.550 ;
        RECT 119.130 38.000 122.930 38.550 ;
        RECT 119.130 37.550 119.430 38.000 ;
        RECT 119.130 37.400 122.980 37.550 ;
        RECT 119.130 36.950 119.430 37.400 ;
        RECT 119.130 36.800 122.980 36.950 ;
        RECT 119.130 36.350 119.430 36.800 ;
        RECT 119.130 36.200 122.980 36.350 ;
        RECT 119.130 35.750 119.430 36.200 ;
        RECT 119.130 35.600 122.980 35.750 ;
        RECT 119.130 35.150 119.430 35.600 ;
        RECT 119.130 35.000 122.980 35.150 ;
        RECT 119.130 34.550 119.430 35.000 ;
        RECT 119.130 34.400 122.980 34.550 ;
        RECT 119.130 33.950 119.430 34.400 ;
        RECT 119.130 33.800 122.980 33.950 ;
        RECT 119.130 33.350 119.430 33.800 ;
        RECT 119.130 33.200 122.980 33.350 ;
        RECT 119.130 32.750 119.430 33.200 ;
        RECT 119.130 32.600 122.980 32.750 ;
        RECT 119.130 32.150 119.430 32.600 ;
        RECT 119.130 32.000 122.980 32.150 ;
        RECT 119.130 31.550 119.430 32.000 ;
        RECT 119.130 31.400 122.980 31.550 ;
        RECT 119.130 30.950 119.430 31.400 ;
        RECT 119.130 30.800 122.980 30.950 ;
        RECT 119.130 30.350 119.430 30.800 ;
        RECT 115.530 21.450 115.680 29.650 ;
        RECT 116.130 21.450 116.280 29.650 ;
        RECT 116.730 21.450 116.880 29.650 ;
        RECT 117.330 21.450 117.480 29.650 ;
        RECT 117.930 21.450 118.080 29.650 ;
        RECT 118.530 21.450 118.680 29.650 ;
        RECT 119.130 29.200 119.430 29.650 ;
        RECT 119.130 29.050 122.980 29.200 ;
        RECT 119.130 28.600 119.430 29.050 ;
        RECT 119.130 28.450 122.980 28.600 ;
        RECT 119.130 28.000 119.430 28.450 ;
        RECT 119.130 27.850 122.980 28.000 ;
        RECT 119.130 27.400 119.430 27.850 ;
        RECT 119.130 27.250 122.980 27.400 ;
        RECT 119.130 26.800 119.430 27.250 ;
        RECT 123.830 26.800 124.730 33.200 ;
        RECT 129.850 30.310 131.850 31.585 ;
        RECT 119.130 26.650 122.980 26.800 ;
        RECT 119.130 26.200 119.430 26.650 ;
        RECT 119.130 26.050 122.980 26.200 ;
        RECT 119.130 25.600 119.430 26.050 ;
        RECT 119.130 25.450 122.980 25.600 ;
        RECT 119.130 25.000 119.430 25.450 ;
        RECT 119.130 24.850 122.980 25.000 ;
        RECT 119.130 24.400 119.430 24.850 ;
        RECT 119.130 24.250 122.980 24.400 ;
        RECT 119.130 23.800 119.430 24.250 ;
        RECT 119.130 23.650 122.980 23.800 ;
        RECT 119.130 23.200 119.430 23.650 ;
        RECT 119.130 23.050 122.980 23.200 ;
        RECT 119.130 22.600 119.430 23.050 ;
        RECT 119.130 22.450 122.980 22.600 ;
        RECT 119.130 22.000 119.430 22.450 ;
        RECT 119.130 21.450 122.930 22.000 ;
        RECT 106.530 21.400 122.930 21.450 ;
        RECT 9.630 20.900 19.830 21.400 ;
        RECT 29.630 20.900 39.830 21.400 ;
        RECT 49.630 20.900 59.830 21.400 ;
        RECT 69.630 20.900 79.830 21.400 ;
        RECT 89.630 20.900 99.830 21.400 ;
        RECT 109.630 20.900 119.830 21.400 ;
        RECT 11.530 19.100 17.930 20.900 ;
        RECT 31.530 19.100 37.930 20.900 ;
        RECT 51.530 19.100 57.930 20.900 ;
        RECT 71.530 19.100 77.930 20.900 ;
        RECT 91.530 19.100 97.930 20.900 ;
        RECT 111.530 19.100 117.930 20.900 ;
        RECT 9.630 18.600 19.830 19.100 ;
        RECT 29.630 18.600 39.830 19.100 ;
        RECT 49.630 18.600 59.830 19.100 ;
        RECT 69.630 18.600 79.830 19.100 ;
        RECT 89.630 18.600 99.830 19.100 ;
        RECT 109.630 18.600 119.830 19.100 ;
        RECT 6.530 18.550 22.930 18.600 ;
        RECT 6.530 18.000 10.330 18.550 ;
        RECT 10.030 17.550 10.330 18.000 ;
        RECT 6.480 17.400 10.330 17.550 ;
        RECT 10.030 16.950 10.330 17.400 ;
        RECT 6.480 16.800 10.330 16.950 ;
        RECT 10.030 16.350 10.330 16.800 ;
        RECT 6.480 16.200 10.330 16.350 ;
        RECT 10.030 15.750 10.330 16.200 ;
        RECT 6.480 15.600 10.330 15.750 ;
        RECT 10.030 15.150 10.330 15.600 ;
        RECT 6.480 15.000 10.330 15.150 ;
        RECT 10.030 14.550 10.330 15.000 ;
        RECT 6.480 14.400 10.330 14.550 ;
        RECT 10.030 13.950 10.330 14.400 ;
        RECT 6.480 13.800 10.330 13.950 ;
        RECT 10.030 13.350 10.330 13.800 ;
        RECT 6.480 13.200 10.330 13.350 ;
        RECT 4.730 6.800 5.630 13.200 ;
        RECT 10.030 12.750 10.330 13.200 ;
        RECT 6.480 12.600 10.330 12.750 ;
        RECT 10.030 12.150 10.330 12.600 ;
        RECT 6.480 12.000 10.330 12.150 ;
        RECT 10.030 11.550 10.330 12.000 ;
        RECT 6.480 11.400 10.330 11.550 ;
        RECT 10.030 10.950 10.330 11.400 ;
        RECT 6.480 10.800 10.330 10.950 ;
        RECT 10.030 10.350 10.330 10.800 ;
        RECT 10.780 10.350 10.930 18.550 ;
        RECT 11.380 10.350 11.530 18.550 ;
        RECT 11.980 10.350 12.130 18.550 ;
        RECT 12.580 10.350 12.730 18.550 ;
        RECT 13.180 10.350 13.330 18.550 ;
        RECT 13.780 10.350 13.930 18.550 ;
        RECT 10.030 9.200 10.330 9.650 ;
        RECT 6.480 9.050 10.330 9.200 ;
        RECT 10.030 8.600 10.330 9.050 ;
        RECT 6.480 8.450 10.330 8.600 ;
        RECT 10.030 8.000 10.330 8.450 ;
        RECT 6.480 7.850 10.330 8.000 ;
        RECT 10.030 7.400 10.330 7.850 ;
        RECT 6.480 7.250 10.330 7.400 ;
        RECT 10.030 6.800 10.330 7.250 ;
        RECT 6.480 6.650 10.330 6.800 ;
        RECT 10.030 6.200 10.330 6.650 ;
        RECT 6.480 6.050 10.330 6.200 ;
        RECT 10.030 5.600 10.330 6.050 ;
        RECT 6.480 5.450 10.330 5.600 ;
        RECT 10.030 5.000 10.330 5.450 ;
        RECT 6.480 4.850 10.330 5.000 ;
        RECT 10.030 4.400 10.330 4.850 ;
        RECT 6.480 4.250 10.330 4.400 ;
        RECT 10.030 3.800 10.330 4.250 ;
        RECT 6.480 3.650 10.330 3.800 ;
        RECT 10.030 3.200 10.330 3.650 ;
        RECT 6.480 3.050 10.330 3.200 ;
        RECT 10.030 2.600 10.330 3.050 ;
        RECT 6.480 2.450 10.330 2.600 ;
        RECT 10.030 2.000 10.330 2.450 ;
        RECT 6.530 1.450 10.330 2.000 ;
        RECT 10.780 1.450 10.930 9.650 ;
        RECT 11.380 1.450 11.530 9.650 ;
        RECT 11.980 1.450 12.130 9.650 ;
        RECT 12.580 1.450 12.730 9.650 ;
        RECT 13.180 1.450 13.330 9.650 ;
        RECT 13.780 1.450 13.930 9.650 ;
        RECT 14.380 1.450 15.080 18.550 ;
        RECT 15.530 10.350 15.680 18.550 ;
        RECT 16.130 10.350 16.280 18.550 ;
        RECT 16.730 10.350 16.880 18.550 ;
        RECT 17.330 10.350 17.480 18.550 ;
        RECT 17.930 10.350 18.080 18.550 ;
        RECT 18.530 10.350 18.680 18.550 ;
        RECT 19.130 18.000 22.930 18.550 ;
        RECT 26.530 18.550 42.930 18.600 ;
        RECT 26.530 18.000 30.330 18.550 ;
        RECT 19.130 17.550 19.430 18.000 ;
        RECT 30.030 17.550 30.330 18.000 ;
        RECT 19.130 17.400 22.980 17.550 ;
        RECT 26.480 17.400 30.330 17.550 ;
        RECT 19.130 16.950 19.430 17.400 ;
        RECT 30.030 16.950 30.330 17.400 ;
        RECT 19.130 16.800 22.980 16.950 ;
        RECT 26.480 16.800 30.330 16.950 ;
        RECT 19.130 16.350 19.430 16.800 ;
        RECT 30.030 16.350 30.330 16.800 ;
        RECT 19.130 16.200 22.980 16.350 ;
        RECT 26.480 16.200 30.330 16.350 ;
        RECT 19.130 15.750 19.430 16.200 ;
        RECT 30.030 15.750 30.330 16.200 ;
        RECT 19.130 15.600 22.980 15.750 ;
        RECT 26.480 15.600 30.330 15.750 ;
        RECT 19.130 15.150 19.430 15.600 ;
        RECT 30.030 15.150 30.330 15.600 ;
        RECT 19.130 15.000 22.980 15.150 ;
        RECT 26.480 15.000 30.330 15.150 ;
        RECT 19.130 14.550 19.430 15.000 ;
        RECT 30.030 14.550 30.330 15.000 ;
        RECT 19.130 14.400 22.980 14.550 ;
        RECT 26.480 14.400 30.330 14.550 ;
        RECT 19.130 13.950 19.430 14.400 ;
        RECT 30.030 13.950 30.330 14.400 ;
        RECT 19.130 13.800 22.980 13.950 ;
        RECT 26.480 13.800 30.330 13.950 ;
        RECT 19.130 13.350 19.430 13.800 ;
        RECT 30.030 13.350 30.330 13.800 ;
        RECT 19.130 13.200 22.980 13.350 ;
        RECT 26.480 13.200 30.330 13.350 ;
        RECT 19.130 12.750 19.430 13.200 ;
        RECT 19.130 12.600 22.980 12.750 ;
        RECT 19.130 12.150 19.430 12.600 ;
        RECT 19.130 12.000 22.980 12.150 ;
        RECT 19.130 11.550 19.430 12.000 ;
        RECT 19.130 11.400 22.980 11.550 ;
        RECT 19.130 10.950 19.430 11.400 ;
        RECT 19.130 10.800 22.980 10.950 ;
        RECT 19.130 10.350 19.430 10.800 ;
        RECT 15.530 1.450 15.680 9.650 ;
        RECT 16.130 1.450 16.280 9.650 ;
        RECT 16.730 1.450 16.880 9.650 ;
        RECT 17.330 1.450 17.480 9.650 ;
        RECT 17.930 1.450 18.080 9.650 ;
        RECT 18.530 1.450 18.680 9.650 ;
        RECT 19.130 9.200 19.430 9.650 ;
        RECT 19.130 9.050 22.980 9.200 ;
        RECT 19.130 8.600 19.430 9.050 ;
        RECT 19.130 8.450 22.980 8.600 ;
        RECT 19.130 8.000 19.430 8.450 ;
        RECT 19.130 7.850 22.980 8.000 ;
        RECT 19.130 7.400 19.430 7.850 ;
        RECT 19.130 7.250 22.980 7.400 ;
        RECT 19.130 6.800 19.430 7.250 ;
        RECT 23.830 6.800 25.630 13.200 ;
        RECT 30.030 12.750 30.330 13.200 ;
        RECT 26.480 12.600 30.330 12.750 ;
        RECT 30.030 12.150 30.330 12.600 ;
        RECT 26.480 12.000 30.330 12.150 ;
        RECT 30.030 11.550 30.330 12.000 ;
        RECT 26.480 11.400 30.330 11.550 ;
        RECT 30.030 10.950 30.330 11.400 ;
        RECT 26.480 10.800 30.330 10.950 ;
        RECT 30.030 10.350 30.330 10.800 ;
        RECT 30.780 10.350 30.930 18.550 ;
        RECT 31.380 10.350 31.530 18.550 ;
        RECT 31.980 10.350 32.130 18.550 ;
        RECT 32.580 10.350 32.730 18.550 ;
        RECT 33.180 10.350 33.330 18.550 ;
        RECT 33.780 10.350 33.930 18.550 ;
        RECT 30.030 9.200 30.330 9.650 ;
        RECT 26.480 9.050 30.330 9.200 ;
        RECT 30.030 8.600 30.330 9.050 ;
        RECT 26.480 8.450 30.330 8.600 ;
        RECT 30.030 8.000 30.330 8.450 ;
        RECT 26.480 7.850 30.330 8.000 ;
        RECT 30.030 7.400 30.330 7.850 ;
        RECT 26.480 7.250 30.330 7.400 ;
        RECT 30.030 6.800 30.330 7.250 ;
        RECT 19.130 6.650 22.980 6.800 ;
        RECT 26.480 6.650 30.330 6.800 ;
        RECT 19.130 6.200 19.430 6.650 ;
        RECT 30.030 6.200 30.330 6.650 ;
        RECT 19.130 6.050 22.980 6.200 ;
        RECT 26.480 6.050 30.330 6.200 ;
        RECT 19.130 5.600 19.430 6.050 ;
        RECT 30.030 5.600 30.330 6.050 ;
        RECT 19.130 5.450 22.980 5.600 ;
        RECT 26.480 5.450 30.330 5.600 ;
        RECT 19.130 5.000 19.430 5.450 ;
        RECT 30.030 5.000 30.330 5.450 ;
        RECT 19.130 4.850 22.980 5.000 ;
        RECT 26.480 4.850 30.330 5.000 ;
        RECT 19.130 4.400 19.430 4.850 ;
        RECT 30.030 4.400 30.330 4.850 ;
        RECT 19.130 4.250 22.980 4.400 ;
        RECT 26.480 4.250 30.330 4.400 ;
        RECT 19.130 3.800 19.430 4.250 ;
        RECT 30.030 3.800 30.330 4.250 ;
        RECT 19.130 3.650 22.980 3.800 ;
        RECT 26.480 3.650 30.330 3.800 ;
        RECT 19.130 3.200 19.430 3.650 ;
        RECT 30.030 3.200 30.330 3.650 ;
        RECT 19.130 3.050 22.980 3.200 ;
        RECT 26.480 3.050 30.330 3.200 ;
        RECT 19.130 2.600 19.430 3.050 ;
        RECT 30.030 2.600 30.330 3.050 ;
        RECT 19.130 2.450 22.980 2.600 ;
        RECT 26.480 2.450 30.330 2.600 ;
        RECT 19.130 2.000 19.430 2.450 ;
        RECT 30.030 2.000 30.330 2.450 ;
        RECT 19.130 1.450 22.930 2.000 ;
        RECT 6.530 1.400 22.930 1.450 ;
        RECT 26.530 1.450 30.330 2.000 ;
        RECT 30.780 1.450 30.930 9.650 ;
        RECT 31.380 1.450 31.530 9.650 ;
        RECT 31.980 1.450 32.130 9.650 ;
        RECT 32.580 1.450 32.730 9.650 ;
        RECT 33.180 1.450 33.330 9.650 ;
        RECT 33.780 1.450 33.930 9.650 ;
        RECT 34.380 1.450 35.080 18.550 ;
        RECT 35.530 10.350 35.680 18.550 ;
        RECT 36.130 10.350 36.280 18.550 ;
        RECT 36.730 10.350 36.880 18.550 ;
        RECT 37.330 10.350 37.480 18.550 ;
        RECT 37.930 10.350 38.080 18.550 ;
        RECT 38.530 10.350 38.680 18.550 ;
        RECT 39.130 18.000 42.930 18.550 ;
        RECT 46.530 18.550 62.930 18.600 ;
        RECT 46.530 18.000 50.330 18.550 ;
        RECT 39.130 17.550 39.430 18.000 ;
        RECT 50.030 17.550 50.330 18.000 ;
        RECT 39.130 17.400 42.980 17.550 ;
        RECT 46.480 17.400 50.330 17.550 ;
        RECT 39.130 16.950 39.430 17.400 ;
        RECT 50.030 16.950 50.330 17.400 ;
        RECT 39.130 16.800 42.980 16.950 ;
        RECT 46.480 16.800 50.330 16.950 ;
        RECT 39.130 16.350 39.430 16.800 ;
        RECT 50.030 16.350 50.330 16.800 ;
        RECT 39.130 16.200 42.980 16.350 ;
        RECT 46.480 16.200 50.330 16.350 ;
        RECT 39.130 15.750 39.430 16.200 ;
        RECT 50.030 15.750 50.330 16.200 ;
        RECT 39.130 15.600 42.980 15.750 ;
        RECT 46.480 15.600 50.330 15.750 ;
        RECT 39.130 15.150 39.430 15.600 ;
        RECT 50.030 15.150 50.330 15.600 ;
        RECT 39.130 15.000 42.980 15.150 ;
        RECT 46.480 15.000 50.330 15.150 ;
        RECT 39.130 14.550 39.430 15.000 ;
        RECT 50.030 14.550 50.330 15.000 ;
        RECT 39.130 14.400 42.980 14.550 ;
        RECT 46.480 14.400 50.330 14.550 ;
        RECT 39.130 13.950 39.430 14.400 ;
        RECT 50.030 13.950 50.330 14.400 ;
        RECT 39.130 13.800 42.980 13.950 ;
        RECT 46.480 13.800 50.330 13.950 ;
        RECT 39.130 13.350 39.430 13.800 ;
        RECT 50.030 13.350 50.330 13.800 ;
        RECT 39.130 13.200 42.980 13.350 ;
        RECT 46.480 13.200 50.330 13.350 ;
        RECT 39.130 12.750 39.430 13.200 ;
        RECT 39.130 12.600 42.980 12.750 ;
        RECT 39.130 12.150 39.430 12.600 ;
        RECT 39.130 12.000 42.980 12.150 ;
        RECT 39.130 11.550 39.430 12.000 ;
        RECT 39.130 11.400 42.980 11.550 ;
        RECT 39.130 10.950 39.430 11.400 ;
        RECT 39.130 10.800 42.980 10.950 ;
        RECT 39.130 10.350 39.430 10.800 ;
        RECT 35.530 1.450 35.680 9.650 ;
        RECT 36.130 1.450 36.280 9.650 ;
        RECT 36.730 1.450 36.880 9.650 ;
        RECT 37.330 1.450 37.480 9.650 ;
        RECT 37.930 1.450 38.080 9.650 ;
        RECT 38.530 1.450 38.680 9.650 ;
        RECT 39.130 9.200 39.430 9.650 ;
        RECT 39.130 9.050 42.980 9.200 ;
        RECT 39.130 8.600 39.430 9.050 ;
        RECT 39.130 8.450 42.980 8.600 ;
        RECT 39.130 8.000 39.430 8.450 ;
        RECT 39.130 7.850 42.980 8.000 ;
        RECT 39.130 7.400 39.430 7.850 ;
        RECT 39.130 7.250 42.980 7.400 ;
        RECT 39.130 6.800 39.430 7.250 ;
        RECT 43.830 6.800 45.630 13.200 ;
        RECT 50.030 12.750 50.330 13.200 ;
        RECT 46.480 12.600 50.330 12.750 ;
        RECT 50.030 12.150 50.330 12.600 ;
        RECT 46.480 12.000 50.330 12.150 ;
        RECT 50.030 11.550 50.330 12.000 ;
        RECT 46.480 11.400 50.330 11.550 ;
        RECT 50.030 10.950 50.330 11.400 ;
        RECT 46.480 10.800 50.330 10.950 ;
        RECT 50.030 10.350 50.330 10.800 ;
        RECT 50.780 10.350 50.930 18.550 ;
        RECT 51.380 10.350 51.530 18.550 ;
        RECT 51.980 10.350 52.130 18.550 ;
        RECT 52.580 10.350 52.730 18.550 ;
        RECT 53.180 10.350 53.330 18.550 ;
        RECT 53.780 10.350 53.930 18.550 ;
        RECT 50.030 9.200 50.330 9.650 ;
        RECT 46.480 9.050 50.330 9.200 ;
        RECT 50.030 8.600 50.330 9.050 ;
        RECT 46.480 8.450 50.330 8.600 ;
        RECT 50.030 8.000 50.330 8.450 ;
        RECT 46.480 7.850 50.330 8.000 ;
        RECT 50.030 7.400 50.330 7.850 ;
        RECT 46.480 7.250 50.330 7.400 ;
        RECT 50.030 6.800 50.330 7.250 ;
        RECT 39.130 6.650 42.980 6.800 ;
        RECT 46.480 6.650 50.330 6.800 ;
        RECT 39.130 6.200 39.430 6.650 ;
        RECT 50.030 6.200 50.330 6.650 ;
        RECT 39.130 6.050 42.980 6.200 ;
        RECT 46.480 6.050 50.330 6.200 ;
        RECT 39.130 5.600 39.430 6.050 ;
        RECT 50.030 5.600 50.330 6.050 ;
        RECT 39.130 5.450 42.980 5.600 ;
        RECT 46.480 5.450 50.330 5.600 ;
        RECT 39.130 5.000 39.430 5.450 ;
        RECT 50.030 5.000 50.330 5.450 ;
        RECT 39.130 4.850 42.980 5.000 ;
        RECT 46.480 4.850 50.330 5.000 ;
        RECT 39.130 4.400 39.430 4.850 ;
        RECT 50.030 4.400 50.330 4.850 ;
        RECT 39.130 4.250 42.980 4.400 ;
        RECT 46.480 4.250 50.330 4.400 ;
        RECT 39.130 3.800 39.430 4.250 ;
        RECT 50.030 3.800 50.330 4.250 ;
        RECT 39.130 3.650 42.980 3.800 ;
        RECT 46.480 3.650 50.330 3.800 ;
        RECT 39.130 3.200 39.430 3.650 ;
        RECT 50.030 3.200 50.330 3.650 ;
        RECT 39.130 3.050 42.980 3.200 ;
        RECT 46.480 3.050 50.330 3.200 ;
        RECT 39.130 2.600 39.430 3.050 ;
        RECT 50.030 2.600 50.330 3.050 ;
        RECT 39.130 2.450 42.980 2.600 ;
        RECT 46.480 2.450 50.330 2.600 ;
        RECT 39.130 2.000 39.430 2.450 ;
        RECT 50.030 2.000 50.330 2.450 ;
        RECT 39.130 1.450 42.930 2.000 ;
        RECT 26.530 1.400 42.930 1.450 ;
        RECT 46.530 1.450 50.330 2.000 ;
        RECT 50.780 1.450 50.930 9.650 ;
        RECT 51.380 1.450 51.530 9.650 ;
        RECT 51.980 1.450 52.130 9.650 ;
        RECT 52.580 1.450 52.730 9.650 ;
        RECT 53.180 1.450 53.330 9.650 ;
        RECT 53.780 1.450 53.930 9.650 ;
        RECT 54.380 1.450 55.080 18.550 ;
        RECT 55.530 10.350 55.680 18.550 ;
        RECT 56.130 10.350 56.280 18.550 ;
        RECT 56.730 10.350 56.880 18.550 ;
        RECT 57.330 10.350 57.480 18.550 ;
        RECT 57.930 10.350 58.080 18.550 ;
        RECT 58.530 10.350 58.680 18.550 ;
        RECT 59.130 18.000 62.930 18.550 ;
        RECT 66.530 18.550 82.930 18.600 ;
        RECT 66.530 18.000 70.330 18.550 ;
        RECT 59.130 17.550 59.430 18.000 ;
        RECT 70.030 17.550 70.330 18.000 ;
        RECT 59.130 17.400 62.980 17.550 ;
        RECT 66.480 17.400 70.330 17.550 ;
        RECT 59.130 16.950 59.430 17.400 ;
        RECT 70.030 16.950 70.330 17.400 ;
        RECT 59.130 16.800 62.980 16.950 ;
        RECT 66.480 16.800 70.330 16.950 ;
        RECT 59.130 16.350 59.430 16.800 ;
        RECT 70.030 16.350 70.330 16.800 ;
        RECT 59.130 16.200 62.980 16.350 ;
        RECT 66.480 16.200 70.330 16.350 ;
        RECT 59.130 15.750 59.430 16.200 ;
        RECT 70.030 15.750 70.330 16.200 ;
        RECT 59.130 15.600 62.980 15.750 ;
        RECT 66.480 15.600 70.330 15.750 ;
        RECT 59.130 15.150 59.430 15.600 ;
        RECT 70.030 15.150 70.330 15.600 ;
        RECT 59.130 15.000 62.980 15.150 ;
        RECT 66.480 15.000 70.330 15.150 ;
        RECT 59.130 14.550 59.430 15.000 ;
        RECT 70.030 14.550 70.330 15.000 ;
        RECT 59.130 14.400 62.980 14.550 ;
        RECT 66.480 14.400 70.330 14.550 ;
        RECT 59.130 13.950 59.430 14.400 ;
        RECT 70.030 13.950 70.330 14.400 ;
        RECT 59.130 13.800 62.980 13.950 ;
        RECT 66.480 13.800 70.330 13.950 ;
        RECT 59.130 13.350 59.430 13.800 ;
        RECT 70.030 13.350 70.330 13.800 ;
        RECT 59.130 13.200 62.980 13.350 ;
        RECT 66.480 13.200 70.330 13.350 ;
        RECT 59.130 12.750 59.430 13.200 ;
        RECT 59.130 12.600 62.980 12.750 ;
        RECT 59.130 12.150 59.430 12.600 ;
        RECT 59.130 12.000 62.980 12.150 ;
        RECT 59.130 11.550 59.430 12.000 ;
        RECT 59.130 11.400 62.980 11.550 ;
        RECT 59.130 10.950 59.430 11.400 ;
        RECT 59.130 10.800 62.980 10.950 ;
        RECT 59.130 10.350 59.430 10.800 ;
        RECT 55.530 1.450 55.680 9.650 ;
        RECT 56.130 1.450 56.280 9.650 ;
        RECT 56.730 1.450 56.880 9.650 ;
        RECT 57.330 1.450 57.480 9.650 ;
        RECT 57.930 1.450 58.080 9.650 ;
        RECT 58.530 1.450 58.680 9.650 ;
        RECT 59.130 9.200 59.430 9.650 ;
        RECT 59.130 9.050 62.980 9.200 ;
        RECT 59.130 8.600 59.430 9.050 ;
        RECT 59.130 8.450 62.980 8.600 ;
        RECT 59.130 8.000 59.430 8.450 ;
        RECT 59.130 7.850 62.980 8.000 ;
        RECT 59.130 7.400 59.430 7.850 ;
        RECT 59.130 7.250 62.980 7.400 ;
        RECT 59.130 6.800 59.430 7.250 ;
        RECT 63.830 6.800 65.630 13.200 ;
        RECT 70.030 12.750 70.330 13.200 ;
        RECT 66.480 12.600 70.330 12.750 ;
        RECT 70.030 12.150 70.330 12.600 ;
        RECT 66.480 12.000 70.330 12.150 ;
        RECT 70.030 11.550 70.330 12.000 ;
        RECT 66.480 11.400 70.330 11.550 ;
        RECT 70.030 10.950 70.330 11.400 ;
        RECT 66.480 10.800 70.330 10.950 ;
        RECT 70.030 10.350 70.330 10.800 ;
        RECT 70.780 10.350 70.930 18.550 ;
        RECT 71.380 10.350 71.530 18.550 ;
        RECT 71.980 10.350 72.130 18.550 ;
        RECT 72.580 10.350 72.730 18.550 ;
        RECT 73.180 10.350 73.330 18.550 ;
        RECT 73.780 10.350 73.930 18.550 ;
        RECT 70.030 9.200 70.330 9.650 ;
        RECT 66.480 9.050 70.330 9.200 ;
        RECT 70.030 8.600 70.330 9.050 ;
        RECT 66.480 8.450 70.330 8.600 ;
        RECT 70.030 8.000 70.330 8.450 ;
        RECT 66.480 7.850 70.330 8.000 ;
        RECT 70.030 7.400 70.330 7.850 ;
        RECT 66.480 7.250 70.330 7.400 ;
        RECT 70.030 6.800 70.330 7.250 ;
        RECT 59.130 6.650 62.980 6.800 ;
        RECT 66.480 6.650 70.330 6.800 ;
        RECT 59.130 6.200 59.430 6.650 ;
        RECT 70.030 6.200 70.330 6.650 ;
        RECT 59.130 6.050 62.980 6.200 ;
        RECT 66.480 6.050 70.330 6.200 ;
        RECT 59.130 5.600 59.430 6.050 ;
        RECT 70.030 5.600 70.330 6.050 ;
        RECT 59.130 5.450 62.980 5.600 ;
        RECT 66.480 5.450 70.330 5.600 ;
        RECT 59.130 5.000 59.430 5.450 ;
        RECT 70.030 5.000 70.330 5.450 ;
        RECT 59.130 4.850 62.980 5.000 ;
        RECT 66.480 4.850 70.330 5.000 ;
        RECT 59.130 4.400 59.430 4.850 ;
        RECT 70.030 4.400 70.330 4.850 ;
        RECT 59.130 4.250 62.980 4.400 ;
        RECT 66.480 4.250 70.330 4.400 ;
        RECT 59.130 3.800 59.430 4.250 ;
        RECT 70.030 3.800 70.330 4.250 ;
        RECT 59.130 3.650 62.980 3.800 ;
        RECT 66.480 3.650 70.330 3.800 ;
        RECT 59.130 3.200 59.430 3.650 ;
        RECT 70.030 3.200 70.330 3.650 ;
        RECT 59.130 3.050 62.980 3.200 ;
        RECT 66.480 3.050 70.330 3.200 ;
        RECT 59.130 2.600 59.430 3.050 ;
        RECT 70.030 2.600 70.330 3.050 ;
        RECT 59.130 2.450 62.980 2.600 ;
        RECT 66.480 2.450 70.330 2.600 ;
        RECT 59.130 2.000 59.430 2.450 ;
        RECT 70.030 2.000 70.330 2.450 ;
        RECT 59.130 1.450 62.930 2.000 ;
        RECT 46.530 1.400 62.930 1.450 ;
        RECT 66.530 1.450 70.330 2.000 ;
        RECT 70.780 1.450 70.930 9.650 ;
        RECT 71.380 1.450 71.530 9.650 ;
        RECT 71.980 1.450 72.130 9.650 ;
        RECT 72.580 1.450 72.730 9.650 ;
        RECT 73.180 1.450 73.330 9.650 ;
        RECT 73.780 1.450 73.930 9.650 ;
        RECT 74.380 1.450 75.080 18.550 ;
        RECT 75.530 10.350 75.680 18.550 ;
        RECT 76.130 10.350 76.280 18.550 ;
        RECT 76.730 10.350 76.880 18.550 ;
        RECT 77.330 10.350 77.480 18.550 ;
        RECT 77.930 10.350 78.080 18.550 ;
        RECT 78.530 10.350 78.680 18.550 ;
        RECT 79.130 18.000 82.930 18.550 ;
        RECT 86.530 18.550 102.930 18.600 ;
        RECT 86.530 18.000 90.330 18.550 ;
        RECT 79.130 17.550 79.430 18.000 ;
        RECT 90.030 17.550 90.330 18.000 ;
        RECT 79.130 17.400 82.980 17.550 ;
        RECT 86.480 17.400 90.330 17.550 ;
        RECT 79.130 16.950 79.430 17.400 ;
        RECT 90.030 16.950 90.330 17.400 ;
        RECT 79.130 16.800 82.980 16.950 ;
        RECT 86.480 16.800 90.330 16.950 ;
        RECT 79.130 16.350 79.430 16.800 ;
        RECT 90.030 16.350 90.330 16.800 ;
        RECT 79.130 16.200 82.980 16.350 ;
        RECT 86.480 16.200 90.330 16.350 ;
        RECT 79.130 15.750 79.430 16.200 ;
        RECT 90.030 15.750 90.330 16.200 ;
        RECT 79.130 15.600 82.980 15.750 ;
        RECT 86.480 15.600 90.330 15.750 ;
        RECT 79.130 15.150 79.430 15.600 ;
        RECT 90.030 15.150 90.330 15.600 ;
        RECT 79.130 15.000 82.980 15.150 ;
        RECT 86.480 15.000 90.330 15.150 ;
        RECT 79.130 14.550 79.430 15.000 ;
        RECT 90.030 14.550 90.330 15.000 ;
        RECT 79.130 14.400 82.980 14.550 ;
        RECT 86.480 14.400 90.330 14.550 ;
        RECT 79.130 13.950 79.430 14.400 ;
        RECT 90.030 13.950 90.330 14.400 ;
        RECT 79.130 13.800 82.980 13.950 ;
        RECT 86.480 13.800 90.330 13.950 ;
        RECT 79.130 13.350 79.430 13.800 ;
        RECT 90.030 13.350 90.330 13.800 ;
        RECT 79.130 13.200 82.980 13.350 ;
        RECT 86.480 13.200 90.330 13.350 ;
        RECT 79.130 12.750 79.430 13.200 ;
        RECT 79.130 12.600 82.980 12.750 ;
        RECT 79.130 12.150 79.430 12.600 ;
        RECT 79.130 12.000 82.980 12.150 ;
        RECT 79.130 11.550 79.430 12.000 ;
        RECT 79.130 11.400 82.980 11.550 ;
        RECT 79.130 10.950 79.430 11.400 ;
        RECT 79.130 10.800 82.980 10.950 ;
        RECT 79.130 10.350 79.430 10.800 ;
        RECT 75.530 1.450 75.680 9.650 ;
        RECT 76.130 1.450 76.280 9.650 ;
        RECT 76.730 1.450 76.880 9.650 ;
        RECT 77.330 1.450 77.480 9.650 ;
        RECT 77.930 1.450 78.080 9.650 ;
        RECT 78.530 1.450 78.680 9.650 ;
        RECT 79.130 9.200 79.430 9.650 ;
        RECT 79.130 9.050 82.980 9.200 ;
        RECT 79.130 8.600 79.430 9.050 ;
        RECT 79.130 8.450 82.980 8.600 ;
        RECT 79.130 8.000 79.430 8.450 ;
        RECT 79.130 7.850 82.980 8.000 ;
        RECT 79.130 7.400 79.430 7.850 ;
        RECT 79.130 7.250 82.980 7.400 ;
        RECT 79.130 6.800 79.430 7.250 ;
        RECT 83.830 6.800 85.630 13.200 ;
        RECT 90.030 12.750 90.330 13.200 ;
        RECT 86.480 12.600 90.330 12.750 ;
        RECT 90.030 12.150 90.330 12.600 ;
        RECT 86.480 12.000 90.330 12.150 ;
        RECT 90.030 11.550 90.330 12.000 ;
        RECT 86.480 11.400 90.330 11.550 ;
        RECT 90.030 10.950 90.330 11.400 ;
        RECT 86.480 10.800 90.330 10.950 ;
        RECT 90.030 10.350 90.330 10.800 ;
        RECT 90.780 10.350 90.930 18.550 ;
        RECT 91.380 10.350 91.530 18.550 ;
        RECT 91.980 10.350 92.130 18.550 ;
        RECT 92.580 10.350 92.730 18.550 ;
        RECT 93.180 10.350 93.330 18.550 ;
        RECT 93.780 10.350 93.930 18.550 ;
        RECT 90.030 9.200 90.330 9.650 ;
        RECT 86.480 9.050 90.330 9.200 ;
        RECT 90.030 8.600 90.330 9.050 ;
        RECT 86.480 8.450 90.330 8.600 ;
        RECT 90.030 8.000 90.330 8.450 ;
        RECT 86.480 7.850 90.330 8.000 ;
        RECT 90.030 7.400 90.330 7.850 ;
        RECT 86.480 7.250 90.330 7.400 ;
        RECT 90.030 6.800 90.330 7.250 ;
        RECT 79.130 6.650 82.980 6.800 ;
        RECT 86.480 6.650 90.330 6.800 ;
        RECT 79.130 6.200 79.430 6.650 ;
        RECT 90.030 6.200 90.330 6.650 ;
        RECT 79.130 6.050 82.980 6.200 ;
        RECT 86.480 6.050 90.330 6.200 ;
        RECT 79.130 5.600 79.430 6.050 ;
        RECT 90.030 5.600 90.330 6.050 ;
        RECT 79.130 5.450 82.980 5.600 ;
        RECT 86.480 5.450 90.330 5.600 ;
        RECT 79.130 5.000 79.430 5.450 ;
        RECT 90.030 5.000 90.330 5.450 ;
        RECT 79.130 4.850 82.980 5.000 ;
        RECT 86.480 4.850 90.330 5.000 ;
        RECT 79.130 4.400 79.430 4.850 ;
        RECT 90.030 4.400 90.330 4.850 ;
        RECT 79.130 4.250 82.980 4.400 ;
        RECT 86.480 4.250 90.330 4.400 ;
        RECT 79.130 3.800 79.430 4.250 ;
        RECT 90.030 3.800 90.330 4.250 ;
        RECT 79.130 3.650 82.980 3.800 ;
        RECT 86.480 3.650 90.330 3.800 ;
        RECT 79.130 3.200 79.430 3.650 ;
        RECT 90.030 3.200 90.330 3.650 ;
        RECT 79.130 3.050 82.980 3.200 ;
        RECT 86.480 3.050 90.330 3.200 ;
        RECT 79.130 2.600 79.430 3.050 ;
        RECT 90.030 2.600 90.330 3.050 ;
        RECT 79.130 2.450 82.980 2.600 ;
        RECT 86.480 2.450 90.330 2.600 ;
        RECT 79.130 2.000 79.430 2.450 ;
        RECT 90.030 2.000 90.330 2.450 ;
        RECT 79.130 1.450 82.930 2.000 ;
        RECT 66.530 1.400 82.930 1.450 ;
        RECT 86.530 1.450 90.330 2.000 ;
        RECT 90.780 1.450 90.930 9.650 ;
        RECT 91.380 1.450 91.530 9.650 ;
        RECT 91.980 1.450 92.130 9.650 ;
        RECT 92.580 1.450 92.730 9.650 ;
        RECT 93.180 1.450 93.330 9.650 ;
        RECT 93.780 1.450 93.930 9.650 ;
        RECT 94.380 1.450 95.080 18.550 ;
        RECT 95.530 10.350 95.680 18.550 ;
        RECT 96.130 10.350 96.280 18.550 ;
        RECT 96.730 10.350 96.880 18.550 ;
        RECT 97.330 10.350 97.480 18.550 ;
        RECT 97.930 10.350 98.080 18.550 ;
        RECT 98.530 10.350 98.680 18.550 ;
        RECT 99.130 18.000 102.930 18.550 ;
        RECT 106.530 18.550 122.930 18.600 ;
        RECT 106.530 18.000 110.330 18.550 ;
        RECT 99.130 17.550 99.430 18.000 ;
        RECT 110.030 17.550 110.330 18.000 ;
        RECT 99.130 17.400 102.980 17.550 ;
        RECT 106.480 17.400 110.330 17.550 ;
        RECT 99.130 16.950 99.430 17.400 ;
        RECT 110.030 16.950 110.330 17.400 ;
        RECT 99.130 16.800 102.980 16.950 ;
        RECT 106.480 16.800 110.330 16.950 ;
        RECT 99.130 16.350 99.430 16.800 ;
        RECT 110.030 16.350 110.330 16.800 ;
        RECT 99.130 16.200 102.980 16.350 ;
        RECT 106.480 16.200 110.330 16.350 ;
        RECT 99.130 15.750 99.430 16.200 ;
        RECT 110.030 15.750 110.330 16.200 ;
        RECT 99.130 15.600 102.980 15.750 ;
        RECT 106.480 15.600 110.330 15.750 ;
        RECT 99.130 15.150 99.430 15.600 ;
        RECT 110.030 15.150 110.330 15.600 ;
        RECT 99.130 15.000 102.980 15.150 ;
        RECT 106.480 15.000 110.330 15.150 ;
        RECT 99.130 14.550 99.430 15.000 ;
        RECT 110.030 14.550 110.330 15.000 ;
        RECT 99.130 14.400 102.980 14.550 ;
        RECT 106.480 14.400 110.330 14.550 ;
        RECT 99.130 13.950 99.430 14.400 ;
        RECT 110.030 13.950 110.330 14.400 ;
        RECT 99.130 13.800 102.980 13.950 ;
        RECT 106.480 13.800 110.330 13.950 ;
        RECT 99.130 13.350 99.430 13.800 ;
        RECT 110.030 13.350 110.330 13.800 ;
        RECT 99.130 13.200 102.980 13.350 ;
        RECT 106.480 13.200 110.330 13.350 ;
        RECT 99.130 12.750 99.430 13.200 ;
        RECT 99.130 12.600 102.980 12.750 ;
        RECT 99.130 12.150 99.430 12.600 ;
        RECT 99.130 12.000 102.980 12.150 ;
        RECT 99.130 11.550 99.430 12.000 ;
        RECT 99.130 11.400 102.980 11.550 ;
        RECT 99.130 10.950 99.430 11.400 ;
        RECT 99.130 10.800 102.980 10.950 ;
        RECT 99.130 10.350 99.430 10.800 ;
        RECT 95.530 1.450 95.680 9.650 ;
        RECT 96.130 1.450 96.280 9.650 ;
        RECT 96.730 1.450 96.880 9.650 ;
        RECT 97.330 1.450 97.480 9.650 ;
        RECT 97.930 1.450 98.080 9.650 ;
        RECT 98.530 1.450 98.680 9.650 ;
        RECT 99.130 9.200 99.430 9.650 ;
        RECT 99.130 9.050 102.980 9.200 ;
        RECT 99.130 8.600 99.430 9.050 ;
        RECT 99.130 8.450 102.980 8.600 ;
        RECT 99.130 8.000 99.430 8.450 ;
        RECT 99.130 7.850 102.980 8.000 ;
        RECT 99.130 7.400 99.430 7.850 ;
        RECT 99.130 7.250 102.980 7.400 ;
        RECT 99.130 6.800 99.430 7.250 ;
        RECT 103.830 6.800 105.630 13.200 ;
        RECT 110.030 12.750 110.330 13.200 ;
        RECT 106.480 12.600 110.330 12.750 ;
        RECT 110.030 12.150 110.330 12.600 ;
        RECT 106.480 12.000 110.330 12.150 ;
        RECT 110.030 11.550 110.330 12.000 ;
        RECT 106.480 11.400 110.330 11.550 ;
        RECT 110.030 10.950 110.330 11.400 ;
        RECT 106.480 10.800 110.330 10.950 ;
        RECT 110.030 10.350 110.330 10.800 ;
        RECT 110.780 10.350 110.930 18.550 ;
        RECT 111.380 10.350 111.530 18.550 ;
        RECT 111.980 10.350 112.130 18.550 ;
        RECT 112.580 10.350 112.730 18.550 ;
        RECT 113.180 10.350 113.330 18.550 ;
        RECT 113.780 10.350 113.930 18.550 ;
        RECT 110.030 9.200 110.330 9.650 ;
        RECT 106.480 9.050 110.330 9.200 ;
        RECT 110.030 8.600 110.330 9.050 ;
        RECT 106.480 8.450 110.330 8.600 ;
        RECT 110.030 8.000 110.330 8.450 ;
        RECT 106.480 7.850 110.330 8.000 ;
        RECT 110.030 7.400 110.330 7.850 ;
        RECT 106.480 7.250 110.330 7.400 ;
        RECT 110.030 6.800 110.330 7.250 ;
        RECT 99.130 6.650 102.980 6.800 ;
        RECT 106.480 6.650 110.330 6.800 ;
        RECT 99.130 6.200 99.430 6.650 ;
        RECT 110.030 6.200 110.330 6.650 ;
        RECT 99.130 6.050 102.980 6.200 ;
        RECT 106.480 6.050 110.330 6.200 ;
        RECT 99.130 5.600 99.430 6.050 ;
        RECT 110.030 5.600 110.330 6.050 ;
        RECT 99.130 5.450 102.980 5.600 ;
        RECT 106.480 5.450 110.330 5.600 ;
        RECT 99.130 5.000 99.430 5.450 ;
        RECT 110.030 5.000 110.330 5.450 ;
        RECT 99.130 4.850 102.980 5.000 ;
        RECT 106.480 4.850 110.330 5.000 ;
        RECT 99.130 4.400 99.430 4.850 ;
        RECT 110.030 4.400 110.330 4.850 ;
        RECT 99.130 4.250 102.980 4.400 ;
        RECT 106.480 4.250 110.330 4.400 ;
        RECT 99.130 3.800 99.430 4.250 ;
        RECT 110.030 3.800 110.330 4.250 ;
        RECT 99.130 3.650 102.980 3.800 ;
        RECT 106.480 3.650 110.330 3.800 ;
        RECT 99.130 3.200 99.430 3.650 ;
        RECT 110.030 3.200 110.330 3.650 ;
        RECT 99.130 3.050 102.980 3.200 ;
        RECT 106.480 3.050 110.330 3.200 ;
        RECT 99.130 2.600 99.430 3.050 ;
        RECT 110.030 2.600 110.330 3.050 ;
        RECT 99.130 2.450 102.980 2.600 ;
        RECT 106.480 2.450 110.330 2.600 ;
        RECT 99.130 2.000 99.430 2.450 ;
        RECT 110.030 2.000 110.330 2.450 ;
        RECT 99.130 1.450 102.930 2.000 ;
        RECT 86.530 1.400 102.930 1.450 ;
        RECT 106.530 1.450 110.330 2.000 ;
        RECT 110.780 1.450 110.930 9.650 ;
        RECT 111.380 1.450 111.530 9.650 ;
        RECT 111.980 1.450 112.130 9.650 ;
        RECT 112.580 1.450 112.730 9.650 ;
        RECT 113.180 1.450 113.330 9.650 ;
        RECT 113.780 1.450 113.930 9.650 ;
        RECT 114.380 1.450 115.080 18.550 ;
        RECT 115.530 10.350 115.680 18.550 ;
        RECT 116.130 10.350 116.280 18.550 ;
        RECT 116.730 10.350 116.880 18.550 ;
        RECT 117.330 10.350 117.480 18.550 ;
        RECT 117.930 10.350 118.080 18.550 ;
        RECT 118.530 10.350 118.680 18.550 ;
        RECT 119.130 18.000 122.930 18.550 ;
        RECT 119.130 17.550 119.430 18.000 ;
        RECT 119.130 17.400 122.980 17.550 ;
        RECT 119.130 16.950 119.430 17.400 ;
        RECT 119.130 16.800 122.980 16.950 ;
        RECT 119.130 16.350 119.430 16.800 ;
        RECT 119.130 16.200 122.980 16.350 ;
        RECT 119.130 15.750 119.430 16.200 ;
        RECT 119.130 15.600 122.980 15.750 ;
        RECT 119.130 15.150 119.430 15.600 ;
        RECT 119.130 15.000 122.980 15.150 ;
        RECT 119.130 14.550 119.430 15.000 ;
        RECT 119.130 14.400 122.980 14.550 ;
        RECT 119.130 13.950 119.430 14.400 ;
        RECT 119.130 13.800 122.980 13.950 ;
        RECT 119.130 13.350 119.430 13.800 ;
        RECT 119.130 13.200 122.980 13.350 ;
        RECT 119.130 12.750 119.430 13.200 ;
        RECT 119.130 12.600 122.980 12.750 ;
        RECT 119.130 12.150 119.430 12.600 ;
        RECT 119.130 12.000 122.980 12.150 ;
        RECT 119.130 11.550 119.430 12.000 ;
        RECT 119.130 11.400 122.980 11.550 ;
        RECT 119.130 10.950 119.430 11.400 ;
        RECT 119.130 10.800 122.980 10.950 ;
        RECT 119.130 10.350 119.430 10.800 ;
        RECT 115.530 1.450 115.680 9.650 ;
        RECT 116.130 1.450 116.280 9.650 ;
        RECT 116.730 1.450 116.880 9.650 ;
        RECT 117.330 1.450 117.480 9.650 ;
        RECT 117.930 1.450 118.080 9.650 ;
        RECT 118.530 1.450 118.680 9.650 ;
        RECT 119.130 9.200 119.430 9.650 ;
        RECT 119.130 9.050 122.980 9.200 ;
        RECT 119.130 8.600 119.430 9.050 ;
        RECT 119.130 8.450 122.980 8.600 ;
        RECT 119.130 8.000 119.430 8.450 ;
        RECT 119.130 7.850 122.980 8.000 ;
        RECT 119.130 7.400 119.430 7.850 ;
        RECT 119.130 7.250 122.980 7.400 ;
        RECT 119.130 6.800 119.430 7.250 ;
        RECT 123.830 6.800 124.730 13.200 ;
        RECT 129.850 10.250 131.850 11.525 ;
        RECT 119.130 6.650 122.980 6.800 ;
        RECT 119.130 6.200 119.430 6.650 ;
        RECT 119.130 6.050 122.980 6.200 ;
        RECT 119.130 5.600 119.430 6.050 ;
        RECT 119.130 5.450 122.980 5.600 ;
        RECT 119.130 5.000 119.430 5.450 ;
        RECT 119.130 4.850 122.980 5.000 ;
        RECT 119.130 4.400 119.430 4.850 ;
        RECT 119.130 4.250 122.980 4.400 ;
        RECT 119.130 3.800 119.430 4.250 ;
        RECT 119.130 3.650 122.980 3.800 ;
        RECT 119.130 3.200 119.430 3.650 ;
        RECT 119.130 3.050 122.980 3.200 ;
        RECT 119.130 2.600 119.430 3.050 ;
        RECT 119.130 2.450 122.980 2.600 ;
        RECT 119.130 2.000 119.430 2.450 ;
        RECT 119.130 1.450 122.930 2.000 ;
        RECT 106.530 1.400 122.930 1.450 ;
        RECT 9.630 0.900 19.830 1.400 ;
        RECT 29.630 0.900 39.830 1.400 ;
        RECT 49.630 0.900 59.830 1.400 ;
        RECT 69.630 0.900 79.830 1.400 ;
        RECT 89.630 0.900 99.830 1.400 ;
        RECT 109.630 0.900 119.830 1.400 ;
        RECT 11.530 0.000 17.930 0.900 ;
        RECT 31.530 0.000 37.930 0.900 ;
        RECT 51.530 0.000 57.930 0.900 ;
        RECT 71.530 0.000 77.930 0.900 ;
        RECT 91.530 0.000 97.930 0.900 ;
        RECT 111.530 0.000 117.930 0.900 ;
      LAYER via2 ;
        RECT 130.050 329.975 130.410 330.355 ;
        RECT 130.680 329.975 131.040 330.355 ;
        RECT 131.280 329.975 131.640 330.355 ;
        RECT 130.050 329.385 130.410 329.765 ;
        RECT 130.680 329.385 131.040 329.765 ;
        RECT 131.280 329.385 131.640 329.765 ;
        RECT 130.050 309.910 130.410 310.290 ;
        RECT 130.680 309.910 131.040 310.290 ;
        RECT 131.280 309.910 131.640 310.290 ;
        RECT 130.050 309.320 130.410 309.700 ;
        RECT 130.680 309.320 131.040 309.700 ;
        RECT 131.280 309.320 131.640 309.700 ;
        RECT 130.050 289.905 130.410 290.285 ;
        RECT 130.680 289.905 131.040 290.285 ;
        RECT 131.280 289.905 131.640 290.285 ;
        RECT 130.050 289.315 130.410 289.695 ;
        RECT 130.680 289.315 131.040 289.695 ;
        RECT 131.280 289.315 131.640 289.695 ;
        RECT 130.050 270.100 130.410 270.480 ;
        RECT 130.680 270.100 131.040 270.480 ;
        RECT 131.280 270.100 131.640 270.480 ;
        RECT 130.050 269.510 130.410 269.890 ;
        RECT 130.680 269.510 131.040 269.890 ;
        RECT 131.280 269.510 131.640 269.890 ;
        RECT 130.050 250.015 130.410 250.395 ;
        RECT 130.680 250.015 131.040 250.395 ;
        RECT 131.280 250.015 131.640 250.395 ;
        RECT 130.050 249.425 130.410 249.805 ;
        RECT 130.680 249.425 131.040 249.805 ;
        RECT 131.280 249.425 131.640 249.805 ;
        RECT 130.050 230.410 130.410 230.790 ;
        RECT 130.680 230.410 131.040 230.790 ;
        RECT 131.280 230.410 131.640 230.790 ;
        RECT 130.050 229.820 130.410 230.200 ;
        RECT 130.680 229.820 131.040 230.200 ;
        RECT 131.280 229.820 131.640 230.200 ;
        RECT 130.050 209.120 130.410 209.500 ;
        RECT 130.680 209.120 131.040 209.500 ;
        RECT 131.280 209.120 131.640 209.500 ;
        RECT 130.050 208.530 130.410 208.910 ;
        RECT 130.680 208.530 131.040 208.910 ;
        RECT 131.280 208.530 131.640 208.910 ;
        RECT 130.050 130.270 130.410 130.650 ;
        RECT 130.680 130.270 131.040 130.650 ;
        RECT 131.280 130.270 131.640 130.650 ;
        RECT 130.050 129.680 130.410 130.060 ;
        RECT 130.680 129.680 131.040 130.060 ;
        RECT 131.280 129.680 131.640 130.060 ;
        RECT 130.050 109.475 130.410 109.855 ;
        RECT 130.680 109.475 131.040 109.855 ;
        RECT 131.280 109.475 131.640 109.855 ;
        RECT 130.050 108.885 130.410 109.265 ;
        RECT 130.680 108.885 131.040 109.265 ;
        RECT 131.280 108.885 131.640 109.265 ;
        RECT 130.050 90.525 130.410 90.905 ;
        RECT 130.680 90.525 131.040 90.905 ;
        RECT 131.280 90.525 131.640 90.905 ;
        RECT 130.050 89.935 130.410 90.315 ;
        RECT 130.680 89.935 131.040 90.315 ;
        RECT 131.280 89.935 131.640 90.315 ;
        RECT 130.050 69.990 130.410 70.370 ;
        RECT 130.680 69.990 131.040 70.370 ;
        RECT 131.280 69.990 131.640 70.370 ;
        RECT 130.050 69.400 130.410 69.780 ;
        RECT 130.680 69.400 131.040 69.780 ;
        RECT 131.280 69.400 131.640 69.780 ;
        RECT 130.050 50.900 130.410 51.280 ;
        RECT 130.680 50.900 131.040 51.280 ;
        RECT 131.280 50.900 131.640 51.280 ;
        RECT 130.050 50.310 130.410 50.690 ;
        RECT 130.680 50.310 131.040 50.690 ;
        RECT 131.280 50.310 131.640 50.690 ;
        RECT 130.050 31.080 130.410 31.460 ;
        RECT 130.680 31.080 131.040 31.460 ;
        RECT 131.280 31.080 131.640 31.460 ;
        RECT 130.050 30.490 130.410 30.870 ;
        RECT 130.680 30.490 131.040 30.870 ;
        RECT 131.280 30.490 131.640 30.870 ;
        RECT 130.050 11.020 130.410 11.400 ;
        RECT 130.680 11.020 131.040 11.400 ;
        RECT 131.280 11.020 131.640 11.400 ;
        RECT 130.050 10.430 130.410 10.810 ;
        RECT 130.680 10.430 131.040 10.810 ;
        RECT 131.280 10.430 131.640 10.810 ;
      LAYER met3 ;
        RECT 129.850 329.205 131.850 330.480 ;
        RECT 129.850 309.140 131.850 310.415 ;
        RECT 129.850 289.135 131.850 290.410 ;
        RECT 129.850 269.330 131.850 270.605 ;
        RECT 129.850 249.245 131.850 250.520 ;
        RECT 129.850 229.640 131.850 230.915 ;
        RECT 129.850 208.350 131.850 209.625 ;
        RECT 129.850 129.500 131.850 130.775 ;
        RECT 129.850 108.705 131.850 109.980 ;
        RECT 129.850 89.755 131.850 91.030 ;
        RECT 129.850 69.220 131.850 70.495 ;
        RECT 129.850 50.130 131.850 51.405 ;
        RECT 129.850 30.310 131.850 31.585 ;
        RECT 129.850 10.250 131.850 11.525 ;
      LAYER via3 ;
        RECT 130.050 329.975 130.410 330.355 ;
        RECT 130.680 329.975 131.040 330.355 ;
        RECT 131.280 329.975 131.640 330.355 ;
        RECT 130.050 329.385 130.410 329.765 ;
        RECT 130.680 329.385 131.040 329.765 ;
        RECT 131.280 329.385 131.640 329.765 ;
        RECT 130.050 309.910 130.410 310.290 ;
        RECT 130.680 309.910 131.040 310.290 ;
        RECT 131.280 309.910 131.640 310.290 ;
        RECT 130.050 309.320 130.410 309.700 ;
        RECT 130.680 309.320 131.040 309.700 ;
        RECT 131.280 309.320 131.640 309.700 ;
        RECT 130.050 289.905 130.410 290.285 ;
        RECT 130.680 289.905 131.040 290.285 ;
        RECT 131.280 289.905 131.640 290.285 ;
        RECT 130.050 289.315 130.410 289.695 ;
        RECT 130.680 289.315 131.040 289.695 ;
        RECT 131.280 289.315 131.640 289.695 ;
        RECT 130.050 270.100 130.410 270.480 ;
        RECT 130.680 270.100 131.040 270.480 ;
        RECT 131.280 270.100 131.640 270.480 ;
        RECT 130.050 269.510 130.410 269.890 ;
        RECT 130.680 269.510 131.040 269.890 ;
        RECT 131.280 269.510 131.640 269.890 ;
        RECT 130.050 250.015 130.410 250.395 ;
        RECT 130.680 250.015 131.040 250.395 ;
        RECT 131.280 250.015 131.640 250.395 ;
        RECT 130.050 249.425 130.410 249.805 ;
        RECT 130.680 249.425 131.040 249.805 ;
        RECT 131.280 249.425 131.640 249.805 ;
        RECT 130.050 230.410 130.410 230.790 ;
        RECT 130.680 230.410 131.040 230.790 ;
        RECT 131.280 230.410 131.640 230.790 ;
        RECT 130.050 229.820 130.410 230.200 ;
        RECT 130.680 229.820 131.040 230.200 ;
        RECT 131.280 229.820 131.640 230.200 ;
        RECT 130.050 209.120 130.410 209.500 ;
        RECT 130.680 209.120 131.040 209.500 ;
        RECT 131.280 209.120 131.640 209.500 ;
        RECT 130.050 208.530 130.410 208.910 ;
        RECT 130.680 208.530 131.040 208.910 ;
        RECT 131.280 208.530 131.640 208.910 ;
        RECT 130.050 130.270 130.410 130.650 ;
        RECT 130.680 130.270 131.040 130.650 ;
        RECT 131.280 130.270 131.640 130.650 ;
        RECT 130.050 129.680 130.410 130.060 ;
        RECT 130.680 129.680 131.040 130.060 ;
        RECT 131.280 129.680 131.640 130.060 ;
        RECT 130.050 109.475 130.410 109.855 ;
        RECT 130.680 109.475 131.040 109.855 ;
        RECT 131.280 109.475 131.640 109.855 ;
        RECT 130.050 108.885 130.410 109.265 ;
        RECT 130.680 108.885 131.040 109.265 ;
        RECT 131.280 108.885 131.640 109.265 ;
        RECT 130.050 90.525 130.410 90.905 ;
        RECT 130.680 90.525 131.040 90.905 ;
        RECT 131.280 90.525 131.640 90.905 ;
        RECT 130.050 89.935 130.410 90.315 ;
        RECT 130.680 89.935 131.040 90.315 ;
        RECT 131.280 89.935 131.640 90.315 ;
        RECT 130.050 69.990 130.410 70.370 ;
        RECT 130.680 69.990 131.040 70.370 ;
        RECT 131.280 69.990 131.640 70.370 ;
        RECT 130.050 69.400 130.410 69.780 ;
        RECT 130.680 69.400 131.040 69.780 ;
        RECT 131.280 69.400 131.640 69.780 ;
        RECT 130.050 50.900 130.410 51.280 ;
        RECT 130.680 50.900 131.040 51.280 ;
        RECT 131.280 50.900 131.640 51.280 ;
        RECT 130.050 50.310 130.410 50.690 ;
        RECT 130.680 50.310 131.040 50.690 ;
        RECT 131.280 50.310 131.640 50.690 ;
        RECT 130.050 31.080 130.410 31.460 ;
        RECT 130.680 31.080 131.040 31.460 ;
        RECT 131.280 31.080 131.640 31.460 ;
        RECT 130.050 30.490 130.410 30.870 ;
        RECT 130.680 30.490 131.040 30.870 ;
        RECT 131.280 30.490 131.640 30.870 ;
        RECT 130.050 11.020 130.410 11.400 ;
        RECT 130.680 11.020 131.040 11.400 ;
        RECT 131.280 11.020 131.640 11.400 ;
        RECT 130.050 10.430 130.410 10.810 ;
        RECT 130.680 10.430 131.040 10.810 ;
        RECT 131.280 10.430 131.640 10.810 ;
      LAYER met4 ;
        RECT 129.850 0.000 131.850 340.000 ;
    END
  END vcm
  OBS
      LAYER pwell ;
        RECT 17.765 175.350 17.935 175.540 ;
        RECT 20.525 175.350 20.695 175.540 ;
        RECT 21.910 175.370 22.080 175.540 ;
        RECT 23.290 175.370 23.460 175.540 ;
        RECT 21.910 175.350 22.015 175.370 ;
        RECT 23.290 175.350 23.395 175.370 ;
        RECT 15.470 174.440 18.080 175.350 ;
        RECT 18.230 174.440 20.840 175.350 ;
        RECT 21.085 174.440 22.015 175.350 ;
        RECT 22.465 174.440 23.395 175.350 ;
        RECT 8.430 170.120 9.780 171.030 ;
        RECT 10.475 170.800 14.225 171.030 ;
        RECT 15.075 170.800 18.825 171.030 ;
        RECT 19.675 170.800 23.425 171.030 ;
        RECT 9.990 170.120 14.225 170.800 ;
        RECT 14.590 170.120 18.825 170.800 ;
        RECT 19.190 170.120 23.425 170.800 ;
        RECT 7.190 169.930 7.360 170.100 ;
        RECT 7.255 169.910 7.360 169.930 ;
        RECT 8.565 169.910 8.735 170.100 ;
        RECT 9.495 169.930 9.665 170.120 ;
        RECT 9.990 170.100 10.100 170.120 ;
        RECT 14.590 170.100 14.700 170.120 ;
        RECT 19.190 170.100 19.300 170.120 ;
        RECT 9.930 169.930 10.100 170.100 ;
        RECT 14.530 169.930 14.700 170.100 ;
        RECT 19.130 169.930 19.300 170.100 ;
        RECT 9.990 169.910 10.100 169.930 ;
        RECT 14.590 169.910 14.700 169.930 ;
        RECT 19.190 169.910 19.300 169.930 ;
        RECT 7.255 169.000 8.185 169.910 ;
        RECT 8.450 169.000 9.800 169.910 ;
        RECT 9.990 169.230 14.225 169.910 ;
        RECT 14.590 169.230 18.825 169.910 ;
        RECT 19.190 169.230 23.425 169.910 ;
        RECT 10.475 169.000 14.225 169.230 ;
        RECT 15.075 169.000 18.825 169.230 ;
        RECT 19.675 169.000 23.425 169.230 ;
        RECT 15.470 164.680 18.080 165.590 ;
        RECT 18.230 164.680 20.840 165.590 ;
        RECT 21.085 164.680 22.015 165.590 ;
        RECT 22.465 164.680 23.395 165.590 ;
        RECT 17.765 164.490 17.935 164.680 ;
        RECT 20.525 164.490 20.695 164.680 ;
        RECT 21.910 164.660 22.015 164.680 ;
        RECT 23.290 164.660 23.395 164.680 ;
        RECT 21.910 164.490 22.080 164.660 ;
        RECT 23.290 164.490 23.460 164.660 ;
      LAYER li1 ;
        RECT 8.250 176.115 8.980 176.645 ;
        RECT 10.960 176.115 11.135 176.185 ;
        RECT 8.250 175.945 11.135 176.115 ;
        RECT 12.695 175.980 13.425 176.680 ;
        RECT 8.810 173.450 8.980 175.450 ;
        RECT 10.960 175.390 11.135 175.945 ;
        RECT 10.965 173.440 11.135 175.390 ;
        RECT 13.190 173.445 13.360 175.980 ;
        RECT 14.425 174.730 14.755 174.910 ;
        RECT 16.060 174.720 16.230 175.200 ;
        RECT 16.900 174.720 17.070 175.200 ;
        RECT 17.740 174.720 17.910 175.200 ;
        RECT 16.060 174.550 17.070 174.720 ;
        RECT 17.275 174.550 17.910 174.720 ;
        RECT 18.820 174.720 18.990 175.200 ;
        RECT 19.660 174.720 19.830 175.200 ;
        RECT 20.500 174.720 20.670 175.200 ;
        RECT 18.820 174.550 19.830 174.720 ;
        RECT 20.035 174.550 20.670 174.720 ;
        RECT 21.175 174.570 21.505 175.200 ;
        RECT 22.555 174.570 22.885 175.200 ;
        RECT 14.500 174.180 14.865 174.350 ;
        RECT 16.060 174.010 16.555 174.550 ;
        RECT 17.275 174.380 17.445 174.550 ;
        RECT 16.945 174.210 17.445 174.380 ;
        RECT 16.060 173.840 17.070 174.010 ;
        RECT 16.060 172.990 16.230 173.840 ;
        RECT 16.900 172.990 17.070 173.840 ;
        RECT 17.275 173.970 17.445 174.210 ;
        RECT 17.615 174.140 17.995 174.380 ;
        RECT 18.820 174.010 19.315 174.550 ;
        RECT 20.035 174.380 20.205 174.550 ;
        RECT 19.705 174.210 20.205 174.380 ;
        RECT 17.275 173.800 17.990 173.970 ;
        RECT 17.660 172.990 17.990 173.800 ;
        RECT 18.820 173.840 19.830 174.010 ;
        RECT 18.820 172.990 18.990 173.840 ;
        RECT 19.660 172.990 19.830 173.840 ;
        RECT 20.035 173.970 20.205 174.210 ;
        RECT 20.375 174.140 20.755 174.380 ;
        RECT 21.175 173.970 21.405 174.570 ;
        RECT 22.555 174.380 22.785 174.570 ;
        RECT 21.575 174.140 22.785 174.380 ;
        RECT 22.955 174.145 23.315 174.380 ;
        RECT 22.955 174.140 23.285 174.145 ;
        RECT 22.555 173.970 22.785 174.140 ;
        RECT 20.035 173.800 20.750 173.970 ;
        RECT 20.420 172.990 20.750 173.800 ;
        RECT 21.175 172.990 21.505 173.970 ;
        RECT 22.555 172.990 22.885 173.970 ;
        RECT 8.940 171.500 9.270 172.480 ;
        RECT 9.890 172.055 10.330 172.480 ;
        RECT 9.890 171.885 10.885 172.055 ;
        RECT 9.035 170.900 9.205 171.500 ;
        RECT 9.375 171.070 9.710 171.340 ;
        RECT 9.890 171.010 10.380 171.715 ;
        RECT 10.550 171.340 10.885 171.885 ;
        RECT 11.055 171.690 11.325 172.480 ;
        RECT 11.495 172.055 11.745 172.480 ;
        RECT 11.495 171.860 12.300 172.055 ;
        RECT 11.055 171.510 11.780 171.690 ;
        RECT 10.550 171.010 10.960 171.340 ;
        RECT 11.130 171.010 11.780 171.510 ;
        RECT 11.950 171.340 12.300 171.860 ;
        RECT 12.470 171.690 12.720 172.480 ;
        RECT 12.890 172.055 13.160 172.480 ;
        RECT 12.890 171.860 13.715 172.055 ;
        RECT 12.470 171.510 13.195 171.690 ;
        RECT 11.950 171.010 12.375 171.340 ;
        RECT 12.545 171.010 13.195 171.510 ;
        RECT 13.365 171.340 13.715 171.860 ;
        RECT 13.885 171.715 14.320 172.480 ;
        RECT 14.490 172.055 14.930 172.480 ;
        RECT 14.490 171.885 15.485 172.055 ;
        RECT 13.885 171.510 14.980 171.715 ;
        RECT 13.365 171.010 13.790 171.340 ;
        RECT 13.960 171.010 14.980 171.510 ;
        RECT 15.150 171.340 15.485 171.885 ;
        RECT 15.655 171.690 15.925 172.480 ;
        RECT 16.095 172.055 16.345 172.480 ;
        RECT 16.095 171.860 16.900 172.055 ;
        RECT 15.655 171.510 16.380 171.690 ;
        RECT 15.150 171.010 15.560 171.340 ;
        RECT 15.730 171.010 16.380 171.510 ;
        RECT 16.550 171.340 16.900 171.860 ;
        RECT 17.070 171.690 17.320 172.480 ;
        RECT 17.490 172.055 17.760 172.480 ;
        RECT 17.490 171.860 18.315 172.055 ;
        RECT 17.070 171.510 17.795 171.690 ;
        RECT 16.550 171.010 16.975 171.340 ;
        RECT 17.145 171.010 17.795 171.510 ;
        RECT 17.965 171.340 18.315 171.860 ;
        RECT 18.485 171.715 18.920 172.480 ;
        RECT 19.090 172.055 19.530 172.480 ;
        RECT 19.090 171.885 20.085 172.055 ;
        RECT 18.485 171.510 19.580 171.715 ;
        RECT 17.965 171.010 18.390 171.340 ;
        RECT 18.560 171.010 19.580 171.510 ;
        RECT 19.750 171.340 20.085 171.885 ;
        RECT 20.255 171.690 20.525 172.480 ;
        RECT 20.695 172.055 20.945 172.480 ;
        RECT 20.695 171.860 21.500 172.055 ;
        RECT 20.255 171.510 20.980 171.690 ;
        RECT 19.750 171.010 20.160 171.340 ;
        RECT 20.330 171.010 20.980 171.510 ;
        RECT 21.150 171.340 21.500 171.860 ;
        RECT 21.670 171.690 21.920 172.480 ;
        RECT 22.090 172.055 22.360 172.480 ;
        RECT 22.090 171.860 22.915 172.055 ;
        RECT 21.670 171.510 22.395 171.690 ;
        RECT 21.150 171.010 21.575 171.340 ;
        RECT 21.745 171.010 22.395 171.510 ;
        RECT 22.565 171.340 22.915 171.860 ;
        RECT 23.085 171.510 23.520 172.480 ;
        RECT 22.565 171.010 22.990 171.340 ;
        RECT 8.510 170.270 9.205 170.900 ;
        RECT 10.550 170.840 10.885 171.010 ;
        RECT 11.130 170.840 11.325 171.010 ;
        RECT 11.950 170.840 12.300 171.010 ;
        RECT 12.545 170.840 12.720 171.010 ;
        RECT 13.365 170.840 13.715 171.010 ;
        RECT 13.960 170.840 14.320 171.010 ;
        RECT 15.150 170.840 15.485 171.010 ;
        RECT 15.730 170.840 15.925 171.010 ;
        RECT 16.550 170.840 16.900 171.010 ;
        RECT 17.145 170.840 17.320 171.010 ;
        RECT 17.965 170.840 18.315 171.010 ;
        RECT 18.560 170.840 18.920 171.010 ;
        RECT 19.750 170.840 20.085 171.010 ;
        RECT 20.330 170.840 20.525 171.010 ;
        RECT 21.150 170.840 21.500 171.010 ;
        RECT 21.745 170.840 21.920 171.010 ;
        RECT 22.565 170.840 22.915 171.010 ;
        RECT 23.160 170.840 23.520 171.510 ;
        RECT 9.890 170.670 10.885 170.840 ;
        RECT 9.890 170.270 10.330 170.670 ;
        RECT 11.055 170.270 11.325 170.840 ;
        RECT 11.495 170.670 12.300 170.840 ;
        RECT 11.495 170.270 11.745 170.670 ;
        RECT 12.470 170.270 12.720 170.840 ;
        RECT 12.890 170.670 13.715 170.840 ;
        RECT 12.890 170.270 13.160 170.670 ;
        RECT 13.885 170.270 14.320 170.840 ;
        RECT 14.490 170.670 15.485 170.840 ;
        RECT 14.490 170.270 14.930 170.670 ;
        RECT 15.655 170.270 15.925 170.840 ;
        RECT 16.095 170.670 16.900 170.840 ;
        RECT 16.095 170.270 16.345 170.670 ;
        RECT 17.070 170.270 17.320 170.840 ;
        RECT 17.490 170.670 18.315 170.840 ;
        RECT 17.490 170.270 17.760 170.670 ;
        RECT 18.485 170.270 18.920 170.840 ;
        RECT 19.090 170.670 20.085 170.840 ;
        RECT 19.090 170.270 19.530 170.670 ;
        RECT 20.255 170.270 20.525 170.840 ;
        RECT 20.695 170.670 21.500 170.840 ;
        RECT 20.695 170.270 20.945 170.670 ;
        RECT 21.670 170.270 21.920 170.840 ;
        RECT 22.090 170.670 22.915 170.840 ;
        RECT 22.090 170.270 22.360 170.670 ;
        RECT 23.085 170.270 23.520 170.840 ;
        RECT 7.765 169.130 8.095 169.760 ;
        RECT 7.865 168.940 8.095 169.130 ;
        RECT 9.025 169.130 9.720 169.760 ;
        RECT 9.890 169.360 10.330 169.760 ;
        RECT 9.890 169.190 10.885 169.360 ;
        RECT 11.055 169.190 11.325 169.760 ;
        RECT 11.495 169.360 11.745 169.760 ;
        RECT 11.495 169.190 12.300 169.360 ;
        RECT 12.470 169.190 12.720 169.760 ;
        RECT 12.890 169.360 13.160 169.760 ;
        RECT 12.890 169.190 13.715 169.360 ;
        RECT 13.885 169.190 14.320 169.760 ;
        RECT 14.490 169.360 14.930 169.760 ;
        RECT 14.490 169.190 15.485 169.360 ;
        RECT 15.655 169.190 15.925 169.760 ;
        RECT 16.095 169.360 16.345 169.760 ;
        RECT 16.095 169.190 16.900 169.360 ;
        RECT 17.070 169.190 17.320 169.760 ;
        RECT 17.490 169.360 17.760 169.760 ;
        RECT 17.490 169.190 18.315 169.360 ;
        RECT 18.485 169.190 18.920 169.760 ;
        RECT 19.090 169.360 19.530 169.760 ;
        RECT 19.090 169.190 20.085 169.360 ;
        RECT 20.255 169.190 20.525 169.760 ;
        RECT 20.695 169.360 20.945 169.760 ;
        RECT 20.695 169.190 21.500 169.360 ;
        RECT 21.670 169.190 21.920 169.760 ;
        RECT 22.090 169.360 22.360 169.760 ;
        RECT 22.090 169.190 22.915 169.360 ;
        RECT 23.085 169.190 23.520 169.760 ;
        RECT 8.520 168.940 8.855 168.960 ;
        RECT 7.865 168.725 8.855 168.940 ;
        RECT 7.865 168.530 8.095 168.725 ;
        RECT 8.520 168.690 8.855 168.725 ;
        RECT 9.025 168.530 9.195 169.130 ;
        RECT 10.550 169.020 10.885 169.190 ;
        RECT 11.130 169.020 11.325 169.190 ;
        RECT 11.950 169.020 12.300 169.190 ;
        RECT 12.545 169.020 12.720 169.190 ;
        RECT 13.365 169.020 13.715 169.190 ;
        RECT 13.960 169.020 14.320 169.190 ;
        RECT 15.150 169.020 15.485 169.190 ;
        RECT 15.730 169.020 15.925 169.190 ;
        RECT 16.550 169.020 16.900 169.190 ;
        RECT 17.145 169.020 17.320 169.190 ;
        RECT 17.965 169.020 18.315 169.190 ;
        RECT 18.560 169.020 18.920 169.190 ;
        RECT 19.750 169.020 20.085 169.190 ;
        RECT 20.330 169.020 20.525 169.190 ;
        RECT 21.150 169.020 21.500 169.190 ;
        RECT 21.745 169.020 21.920 169.190 ;
        RECT 22.565 169.020 22.915 169.190 ;
        RECT 9.365 168.690 9.700 168.940 ;
        RECT 7.765 167.550 8.095 168.530 ;
        RECT 8.960 167.550 9.290 168.530 ;
        RECT 9.890 168.315 10.380 169.020 ;
        RECT 10.550 168.690 10.960 169.020 ;
        RECT 10.550 168.145 10.885 168.690 ;
        RECT 11.130 168.520 11.780 169.020 ;
        RECT 9.890 167.975 10.885 168.145 ;
        RECT 11.055 168.340 11.780 168.520 ;
        RECT 11.950 168.690 12.375 169.020 ;
        RECT 9.890 167.550 10.330 167.975 ;
        RECT 11.055 167.550 11.325 168.340 ;
        RECT 11.950 168.170 12.300 168.690 ;
        RECT 12.545 168.520 13.195 169.020 ;
        RECT 11.495 167.975 12.300 168.170 ;
        RECT 12.470 168.340 13.195 168.520 ;
        RECT 13.365 168.690 13.790 169.020 ;
        RECT 11.495 167.550 11.745 167.975 ;
        RECT 12.470 167.550 12.720 168.340 ;
        RECT 13.365 168.170 13.715 168.690 ;
        RECT 13.960 168.520 14.980 169.020 ;
        RECT 12.890 167.975 13.715 168.170 ;
        RECT 13.885 168.315 14.980 168.520 ;
        RECT 15.150 168.690 15.560 169.020 ;
        RECT 12.890 167.550 13.160 167.975 ;
        RECT 13.885 167.550 14.320 168.315 ;
        RECT 15.150 168.145 15.485 168.690 ;
        RECT 15.730 168.520 16.380 169.020 ;
        RECT 14.490 167.975 15.485 168.145 ;
        RECT 15.655 168.340 16.380 168.520 ;
        RECT 16.550 168.690 16.975 169.020 ;
        RECT 14.490 167.550 14.930 167.975 ;
        RECT 15.655 167.550 15.925 168.340 ;
        RECT 16.550 168.170 16.900 168.690 ;
        RECT 17.145 168.520 17.795 169.020 ;
        RECT 16.095 167.975 16.900 168.170 ;
        RECT 17.070 168.340 17.795 168.520 ;
        RECT 17.965 168.690 18.390 169.020 ;
        RECT 16.095 167.550 16.345 167.975 ;
        RECT 17.070 167.550 17.320 168.340 ;
        RECT 17.965 168.170 18.315 168.690 ;
        RECT 18.560 168.520 19.580 169.020 ;
        RECT 17.490 167.975 18.315 168.170 ;
        RECT 18.485 168.315 19.580 168.520 ;
        RECT 19.750 168.690 20.160 169.020 ;
        RECT 17.490 167.550 17.760 167.975 ;
        RECT 18.485 167.550 18.920 168.315 ;
        RECT 19.750 168.145 20.085 168.690 ;
        RECT 20.330 168.520 20.980 169.020 ;
        RECT 19.090 167.975 20.085 168.145 ;
        RECT 20.255 168.340 20.980 168.520 ;
        RECT 21.150 168.690 21.575 169.020 ;
        RECT 19.090 167.550 19.530 167.975 ;
        RECT 20.255 167.550 20.525 168.340 ;
        RECT 21.150 168.170 21.500 168.690 ;
        RECT 21.745 168.520 22.395 169.020 ;
        RECT 20.695 167.975 21.500 168.170 ;
        RECT 21.670 168.340 22.395 168.520 ;
        RECT 22.565 168.690 22.990 169.020 ;
        RECT 20.695 167.550 20.945 167.975 ;
        RECT 21.670 167.550 21.920 168.340 ;
        RECT 22.565 168.170 22.915 168.690 ;
        RECT 23.160 168.520 23.520 169.190 ;
        RECT 22.090 167.975 22.915 168.170 ;
        RECT 22.090 167.550 22.360 167.975 ;
        RECT 23.085 167.550 23.520 168.520 ;
        RECT 8.400 165.935 8.695 166.875 ;
        RECT 9.785 165.145 9.955 166.585 ;
        RECT 9.730 164.605 9.955 165.145 ;
        RECT 11.365 165.145 11.535 166.585 ;
        RECT 12.185 166.275 12.355 166.585 ;
        RECT 12.180 165.145 12.355 166.275 ;
        RECT 11.365 164.605 11.590 165.145 ;
        RECT 12.115 164.605 12.355 165.145 ;
        RECT 12.975 164.190 13.145 166.585 ;
        RECT 13.765 165.145 13.935 166.585 ;
        RECT 16.060 166.190 16.230 167.040 ;
        RECT 16.900 166.190 17.070 167.040 ;
        RECT 17.660 166.230 17.990 167.040 ;
        RECT 16.060 166.020 17.070 166.190 ;
        RECT 17.275 166.060 17.990 166.230 ;
        RECT 18.820 166.190 18.990 167.040 ;
        RECT 19.660 166.190 19.830 167.040 ;
        RECT 20.420 166.230 20.750 167.040 ;
        RECT 14.720 165.690 15.060 165.860 ;
        RECT 16.060 165.480 16.555 166.020 ;
        RECT 17.275 165.820 17.445 166.060 ;
        RECT 18.820 166.020 19.830 166.190 ;
        RECT 20.035 166.060 20.750 166.230 ;
        RECT 21.175 166.060 21.505 167.040 ;
        RECT 22.555 166.060 22.885 167.040 ;
        RECT 16.945 165.650 17.445 165.820 ;
        RECT 17.615 165.650 17.995 165.890 ;
        RECT 17.275 165.480 17.445 165.650 ;
        RECT 18.820 165.480 19.315 166.020 ;
        RECT 20.035 165.820 20.205 166.060 ;
        RECT 19.705 165.650 20.205 165.820 ;
        RECT 20.375 165.650 20.755 165.890 ;
        RECT 20.035 165.480 20.205 165.650 ;
        RECT 16.060 165.310 17.070 165.480 ;
        RECT 17.275 165.310 17.910 165.480 ;
        RECT 13.765 164.640 14.000 165.145 ;
        RECT 14.565 164.935 14.780 165.290 ;
        RECT 16.060 164.830 16.230 165.310 ;
        RECT 16.900 164.830 17.070 165.310 ;
        RECT 17.740 164.830 17.910 165.310 ;
        RECT 18.820 165.310 19.830 165.480 ;
        RECT 20.035 165.310 20.670 165.480 ;
        RECT 18.820 164.830 18.990 165.310 ;
        RECT 19.660 164.830 19.830 165.310 ;
        RECT 20.500 164.830 20.670 165.310 ;
        RECT 21.175 165.460 21.405 166.060 ;
        RECT 22.555 165.890 22.785 166.060 ;
        RECT 21.575 165.650 22.785 165.890 ;
        RECT 22.955 165.655 23.305 165.890 ;
        RECT 22.955 165.650 23.285 165.655 ;
        RECT 22.555 165.460 22.785 165.650 ;
        RECT 21.175 164.830 21.505 165.460 ;
        RECT 22.555 164.830 22.885 165.460 ;
        RECT 13.765 164.190 14.395 164.640 ;
        RECT 12.690 163.515 13.425 164.190 ;
        RECT 13.760 163.535 14.495 164.190 ;
      LAYER mcon ;
        RECT 8.310 176.395 8.520 176.605 ;
        RECT 8.710 176.395 8.920 176.605 ;
        RECT 8.310 175.995 8.520 176.205 ;
        RECT 8.710 175.995 8.920 176.205 ;
        RECT 12.755 176.430 12.965 176.640 ;
        RECT 13.155 176.430 13.365 176.640 ;
        RECT 10.960 175.955 11.135 176.150 ;
        RECT 12.755 176.030 12.965 176.240 ;
        RECT 13.155 176.030 13.365 176.240 ;
        RECT 8.810 173.530 8.980 173.910 ;
        RECT 14.505 174.735 14.675 174.905 ;
        RECT 21.255 174.630 21.425 174.800 ;
        RECT 14.605 174.180 14.775 174.350 ;
        RECT 16.265 174.180 16.440 174.350 ;
        RECT 17.765 174.180 17.935 174.350 ;
        RECT 19.000 173.895 19.175 174.065 ;
        RECT 20.525 174.180 20.695 174.350 ;
        RECT 21.695 174.180 21.865 174.350 ;
        RECT 23.075 174.180 23.250 174.355 ;
        RECT 9.035 171.135 9.205 171.305 ;
        RECT 9.495 171.120 9.665 171.290 ;
        RECT 10.145 171.090 10.315 171.260 ;
        RECT 23.310 171.120 23.480 171.290 ;
        RECT 9.025 168.765 9.195 168.935 ;
        RECT 9.445 168.770 9.615 168.940 ;
        RECT 9.930 168.740 10.100 168.910 ;
        RECT 23.310 168.740 23.480 168.910 ;
        RECT 8.430 166.550 8.660 166.790 ;
        RECT 8.430 166.000 8.660 166.225 ;
        RECT 9.785 165.450 9.955 165.720 ;
        RECT 11.365 165.445 11.535 165.715 ;
        RECT 12.180 165.475 12.355 165.730 ;
        RECT 13.765 165.460 13.935 165.715 ;
        RECT 14.810 165.690 14.980 165.860 ;
        RECT 16.185 165.685 16.355 165.855 ;
        RECT 19.035 165.965 19.205 166.135 ;
        RECT 17.765 165.680 17.935 165.850 ;
        RECT 20.525 165.680 20.695 165.850 ;
        RECT 14.580 165.015 14.765 165.190 ;
        RECT 22.615 165.680 22.785 165.850 ;
        RECT 23.075 165.680 23.245 165.850 ;
        RECT 21.255 165.230 21.425 165.400 ;
        RECT 12.755 163.940 12.965 164.150 ;
        RECT 13.155 163.940 13.365 164.150 ;
        RECT 12.755 163.555 12.965 163.750 ;
        RECT 13.155 163.555 13.365 163.750 ;
        RECT 13.825 163.940 14.035 164.150 ;
        RECT 14.225 163.940 14.435 164.150 ;
        RECT 13.825 163.565 14.035 163.735 ;
        RECT 14.225 163.565 14.435 163.735 ;
      LAYER met1 ;
        RECT 8.250 176.165 8.980 176.645 ;
        RECT 10.835 176.165 11.195 176.180 ;
        RECT 8.250 175.945 11.195 176.165 ;
        RECT 12.695 175.980 13.425 176.680 ;
        RECT 10.835 175.925 11.195 175.945 ;
        RECT 14.445 174.910 14.750 174.935 ;
        RECT 14.445 174.730 16.850 174.910 ;
        RECT 14.445 174.705 14.750 174.730 ;
        RECT 14.500 174.145 16.505 174.380 ;
        RECT 7.475 173.850 7.845 173.905 ;
        RECT 8.775 173.850 9.010 173.970 ;
        RECT 16.710 173.860 16.850 174.730 ;
        RECT 18.075 174.600 21.485 174.830 ;
        RECT 17.615 174.380 17.935 174.400 ;
        RECT 18.075 174.380 18.250 174.600 ;
        RECT 20.460 174.380 20.780 174.390 ;
        RECT 23.050 174.385 23.310 174.425 ;
        RECT 17.615 174.150 18.250 174.380 ;
        RECT 20.375 174.150 21.925 174.380 ;
        RECT 17.615 174.140 17.935 174.150 ;
        RECT 20.460 174.130 20.780 174.150 ;
        RECT 23.040 174.145 23.310 174.385 ;
        RECT 18.960 173.860 19.205 174.125 ;
        RECT 23.050 174.105 23.310 174.145 ;
        RECT 7.475 173.585 9.010 173.850 ;
        RECT 16.705 173.685 19.205 173.860 ;
        RECT 8.775 173.470 9.010 173.585 ;
        RECT 18.040 171.670 18.300 171.770 ;
        RECT 9.465 171.525 18.300 171.670 ;
        RECT 9.005 171.050 9.235 171.375 ;
        RECT 9.465 171.060 9.705 171.525 ;
        RECT 18.040 171.450 18.300 171.525 ;
        RECT 9.025 170.920 9.235 171.050 ;
        RECT 10.095 171.010 10.380 171.375 ;
        RECT 23.260 171.045 23.520 171.365 ;
        RECT 10.095 170.920 10.315 171.010 ;
        RECT 9.025 170.775 10.315 170.920 ;
        RECT 17.585 169.445 17.905 169.485 ;
        RECT 9.370 169.270 17.905 169.445 ;
        RECT 8.995 168.540 9.225 169.255 ;
        RECT 9.370 168.690 9.700 169.270 ;
        RECT 17.585 169.225 17.905 169.270 ;
        RECT 9.900 168.540 10.160 168.975 ;
        RECT 23.260 168.665 23.520 168.985 ;
        RECT 8.995 168.400 10.160 168.540 ;
        RECT 8.400 165.750 8.695 166.875 ;
        RECT 16.660 166.325 19.205 166.500 ;
        RECT 8.400 165.420 11.600 165.750 ;
        RECT 12.080 165.425 14.020 165.760 ;
        RECT 14.635 165.655 16.475 165.890 ;
        RECT 8.400 165.415 8.695 165.420 ;
        RECT 9.725 165.415 11.600 165.420 ;
        RECT 16.660 165.345 16.875 166.325 ;
        RECT 19.030 166.165 19.205 166.325 ;
        RECT 17.735 165.880 18.230 165.910 ;
        RECT 19.005 165.905 19.240 166.165 ;
        RECT 17.615 165.650 18.230 165.880 ;
        RECT 14.845 165.290 16.875 165.345 ;
        RECT 14.550 165.170 16.875 165.290 ;
        RECT 18.050 165.430 18.230 165.650 ;
        RECT 20.375 165.890 20.780 165.900 ;
        RECT 20.375 165.650 22.845 165.890 ;
        RECT 20.375 165.640 20.780 165.650 ;
        RECT 23.045 165.615 23.305 165.935 ;
        RECT 18.050 165.190 21.485 165.430 ;
        RECT 14.550 165.115 14.935 165.170 ;
        RECT 14.550 164.955 14.795 165.115 ;
        RECT 12.690 163.245 13.425 164.190 ;
        RECT 13.760 163.535 14.495 164.190 ;
      LAYER via ;
        RECT 8.310 176.345 8.570 176.605 ;
        RECT 8.660 176.345 8.920 176.605 ;
        RECT 8.310 175.995 8.570 176.255 ;
        RECT 8.660 175.995 8.920 176.255 ;
        RECT 12.755 176.380 13.015 176.640 ;
        RECT 13.105 176.380 13.365 176.640 ;
        RECT 12.755 176.030 13.015 176.290 ;
        RECT 13.105 176.030 13.365 176.290 ;
        RECT 7.515 173.610 7.815 173.870 ;
        RECT 17.645 174.140 17.905 174.400 ;
        RECT 23.050 174.135 23.310 174.395 ;
        RECT 18.040 171.480 18.300 171.740 ;
        RECT 23.260 171.075 23.520 171.335 ;
        RECT 17.615 169.225 17.875 169.485 ;
        RECT 23.260 168.695 23.520 168.955 ;
        RECT 8.415 166.530 8.675 166.790 ;
        RECT 8.415 166.000 8.675 166.260 ;
        RECT 17.765 165.650 18.025 165.910 ;
        RECT 23.045 165.645 23.305 165.905 ;
        RECT 12.755 163.890 13.015 164.150 ;
        RECT 13.105 163.890 13.365 164.150 ;
        RECT 12.755 163.555 13.015 163.815 ;
        RECT 13.105 163.555 13.365 163.815 ;
        RECT 13.825 163.890 14.085 164.150 ;
        RECT 14.175 163.890 14.435 164.150 ;
        RECT 13.825 163.565 14.085 163.825 ;
        RECT 14.175 163.565 14.435 163.825 ;
      LAYER met2 ;
        RECT 8.250 178.880 11.990 179.700 ;
        RECT 8.250 178.870 11.980 178.880 ;
        RECT 7.055 175.845 7.845 176.665 ;
        RECT 8.250 175.945 8.980 178.870 ;
        RECT 16.760 178.775 17.510 179.595 ;
        RECT 16.760 178.770 17.500 178.775 ;
        RECT 7.475 173.585 7.845 175.845 ;
        RECT 8.400 165.935 8.695 175.945 ;
        RECT 12.690 162.380 13.425 176.680 ;
        RECT 13.755 176.265 14.495 176.660 ;
        RECT 13.760 163.535 14.495 176.265 ;
        RECT 16.760 175.845 17.495 178.770 ;
        RECT 17.615 174.140 17.935 174.400 ;
        RECT 17.685 169.485 17.840 174.140 ;
        RECT 23.050 174.105 23.520 174.425 ;
        RECT 18.040 171.450 18.300 171.770 ;
        RECT 17.585 169.225 17.905 169.485 ;
        RECT 18.100 165.925 18.245 171.450 ;
        RECT 23.260 171.045 23.520 174.105 ;
        RECT 23.260 165.935 23.520 168.985 ;
        RECT 17.680 165.630 18.245 165.925 ;
        RECT 23.045 165.615 23.520 165.935 ;
        RECT 12.675 162.375 13.425 162.380 ;
        RECT 12.675 161.955 13.445 162.375 ;
      LAYER via2 ;
        RECT 11.285 179.345 11.565 179.625 ;
        RECT 11.685 179.345 11.965 179.625 ;
        RECT 11.285 178.945 11.565 179.225 ;
        RECT 11.685 178.945 11.965 179.225 ;
        RECT 16.805 179.240 17.085 179.520 ;
        RECT 17.205 179.240 17.485 179.520 ;
        RECT 7.080 176.315 7.360 176.595 ;
        RECT 7.490 176.320 7.770 176.600 ;
        RECT 7.085 175.915 7.365 176.195 ;
        RECT 7.495 175.920 7.775 176.200 ;
        RECT 16.805 178.840 17.085 179.120 ;
        RECT 17.205 178.840 17.485 179.120 ;
        RECT 13.800 176.310 14.080 176.590 ;
        RECT 14.200 176.305 14.480 176.585 ;
        RECT 13.805 175.905 14.085 176.185 ;
        RECT 14.205 175.905 14.485 176.185 ;
        RECT 16.800 176.305 17.080 176.585 ;
        RECT 17.200 176.300 17.480 176.580 ;
        RECT 16.805 175.900 17.085 176.180 ;
        RECT 17.205 175.900 17.485 176.180 ;
        RECT 12.720 162.005 13.000 162.315 ;
        RECT 13.120 162.005 13.400 162.315 ;
      LAYER met3 ;
        RECT 4.730 338.750 9.130 340.000 ;
        RECT 11.530 339.150 17.930 340.000 ;
        RECT 20.330 338.750 29.130 340.000 ;
        RECT 31.530 339.150 37.930 340.000 ;
        RECT 40.330 338.750 49.130 340.000 ;
        RECT 51.530 339.150 57.930 340.000 ;
        RECT 60.330 338.750 69.130 340.000 ;
        RECT 71.530 339.150 77.930 340.000 ;
        RECT 80.330 338.750 89.130 340.000 ;
        RECT 91.530 339.150 97.930 340.000 ;
        RECT 100.330 338.750 109.130 340.000 ;
        RECT 111.530 339.150 117.930 340.000 ;
        RECT 120.330 338.750 124.730 340.000 ;
        RECT 4.730 335.600 124.730 338.750 ;
        RECT 4.730 326.800 5.580 333.200 ;
        RECT 5.980 324.400 23.480 335.600 ;
        RECT 23.880 326.800 25.580 333.200 ;
        RECT 25.980 324.400 43.480 335.600 ;
        RECT 43.880 326.800 45.580 333.200 ;
        RECT 45.980 324.400 63.480 335.600 ;
        RECT 63.880 326.800 65.580 333.200 ;
        RECT 65.980 324.400 83.480 335.600 ;
        RECT 83.880 326.800 85.580 333.200 ;
        RECT 85.980 324.400 103.480 335.600 ;
        RECT 103.880 326.800 105.580 333.200 ;
        RECT 105.980 324.400 123.480 335.600 ;
        RECT 123.880 326.800 124.730 333.200 ;
        RECT 4.730 321.250 124.730 324.400 ;
        RECT 4.730 318.750 9.130 321.250 ;
        RECT 11.530 319.150 17.930 320.850 ;
        RECT 20.330 318.750 29.130 321.250 ;
        RECT 31.530 319.150 37.930 320.850 ;
        RECT 40.330 318.750 49.130 321.250 ;
        RECT 51.530 319.150 57.930 320.850 ;
        RECT 60.330 318.750 69.130 321.250 ;
        RECT 71.530 319.150 77.930 320.850 ;
        RECT 80.330 318.750 89.130 321.250 ;
        RECT 91.530 319.150 97.930 320.850 ;
        RECT 100.330 318.750 109.130 321.250 ;
        RECT 111.530 319.150 117.930 320.850 ;
        RECT 120.330 318.750 124.730 321.250 ;
        RECT 4.730 315.600 124.730 318.750 ;
        RECT 4.730 306.800 5.580 313.200 ;
        RECT 5.980 304.400 23.480 315.600 ;
        RECT 23.880 306.800 25.580 313.200 ;
        RECT 25.980 304.400 43.480 315.600 ;
        RECT 43.880 306.800 45.580 313.200 ;
        RECT 45.980 304.400 63.480 315.600 ;
        RECT 63.880 306.800 65.580 313.200 ;
        RECT 65.980 304.400 83.480 315.600 ;
        RECT 83.880 306.800 85.580 313.200 ;
        RECT 85.980 304.400 103.480 315.600 ;
        RECT 103.880 306.800 105.580 313.200 ;
        RECT 105.980 304.400 123.480 315.600 ;
        RECT 123.880 306.800 124.730 313.200 ;
        RECT 4.730 301.250 124.730 304.400 ;
        RECT 4.730 298.750 9.130 301.250 ;
        RECT 11.530 299.150 17.930 300.850 ;
        RECT 20.330 298.750 29.130 301.250 ;
        RECT 31.530 299.150 37.930 300.850 ;
        RECT 40.330 298.750 49.130 301.250 ;
        RECT 51.530 299.150 57.930 300.850 ;
        RECT 60.330 298.750 69.130 301.250 ;
        RECT 71.530 299.150 77.930 300.850 ;
        RECT 80.330 298.750 89.130 301.250 ;
        RECT 91.530 299.150 97.930 300.850 ;
        RECT 100.330 298.750 109.130 301.250 ;
        RECT 111.530 299.150 117.930 300.850 ;
        RECT 120.330 298.750 124.730 301.250 ;
        RECT 4.730 295.600 124.730 298.750 ;
        RECT 4.730 286.800 5.580 293.200 ;
        RECT 5.980 284.400 23.480 295.600 ;
        RECT 23.880 286.800 25.580 293.200 ;
        RECT 25.980 284.400 43.480 295.600 ;
        RECT 43.880 286.800 45.580 293.200 ;
        RECT 45.980 284.400 63.480 295.600 ;
        RECT 63.880 286.800 65.580 293.200 ;
        RECT 65.980 284.400 83.480 295.600 ;
        RECT 83.880 286.800 85.580 293.200 ;
        RECT 85.980 284.400 103.480 295.600 ;
        RECT 103.880 286.800 105.580 293.200 ;
        RECT 105.980 284.400 123.480 295.600 ;
        RECT 123.880 286.800 124.730 293.200 ;
        RECT 4.730 281.250 124.730 284.400 ;
        RECT 4.730 278.750 9.130 281.250 ;
        RECT 11.530 279.150 17.930 280.850 ;
        RECT 20.330 278.750 29.130 281.250 ;
        RECT 31.530 279.150 37.930 280.850 ;
        RECT 40.330 278.750 49.130 281.250 ;
        RECT 51.530 279.150 57.930 280.850 ;
        RECT 60.330 278.750 69.130 281.250 ;
        RECT 71.530 279.150 77.930 280.850 ;
        RECT 80.330 278.750 89.130 281.250 ;
        RECT 91.530 279.150 97.930 280.850 ;
        RECT 100.330 278.750 109.130 281.250 ;
        RECT 111.530 279.150 117.930 280.850 ;
        RECT 120.330 278.750 124.730 281.250 ;
        RECT 4.730 275.600 124.730 278.750 ;
        RECT 4.730 266.800 5.580 273.200 ;
        RECT 5.980 264.400 23.480 275.600 ;
        RECT 23.880 266.800 25.580 273.200 ;
        RECT 25.980 264.400 43.480 275.600 ;
        RECT 43.880 266.800 45.580 273.200 ;
        RECT 45.980 264.400 63.480 275.600 ;
        RECT 63.880 266.800 65.580 273.200 ;
        RECT 65.980 264.400 83.480 275.600 ;
        RECT 83.880 266.800 85.580 273.200 ;
        RECT 85.980 264.400 103.480 275.600 ;
        RECT 103.880 266.800 105.580 273.200 ;
        RECT 105.980 264.400 123.480 275.600 ;
        RECT 123.880 266.800 124.730 273.200 ;
        RECT 4.730 261.250 124.730 264.400 ;
        RECT 4.730 258.750 9.130 261.250 ;
        RECT 11.530 259.150 17.930 260.850 ;
        RECT 20.330 258.750 29.130 261.250 ;
        RECT 31.530 259.150 37.930 260.850 ;
        RECT 40.330 258.750 49.130 261.250 ;
        RECT 51.530 259.150 57.930 260.850 ;
        RECT 60.330 258.750 69.130 261.250 ;
        RECT 71.530 259.150 77.930 260.850 ;
        RECT 80.330 258.750 89.130 261.250 ;
        RECT 91.530 259.150 97.930 260.850 ;
        RECT 100.330 258.750 109.130 261.250 ;
        RECT 111.530 259.150 117.930 260.850 ;
        RECT 120.330 258.750 124.730 261.250 ;
        RECT 4.730 255.600 124.730 258.750 ;
        RECT 4.730 246.800 5.580 253.200 ;
        RECT 5.980 244.400 23.480 255.600 ;
        RECT 23.880 246.800 25.580 253.200 ;
        RECT 25.980 244.400 43.480 255.600 ;
        RECT 43.880 246.800 45.580 253.200 ;
        RECT 45.980 244.400 63.480 255.600 ;
        RECT 63.880 246.800 65.580 253.200 ;
        RECT 65.980 244.400 83.480 255.600 ;
        RECT 83.880 246.800 85.580 253.200 ;
        RECT 85.980 244.400 103.480 255.600 ;
        RECT 103.880 246.800 105.580 253.200 ;
        RECT 105.980 244.400 123.480 255.600 ;
        RECT 123.880 246.800 124.730 253.200 ;
        RECT 4.730 241.250 124.730 244.400 ;
        RECT 4.730 238.750 9.130 241.250 ;
        RECT 11.530 239.150 17.930 240.850 ;
        RECT 20.330 238.750 29.130 241.250 ;
        RECT 31.530 239.150 37.930 240.850 ;
        RECT 40.330 238.750 49.130 241.250 ;
        RECT 51.530 239.150 57.930 240.850 ;
        RECT 60.330 238.750 69.130 241.250 ;
        RECT 71.530 239.150 77.930 240.850 ;
        RECT 80.330 238.750 89.130 241.250 ;
        RECT 91.530 239.150 97.930 240.850 ;
        RECT 100.330 238.750 109.130 241.250 ;
        RECT 111.530 239.150 117.930 240.850 ;
        RECT 120.330 238.750 124.730 241.250 ;
        RECT 4.730 235.600 124.730 238.750 ;
        RECT 4.730 226.800 5.580 233.200 ;
        RECT 5.980 224.400 23.480 235.600 ;
        RECT 23.880 226.800 25.580 233.200 ;
        RECT 25.980 224.400 43.480 235.600 ;
        RECT 43.880 226.800 45.580 233.200 ;
        RECT 45.980 224.400 63.480 235.600 ;
        RECT 63.880 226.800 65.580 233.200 ;
        RECT 65.980 224.400 83.480 235.600 ;
        RECT 83.880 226.800 85.580 233.200 ;
        RECT 85.980 224.400 103.480 235.600 ;
        RECT 103.880 226.800 105.580 233.200 ;
        RECT 105.980 224.400 123.480 235.600 ;
        RECT 123.880 226.800 124.730 233.200 ;
        RECT 4.730 221.250 124.730 224.400 ;
        RECT 4.730 218.750 9.130 221.250 ;
        RECT 11.530 219.150 17.930 220.850 ;
        RECT 20.330 218.750 29.130 221.250 ;
        RECT 31.530 219.150 37.930 220.850 ;
        RECT 40.330 218.750 49.130 221.250 ;
        RECT 51.530 219.150 57.930 220.850 ;
        RECT 60.330 218.750 69.130 221.250 ;
        RECT 71.530 219.150 77.930 220.850 ;
        RECT 80.330 218.750 89.130 221.250 ;
        RECT 91.530 219.150 97.930 220.850 ;
        RECT 100.330 218.750 109.130 221.250 ;
        RECT 111.530 219.150 117.930 220.850 ;
        RECT 120.330 218.750 124.730 221.250 ;
        RECT 4.730 215.600 124.730 218.750 ;
        RECT 4.730 206.800 5.580 213.200 ;
        RECT 5.980 204.400 23.480 215.600 ;
        RECT 23.880 206.800 25.580 213.200 ;
        RECT 25.980 204.400 43.480 215.600 ;
        RECT 43.880 206.800 45.580 213.200 ;
        RECT 45.980 204.400 63.480 215.600 ;
        RECT 63.880 206.800 65.580 213.200 ;
        RECT 65.980 204.400 83.480 215.600 ;
        RECT 83.880 206.800 85.580 213.200 ;
        RECT 85.980 204.400 103.480 215.600 ;
        RECT 103.880 206.800 105.580 213.200 ;
        RECT 105.980 204.400 123.480 215.600 ;
        RECT 123.880 206.800 124.730 213.200 ;
        RECT 4.730 201.250 124.730 204.400 ;
        RECT 4.730 200.000 9.130 201.250 ;
        RECT 11.530 200.000 17.930 200.850 ;
        RECT 20.330 200.000 29.130 201.250 ;
        RECT 31.530 200.000 37.930 200.850 ;
        RECT 40.330 200.000 49.130 201.250 ;
        RECT 51.530 200.000 57.930 200.850 ;
        RECT 60.330 200.000 69.130 201.250 ;
        RECT 71.530 200.000 77.930 200.850 ;
        RECT 80.330 200.000 89.130 201.250 ;
        RECT 91.530 200.000 97.930 200.850 ;
        RECT 100.330 200.000 109.130 201.250 ;
        RECT 111.530 200.000 117.930 200.850 ;
        RECT 120.330 200.000 124.730 201.250 ;
        RECT 11.240 178.875 12.005 179.700 ;
        RECT 16.760 178.770 21.725 179.600 ;
        RECT 13.445 176.665 17.510 176.670 ;
        RECT 7.055 175.845 17.510 176.665 ;
        RECT 12.675 162.375 13.440 162.380 ;
        RECT 12.675 161.955 13.445 162.375 ;
        RECT 11.530 139.150 17.930 140.000 ;
        RECT 31.530 139.150 37.930 140.000 ;
        RECT 51.530 139.150 57.930 140.000 ;
        RECT 71.530 139.150 77.930 140.000 ;
        RECT 91.530 139.150 97.930 140.000 ;
        RECT 111.530 139.150 117.930 140.000 ;
        RECT 4.730 126.800 5.580 133.200 ;
        RECT 23.880 126.800 25.580 133.200 ;
        RECT 43.880 126.800 45.580 133.200 ;
        RECT 63.880 126.800 65.580 133.200 ;
        RECT 83.880 126.800 85.580 133.200 ;
        RECT 103.880 126.800 105.580 133.200 ;
        RECT 123.880 126.800 124.730 133.200 ;
        RECT 11.530 119.150 17.930 120.850 ;
        RECT 31.530 119.150 37.930 120.850 ;
        RECT 51.530 119.150 57.930 120.850 ;
        RECT 71.530 119.150 77.930 120.850 ;
        RECT 91.530 119.150 97.930 120.850 ;
        RECT 111.530 119.150 117.930 120.850 ;
        RECT 4.730 106.800 5.580 113.200 ;
        RECT 23.880 106.800 25.580 113.200 ;
        RECT 43.880 106.800 45.580 113.200 ;
        RECT 63.880 106.800 65.580 113.200 ;
        RECT 83.880 106.800 85.580 113.200 ;
        RECT 103.880 106.800 105.580 113.200 ;
        RECT 123.880 106.800 124.730 113.200 ;
        RECT 11.530 99.150 17.930 100.850 ;
        RECT 31.530 99.150 37.930 100.850 ;
        RECT 51.530 99.150 57.930 100.850 ;
        RECT 71.530 99.150 77.930 100.850 ;
        RECT 91.530 99.150 97.930 100.850 ;
        RECT 111.530 99.150 117.930 100.850 ;
        RECT 4.730 86.800 5.580 93.200 ;
        RECT 23.880 86.800 25.580 93.200 ;
        RECT 43.880 86.800 45.580 93.200 ;
        RECT 63.880 86.800 65.580 93.200 ;
        RECT 83.880 86.800 85.580 93.200 ;
        RECT 103.880 86.800 105.580 93.200 ;
        RECT 123.880 86.800 124.730 93.200 ;
        RECT 11.530 79.150 17.930 80.850 ;
        RECT 31.530 79.150 37.930 80.850 ;
        RECT 51.530 79.150 57.930 80.850 ;
        RECT 71.530 79.150 77.930 80.850 ;
        RECT 91.530 79.150 97.930 80.850 ;
        RECT 111.530 79.150 117.930 80.850 ;
        RECT 4.730 66.800 5.580 73.200 ;
        RECT 23.880 66.800 25.580 73.200 ;
        RECT 43.880 66.800 45.580 73.200 ;
        RECT 63.880 66.800 65.580 73.200 ;
        RECT 83.880 66.800 85.580 73.200 ;
        RECT 103.880 66.800 105.580 73.200 ;
        RECT 123.880 66.800 124.730 73.200 ;
        RECT 11.530 59.150 17.930 60.850 ;
        RECT 31.530 59.150 37.930 60.850 ;
        RECT 51.530 59.150 57.930 60.850 ;
        RECT 71.530 59.150 77.930 60.850 ;
        RECT 91.530 59.150 97.930 60.850 ;
        RECT 111.530 59.150 117.930 60.850 ;
        RECT 4.730 46.800 5.580 53.200 ;
        RECT 23.880 46.800 25.580 53.200 ;
        RECT 43.880 46.800 45.580 53.200 ;
        RECT 63.880 46.800 65.580 53.200 ;
        RECT 83.880 46.800 85.580 53.200 ;
        RECT 103.880 46.800 105.580 53.200 ;
        RECT 123.880 46.800 124.730 53.200 ;
        RECT 11.530 39.150 17.930 40.850 ;
        RECT 31.530 39.150 37.930 40.850 ;
        RECT 51.530 39.150 57.930 40.850 ;
        RECT 71.530 39.150 77.930 40.850 ;
        RECT 91.530 39.150 97.930 40.850 ;
        RECT 111.530 39.150 117.930 40.850 ;
        RECT 4.730 26.800 5.580 33.200 ;
        RECT 23.880 26.800 25.580 33.200 ;
        RECT 43.880 26.800 45.580 33.200 ;
        RECT 63.880 26.800 65.580 33.200 ;
        RECT 83.880 26.800 85.580 33.200 ;
        RECT 103.880 26.800 105.580 33.200 ;
        RECT 123.880 26.800 124.730 33.200 ;
        RECT 11.530 19.150 17.930 20.850 ;
        RECT 31.530 19.150 37.930 20.850 ;
        RECT 51.530 19.150 57.930 20.850 ;
        RECT 71.530 19.150 77.930 20.850 ;
        RECT 91.530 19.150 97.930 20.850 ;
        RECT 111.530 19.150 117.930 20.850 ;
        RECT 4.730 6.800 5.580 13.200 ;
        RECT 23.880 6.800 25.580 13.200 ;
        RECT 43.880 6.800 45.580 13.200 ;
        RECT 63.880 6.800 65.580 13.200 ;
        RECT 83.880 6.800 85.580 13.200 ;
        RECT 103.880 6.800 105.580 13.200 ;
        RECT 123.880 6.800 124.730 13.200 ;
        RECT 11.530 0.000 17.930 0.850 ;
        RECT 31.530 0.000 37.930 0.850 ;
        RECT 51.530 0.000 57.930 0.850 ;
        RECT 71.530 0.000 77.930 0.850 ;
        RECT 91.530 0.000 97.930 0.850 ;
        RECT 111.530 0.000 117.930 0.850 ;
      LAYER via3 ;
        RECT 4.830 339.050 5.680 339.900 ;
        RECT 5.780 339.050 6.630 339.900 ;
        RECT 7.230 339.050 8.080 339.900 ;
        RECT 8.180 339.050 9.030 339.900 ;
        RECT 11.630 339.250 12.280 339.900 ;
        RECT 12.430 339.250 13.080 339.900 ;
        RECT 13.230 339.250 13.880 339.900 ;
        RECT 15.580 339.250 16.230 339.900 ;
        RECT 16.380 339.250 17.030 339.900 ;
        RECT 17.180 339.250 17.830 339.900 ;
        RECT 4.830 338.100 5.680 338.950 ;
        RECT 20.430 339.050 21.280 339.900 ;
        RECT 21.380 339.050 22.230 339.900 ;
        RECT 22.830 339.050 23.680 339.900 ;
        RECT 23.780 339.050 24.630 339.900 ;
        RECT 24.830 339.050 25.680 339.900 ;
        RECT 25.780 339.050 26.630 339.900 ;
        RECT 27.230 339.050 28.080 339.900 ;
        RECT 28.180 339.050 29.030 339.900 ;
        RECT 31.630 339.250 32.280 339.900 ;
        RECT 32.430 339.250 33.080 339.900 ;
        RECT 33.230 339.250 33.880 339.900 ;
        RECT 35.580 339.250 36.230 339.900 ;
        RECT 36.380 339.250 37.030 339.900 ;
        RECT 37.180 339.250 37.830 339.900 ;
        RECT 23.780 338.100 24.630 338.950 ;
        RECT 24.830 338.100 25.680 338.950 ;
        RECT 40.430 339.050 41.280 339.900 ;
        RECT 41.380 339.050 42.230 339.900 ;
        RECT 42.830 339.050 43.680 339.900 ;
        RECT 43.780 339.050 44.630 339.900 ;
        RECT 44.830 339.050 45.680 339.900 ;
        RECT 45.780 339.050 46.630 339.900 ;
        RECT 47.230 339.050 48.080 339.900 ;
        RECT 48.180 339.050 49.030 339.900 ;
        RECT 51.630 339.250 52.280 339.900 ;
        RECT 52.430 339.250 53.080 339.900 ;
        RECT 53.230 339.250 53.880 339.900 ;
        RECT 55.580 339.250 56.230 339.900 ;
        RECT 56.380 339.250 57.030 339.900 ;
        RECT 57.180 339.250 57.830 339.900 ;
        RECT 43.780 338.100 44.630 338.950 ;
        RECT 44.830 338.100 45.680 338.950 ;
        RECT 60.430 339.050 61.280 339.900 ;
        RECT 61.380 339.050 62.230 339.900 ;
        RECT 62.830 339.050 63.680 339.900 ;
        RECT 63.780 339.050 64.630 339.900 ;
        RECT 64.830 339.050 65.680 339.900 ;
        RECT 65.780 339.050 66.630 339.900 ;
        RECT 67.230 339.050 68.080 339.900 ;
        RECT 68.180 339.050 69.030 339.900 ;
        RECT 71.630 339.250 72.280 339.900 ;
        RECT 72.430 339.250 73.080 339.900 ;
        RECT 73.230 339.250 73.880 339.900 ;
        RECT 75.580 339.250 76.230 339.900 ;
        RECT 76.380 339.250 77.030 339.900 ;
        RECT 77.180 339.250 77.830 339.900 ;
        RECT 63.780 338.100 64.630 338.950 ;
        RECT 64.830 338.100 65.680 338.950 ;
        RECT 80.430 339.050 81.280 339.900 ;
        RECT 81.380 339.050 82.230 339.900 ;
        RECT 82.830 339.050 83.680 339.900 ;
        RECT 83.780 339.050 84.630 339.900 ;
        RECT 84.830 339.050 85.680 339.900 ;
        RECT 85.780 339.050 86.630 339.900 ;
        RECT 87.230 339.050 88.080 339.900 ;
        RECT 88.180 339.050 89.030 339.900 ;
        RECT 91.630 339.250 92.280 339.900 ;
        RECT 92.430 339.250 93.080 339.900 ;
        RECT 93.230 339.250 93.880 339.900 ;
        RECT 95.580 339.250 96.230 339.900 ;
        RECT 96.380 339.250 97.030 339.900 ;
        RECT 97.180 339.250 97.830 339.900 ;
        RECT 83.780 338.100 84.630 338.950 ;
        RECT 84.830 338.100 85.680 338.950 ;
        RECT 100.430 339.050 101.280 339.900 ;
        RECT 101.380 339.050 102.230 339.900 ;
        RECT 102.830 339.050 103.680 339.900 ;
        RECT 103.780 339.050 104.630 339.900 ;
        RECT 104.830 339.050 105.680 339.900 ;
        RECT 105.780 339.050 106.630 339.900 ;
        RECT 107.230 339.050 108.080 339.900 ;
        RECT 108.180 339.050 109.030 339.900 ;
        RECT 111.630 339.250 112.280 339.900 ;
        RECT 112.430 339.250 113.080 339.900 ;
        RECT 113.230 339.250 113.880 339.900 ;
        RECT 115.580 339.250 116.230 339.900 ;
        RECT 116.380 339.250 117.030 339.900 ;
        RECT 117.180 339.250 117.830 339.900 ;
        RECT 103.780 338.100 104.630 338.950 ;
        RECT 104.830 338.100 105.680 338.950 ;
        RECT 120.430 339.050 121.280 339.900 ;
        RECT 121.380 339.050 122.230 339.900 ;
        RECT 122.830 339.050 123.680 339.900 ;
        RECT 123.780 339.050 124.630 339.900 ;
        RECT 123.780 338.100 124.630 338.950 ;
        RECT 4.830 336.650 5.680 337.500 ;
        RECT 23.780 336.650 24.630 337.500 ;
        RECT 24.830 336.650 25.680 337.500 ;
        RECT 43.780 336.650 44.630 337.500 ;
        RECT 44.830 336.650 45.680 337.500 ;
        RECT 63.780 336.650 64.630 337.500 ;
        RECT 64.830 336.650 65.680 337.500 ;
        RECT 83.780 336.650 84.630 337.500 ;
        RECT 84.830 336.650 85.680 337.500 ;
        RECT 103.780 336.650 104.630 337.500 ;
        RECT 104.830 336.650 105.680 337.500 ;
        RECT 123.780 336.650 124.630 337.500 ;
        RECT 4.830 335.700 5.680 336.550 ;
        RECT 23.780 335.700 24.630 336.550 ;
        RECT 24.830 335.700 25.680 336.550 ;
        RECT 43.780 335.700 44.630 336.550 ;
        RECT 44.830 335.700 45.680 336.550 ;
        RECT 63.780 335.700 64.630 336.550 ;
        RECT 64.830 335.700 65.680 336.550 ;
        RECT 83.780 335.700 84.630 336.550 ;
        RECT 84.830 335.700 85.680 336.550 ;
        RECT 103.780 335.700 104.630 336.550 ;
        RECT 104.830 335.700 105.680 336.550 ;
        RECT 123.780 335.700 124.630 336.550 ;
        RECT 4.830 332.450 5.480 333.100 ;
        RECT 4.830 331.650 5.480 332.300 ;
        RECT 4.830 330.850 5.480 331.500 ;
        RECT 4.830 328.500 5.480 329.150 ;
        RECT 4.830 327.700 5.480 328.350 ;
        RECT 4.830 326.900 5.480 327.550 ;
        RECT 23.980 332.450 24.630 333.100 ;
        RECT 24.830 332.450 25.480 333.100 ;
        RECT 23.980 331.650 24.630 332.300 ;
        RECT 24.830 331.650 25.480 332.300 ;
        RECT 23.980 330.850 24.630 331.500 ;
        RECT 24.830 330.850 25.480 331.500 ;
        RECT 23.980 328.500 24.630 329.150 ;
        RECT 24.830 328.500 25.480 329.150 ;
        RECT 23.980 327.700 24.630 328.350 ;
        RECT 24.830 327.700 25.480 328.350 ;
        RECT 23.980 326.900 24.630 327.550 ;
        RECT 24.830 326.900 25.480 327.550 ;
        RECT 43.980 332.450 44.630 333.100 ;
        RECT 44.830 332.450 45.480 333.100 ;
        RECT 43.980 331.650 44.630 332.300 ;
        RECT 44.830 331.650 45.480 332.300 ;
        RECT 43.980 330.850 44.630 331.500 ;
        RECT 44.830 330.850 45.480 331.500 ;
        RECT 43.980 328.500 44.630 329.150 ;
        RECT 44.830 328.500 45.480 329.150 ;
        RECT 43.980 327.700 44.630 328.350 ;
        RECT 44.830 327.700 45.480 328.350 ;
        RECT 43.980 326.900 44.630 327.550 ;
        RECT 44.830 326.900 45.480 327.550 ;
        RECT 63.980 332.450 64.630 333.100 ;
        RECT 64.830 332.450 65.480 333.100 ;
        RECT 63.980 331.650 64.630 332.300 ;
        RECT 64.830 331.650 65.480 332.300 ;
        RECT 63.980 330.850 64.630 331.500 ;
        RECT 64.830 330.850 65.480 331.500 ;
        RECT 63.980 328.500 64.630 329.150 ;
        RECT 64.830 328.500 65.480 329.150 ;
        RECT 63.980 327.700 64.630 328.350 ;
        RECT 64.830 327.700 65.480 328.350 ;
        RECT 63.980 326.900 64.630 327.550 ;
        RECT 64.830 326.900 65.480 327.550 ;
        RECT 83.980 332.450 84.630 333.100 ;
        RECT 84.830 332.450 85.480 333.100 ;
        RECT 83.980 331.650 84.630 332.300 ;
        RECT 84.830 331.650 85.480 332.300 ;
        RECT 83.980 330.850 84.630 331.500 ;
        RECT 84.830 330.850 85.480 331.500 ;
        RECT 83.980 328.500 84.630 329.150 ;
        RECT 84.830 328.500 85.480 329.150 ;
        RECT 83.980 327.700 84.630 328.350 ;
        RECT 84.830 327.700 85.480 328.350 ;
        RECT 83.980 326.900 84.630 327.550 ;
        RECT 84.830 326.900 85.480 327.550 ;
        RECT 103.980 332.450 104.630 333.100 ;
        RECT 104.830 332.450 105.480 333.100 ;
        RECT 103.980 331.650 104.630 332.300 ;
        RECT 104.830 331.650 105.480 332.300 ;
        RECT 103.980 330.850 104.630 331.500 ;
        RECT 104.830 330.850 105.480 331.500 ;
        RECT 103.980 328.500 104.630 329.150 ;
        RECT 104.830 328.500 105.480 329.150 ;
        RECT 103.980 327.700 104.630 328.350 ;
        RECT 104.830 327.700 105.480 328.350 ;
        RECT 103.980 326.900 104.630 327.550 ;
        RECT 104.830 326.900 105.480 327.550 ;
        RECT 123.980 332.450 124.630 333.100 ;
        RECT 123.980 331.650 124.630 332.300 ;
        RECT 123.980 330.850 124.630 331.500 ;
        RECT 123.980 328.500 124.630 329.150 ;
        RECT 123.980 327.700 124.630 328.350 ;
        RECT 123.980 326.900 124.630 327.550 ;
        RECT 4.830 323.450 5.680 324.300 ;
        RECT 23.780 323.450 24.630 324.300 ;
        RECT 24.830 323.450 25.680 324.300 ;
        RECT 43.780 323.450 44.630 324.300 ;
        RECT 44.830 323.450 45.680 324.300 ;
        RECT 63.780 323.450 64.630 324.300 ;
        RECT 64.830 323.450 65.680 324.300 ;
        RECT 83.780 323.450 84.630 324.300 ;
        RECT 84.830 323.450 85.680 324.300 ;
        RECT 103.780 323.450 104.630 324.300 ;
        RECT 104.830 323.450 105.680 324.300 ;
        RECT 123.780 323.450 124.630 324.300 ;
        RECT 4.830 322.500 5.680 323.350 ;
        RECT 23.780 322.500 24.630 323.350 ;
        RECT 24.830 322.500 25.680 323.350 ;
        RECT 43.780 322.500 44.630 323.350 ;
        RECT 44.830 322.500 45.680 323.350 ;
        RECT 63.780 322.500 64.630 323.350 ;
        RECT 64.830 322.500 65.680 323.350 ;
        RECT 83.780 322.500 84.630 323.350 ;
        RECT 84.830 322.500 85.680 323.350 ;
        RECT 103.780 322.500 104.630 323.350 ;
        RECT 104.830 322.500 105.680 323.350 ;
        RECT 123.780 322.500 124.630 323.350 ;
        RECT 4.830 321.050 5.680 321.900 ;
        RECT 4.830 320.100 5.680 320.950 ;
        RECT 5.780 320.100 6.630 320.950 ;
        RECT 7.230 320.100 8.080 320.950 ;
        RECT 8.180 320.100 9.030 320.950 ;
        RECT 23.780 321.050 24.630 321.900 ;
        RECT 24.830 321.050 25.680 321.900 ;
        RECT 4.830 319.050 5.680 319.900 ;
        RECT 5.780 319.050 6.630 319.900 ;
        RECT 7.230 319.050 8.080 319.900 ;
        RECT 8.180 319.050 9.030 319.900 ;
        RECT 11.630 320.100 12.280 320.750 ;
        RECT 12.430 320.100 13.080 320.750 ;
        RECT 13.230 320.100 13.880 320.750 ;
        RECT 15.580 320.100 16.230 320.750 ;
        RECT 16.380 320.100 17.030 320.750 ;
        RECT 17.180 320.100 17.830 320.750 ;
        RECT 11.630 319.250 12.280 319.900 ;
        RECT 12.430 319.250 13.080 319.900 ;
        RECT 13.230 319.250 13.880 319.900 ;
        RECT 15.580 319.250 16.230 319.900 ;
        RECT 16.380 319.250 17.030 319.900 ;
        RECT 17.180 319.250 17.830 319.900 ;
        RECT 20.430 320.100 21.280 320.950 ;
        RECT 21.380 320.100 22.230 320.950 ;
        RECT 22.830 320.100 23.680 320.950 ;
        RECT 23.780 320.100 24.630 320.950 ;
        RECT 24.830 320.100 25.680 320.950 ;
        RECT 25.780 320.100 26.630 320.950 ;
        RECT 27.230 320.100 28.080 320.950 ;
        RECT 28.180 320.100 29.030 320.950 ;
        RECT 43.780 321.050 44.630 321.900 ;
        RECT 44.830 321.050 45.680 321.900 ;
        RECT 4.830 318.100 5.680 318.950 ;
        RECT 20.430 319.050 21.280 319.900 ;
        RECT 21.380 319.050 22.230 319.900 ;
        RECT 22.830 319.050 23.680 319.900 ;
        RECT 23.780 319.050 24.630 319.900 ;
        RECT 24.830 319.050 25.680 319.900 ;
        RECT 25.780 319.050 26.630 319.900 ;
        RECT 27.230 319.050 28.080 319.900 ;
        RECT 28.180 319.050 29.030 319.900 ;
        RECT 31.630 320.100 32.280 320.750 ;
        RECT 32.430 320.100 33.080 320.750 ;
        RECT 33.230 320.100 33.880 320.750 ;
        RECT 35.580 320.100 36.230 320.750 ;
        RECT 36.380 320.100 37.030 320.750 ;
        RECT 37.180 320.100 37.830 320.750 ;
        RECT 31.630 319.250 32.280 319.900 ;
        RECT 32.430 319.250 33.080 319.900 ;
        RECT 33.230 319.250 33.880 319.900 ;
        RECT 35.580 319.250 36.230 319.900 ;
        RECT 36.380 319.250 37.030 319.900 ;
        RECT 37.180 319.250 37.830 319.900 ;
        RECT 40.430 320.100 41.280 320.950 ;
        RECT 41.380 320.100 42.230 320.950 ;
        RECT 42.830 320.100 43.680 320.950 ;
        RECT 43.780 320.100 44.630 320.950 ;
        RECT 44.830 320.100 45.680 320.950 ;
        RECT 45.780 320.100 46.630 320.950 ;
        RECT 47.230 320.100 48.080 320.950 ;
        RECT 48.180 320.100 49.030 320.950 ;
        RECT 63.780 321.050 64.630 321.900 ;
        RECT 64.830 321.050 65.680 321.900 ;
        RECT 23.780 318.100 24.630 318.950 ;
        RECT 24.830 318.100 25.680 318.950 ;
        RECT 40.430 319.050 41.280 319.900 ;
        RECT 41.380 319.050 42.230 319.900 ;
        RECT 42.830 319.050 43.680 319.900 ;
        RECT 43.780 319.050 44.630 319.900 ;
        RECT 44.830 319.050 45.680 319.900 ;
        RECT 45.780 319.050 46.630 319.900 ;
        RECT 47.230 319.050 48.080 319.900 ;
        RECT 48.180 319.050 49.030 319.900 ;
        RECT 51.630 320.100 52.280 320.750 ;
        RECT 52.430 320.100 53.080 320.750 ;
        RECT 53.230 320.100 53.880 320.750 ;
        RECT 55.580 320.100 56.230 320.750 ;
        RECT 56.380 320.100 57.030 320.750 ;
        RECT 57.180 320.100 57.830 320.750 ;
        RECT 51.630 319.250 52.280 319.900 ;
        RECT 52.430 319.250 53.080 319.900 ;
        RECT 53.230 319.250 53.880 319.900 ;
        RECT 55.580 319.250 56.230 319.900 ;
        RECT 56.380 319.250 57.030 319.900 ;
        RECT 57.180 319.250 57.830 319.900 ;
        RECT 60.430 320.100 61.280 320.950 ;
        RECT 61.380 320.100 62.230 320.950 ;
        RECT 62.830 320.100 63.680 320.950 ;
        RECT 63.780 320.100 64.630 320.950 ;
        RECT 64.830 320.100 65.680 320.950 ;
        RECT 65.780 320.100 66.630 320.950 ;
        RECT 67.230 320.100 68.080 320.950 ;
        RECT 68.180 320.100 69.030 320.950 ;
        RECT 83.780 321.050 84.630 321.900 ;
        RECT 84.830 321.050 85.680 321.900 ;
        RECT 43.780 318.100 44.630 318.950 ;
        RECT 44.830 318.100 45.680 318.950 ;
        RECT 60.430 319.050 61.280 319.900 ;
        RECT 61.380 319.050 62.230 319.900 ;
        RECT 62.830 319.050 63.680 319.900 ;
        RECT 63.780 319.050 64.630 319.900 ;
        RECT 64.830 319.050 65.680 319.900 ;
        RECT 65.780 319.050 66.630 319.900 ;
        RECT 67.230 319.050 68.080 319.900 ;
        RECT 68.180 319.050 69.030 319.900 ;
        RECT 71.630 320.100 72.280 320.750 ;
        RECT 72.430 320.100 73.080 320.750 ;
        RECT 73.230 320.100 73.880 320.750 ;
        RECT 75.580 320.100 76.230 320.750 ;
        RECT 76.380 320.100 77.030 320.750 ;
        RECT 77.180 320.100 77.830 320.750 ;
        RECT 71.630 319.250 72.280 319.900 ;
        RECT 72.430 319.250 73.080 319.900 ;
        RECT 73.230 319.250 73.880 319.900 ;
        RECT 75.580 319.250 76.230 319.900 ;
        RECT 76.380 319.250 77.030 319.900 ;
        RECT 77.180 319.250 77.830 319.900 ;
        RECT 80.430 320.100 81.280 320.950 ;
        RECT 81.380 320.100 82.230 320.950 ;
        RECT 82.830 320.100 83.680 320.950 ;
        RECT 83.780 320.100 84.630 320.950 ;
        RECT 84.830 320.100 85.680 320.950 ;
        RECT 85.780 320.100 86.630 320.950 ;
        RECT 87.230 320.100 88.080 320.950 ;
        RECT 88.180 320.100 89.030 320.950 ;
        RECT 103.780 321.050 104.630 321.900 ;
        RECT 104.830 321.050 105.680 321.900 ;
        RECT 63.780 318.100 64.630 318.950 ;
        RECT 64.830 318.100 65.680 318.950 ;
        RECT 80.430 319.050 81.280 319.900 ;
        RECT 81.380 319.050 82.230 319.900 ;
        RECT 82.830 319.050 83.680 319.900 ;
        RECT 83.780 319.050 84.630 319.900 ;
        RECT 84.830 319.050 85.680 319.900 ;
        RECT 85.780 319.050 86.630 319.900 ;
        RECT 87.230 319.050 88.080 319.900 ;
        RECT 88.180 319.050 89.030 319.900 ;
        RECT 91.630 320.100 92.280 320.750 ;
        RECT 92.430 320.100 93.080 320.750 ;
        RECT 93.230 320.100 93.880 320.750 ;
        RECT 95.580 320.100 96.230 320.750 ;
        RECT 96.380 320.100 97.030 320.750 ;
        RECT 97.180 320.100 97.830 320.750 ;
        RECT 91.630 319.250 92.280 319.900 ;
        RECT 92.430 319.250 93.080 319.900 ;
        RECT 93.230 319.250 93.880 319.900 ;
        RECT 95.580 319.250 96.230 319.900 ;
        RECT 96.380 319.250 97.030 319.900 ;
        RECT 97.180 319.250 97.830 319.900 ;
        RECT 100.430 320.100 101.280 320.950 ;
        RECT 101.380 320.100 102.230 320.950 ;
        RECT 102.830 320.100 103.680 320.950 ;
        RECT 103.780 320.100 104.630 320.950 ;
        RECT 104.830 320.100 105.680 320.950 ;
        RECT 105.780 320.100 106.630 320.950 ;
        RECT 107.230 320.100 108.080 320.950 ;
        RECT 108.180 320.100 109.030 320.950 ;
        RECT 123.780 321.050 124.630 321.900 ;
        RECT 83.780 318.100 84.630 318.950 ;
        RECT 84.830 318.100 85.680 318.950 ;
        RECT 100.430 319.050 101.280 319.900 ;
        RECT 101.380 319.050 102.230 319.900 ;
        RECT 102.830 319.050 103.680 319.900 ;
        RECT 103.780 319.050 104.630 319.900 ;
        RECT 104.830 319.050 105.680 319.900 ;
        RECT 105.780 319.050 106.630 319.900 ;
        RECT 107.230 319.050 108.080 319.900 ;
        RECT 108.180 319.050 109.030 319.900 ;
        RECT 111.630 320.100 112.280 320.750 ;
        RECT 112.430 320.100 113.080 320.750 ;
        RECT 113.230 320.100 113.880 320.750 ;
        RECT 115.580 320.100 116.230 320.750 ;
        RECT 116.380 320.100 117.030 320.750 ;
        RECT 117.180 320.100 117.830 320.750 ;
        RECT 111.630 319.250 112.280 319.900 ;
        RECT 112.430 319.250 113.080 319.900 ;
        RECT 113.230 319.250 113.880 319.900 ;
        RECT 115.580 319.250 116.230 319.900 ;
        RECT 116.380 319.250 117.030 319.900 ;
        RECT 117.180 319.250 117.830 319.900 ;
        RECT 120.430 320.100 121.280 320.950 ;
        RECT 121.380 320.100 122.230 320.950 ;
        RECT 122.830 320.100 123.680 320.950 ;
        RECT 123.780 320.100 124.630 320.950 ;
        RECT 103.780 318.100 104.630 318.950 ;
        RECT 104.830 318.100 105.680 318.950 ;
        RECT 120.430 319.050 121.280 319.900 ;
        RECT 121.380 319.050 122.230 319.900 ;
        RECT 122.830 319.050 123.680 319.900 ;
        RECT 123.780 319.050 124.630 319.900 ;
        RECT 123.780 318.100 124.630 318.950 ;
        RECT 4.830 316.650 5.680 317.500 ;
        RECT 23.780 316.650 24.630 317.500 ;
        RECT 24.830 316.650 25.680 317.500 ;
        RECT 43.780 316.650 44.630 317.500 ;
        RECT 44.830 316.650 45.680 317.500 ;
        RECT 63.780 316.650 64.630 317.500 ;
        RECT 64.830 316.650 65.680 317.500 ;
        RECT 83.780 316.650 84.630 317.500 ;
        RECT 84.830 316.650 85.680 317.500 ;
        RECT 103.780 316.650 104.630 317.500 ;
        RECT 104.830 316.650 105.680 317.500 ;
        RECT 123.780 316.650 124.630 317.500 ;
        RECT 4.830 315.700 5.680 316.550 ;
        RECT 23.780 315.700 24.630 316.550 ;
        RECT 24.830 315.700 25.680 316.550 ;
        RECT 43.780 315.700 44.630 316.550 ;
        RECT 44.830 315.700 45.680 316.550 ;
        RECT 63.780 315.700 64.630 316.550 ;
        RECT 64.830 315.700 65.680 316.550 ;
        RECT 83.780 315.700 84.630 316.550 ;
        RECT 84.830 315.700 85.680 316.550 ;
        RECT 103.780 315.700 104.630 316.550 ;
        RECT 104.830 315.700 105.680 316.550 ;
        RECT 123.780 315.700 124.630 316.550 ;
        RECT 4.830 312.450 5.480 313.100 ;
        RECT 4.830 311.650 5.480 312.300 ;
        RECT 4.830 310.850 5.480 311.500 ;
        RECT 4.830 308.500 5.480 309.150 ;
        RECT 4.830 307.700 5.480 308.350 ;
        RECT 4.830 306.900 5.480 307.550 ;
        RECT 23.980 312.450 24.630 313.100 ;
        RECT 24.830 312.450 25.480 313.100 ;
        RECT 23.980 311.650 24.630 312.300 ;
        RECT 24.830 311.650 25.480 312.300 ;
        RECT 23.980 310.850 24.630 311.500 ;
        RECT 24.830 310.850 25.480 311.500 ;
        RECT 23.980 308.500 24.630 309.150 ;
        RECT 24.830 308.500 25.480 309.150 ;
        RECT 23.980 307.700 24.630 308.350 ;
        RECT 24.830 307.700 25.480 308.350 ;
        RECT 23.980 306.900 24.630 307.550 ;
        RECT 24.830 306.900 25.480 307.550 ;
        RECT 43.980 312.450 44.630 313.100 ;
        RECT 44.830 312.450 45.480 313.100 ;
        RECT 43.980 311.650 44.630 312.300 ;
        RECT 44.830 311.650 45.480 312.300 ;
        RECT 43.980 310.850 44.630 311.500 ;
        RECT 44.830 310.850 45.480 311.500 ;
        RECT 43.980 308.500 44.630 309.150 ;
        RECT 44.830 308.500 45.480 309.150 ;
        RECT 43.980 307.700 44.630 308.350 ;
        RECT 44.830 307.700 45.480 308.350 ;
        RECT 43.980 306.900 44.630 307.550 ;
        RECT 44.830 306.900 45.480 307.550 ;
        RECT 63.980 312.450 64.630 313.100 ;
        RECT 64.830 312.450 65.480 313.100 ;
        RECT 63.980 311.650 64.630 312.300 ;
        RECT 64.830 311.650 65.480 312.300 ;
        RECT 63.980 310.850 64.630 311.500 ;
        RECT 64.830 310.850 65.480 311.500 ;
        RECT 63.980 308.500 64.630 309.150 ;
        RECT 64.830 308.500 65.480 309.150 ;
        RECT 63.980 307.700 64.630 308.350 ;
        RECT 64.830 307.700 65.480 308.350 ;
        RECT 63.980 306.900 64.630 307.550 ;
        RECT 64.830 306.900 65.480 307.550 ;
        RECT 83.980 312.450 84.630 313.100 ;
        RECT 84.830 312.450 85.480 313.100 ;
        RECT 83.980 311.650 84.630 312.300 ;
        RECT 84.830 311.650 85.480 312.300 ;
        RECT 83.980 310.850 84.630 311.500 ;
        RECT 84.830 310.850 85.480 311.500 ;
        RECT 83.980 308.500 84.630 309.150 ;
        RECT 84.830 308.500 85.480 309.150 ;
        RECT 83.980 307.700 84.630 308.350 ;
        RECT 84.830 307.700 85.480 308.350 ;
        RECT 83.980 306.900 84.630 307.550 ;
        RECT 84.830 306.900 85.480 307.550 ;
        RECT 103.980 312.450 104.630 313.100 ;
        RECT 104.830 312.450 105.480 313.100 ;
        RECT 103.980 311.650 104.630 312.300 ;
        RECT 104.830 311.650 105.480 312.300 ;
        RECT 103.980 310.850 104.630 311.500 ;
        RECT 104.830 310.850 105.480 311.500 ;
        RECT 103.980 308.500 104.630 309.150 ;
        RECT 104.830 308.500 105.480 309.150 ;
        RECT 103.980 307.700 104.630 308.350 ;
        RECT 104.830 307.700 105.480 308.350 ;
        RECT 103.980 306.900 104.630 307.550 ;
        RECT 104.830 306.900 105.480 307.550 ;
        RECT 123.980 312.450 124.630 313.100 ;
        RECT 123.980 311.650 124.630 312.300 ;
        RECT 123.980 310.850 124.630 311.500 ;
        RECT 123.980 308.500 124.630 309.150 ;
        RECT 123.980 307.700 124.630 308.350 ;
        RECT 123.980 306.900 124.630 307.550 ;
        RECT 4.830 303.450 5.680 304.300 ;
        RECT 23.780 303.450 24.630 304.300 ;
        RECT 24.830 303.450 25.680 304.300 ;
        RECT 43.780 303.450 44.630 304.300 ;
        RECT 44.830 303.450 45.680 304.300 ;
        RECT 63.780 303.450 64.630 304.300 ;
        RECT 64.830 303.450 65.680 304.300 ;
        RECT 83.780 303.450 84.630 304.300 ;
        RECT 84.830 303.450 85.680 304.300 ;
        RECT 103.780 303.450 104.630 304.300 ;
        RECT 104.830 303.450 105.680 304.300 ;
        RECT 123.780 303.450 124.630 304.300 ;
        RECT 4.830 302.500 5.680 303.350 ;
        RECT 23.780 302.500 24.630 303.350 ;
        RECT 24.830 302.500 25.680 303.350 ;
        RECT 43.780 302.500 44.630 303.350 ;
        RECT 44.830 302.500 45.680 303.350 ;
        RECT 63.780 302.500 64.630 303.350 ;
        RECT 64.830 302.500 65.680 303.350 ;
        RECT 83.780 302.500 84.630 303.350 ;
        RECT 84.830 302.500 85.680 303.350 ;
        RECT 103.780 302.500 104.630 303.350 ;
        RECT 104.830 302.500 105.680 303.350 ;
        RECT 123.780 302.500 124.630 303.350 ;
        RECT 4.830 301.050 5.680 301.900 ;
        RECT 4.830 300.100 5.680 300.950 ;
        RECT 5.780 300.100 6.630 300.950 ;
        RECT 7.230 300.100 8.080 300.950 ;
        RECT 8.180 300.100 9.030 300.950 ;
        RECT 23.780 301.050 24.630 301.900 ;
        RECT 24.830 301.050 25.680 301.900 ;
        RECT 4.830 299.050 5.680 299.900 ;
        RECT 5.780 299.050 6.630 299.900 ;
        RECT 7.230 299.050 8.080 299.900 ;
        RECT 8.180 299.050 9.030 299.900 ;
        RECT 11.630 300.100 12.280 300.750 ;
        RECT 12.430 300.100 13.080 300.750 ;
        RECT 13.230 300.100 13.880 300.750 ;
        RECT 15.580 300.100 16.230 300.750 ;
        RECT 16.380 300.100 17.030 300.750 ;
        RECT 17.180 300.100 17.830 300.750 ;
        RECT 11.630 299.250 12.280 299.900 ;
        RECT 12.430 299.250 13.080 299.900 ;
        RECT 13.230 299.250 13.880 299.900 ;
        RECT 15.580 299.250 16.230 299.900 ;
        RECT 16.380 299.250 17.030 299.900 ;
        RECT 17.180 299.250 17.830 299.900 ;
        RECT 20.430 300.100 21.280 300.950 ;
        RECT 21.380 300.100 22.230 300.950 ;
        RECT 22.830 300.100 23.680 300.950 ;
        RECT 23.780 300.100 24.630 300.950 ;
        RECT 24.830 300.100 25.680 300.950 ;
        RECT 25.780 300.100 26.630 300.950 ;
        RECT 27.230 300.100 28.080 300.950 ;
        RECT 28.180 300.100 29.030 300.950 ;
        RECT 43.780 301.050 44.630 301.900 ;
        RECT 44.830 301.050 45.680 301.900 ;
        RECT 4.830 298.100 5.680 298.950 ;
        RECT 20.430 299.050 21.280 299.900 ;
        RECT 21.380 299.050 22.230 299.900 ;
        RECT 22.830 299.050 23.680 299.900 ;
        RECT 23.780 299.050 24.630 299.900 ;
        RECT 24.830 299.050 25.680 299.900 ;
        RECT 25.780 299.050 26.630 299.900 ;
        RECT 27.230 299.050 28.080 299.900 ;
        RECT 28.180 299.050 29.030 299.900 ;
        RECT 31.630 300.100 32.280 300.750 ;
        RECT 32.430 300.100 33.080 300.750 ;
        RECT 33.230 300.100 33.880 300.750 ;
        RECT 35.580 300.100 36.230 300.750 ;
        RECT 36.380 300.100 37.030 300.750 ;
        RECT 37.180 300.100 37.830 300.750 ;
        RECT 31.630 299.250 32.280 299.900 ;
        RECT 32.430 299.250 33.080 299.900 ;
        RECT 33.230 299.250 33.880 299.900 ;
        RECT 35.580 299.250 36.230 299.900 ;
        RECT 36.380 299.250 37.030 299.900 ;
        RECT 37.180 299.250 37.830 299.900 ;
        RECT 40.430 300.100 41.280 300.950 ;
        RECT 41.380 300.100 42.230 300.950 ;
        RECT 42.830 300.100 43.680 300.950 ;
        RECT 43.780 300.100 44.630 300.950 ;
        RECT 44.830 300.100 45.680 300.950 ;
        RECT 45.780 300.100 46.630 300.950 ;
        RECT 47.230 300.100 48.080 300.950 ;
        RECT 48.180 300.100 49.030 300.950 ;
        RECT 63.780 301.050 64.630 301.900 ;
        RECT 64.830 301.050 65.680 301.900 ;
        RECT 23.780 298.100 24.630 298.950 ;
        RECT 24.830 298.100 25.680 298.950 ;
        RECT 40.430 299.050 41.280 299.900 ;
        RECT 41.380 299.050 42.230 299.900 ;
        RECT 42.830 299.050 43.680 299.900 ;
        RECT 43.780 299.050 44.630 299.900 ;
        RECT 44.830 299.050 45.680 299.900 ;
        RECT 45.780 299.050 46.630 299.900 ;
        RECT 47.230 299.050 48.080 299.900 ;
        RECT 48.180 299.050 49.030 299.900 ;
        RECT 51.630 300.100 52.280 300.750 ;
        RECT 52.430 300.100 53.080 300.750 ;
        RECT 53.230 300.100 53.880 300.750 ;
        RECT 55.580 300.100 56.230 300.750 ;
        RECT 56.380 300.100 57.030 300.750 ;
        RECT 57.180 300.100 57.830 300.750 ;
        RECT 51.630 299.250 52.280 299.900 ;
        RECT 52.430 299.250 53.080 299.900 ;
        RECT 53.230 299.250 53.880 299.900 ;
        RECT 55.580 299.250 56.230 299.900 ;
        RECT 56.380 299.250 57.030 299.900 ;
        RECT 57.180 299.250 57.830 299.900 ;
        RECT 60.430 300.100 61.280 300.950 ;
        RECT 61.380 300.100 62.230 300.950 ;
        RECT 62.830 300.100 63.680 300.950 ;
        RECT 63.780 300.100 64.630 300.950 ;
        RECT 64.830 300.100 65.680 300.950 ;
        RECT 65.780 300.100 66.630 300.950 ;
        RECT 67.230 300.100 68.080 300.950 ;
        RECT 68.180 300.100 69.030 300.950 ;
        RECT 83.780 301.050 84.630 301.900 ;
        RECT 84.830 301.050 85.680 301.900 ;
        RECT 43.780 298.100 44.630 298.950 ;
        RECT 44.830 298.100 45.680 298.950 ;
        RECT 60.430 299.050 61.280 299.900 ;
        RECT 61.380 299.050 62.230 299.900 ;
        RECT 62.830 299.050 63.680 299.900 ;
        RECT 63.780 299.050 64.630 299.900 ;
        RECT 64.830 299.050 65.680 299.900 ;
        RECT 65.780 299.050 66.630 299.900 ;
        RECT 67.230 299.050 68.080 299.900 ;
        RECT 68.180 299.050 69.030 299.900 ;
        RECT 71.630 300.100 72.280 300.750 ;
        RECT 72.430 300.100 73.080 300.750 ;
        RECT 73.230 300.100 73.880 300.750 ;
        RECT 75.580 300.100 76.230 300.750 ;
        RECT 76.380 300.100 77.030 300.750 ;
        RECT 77.180 300.100 77.830 300.750 ;
        RECT 71.630 299.250 72.280 299.900 ;
        RECT 72.430 299.250 73.080 299.900 ;
        RECT 73.230 299.250 73.880 299.900 ;
        RECT 75.580 299.250 76.230 299.900 ;
        RECT 76.380 299.250 77.030 299.900 ;
        RECT 77.180 299.250 77.830 299.900 ;
        RECT 80.430 300.100 81.280 300.950 ;
        RECT 81.380 300.100 82.230 300.950 ;
        RECT 82.830 300.100 83.680 300.950 ;
        RECT 83.780 300.100 84.630 300.950 ;
        RECT 84.830 300.100 85.680 300.950 ;
        RECT 85.780 300.100 86.630 300.950 ;
        RECT 87.230 300.100 88.080 300.950 ;
        RECT 88.180 300.100 89.030 300.950 ;
        RECT 103.780 301.050 104.630 301.900 ;
        RECT 104.830 301.050 105.680 301.900 ;
        RECT 63.780 298.100 64.630 298.950 ;
        RECT 64.830 298.100 65.680 298.950 ;
        RECT 80.430 299.050 81.280 299.900 ;
        RECT 81.380 299.050 82.230 299.900 ;
        RECT 82.830 299.050 83.680 299.900 ;
        RECT 83.780 299.050 84.630 299.900 ;
        RECT 84.830 299.050 85.680 299.900 ;
        RECT 85.780 299.050 86.630 299.900 ;
        RECT 87.230 299.050 88.080 299.900 ;
        RECT 88.180 299.050 89.030 299.900 ;
        RECT 91.630 300.100 92.280 300.750 ;
        RECT 92.430 300.100 93.080 300.750 ;
        RECT 93.230 300.100 93.880 300.750 ;
        RECT 95.580 300.100 96.230 300.750 ;
        RECT 96.380 300.100 97.030 300.750 ;
        RECT 97.180 300.100 97.830 300.750 ;
        RECT 91.630 299.250 92.280 299.900 ;
        RECT 92.430 299.250 93.080 299.900 ;
        RECT 93.230 299.250 93.880 299.900 ;
        RECT 95.580 299.250 96.230 299.900 ;
        RECT 96.380 299.250 97.030 299.900 ;
        RECT 97.180 299.250 97.830 299.900 ;
        RECT 100.430 300.100 101.280 300.950 ;
        RECT 101.380 300.100 102.230 300.950 ;
        RECT 102.830 300.100 103.680 300.950 ;
        RECT 103.780 300.100 104.630 300.950 ;
        RECT 104.830 300.100 105.680 300.950 ;
        RECT 105.780 300.100 106.630 300.950 ;
        RECT 107.230 300.100 108.080 300.950 ;
        RECT 108.180 300.100 109.030 300.950 ;
        RECT 123.780 301.050 124.630 301.900 ;
        RECT 83.780 298.100 84.630 298.950 ;
        RECT 84.830 298.100 85.680 298.950 ;
        RECT 100.430 299.050 101.280 299.900 ;
        RECT 101.380 299.050 102.230 299.900 ;
        RECT 102.830 299.050 103.680 299.900 ;
        RECT 103.780 299.050 104.630 299.900 ;
        RECT 104.830 299.050 105.680 299.900 ;
        RECT 105.780 299.050 106.630 299.900 ;
        RECT 107.230 299.050 108.080 299.900 ;
        RECT 108.180 299.050 109.030 299.900 ;
        RECT 111.630 300.100 112.280 300.750 ;
        RECT 112.430 300.100 113.080 300.750 ;
        RECT 113.230 300.100 113.880 300.750 ;
        RECT 115.580 300.100 116.230 300.750 ;
        RECT 116.380 300.100 117.030 300.750 ;
        RECT 117.180 300.100 117.830 300.750 ;
        RECT 111.630 299.250 112.280 299.900 ;
        RECT 112.430 299.250 113.080 299.900 ;
        RECT 113.230 299.250 113.880 299.900 ;
        RECT 115.580 299.250 116.230 299.900 ;
        RECT 116.380 299.250 117.030 299.900 ;
        RECT 117.180 299.250 117.830 299.900 ;
        RECT 120.430 300.100 121.280 300.950 ;
        RECT 121.380 300.100 122.230 300.950 ;
        RECT 122.830 300.100 123.680 300.950 ;
        RECT 123.780 300.100 124.630 300.950 ;
        RECT 103.780 298.100 104.630 298.950 ;
        RECT 104.830 298.100 105.680 298.950 ;
        RECT 120.430 299.050 121.280 299.900 ;
        RECT 121.380 299.050 122.230 299.900 ;
        RECT 122.830 299.050 123.680 299.900 ;
        RECT 123.780 299.050 124.630 299.900 ;
        RECT 123.780 298.100 124.630 298.950 ;
        RECT 4.830 296.650 5.680 297.500 ;
        RECT 23.780 296.650 24.630 297.500 ;
        RECT 24.830 296.650 25.680 297.500 ;
        RECT 43.780 296.650 44.630 297.500 ;
        RECT 44.830 296.650 45.680 297.500 ;
        RECT 63.780 296.650 64.630 297.500 ;
        RECT 64.830 296.650 65.680 297.500 ;
        RECT 83.780 296.650 84.630 297.500 ;
        RECT 84.830 296.650 85.680 297.500 ;
        RECT 103.780 296.650 104.630 297.500 ;
        RECT 104.830 296.650 105.680 297.500 ;
        RECT 123.780 296.650 124.630 297.500 ;
        RECT 4.830 295.700 5.680 296.550 ;
        RECT 23.780 295.700 24.630 296.550 ;
        RECT 24.830 295.700 25.680 296.550 ;
        RECT 43.780 295.700 44.630 296.550 ;
        RECT 44.830 295.700 45.680 296.550 ;
        RECT 63.780 295.700 64.630 296.550 ;
        RECT 64.830 295.700 65.680 296.550 ;
        RECT 83.780 295.700 84.630 296.550 ;
        RECT 84.830 295.700 85.680 296.550 ;
        RECT 103.780 295.700 104.630 296.550 ;
        RECT 104.830 295.700 105.680 296.550 ;
        RECT 123.780 295.700 124.630 296.550 ;
        RECT 4.830 292.450 5.480 293.100 ;
        RECT 4.830 291.650 5.480 292.300 ;
        RECT 4.830 290.850 5.480 291.500 ;
        RECT 4.830 288.500 5.480 289.150 ;
        RECT 4.830 287.700 5.480 288.350 ;
        RECT 4.830 286.900 5.480 287.550 ;
        RECT 23.980 292.450 24.630 293.100 ;
        RECT 24.830 292.450 25.480 293.100 ;
        RECT 23.980 291.650 24.630 292.300 ;
        RECT 24.830 291.650 25.480 292.300 ;
        RECT 23.980 290.850 24.630 291.500 ;
        RECT 24.830 290.850 25.480 291.500 ;
        RECT 23.980 288.500 24.630 289.150 ;
        RECT 24.830 288.500 25.480 289.150 ;
        RECT 23.980 287.700 24.630 288.350 ;
        RECT 24.830 287.700 25.480 288.350 ;
        RECT 23.980 286.900 24.630 287.550 ;
        RECT 24.830 286.900 25.480 287.550 ;
        RECT 43.980 292.450 44.630 293.100 ;
        RECT 44.830 292.450 45.480 293.100 ;
        RECT 43.980 291.650 44.630 292.300 ;
        RECT 44.830 291.650 45.480 292.300 ;
        RECT 43.980 290.850 44.630 291.500 ;
        RECT 44.830 290.850 45.480 291.500 ;
        RECT 43.980 288.500 44.630 289.150 ;
        RECT 44.830 288.500 45.480 289.150 ;
        RECT 43.980 287.700 44.630 288.350 ;
        RECT 44.830 287.700 45.480 288.350 ;
        RECT 43.980 286.900 44.630 287.550 ;
        RECT 44.830 286.900 45.480 287.550 ;
        RECT 63.980 292.450 64.630 293.100 ;
        RECT 64.830 292.450 65.480 293.100 ;
        RECT 63.980 291.650 64.630 292.300 ;
        RECT 64.830 291.650 65.480 292.300 ;
        RECT 63.980 290.850 64.630 291.500 ;
        RECT 64.830 290.850 65.480 291.500 ;
        RECT 63.980 288.500 64.630 289.150 ;
        RECT 64.830 288.500 65.480 289.150 ;
        RECT 63.980 287.700 64.630 288.350 ;
        RECT 64.830 287.700 65.480 288.350 ;
        RECT 63.980 286.900 64.630 287.550 ;
        RECT 64.830 286.900 65.480 287.550 ;
        RECT 83.980 292.450 84.630 293.100 ;
        RECT 84.830 292.450 85.480 293.100 ;
        RECT 83.980 291.650 84.630 292.300 ;
        RECT 84.830 291.650 85.480 292.300 ;
        RECT 83.980 290.850 84.630 291.500 ;
        RECT 84.830 290.850 85.480 291.500 ;
        RECT 83.980 288.500 84.630 289.150 ;
        RECT 84.830 288.500 85.480 289.150 ;
        RECT 83.980 287.700 84.630 288.350 ;
        RECT 84.830 287.700 85.480 288.350 ;
        RECT 83.980 286.900 84.630 287.550 ;
        RECT 84.830 286.900 85.480 287.550 ;
        RECT 103.980 292.450 104.630 293.100 ;
        RECT 104.830 292.450 105.480 293.100 ;
        RECT 103.980 291.650 104.630 292.300 ;
        RECT 104.830 291.650 105.480 292.300 ;
        RECT 103.980 290.850 104.630 291.500 ;
        RECT 104.830 290.850 105.480 291.500 ;
        RECT 103.980 288.500 104.630 289.150 ;
        RECT 104.830 288.500 105.480 289.150 ;
        RECT 103.980 287.700 104.630 288.350 ;
        RECT 104.830 287.700 105.480 288.350 ;
        RECT 103.980 286.900 104.630 287.550 ;
        RECT 104.830 286.900 105.480 287.550 ;
        RECT 123.980 292.450 124.630 293.100 ;
        RECT 123.980 291.650 124.630 292.300 ;
        RECT 123.980 290.850 124.630 291.500 ;
        RECT 123.980 288.500 124.630 289.150 ;
        RECT 123.980 287.700 124.630 288.350 ;
        RECT 123.980 286.900 124.630 287.550 ;
        RECT 4.830 283.450 5.680 284.300 ;
        RECT 23.780 283.450 24.630 284.300 ;
        RECT 24.830 283.450 25.680 284.300 ;
        RECT 43.780 283.450 44.630 284.300 ;
        RECT 44.830 283.450 45.680 284.300 ;
        RECT 63.780 283.450 64.630 284.300 ;
        RECT 64.830 283.450 65.680 284.300 ;
        RECT 83.780 283.450 84.630 284.300 ;
        RECT 84.830 283.450 85.680 284.300 ;
        RECT 103.780 283.450 104.630 284.300 ;
        RECT 104.830 283.450 105.680 284.300 ;
        RECT 123.780 283.450 124.630 284.300 ;
        RECT 4.830 282.500 5.680 283.350 ;
        RECT 23.780 282.500 24.630 283.350 ;
        RECT 24.830 282.500 25.680 283.350 ;
        RECT 43.780 282.500 44.630 283.350 ;
        RECT 44.830 282.500 45.680 283.350 ;
        RECT 63.780 282.500 64.630 283.350 ;
        RECT 64.830 282.500 65.680 283.350 ;
        RECT 83.780 282.500 84.630 283.350 ;
        RECT 84.830 282.500 85.680 283.350 ;
        RECT 103.780 282.500 104.630 283.350 ;
        RECT 104.830 282.500 105.680 283.350 ;
        RECT 123.780 282.500 124.630 283.350 ;
        RECT 4.830 281.050 5.680 281.900 ;
        RECT 4.830 280.100 5.680 280.950 ;
        RECT 5.780 280.100 6.630 280.950 ;
        RECT 7.230 280.100 8.080 280.950 ;
        RECT 8.180 280.100 9.030 280.950 ;
        RECT 23.780 281.050 24.630 281.900 ;
        RECT 24.830 281.050 25.680 281.900 ;
        RECT 4.830 279.050 5.680 279.900 ;
        RECT 5.780 279.050 6.630 279.900 ;
        RECT 7.230 279.050 8.080 279.900 ;
        RECT 8.180 279.050 9.030 279.900 ;
        RECT 11.630 280.100 12.280 280.750 ;
        RECT 12.430 280.100 13.080 280.750 ;
        RECT 13.230 280.100 13.880 280.750 ;
        RECT 15.580 280.100 16.230 280.750 ;
        RECT 16.380 280.100 17.030 280.750 ;
        RECT 17.180 280.100 17.830 280.750 ;
        RECT 11.630 279.250 12.280 279.900 ;
        RECT 12.430 279.250 13.080 279.900 ;
        RECT 13.230 279.250 13.880 279.900 ;
        RECT 15.580 279.250 16.230 279.900 ;
        RECT 16.380 279.250 17.030 279.900 ;
        RECT 17.180 279.250 17.830 279.900 ;
        RECT 20.430 280.100 21.280 280.950 ;
        RECT 21.380 280.100 22.230 280.950 ;
        RECT 22.830 280.100 23.680 280.950 ;
        RECT 23.780 280.100 24.630 280.950 ;
        RECT 24.830 280.100 25.680 280.950 ;
        RECT 25.780 280.100 26.630 280.950 ;
        RECT 27.230 280.100 28.080 280.950 ;
        RECT 28.180 280.100 29.030 280.950 ;
        RECT 43.780 281.050 44.630 281.900 ;
        RECT 44.830 281.050 45.680 281.900 ;
        RECT 4.830 278.100 5.680 278.950 ;
        RECT 20.430 279.050 21.280 279.900 ;
        RECT 21.380 279.050 22.230 279.900 ;
        RECT 22.830 279.050 23.680 279.900 ;
        RECT 23.780 279.050 24.630 279.900 ;
        RECT 24.830 279.050 25.680 279.900 ;
        RECT 25.780 279.050 26.630 279.900 ;
        RECT 27.230 279.050 28.080 279.900 ;
        RECT 28.180 279.050 29.030 279.900 ;
        RECT 31.630 280.100 32.280 280.750 ;
        RECT 32.430 280.100 33.080 280.750 ;
        RECT 33.230 280.100 33.880 280.750 ;
        RECT 35.580 280.100 36.230 280.750 ;
        RECT 36.380 280.100 37.030 280.750 ;
        RECT 37.180 280.100 37.830 280.750 ;
        RECT 31.630 279.250 32.280 279.900 ;
        RECT 32.430 279.250 33.080 279.900 ;
        RECT 33.230 279.250 33.880 279.900 ;
        RECT 35.580 279.250 36.230 279.900 ;
        RECT 36.380 279.250 37.030 279.900 ;
        RECT 37.180 279.250 37.830 279.900 ;
        RECT 40.430 280.100 41.280 280.950 ;
        RECT 41.380 280.100 42.230 280.950 ;
        RECT 42.830 280.100 43.680 280.950 ;
        RECT 43.780 280.100 44.630 280.950 ;
        RECT 44.830 280.100 45.680 280.950 ;
        RECT 45.780 280.100 46.630 280.950 ;
        RECT 47.230 280.100 48.080 280.950 ;
        RECT 48.180 280.100 49.030 280.950 ;
        RECT 63.780 281.050 64.630 281.900 ;
        RECT 64.830 281.050 65.680 281.900 ;
        RECT 23.780 278.100 24.630 278.950 ;
        RECT 24.830 278.100 25.680 278.950 ;
        RECT 40.430 279.050 41.280 279.900 ;
        RECT 41.380 279.050 42.230 279.900 ;
        RECT 42.830 279.050 43.680 279.900 ;
        RECT 43.780 279.050 44.630 279.900 ;
        RECT 44.830 279.050 45.680 279.900 ;
        RECT 45.780 279.050 46.630 279.900 ;
        RECT 47.230 279.050 48.080 279.900 ;
        RECT 48.180 279.050 49.030 279.900 ;
        RECT 51.630 280.100 52.280 280.750 ;
        RECT 52.430 280.100 53.080 280.750 ;
        RECT 53.230 280.100 53.880 280.750 ;
        RECT 55.580 280.100 56.230 280.750 ;
        RECT 56.380 280.100 57.030 280.750 ;
        RECT 57.180 280.100 57.830 280.750 ;
        RECT 51.630 279.250 52.280 279.900 ;
        RECT 52.430 279.250 53.080 279.900 ;
        RECT 53.230 279.250 53.880 279.900 ;
        RECT 55.580 279.250 56.230 279.900 ;
        RECT 56.380 279.250 57.030 279.900 ;
        RECT 57.180 279.250 57.830 279.900 ;
        RECT 60.430 280.100 61.280 280.950 ;
        RECT 61.380 280.100 62.230 280.950 ;
        RECT 62.830 280.100 63.680 280.950 ;
        RECT 63.780 280.100 64.630 280.950 ;
        RECT 64.830 280.100 65.680 280.950 ;
        RECT 65.780 280.100 66.630 280.950 ;
        RECT 67.230 280.100 68.080 280.950 ;
        RECT 68.180 280.100 69.030 280.950 ;
        RECT 83.780 281.050 84.630 281.900 ;
        RECT 84.830 281.050 85.680 281.900 ;
        RECT 43.780 278.100 44.630 278.950 ;
        RECT 44.830 278.100 45.680 278.950 ;
        RECT 60.430 279.050 61.280 279.900 ;
        RECT 61.380 279.050 62.230 279.900 ;
        RECT 62.830 279.050 63.680 279.900 ;
        RECT 63.780 279.050 64.630 279.900 ;
        RECT 64.830 279.050 65.680 279.900 ;
        RECT 65.780 279.050 66.630 279.900 ;
        RECT 67.230 279.050 68.080 279.900 ;
        RECT 68.180 279.050 69.030 279.900 ;
        RECT 71.630 280.100 72.280 280.750 ;
        RECT 72.430 280.100 73.080 280.750 ;
        RECT 73.230 280.100 73.880 280.750 ;
        RECT 75.580 280.100 76.230 280.750 ;
        RECT 76.380 280.100 77.030 280.750 ;
        RECT 77.180 280.100 77.830 280.750 ;
        RECT 71.630 279.250 72.280 279.900 ;
        RECT 72.430 279.250 73.080 279.900 ;
        RECT 73.230 279.250 73.880 279.900 ;
        RECT 75.580 279.250 76.230 279.900 ;
        RECT 76.380 279.250 77.030 279.900 ;
        RECT 77.180 279.250 77.830 279.900 ;
        RECT 80.430 280.100 81.280 280.950 ;
        RECT 81.380 280.100 82.230 280.950 ;
        RECT 82.830 280.100 83.680 280.950 ;
        RECT 83.780 280.100 84.630 280.950 ;
        RECT 84.830 280.100 85.680 280.950 ;
        RECT 85.780 280.100 86.630 280.950 ;
        RECT 87.230 280.100 88.080 280.950 ;
        RECT 88.180 280.100 89.030 280.950 ;
        RECT 103.780 281.050 104.630 281.900 ;
        RECT 104.830 281.050 105.680 281.900 ;
        RECT 63.780 278.100 64.630 278.950 ;
        RECT 64.830 278.100 65.680 278.950 ;
        RECT 80.430 279.050 81.280 279.900 ;
        RECT 81.380 279.050 82.230 279.900 ;
        RECT 82.830 279.050 83.680 279.900 ;
        RECT 83.780 279.050 84.630 279.900 ;
        RECT 84.830 279.050 85.680 279.900 ;
        RECT 85.780 279.050 86.630 279.900 ;
        RECT 87.230 279.050 88.080 279.900 ;
        RECT 88.180 279.050 89.030 279.900 ;
        RECT 91.630 280.100 92.280 280.750 ;
        RECT 92.430 280.100 93.080 280.750 ;
        RECT 93.230 280.100 93.880 280.750 ;
        RECT 95.580 280.100 96.230 280.750 ;
        RECT 96.380 280.100 97.030 280.750 ;
        RECT 97.180 280.100 97.830 280.750 ;
        RECT 91.630 279.250 92.280 279.900 ;
        RECT 92.430 279.250 93.080 279.900 ;
        RECT 93.230 279.250 93.880 279.900 ;
        RECT 95.580 279.250 96.230 279.900 ;
        RECT 96.380 279.250 97.030 279.900 ;
        RECT 97.180 279.250 97.830 279.900 ;
        RECT 100.430 280.100 101.280 280.950 ;
        RECT 101.380 280.100 102.230 280.950 ;
        RECT 102.830 280.100 103.680 280.950 ;
        RECT 103.780 280.100 104.630 280.950 ;
        RECT 104.830 280.100 105.680 280.950 ;
        RECT 105.780 280.100 106.630 280.950 ;
        RECT 107.230 280.100 108.080 280.950 ;
        RECT 108.180 280.100 109.030 280.950 ;
        RECT 123.780 281.050 124.630 281.900 ;
        RECT 83.780 278.100 84.630 278.950 ;
        RECT 84.830 278.100 85.680 278.950 ;
        RECT 100.430 279.050 101.280 279.900 ;
        RECT 101.380 279.050 102.230 279.900 ;
        RECT 102.830 279.050 103.680 279.900 ;
        RECT 103.780 279.050 104.630 279.900 ;
        RECT 104.830 279.050 105.680 279.900 ;
        RECT 105.780 279.050 106.630 279.900 ;
        RECT 107.230 279.050 108.080 279.900 ;
        RECT 108.180 279.050 109.030 279.900 ;
        RECT 111.630 280.100 112.280 280.750 ;
        RECT 112.430 280.100 113.080 280.750 ;
        RECT 113.230 280.100 113.880 280.750 ;
        RECT 115.580 280.100 116.230 280.750 ;
        RECT 116.380 280.100 117.030 280.750 ;
        RECT 117.180 280.100 117.830 280.750 ;
        RECT 111.630 279.250 112.280 279.900 ;
        RECT 112.430 279.250 113.080 279.900 ;
        RECT 113.230 279.250 113.880 279.900 ;
        RECT 115.580 279.250 116.230 279.900 ;
        RECT 116.380 279.250 117.030 279.900 ;
        RECT 117.180 279.250 117.830 279.900 ;
        RECT 120.430 280.100 121.280 280.950 ;
        RECT 121.380 280.100 122.230 280.950 ;
        RECT 122.830 280.100 123.680 280.950 ;
        RECT 123.780 280.100 124.630 280.950 ;
        RECT 103.780 278.100 104.630 278.950 ;
        RECT 104.830 278.100 105.680 278.950 ;
        RECT 120.430 279.050 121.280 279.900 ;
        RECT 121.380 279.050 122.230 279.900 ;
        RECT 122.830 279.050 123.680 279.900 ;
        RECT 123.780 279.050 124.630 279.900 ;
        RECT 123.780 278.100 124.630 278.950 ;
        RECT 4.830 276.650 5.680 277.500 ;
        RECT 23.780 276.650 24.630 277.500 ;
        RECT 24.830 276.650 25.680 277.500 ;
        RECT 43.780 276.650 44.630 277.500 ;
        RECT 44.830 276.650 45.680 277.500 ;
        RECT 63.780 276.650 64.630 277.500 ;
        RECT 64.830 276.650 65.680 277.500 ;
        RECT 83.780 276.650 84.630 277.500 ;
        RECT 84.830 276.650 85.680 277.500 ;
        RECT 103.780 276.650 104.630 277.500 ;
        RECT 104.830 276.650 105.680 277.500 ;
        RECT 123.780 276.650 124.630 277.500 ;
        RECT 4.830 275.700 5.680 276.550 ;
        RECT 23.780 275.700 24.630 276.550 ;
        RECT 24.830 275.700 25.680 276.550 ;
        RECT 43.780 275.700 44.630 276.550 ;
        RECT 44.830 275.700 45.680 276.550 ;
        RECT 63.780 275.700 64.630 276.550 ;
        RECT 64.830 275.700 65.680 276.550 ;
        RECT 83.780 275.700 84.630 276.550 ;
        RECT 84.830 275.700 85.680 276.550 ;
        RECT 103.780 275.700 104.630 276.550 ;
        RECT 104.830 275.700 105.680 276.550 ;
        RECT 123.780 275.700 124.630 276.550 ;
        RECT 4.830 272.450 5.480 273.100 ;
        RECT 4.830 271.650 5.480 272.300 ;
        RECT 4.830 270.850 5.480 271.500 ;
        RECT 4.830 268.500 5.480 269.150 ;
        RECT 4.830 267.700 5.480 268.350 ;
        RECT 4.830 266.900 5.480 267.550 ;
        RECT 23.980 272.450 24.630 273.100 ;
        RECT 24.830 272.450 25.480 273.100 ;
        RECT 23.980 271.650 24.630 272.300 ;
        RECT 24.830 271.650 25.480 272.300 ;
        RECT 23.980 270.850 24.630 271.500 ;
        RECT 24.830 270.850 25.480 271.500 ;
        RECT 23.980 268.500 24.630 269.150 ;
        RECT 24.830 268.500 25.480 269.150 ;
        RECT 23.980 267.700 24.630 268.350 ;
        RECT 24.830 267.700 25.480 268.350 ;
        RECT 23.980 266.900 24.630 267.550 ;
        RECT 24.830 266.900 25.480 267.550 ;
        RECT 43.980 272.450 44.630 273.100 ;
        RECT 44.830 272.450 45.480 273.100 ;
        RECT 43.980 271.650 44.630 272.300 ;
        RECT 44.830 271.650 45.480 272.300 ;
        RECT 43.980 270.850 44.630 271.500 ;
        RECT 44.830 270.850 45.480 271.500 ;
        RECT 43.980 268.500 44.630 269.150 ;
        RECT 44.830 268.500 45.480 269.150 ;
        RECT 43.980 267.700 44.630 268.350 ;
        RECT 44.830 267.700 45.480 268.350 ;
        RECT 43.980 266.900 44.630 267.550 ;
        RECT 44.830 266.900 45.480 267.550 ;
        RECT 63.980 272.450 64.630 273.100 ;
        RECT 64.830 272.450 65.480 273.100 ;
        RECT 63.980 271.650 64.630 272.300 ;
        RECT 64.830 271.650 65.480 272.300 ;
        RECT 63.980 270.850 64.630 271.500 ;
        RECT 64.830 270.850 65.480 271.500 ;
        RECT 63.980 268.500 64.630 269.150 ;
        RECT 64.830 268.500 65.480 269.150 ;
        RECT 63.980 267.700 64.630 268.350 ;
        RECT 64.830 267.700 65.480 268.350 ;
        RECT 63.980 266.900 64.630 267.550 ;
        RECT 64.830 266.900 65.480 267.550 ;
        RECT 83.980 272.450 84.630 273.100 ;
        RECT 84.830 272.450 85.480 273.100 ;
        RECT 83.980 271.650 84.630 272.300 ;
        RECT 84.830 271.650 85.480 272.300 ;
        RECT 83.980 270.850 84.630 271.500 ;
        RECT 84.830 270.850 85.480 271.500 ;
        RECT 83.980 268.500 84.630 269.150 ;
        RECT 84.830 268.500 85.480 269.150 ;
        RECT 83.980 267.700 84.630 268.350 ;
        RECT 84.830 267.700 85.480 268.350 ;
        RECT 83.980 266.900 84.630 267.550 ;
        RECT 84.830 266.900 85.480 267.550 ;
        RECT 103.980 272.450 104.630 273.100 ;
        RECT 104.830 272.450 105.480 273.100 ;
        RECT 103.980 271.650 104.630 272.300 ;
        RECT 104.830 271.650 105.480 272.300 ;
        RECT 103.980 270.850 104.630 271.500 ;
        RECT 104.830 270.850 105.480 271.500 ;
        RECT 103.980 268.500 104.630 269.150 ;
        RECT 104.830 268.500 105.480 269.150 ;
        RECT 103.980 267.700 104.630 268.350 ;
        RECT 104.830 267.700 105.480 268.350 ;
        RECT 103.980 266.900 104.630 267.550 ;
        RECT 104.830 266.900 105.480 267.550 ;
        RECT 123.980 272.450 124.630 273.100 ;
        RECT 123.980 271.650 124.630 272.300 ;
        RECT 123.980 270.850 124.630 271.500 ;
        RECT 123.980 268.500 124.630 269.150 ;
        RECT 123.980 267.700 124.630 268.350 ;
        RECT 123.980 266.900 124.630 267.550 ;
        RECT 4.830 263.450 5.680 264.300 ;
        RECT 23.780 263.450 24.630 264.300 ;
        RECT 24.830 263.450 25.680 264.300 ;
        RECT 43.780 263.450 44.630 264.300 ;
        RECT 44.830 263.450 45.680 264.300 ;
        RECT 63.780 263.450 64.630 264.300 ;
        RECT 64.830 263.450 65.680 264.300 ;
        RECT 83.780 263.450 84.630 264.300 ;
        RECT 84.830 263.450 85.680 264.300 ;
        RECT 103.780 263.450 104.630 264.300 ;
        RECT 104.830 263.450 105.680 264.300 ;
        RECT 123.780 263.450 124.630 264.300 ;
        RECT 4.830 262.500 5.680 263.350 ;
        RECT 23.780 262.500 24.630 263.350 ;
        RECT 24.830 262.500 25.680 263.350 ;
        RECT 43.780 262.500 44.630 263.350 ;
        RECT 44.830 262.500 45.680 263.350 ;
        RECT 63.780 262.500 64.630 263.350 ;
        RECT 64.830 262.500 65.680 263.350 ;
        RECT 83.780 262.500 84.630 263.350 ;
        RECT 84.830 262.500 85.680 263.350 ;
        RECT 103.780 262.500 104.630 263.350 ;
        RECT 104.830 262.500 105.680 263.350 ;
        RECT 123.780 262.500 124.630 263.350 ;
        RECT 4.830 261.050 5.680 261.900 ;
        RECT 4.830 260.100 5.680 260.950 ;
        RECT 5.780 260.100 6.630 260.950 ;
        RECT 7.230 260.100 8.080 260.950 ;
        RECT 8.180 260.100 9.030 260.950 ;
        RECT 23.780 261.050 24.630 261.900 ;
        RECT 24.830 261.050 25.680 261.900 ;
        RECT 4.830 259.050 5.680 259.900 ;
        RECT 5.780 259.050 6.630 259.900 ;
        RECT 7.230 259.050 8.080 259.900 ;
        RECT 8.180 259.050 9.030 259.900 ;
        RECT 11.630 260.100 12.280 260.750 ;
        RECT 12.430 260.100 13.080 260.750 ;
        RECT 13.230 260.100 13.880 260.750 ;
        RECT 15.580 260.100 16.230 260.750 ;
        RECT 16.380 260.100 17.030 260.750 ;
        RECT 17.180 260.100 17.830 260.750 ;
        RECT 11.630 259.250 12.280 259.900 ;
        RECT 12.430 259.250 13.080 259.900 ;
        RECT 13.230 259.250 13.880 259.900 ;
        RECT 15.580 259.250 16.230 259.900 ;
        RECT 16.380 259.250 17.030 259.900 ;
        RECT 17.180 259.250 17.830 259.900 ;
        RECT 20.430 260.100 21.280 260.950 ;
        RECT 21.380 260.100 22.230 260.950 ;
        RECT 22.830 260.100 23.680 260.950 ;
        RECT 23.780 260.100 24.630 260.950 ;
        RECT 24.830 260.100 25.680 260.950 ;
        RECT 25.780 260.100 26.630 260.950 ;
        RECT 27.230 260.100 28.080 260.950 ;
        RECT 28.180 260.100 29.030 260.950 ;
        RECT 43.780 261.050 44.630 261.900 ;
        RECT 44.830 261.050 45.680 261.900 ;
        RECT 4.830 258.100 5.680 258.950 ;
        RECT 20.430 259.050 21.280 259.900 ;
        RECT 21.380 259.050 22.230 259.900 ;
        RECT 22.830 259.050 23.680 259.900 ;
        RECT 23.780 259.050 24.630 259.900 ;
        RECT 24.830 259.050 25.680 259.900 ;
        RECT 25.780 259.050 26.630 259.900 ;
        RECT 27.230 259.050 28.080 259.900 ;
        RECT 28.180 259.050 29.030 259.900 ;
        RECT 31.630 260.100 32.280 260.750 ;
        RECT 32.430 260.100 33.080 260.750 ;
        RECT 33.230 260.100 33.880 260.750 ;
        RECT 35.580 260.100 36.230 260.750 ;
        RECT 36.380 260.100 37.030 260.750 ;
        RECT 37.180 260.100 37.830 260.750 ;
        RECT 31.630 259.250 32.280 259.900 ;
        RECT 32.430 259.250 33.080 259.900 ;
        RECT 33.230 259.250 33.880 259.900 ;
        RECT 35.580 259.250 36.230 259.900 ;
        RECT 36.380 259.250 37.030 259.900 ;
        RECT 37.180 259.250 37.830 259.900 ;
        RECT 40.430 260.100 41.280 260.950 ;
        RECT 41.380 260.100 42.230 260.950 ;
        RECT 42.830 260.100 43.680 260.950 ;
        RECT 43.780 260.100 44.630 260.950 ;
        RECT 44.830 260.100 45.680 260.950 ;
        RECT 45.780 260.100 46.630 260.950 ;
        RECT 47.230 260.100 48.080 260.950 ;
        RECT 48.180 260.100 49.030 260.950 ;
        RECT 63.780 261.050 64.630 261.900 ;
        RECT 64.830 261.050 65.680 261.900 ;
        RECT 23.780 258.100 24.630 258.950 ;
        RECT 24.830 258.100 25.680 258.950 ;
        RECT 40.430 259.050 41.280 259.900 ;
        RECT 41.380 259.050 42.230 259.900 ;
        RECT 42.830 259.050 43.680 259.900 ;
        RECT 43.780 259.050 44.630 259.900 ;
        RECT 44.830 259.050 45.680 259.900 ;
        RECT 45.780 259.050 46.630 259.900 ;
        RECT 47.230 259.050 48.080 259.900 ;
        RECT 48.180 259.050 49.030 259.900 ;
        RECT 51.630 260.100 52.280 260.750 ;
        RECT 52.430 260.100 53.080 260.750 ;
        RECT 53.230 260.100 53.880 260.750 ;
        RECT 55.580 260.100 56.230 260.750 ;
        RECT 56.380 260.100 57.030 260.750 ;
        RECT 57.180 260.100 57.830 260.750 ;
        RECT 51.630 259.250 52.280 259.900 ;
        RECT 52.430 259.250 53.080 259.900 ;
        RECT 53.230 259.250 53.880 259.900 ;
        RECT 55.580 259.250 56.230 259.900 ;
        RECT 56.380 259.250 57.030 259.900 ;
        RECT 57.180 259.250 57.830 259.900 ;
        RECT 60.430 260.100 61.280 260.950 ;
        RECT 61.380 260.100 62.230 260.950 ;
        RECT 62.830 260.100 63.680 260.950 ;
        RECT 63.780 260.100 64.630 260.950 ;
        RECT 64.830 260.100 65.680 260.950 ;
        RECT 65.780 260.100 66.630 260.950 ;
        RECT 67.230 260.100 68.080 260.950 ;
        RECT 68.180 260.100 69.030 260.950 ;
        RECT 83.780 261.050 84.630 261.900 ;
        RECT 84.830 261.050 85.680 261.900 ;
        RECT 43.780 258.100 44.630 258.950 ;
        RECT 44.830 258.100 45.680 258.950 ;
        RECT 60.430 259.050 61.280 259.900 ;
        RECT 61.380 259.050 62.230 259.900 ;
        RECT 62.830 259.050 63.680 259.900 ;
        RECT 63.780 259.050 64.630 259.900 ;
        RECT 64.830 259.050 65.680 259.900 ;
        RECT 65.780 259.050 66.630 259.900 ;
        RECT 67.230 259.050 68.080 259.900 ;
        RECT 68.180 259.050 69.030 259.900 ;
        RECT 71.630 260.100 72.280 260.750 ;
        RECT 72.430 260.100 73.080 260.750 ;
        RECT 73.230 260.100 73.880 260.750 ;
        RECT 75.580 260.100 76.230 260.750 ;
        RECT 76.380 260.100 77.030 260.750 ;
        RECT 77.180 260.100 77.830 260.750 ;
        RECT 71.630 259.250 72.280 259.900 ;
        RECT 72.430 259.250 73.080 259.900 ;
        RECT 73.230 259.250 73.880 259.900 ;
        RECT 75.580 259.250 76.230 259.900 ;
        RECT 76.380 259.250 77.030 259.900 ;
        RECT 77.180 259.250 77.830 259.900 ;
        RECT 80.430 260.100 81.280 260.950 ;
        RECT 81.380 260.100 82.230 260.950 ;
        RECT 82.830 260.100 83.680 260.950 ;
        RECT 83.780 260.100 84.630 260.950 ;
        RECT 84.830 260.100 85.680 260.950 ;
        RECT 85.780 260.100 86.630 260.950 ;
        RECT 87.230 260.100 88.080 260.950 ;
        RECT 88.180 260.100 89.030 260.950 ;
        RECT 103.780 261.050 104.630 261.900 ;
        RECT 104.830 261.050 105.680 261.900 ;
        RECT 63.780 258.100 64.630 258.950 ;
        RECT 64.830 258.100 65.680 258.950 ;
        RECT 80.430 259.050 81.280 259.900 ;
        RECT 81.380 259.050 82.230 259.900 ;
        RECT 82.830 259.050 83.680 259.900 ;
        RECT 83.780 259.050 84.630 259.900 ;
        RECT 84.830 259.050 85.680 259.900 ;
        RECT 85.780 259.050 86.630 259.900 ;
        RECT 87.230 259.050 88.080 259.900 ;
        RECT 88.180 259.050 89.030 259.900 ;
        RECT 91.630 260.100 92.280 260.750 ;
        RECT 92.430 260.100 93.080 260.750 ;
        RECT 93.230 260.100 93.880 260.750 ;
        RECT 95.580 260.100 96.230 260.750 ;
        RECT 96.380 260.100 97.030 260.750 ;
        RECT 97.180 260.100 97.830 260.750 ;
        RECT 91.630 259.250 92.280 259.900 ;
        RECT 92.430 259.250 93.080 259.900 ;
        RECT 93.230 259.250 93.880 259.900 ;
        RECT 95.580 259.250 96.230 259.900 ;
        RECT 96.380 259.250 97.030 259.900 ;
        RECT 97.180 259.250 97.830 259.900 ;
        RECT 100.430 260.100 101.280 260.950 ;
        RECT 101.380 260.100 102.230 260.950 ;
        RECT 102.830 260.100 103.680 260.950 ;
        RECT 103.780 260.100 104.630 260.950 ;
        RECT 104.830 260.100 105.680 260.950 ;
        RECT 105.780 260.100 106.630 260.950 ;
        RECT 107.230 260.100 108.080 260.950 ;
        RECT 108.180 260.100 109.030 260.950 ;
        RECT 123.780 261.050 124.630 261.900 ;
        RECT 83.780 258.100 84.630 258.950 ;
        RECT 84.830 258.100 85.680 258.950 ;
        RECT 100.430 259.050 101.280 259.900 ;
        RECT 101.380 259.050 102.230 259.900 ;
        RECT 102.830 259.050 103.680 259.900 ;
        RECT 103.780 259.050 104.630 259.900 ;
        RECT 104.830 259.050 105.680 259.900 ;
        RECT 105.780 259.050 106.630 259.900 ;
        RECT 107.230 259.050 108.080 259.900 ;
        RECT 108.180 259.050 109.030 259.900 ;
        RECT 111.630 260.100 112.280 260.750 ;
        RECT 112.430 260.100 113.080 260.750 ;
        RECT 113.230 260.100 113.880 260.750 ;
        RECT 115.580 260.100 116.230 260.750 ;
        RECT 116.380 260.100 117.030 260.750 ;
        RECT 117.180 260.100 117.830 260.750 ;
        RECT 111.630 259.250 112.280 259.900 ;
        RECT 112.430 259.250 113.080 259.900 ;
        RECT 113.230 259.250 113.880 259.900 ;
        RECT 115.580 259.250 116.230 259.900 ;
        RECT 116.380 259.250 117.030 259.900 ;
        RECT 117.180 259.250 117.830 259.900 ;
        RECT 120.430 260.100 121.280 260.950 ;
        RECT 121.380 260.100 122.230 260.950 ;
        RECT 122.830 260.100 123.680 260.950 ;
        RECT 123.780 260.100 124.630 260.950 ;
        RECT 103.780 258.100 104.630 258.950 ;
        RECT 104.830 258.100 105.680 258.950 ;
        RECT 120.430 259.050 121.280 259.900 ;
        RECT 121.380 259.050 122.230 259.900 ;
        RECT 122.830 259.050 123.680 259.900 ;
        RECT 123.780 259.050 124.630 259.900 ;
        RECT 123.780 258.100 124.630 258.950 ;
        RECT 4.830 256.650 5.680 257.500 ;
        RECT 23.780 256.650 24.630 257.500 ;
        RECT 24.830 256.650 25.680 257.500 ;
        RECT 43.780 256.650 44.630 257.500 ;
        RECT 44.830 256.650 45.680 257.500 ;
        RECT 63.780 256.650 64.630 257.500 ;
        RECT 64.830 256.650 65.680 257.500 ;
        RECT 83.780 256.650 84.630 257.500 ;
        RECT 84.830 256.650 85.680 257.500 ;
        RECT 103.780 256.650 104.630 257.500 ;
        RECT 104.830 256.650 105.680 257.500 ;
        RECT 123.780 256.650 124.630 257.500 ;
        RECT 4.830 255.700 5.680 256.550 ;
        RECT 23.780 255.700 24.630 256.550 ;
        RECT 24.830 255.700 25.680 256.550 ;
        RECT 43.780 255.700 44.630 256.550 ;
        RECT 44.830 255.700 45.680 256.550 ;
        RECT 63.780 255.700 64.630 256.550 ;
        RECT 64.830 255.700 65.680 256.550 ;
        RECT 83.780 255.700 84.630 256.550 ;
        RECT 84.830 255.700 85.680 256.550 ;
        RECT 103.780 255.700 104.630 256.550 ;
        RECT 104.830 255.700 105.680 256.550 ;
        RECT 123.780 255.700 124.630 256.550 ;
        RECT 4.830 252.450 5.480 253.100 ;
        RECT 4.830 251.650 5.480 252.300 ;
        RECT 4.830 250.850 5.480 251.500 ;
        RECT 4.830 248.500 5.480 249.150 ;
        RECT 4.830 247.700 5.480 248.350 ;
        RECT 4.830 246.900 5.480 247.550 ;
        RECT 23.980 252.450 24.630 253.100 ;
        RECT 24.830 252.450 25.480 253.100 ;
        RECT 23.980 251.650 24.630 252.300 ;
        RECT 24.830 251.650 25.480 252.300 ;
        RECT 23.980 250.850 24.630 251.500 ;
        RECT 24.830 250.850 25.480 251.500 ;
        RECT 23.980 248.500 24.630 249.150 ;
        RECT 24.830 248.500 25.480 249.150 ;
        RECT 23.980 247.700 24.630 248.350 ;
        RECT 24.830 247.700 25.480 248.350 ;
        RECT 23.980 246.900 24.630 247.550 ;
        RECT 24.830 246.900 25.480 247.550 ;
        RECT 43.980 252.450 44.630 253.100 ;
        RECT 44.830 252.450 45.480 253.100 ;
        RECT 43.980 251.650 44.630 252.300 ;
        RECT 44.830 251.650 45.480 252.300 ;
        RECT 43.980 250.850 44.630 251.500 ;
        RECT 44.830 250.850 45.480 251.500 ;
        RECT 43.980 248.500 44.630 249.150 ;
        RECT 44.830 248.500 45.480 249.150 ;
        RECT 43.980 247.700 44.630 248.350 ;
        RECT 44.830 247.700 45.480 248.350 ;
        RECT 43.980 246.900 44.630 247.550 ;
        RECT 44.830 246.900 45.480 247.550 ;
        RECT 63.980 252.450 64.630 253.100 ;
        RECT 64.830 252.450 65.480 253.100 ;
        RECT 63.980 251.650 64.630 252.300 ;
        RECT 64.830 251.650 65.480 252.300 ;
        RECT 63.980 250.850 64.630 251.500 ;
        RECT 64.830 250.850 65.480 251.500 ;
        RECT 63.980 248.500 64.630 249.150 ;
        RECT 64.830 248.500 65.480 249.150 ;
        RECT 63.980 247.700 64.630 248.350 ;
        RECT 64.830 247.700 65.480 248.350 ;
        RECT 63.980 246.900 64.630 247.550 ;
        RECT 64.830 246.900 65.480 247.550 ;
        RECT 83.980 252.450 84.630 253.100 ;
        RECT 84.830 252.450 85.480 253.100 ;
        RECT 83.980 251.650 84.630 252.300 ;
        RECT 84.830 251.650 85.480 252.300 ;
        RECT 83.980 250.850 84.630 251.500 ;
        RECT 84.830 250.850 85.480 251.500 ;
        RECT 83.980 248.500 84.630 249.150 ;
        RECT 84.830 248.500 85.480 249.150 ;
        RECT 83.980 247.700 84.630 248.350 ;
        RECT 84.830 247.700 85.480 248.350 ;
        RECT 83.980 246.900 84.630 247.550 ;
        RECT 84.830 246.900 85.480 247.550 ;
        RECT 103.980 252.450 104.630 253.100 ;
        RECT 104.830 252.450 105.480 253.100 ;
        RECT 103.980 251.650 104.630 252.300 ;
        RECT 104.830 251.650 105.480 252.300 ;
        RECT 103.980 250.850 104.630 251.500 ;
        RECT 104.830 250.850 105.480 251.500 ;
        RECT 103.980 248.500 104.630 249.150 ;
        RECT 104.830 248.500 105.480 249.150 ;
        RECT 103.980 247.700 104.630 248.350 ;
        RECT 104.830 247.700 105.480 248.350 ;
        RECT 103.980 246.900 104.630 247.550 ;
        RECT 104.830 246.900 105.480 247.550 ;
        RECT 123.980 252.450 124.630 253.100 ;
        RECT 123.980 251.650 124.630 252.300 ;
        RECT 123.980 250.850 124.630 251.500 ;
        RECT 123.980 248.500 124.630 249.150 ;
        RECT 123.980 247.700 124.630 248.350 ;
        RECT 123.980 246.900 124.630 247.550 ;
        RECT 4.830 243.450 5.680 244.300 ;
        RECT 23.780 243.450 24.630 244.300 ;
        RECT 24.830 243.450 25.680 244.300 ;
        RECT 43.780 243.450 44.630 244.300 ;
        RECT 44.830 243.450 45.680 244.300 ;
        RECT 63.780 243.450 64.630 244.300 ;
        RECT 64.830 243.450 65.680 244.300 ;
        RECT 83.780 243.450 84.630 244.300 ;
        RECT 84.830 243.450 85.680 244.300 ;
        RECT 103.780 243.450 104.630 244.300 ;
        RECT 104.830 243.450 105.680 244.300 ;
        RECT 123.780 243.450 124.630 244.300 ;
        RECT 4.830 242.500 5.680 243.350 ;
        RECT 23.780 242.500 24.630 243.350 ;
        RECT 24.830 242.500 25.680 243.350 ;
        RECT 43.780 242.500 44.630 243.350 ;
        RECT 44.830 242.500 45.680 243.350 ;
        RECT 63.780 242.500 64.630 243.350 ;
        RECT 64.830 242.500 65.680 243.350 ;
        RECT 83.780 242.500 84.630 243.350 ;
        RECT 84.830 242.500 85.680 243.350 ;
        RECT 103.780 242.500 104.630 243.350 ;
        RECT 104.830 242.500 105.680 243.350 ;
        RECT 123.780 242.500 124.630 243.350 ;
        RECT 4.830 241.050 5.680 241.900 ;
        RECT 4.830 240.100 5.680 240.950 ;
        RECT 5.780 240.100 6.630 240.950 ;
        RECT 7.230 240.100 8.080 240.950 ;
        RECT 8.180 240.100 9.030 240.950 ;
        RECT 23.780 241.050 24.630 241.900 ;
        RECT 24.830 241.050 25.680 241.900 ;
        RECT 4.830 239.050 5.680 239.900 ;
        RECT 5.780 239.050 6.630 239.900 ;
        RECT 7.230 239.050 8.080 239.900 ;
        RECT 8.180 239.050 9.030 239.900 ;
        RECT 11.630 240.100 12.280 240.750 ;
        RECT 12.430 240.100 13.080 240.750 ;
        RECT 13.230 240.100 13.880 240.750 ;
        RECT 15.580 240.100 16.230 240.750 ;
        RECT 16.380 240.100 17.030 240.750 ;
        RECT 17.180 240.100 17.830 240.750 ;
        RECT 11.630 239.250 12.280 239.900 ;
        RECT 12.430 239.250 13.080 239.900 ;
        RECT 13.230 239.250 13.880 239.900 ;
        RECT 15.580 239.250 16.230 239.900 ;
        RECT 16.380 239.250 17.030 239.900 ;
        RECT 17.180 239.250 17.830 239.900 ;
        RECT 20.430 240.100 21.280 240.950 ;
        RECT 21.380 240.100 22.230 240.950 ;
        RECT 22.830 240.100 23.680 240.950 ;
        RECT 23.780 240.100 24.630 240.950 ;
        RECT 24.830 240.100 25.680 240.950 ;
        RECT 25.780 240.100 26.630 240.950 ;
        RECT 27.230 240.100 28.080 240.950 ;
        RECT 28.180 240.100 29.030 240.950 ;
        RECT 43.780 241.050 44.630 241.900 ;
        RECT 44.830 241.050 45.680 241.900 ;
        RECT 4.830 238.100 5.680 238.950 ;
        RECT 20.430 239.050 21.280 239.900 ;
        RECT 21.380 239.050 22.230 239.900 ;
        RECT 22.830 239.050 23.680 239.900 ;
        RECT 23.780 239.050 24.630 239.900 ;
        RECT 24.830 239.050 25.680 239.900 ;
        RECT 25.780 239.050 26.630 239.900 ;
        RECT 27.230 239.050 28.080 239.900 ;
        RECT 28.180 239.050 29.030 239.900 ;
        RECT 31.630 240.100 32.280 240.750 ;
        RECT 32.430 240.100 33.080 240.750 ;
        RECT 33.230 240.100 33.880 240.750 ;
        RECT 35.580 240.100 36.230 240.750 ;
        RECT 36.380 240.100 37.030 240.750 ;
        RECT 37.180 240.100 37.830 240.750 ;
        RECT 31.630 239.250 32.280 239.900 ;
        RECT 32.430 239.250 33.080 239.900 ;
        RECT 33.230 239.250 33.880 239.900 ;
        RECT 35.580 239.250 36.230 239.900 ;
        RECT 36.380 239.250 37.030 239.900 ;
        RECT 37.180 239.250 37.830 239.900 ;
        RECT 40.430 240.100 41.280 240.950 ;
        RECT 41.380 240.100 42.230 240.950 ;
        RECT 42.830 240.100 43.680 240.950 ;
        RECT 43.780 240.100 44.630 240.950 ;
        RECT 44.830 240.100 45.680 240.950 ;
        RECT 45.780 240.100 46.630 240.950 ;
        RECT 47.230 240.100 48.080 240.950 ;
        RECT 48.180 240.100 49.030 240.950 ;
        RECT 63.780 241.050 64.630 241.900 ;
        RECT 64.830 241.050 65.680 241.900 ;
        RECT 23.780 238.100 24.630 238.950 ;
        RECT 24.830 238.100 25.680 238.950 ;
        RECT 40.430 239.050 41.280 239.900 ;
        RECT 41.380 239.050 42.230 239.900 ;
        RECT 42.830 239.050 43.680 239.900 ;
        RECT 43.780 239.050 44.630 239.900 ;
        RECT 44.830 239.050 45.680 239.900 ;
        RECT 45.780 239.050 46.630 239.900 ;
        RECT 47.230 239.050 48.080 239.900 ;
        RECT 48.180 239.050 49.030 239.900 ;
        RECT 51.630 240.100 52.280 240.750 ;
        RECT 52.430 240.100 53.080 240.750 ;
        RECT 53.230 240.100 53.880 240.750 ;
        RECT 55.580 240.100 56.230 240.750 ;
        RECT 56.380 240.100 57.030 240.750 ;
        RECT 57.180 240.100 57.830 240.750 ;
        RECT 51.630 239.250 52.280 239.900 ;
        RECT 52.430 239.250 53.080 239.900 ;
        RECT 53.230 239.250 53.880 239.900 ;
        RECT 55.580 239.250 56.230 239.900 ;
        RECT 56.380 239.250 57.030 239.900 ;
        RECT 57.180 239.250 57.830 239.900 ;
        RECT 60.430 240.100 61.280 240.950 ;
        RECT 61.380 240.100 62.230 240.950 ;
        RECT 62.830 240.100 63.680 240.950 ;
        RECT 63.780 240.100 64.630 240.950 ;
        RECT 64.830 240.100 65.680 240.950 ;
        RECT 65.780 240.100 66.630 240.950 ;
        RECT 67.230 240.100 68.080 240.950 ;
        RECT 68.180 240.100 69.030 240.950 ;
        RECT 83.780 241.050 84.630 241.900 ;
        RECT 84.830 241.050 85.680 241.900 ;
        RECT 43.780 238.100 44.630 238.950 ;
        RECT 44.830 238.100 45.680 238.950 ;
        RECT 60.430 239.050 61.280 239.900 ;
        RECT 61.380 239.050 62.230 239.900 ;
        RECT 62.830 239.050 63.680 239.900 ;
        RECT 63.780 239.050 64.630 239.900 ;
        RECT 64.830 239.050 65.680 239.900 ;
        RECT 65.780 239.050 66.630 239.900 ;
        RECT 67.230 239.050 68.080 239.900 ;
        RECT 68.180 239.050 69.030 239.900 ;
        RECT 71.630 240.100 72.280 240.750 ;
        RECT 72.430 240.100 73.080 240.750 ;
        RECT 73.230 240.100 73.880 240.750 ;
        RECT 75.580 240.100 76.230 240.750 ;
        RECT 76.380 240.100 77.030 240.750 ;
        RECT 77.180 240.100 77.830 240.750 ;
        RECT 71.630 239.250 72.280 239.900 ;
        RECT 72.430 239.250 73.080 239.900 ;
        RECT 73.230 239.250 73.880 239.900 ;
        RECT 75.580 239.250 76.230 239.900 ;
        RECT 76.380 239.250 77.030 239.900 ;
        RECT 77.180 239.250 77.830 239.900 ;
        RECT 80.430 240.100 81.280 240.950 ;
        RECT 81.380 240.100 82.230 240.950 ;
        RECT 82.830 240.100 83.680 240.950 ;
        RECT 83.780 240.100 84.630 240.950 ;
        RECT 84.830 240.100 85.680 240.950 ;
        RECT 85.780 240.100 86.630 240.950 ;
        RECT 87.230 240.100 88.080 240.950 ;
        RECT 88.180 240.100 89.030 240.950 ;
        RECT 103.780 241.050 104.630 241.900 ;
        RECT 104.830 241.050 105.680 241.900 ;
        RECT 63.780 238.100 64.630 238.950 ;
        RECT 64.830 238.100 65.680 238.950 ;
        RECT 80.430 239.050 81.280 239.900 ;
        RECT 81.380 239.050 82.230 239.900 ;
        RECT 82.830 239.050 83.680 239.900 ;
        RECT 83.780 239.050 84.630 239.900 ;
        RECT 84.830 239.050 85.680 239.900 ;
        RECT 85.780 239.050 86.630 239.900 ;
        RECT 87.230 239.050 88.080 239.900 ;
        RECT 88.180 239.050 89.030 239.900 ;
        RECT 91.630 240.100 92.280 240.750 ;
        RECT 92.430 240.100 93.080 240.750 ;
        RECT 93.230 240.100 93.880 240.750 ;
        RECT 95.580 240.100 96.230 240.750 ;
        RECT 96.380 240.100 97.030 240.750 ;
        RECT 97.180 240.100 97.830 240.750 ;
        RECT 91.630 239.250 92.280 239.900 ;
        RECT 92.430 239.250 93.080 239.900 ;
        RECT 93.230 239.250 93.880 239.900 ;
        RECT 95.580 239.250 96.230 239.900 ;
        RECT 96.380 239.250 97.030 239.900 ;
        RECT 97.180 239.250 97.830 239.900 ;
        RECT 100.430 240.100 101.280 240.950 ;
        RECT 101.380 240.100 102.230 240.950 ;
        RECT 102.830 240.100 103.680 240.950 ;
        RECT 103.780 240.100 104.630 240.950 ;
        RECT 104.830 240.100 105.680 240.950 ;
        RECT 105.780 240.100 106.630 240.950 ;
        RECT 107.230 240.100 108.080 240.950 ;
        RECT 108.180 240.100 109.030 240.950 ;
        RECT 123.780 241.050 124.630 241.900 ;
        RECT 83.780 238.100 84.630 238.950 ;
        RECT 84.830 238.100 85.680 238.950 ;
        RECT 100.430 239.050 101.280 239.900 ;
        RECT 101.380 239.050 102.230 239.900 ;
        RECT 102.830 239.050 103.680 239.900 ;
        RECT 103.780 239.050 104.630 239.900 ;
        RECT 104.830 239.050 105.680 239.900 ;
        RECT 105.780 239.050 106.630 239.900 ;
        RECT 107.230 239.050 108.080 239.900 ;
        RECT 108.180 239.050 109.030 239.900 ;
        RECT 111.630 240.100 112.280 240.750 ;
        RECT 112.430 240.100 113.080 240.750 ;
        RECT 113.230 240.100 113.880 240.750 ;
        RECT 115.580 240.100 116.230 240.750 ;
        RECT 116.380 240.100 117.030 240.750 ;
        RECT 117.180 240.100 117.830 240.750 ;
        RECT 111.630 239.250 112.280 239.900 ;
        RECT 112.430 239.250 113.080 239.900 ;
        RECT 113.230 239.250 113.880 239.900 ;
        RECT 115.580 239.250 116.230 239.900 ;
        RECT 116.380 239.250 117.030 239.900 ;
        RECT 117.180 239.250 117.830 239.900 ;
        RECT 120.430 240.100 121.280 240.950 ;
        RECT 121.380 240.100 122.230 240.950 ;
        RECT 122.830 240.100 123.680 240.950 ;
        RECT 123.780 240.100 124.630 240.950 ;
        RECT 103.780 238.100 104.630 238.950 ;
        RECT 104.830 238.100 105.680 238.950 ;
        RECT 120.430 239.050 121.280 239.900 ;
        RECT 121.380 239.050 122.230 239.900 ;
        RECT 122.830 239.050 123.680 239.900 ;
        RECT 123.780 239.050 124.630 239.900 ;
        RECT 123.780 238.100 124.630 238.950 ;
        RECT 4.830 236.650 5.680 237.500 ;
        RECT 23.780 236.650 24.630 237.500 ;
        RECT 24.830 236.650 25.680 237.500 ;
        RECT 43.780 236.650 44.630 237.500 ;
        RECT 44.830 236.650 45.680 237.500 ;
        RECT 63.780 236.650 64.630 237.500 ;
        RECT 64.830 236.650 65.680 237.500 ;
        RECT 83.780 236.650 84.630 237.500 ;
        RECT 84.830 236.650 85.680 237.500 ;
        RECT 103.780 236.650 104.630 237.500 ;
        RECT 104.830 236.650 105.680 237.500 ;
        RECT 123.780 236.650 124.630 237.500 ;
        RECT 4.830 235.700 5.680 236.550 ;
        RECT 23.780 235.700 24.630 236.550 ;
        RECT 24.830 235.700 25.680 236.550 ;
        RECT 43.780 235.700 44.630 236.550 ;
        RECT 44.830 235.700 45.680 236.550 ;
        RECT 63.780 235.700 64.630 236.550 ;
        RECT 64.830 235.700 65.680 236.550 ;
        RECT 83.780 235.700 84.630 236.550 ;
        RECT 84.830 235.700 85.680 236.550 ;
        RECT 103.780 235.700 104.630 236.550 ;
        RECT 104.830 235.700 105.680 236.550 ;
        RECT 123.780 235.700 124.630 236.550 ;
        RECT 4.830 232.450 5.480 233.100 ;
        RECT 4.830 231.650 5.480 232.300 ;
        RECT 4.830 230.850 5.480 231.500 ;
        RECT 4.830 228.500 5.480 229.150 ;
        RECT 4.830 227.700 5.480 228.350 ;
        RECT 4.830 226.900 5.480 227.550 ;
        RECT 23.980 232.450 24.630 233.100 ;
        RECT 24.830 232.450 25.480 233.100 ;
        RECT 23.980 231.650 24.630 232.300 ;
        RECT 24.830 231.650 25.480 232.300 ;
        RECT 23.980 230.850 24.630 231.500 ;
        RECT 24.830 230.850 25.480 231.500 ;
        RECT 23.980 228.500 24.630 229.150 ;
        RECT 24.830 228.500 25.480 229.150 ;
        RECT 23.980 227.700 24.630 228.350 ;
        RECT 24.830 227.700 25.480 228.350 ;
        RECT 23.980 226.900 24.630 227.550 ;
        RECT 24.830 226.900 25.480 227.550 ;
        RECT 43.980 232.450 44.630 233.100 ;
        RECT 44.830 232.450 45.480 233.100 ;
        RECT 43.980 231.650 44.630 232.300 ;
        RECT 44.830 231.650 45.480 232.300 ;
        RECT 43.980 230.850 44.630 231.500 ;
        RECT 44.830 230.850 45.480 231.500 ;
        RECT 43.980 228.500 44.630 229.150 ;
        RECT 44.830 228.500 45.480 229.150 ;
        RECT 43.980 227.700 44.630 228.350 ;
        RECT 44.830 227.700 45.480 228.350 ;
        RECT 43.980 226.900 44.630 227.550 ;
        RECT 44.830 226.900 45.480 227.550 ;
        RECT 63.980 232.450 64.630 233.100 ;
        RECT 64.830 232.450 65.480 233.100 ;
        RECT 63.980 231.650 64.630 232.300 ;
        RECT 64.830 231.650 65.480 232.300 ;
        RECT 63.980 230.850 64.630 231.500 ;
        RECT 64.830 230.850 65.480 231.500 ;
        RECT 63.980 228.500 64.630 229.150 ;
        RECT 64.830 228.500 65.480 229.150 ;
        RECT 63.980 227.700 64.630 228.350 ;
        RECT 64.830 227.700 65.480 228.350 ;
        RECT 63.980 226.900 64.630 227.550 ;
        RECT 64.830 226.900 65.480 227.550 ;
        RECT 83.980 232.450 84.630 233.100 ;
        RECT 84.830 232.450 85.480 233.100 ;
        RECT 83.980 231.650 84.630 232.300 ;
        RECT 84.830 231.650 85.480 232.300 ;
        RECT 83.980 230.850 84.630 231.500 ;
        RECT 84.830 230.850 85.480 231.500 ;
        RECT 83.980 228.500 84.630 229.150 ;
        RECT 84.830 228.500 85.480 229.150 ;
        RECT 83.980 227.700 84.630 228.350 ;
        RECT 84.830 227.700 85.480 228.350 ;
        RECT 83.980 226.900 84.630 227.550 ;
        RECT 84.830 226.900 85.480 227.550 ;
        RECT 103.980 232.450 104.630 233.100 ;
        RECT 104.830 232.450 105.480 233.100 ;
        RECT 103.980 231.650 104.630 232.300 ;
        RECT 104.830 231.650 105.480 232.300 ;
        RECT 103.980 230.850 104.630 231.500 ;
        RECT 104.830 230.850 105.480 231.500 ;
        RECT 103.980 228.500 104.630 229.150 ;
        RECT 104.830 228.500 105.480 229.150 ;
        RECT 103.980 227.700 104.630 228.350 ;
        RECT 104.830 227.700 105.480 228.350 ;
        RECT 103.980 226.900 104.630 227.550 ;
        RECT 104.830 226.900 105.480 227.550 ;
        RECT 123.980 232.450 124.630 233.100 ;
        RECT 123.980 231.650 124.630 232.300 ;
        RECT 123.980 230.850 124.630 231.500 ;
        RECT 123.980 228.500 124.630 229.150 ;
        RECT 123.980 227.700 124.630 228.350 ;
        RECT 123.980 226.900 124.630 227.550 ;
        RECT 4.830 223.450 5.680 224.300 ;
        RECT 23.780 223.450 24.630 224.300 ;
        RECT 24.830 223.450 25.680 224.300 ;
        RECT 43.780 223.450 44.630 224.300 ;
        RECT 44.830 223.450 45.680 224.300 ;
        RECT 63.780 223.450 64.630 224.300 ;
        RECT 64.830 223.450 65.680 224.300 ;
        RECT 83.780 223.450 84.630 224.300 ;
        RECT 84.830 223.450 85.680 224.300 ;
        RECT 103.780 223.450 104.630 224.300 ;
        RECT 104.830 223.450 105.680 224.300 ;
        RECT 123.780 223.450 124.630 224.300 ;
        RECT 4.830 222.500 5.680 223.350 ;
        RECT 23.780 222.500 24.630 223.350 ;
        RECT 24.830 222.500 25.680 223.350 ;
        RECT 43.780 222.500 44.630 223.350 ;
        RECT 44.830 222.500 45.680 223.350 ;
        RECT 63.780 222.500 64.630 223.350 ;
        RECT 64.830 222.500 65.680 223.350 ;
        RECT 83.780 222.500 84.630 223.350 ;
        RECT 84.830 222.500 85.680 223.350 ;
        RECT 103.780 222.500 104.630 223.350 ;
        RECT 104.830 222.500 105.680 223.350 ;
        RECT 123.780 222.500 124.630 223.350 ;
        RECT 4.830 221.050 5.680 221.900 ;
        RECT 4.830 220.100 5.680 220.950 ;
        RECT 5.780 220.100 6.630 220.950 ;
        RECT 7.230 220.100 8.080 220.950 ;
        RECT 8.180 220.100 9.030 220.950 ;
        RECT 23.780 221.050 24.630 221.900 ;
        RECT 24.830 221.050 25.680 221.900 ;
        RECT 4.830 219.050 5.680 219.900 ;
        RECT 5.780 219.050 6.630 219.900 ;
        RECT 7.230 219.050 8.080 219.900 ;
        RECT 8.180 219.050 9.030 219.900 ;
        RECT 11.630 220.100 12.280 220.750 ;
        RECT 12.430 220.100 13.080 220.750 ;
        RECT 13.230 220.100 13.880 220.750 ;
        RECT 15.580 220.100 16.230 220.750 ;
        RECT 16.380 220.100 17.030 220.750 ;
        RECT 17.180 220.100 17.830 220.750 ;
        RECT 11.630 219.250 12.280 219.900 ;
        RECT 12.430 219.250 13.080 219.900 ;
        RECT 13.230 219.250 13.880 219.900 ;
        RECT 15.580 219.250 16.230 219.900 ;
        RECT 16.380 219.250 17.030 219.900 ;
        RECT 17.180 219.250 17.830 219.900 ;
        RECT 20.430 220.100 21.280 220.950 ;
        RECT 21.380 220.100 22.230 220.950 ;
        RECT 22.830 220.100 23.680 220.950 ;
        RECT 23.780 220.100 24.630 220.950 ;
        RECT 24.830 220.100 25.680 220.950 ;
        RECT 25.780 220.100 26.630 220.950 ;
        RECT 27.230 220.100 28.080 220.950 ;
        RECT 28.180 220.100 29.030 220.950 ;
        RECT 43.780 221.050 44.630 221.900 ;
        RECT 44.830 221.050 45.680 221.900 ;
        RECT 4.830 218.100 5.680 218.950 ;
        RECT 20.430 219.050 21.280 219.900 ;
        RECT 21.380 219.050 22.230 219.900 ;
        RECT 22.830 219.050 23.680 219.900 ;
        RECT 23.780 219.050 24.630 219.900 ;
        RECT 24.830 219.050 25.680 219.900 ;
        RECT 25.780 219.050 26.630 219.900 ;
        RECT 27.230 219.050 28.080 219.900 ;
        RECT 28.180 219.050 29.030 219.900 ;
        RECT 31.630 220.100 32.280 220.750 ;
        RECT 32.430 220.100 33.080 220.750 ;
        RECT 33.230 220.100 33.880 220.750 ;
        RECT 35.580 220.100 36.230 220.750 ;
        RECT 36.380 220.100 37.030 220.750 ;
        RECT 37.180 220.100 37.830 220.750 ;
        RECT 31.630 219.250 32.280 219.900 ;
        RECT 32.430 219.250 33.080 219.900 ;
        RECT 33.230 219.250 33.880 219.900 ;
        RECT 35.580 219.250 36.230 219.900 ;
        RECT 36.380 219.250 37.030 219.900 ;
        RECT 37.180 219.250 37.830 219.900 ;
        RECT 40.430 220.100 41.280 220.950 ;
        RECT 41.380 220.100 42.230 220.950 ;
        RECT 42.830 220.100 43.680 220.950 ;
        RECT 43.780 220.100 44.630 220.950 ;
        RECT 44.830 220.100 45.680 220.950 ;
        RECT 45.780 220.100 46.630 220.950 ;
        RECT 47.230 220.100 48.080 220.950 ;
        RECT 48.180 220.100 49.030 220.950 ;
        RECT 63.780 221.050 64.630 221.900 ;
        RECT 64.830 221.050 65.680 221.900 ;
        RECT 23.780 218.100 24.630 218.950 ;
        RECT 24.830 218.100 25.680 218.950 ;
        RECT 40.430 219.050 41.280 219.900 ;
        RECT 41.380 219.050 42.230 219.900 ;
        RECT 42.830 219.050 43.680 219.900 ;
        RECT 43.780 219.050 44.630 219.900 ;
        RECT 44.830 219.050 45.680 219.900 ;
        RECT 45.780 219.050 46.630 219.900 ;
        RECT 47.230 219.050 48.080 219.900 ;
        RECT 48.180 219.050 49.030 219.900 ;
        RECT 51.630 220.100 52.280 220.750 ;
        RECT 52.430 220.100 53.080 220.750 ;
        RECT 53.230 220.100 53.880 220.750 ;
        RECT 55.580 220.100 56.230 220.750 ;
        RECT 56.380 220.100 57.030 220.750 ;
        RECT 57.180 220.100 57.830 220.750 ;
        RECT 51.630 219.250 52.280 219.900 ;
        RECT 52.430 219.250 53.080 219.900 ;
        RECT 53.230 219.250 53.880 219.900 ;
        RECT 55.580 219.250 56.230 219.900 ;
        RECT 56.380 219.250 57.030 219.900 ;
        RECT 57.180 219.250 57.830 219.900 ;
        RECT 60.430 220.100 61.280 220.950 ;
        RECT 61.380 220.100 62.230 220.950 ;
        RECT 62.830 220.100 63.680 220.950 ;
        RECT 63.780 220.100 64.630 220.950 ;
        RECT 64.830 220.100 65.680 220.950 ;
        RECT 65.780 220.100 66.630 220.950 ;
        RECT 67.230 220.100 68.080 220.950 ;
        RECT 68.180 220.100 69.030 220.950 ;
        RECT 83.780 221.050 84.630 221.900 ;
        RECT 84.830 221.050 85.680 221.900 ;
        RECT 43.780 218.100 44.630 218.950 ;
        RECT 44.830 218.100 45.680 218.950 ;
        RECT 60.430 219.050 61.280 219.900 ;
        RECT 61.380 219.050 62.230 219.900 ;
        RECT 62.830 219.050 63.680 219.900 ;
        RECT 63.780 219.050 64.630 219.900 ;
        RECT 64.830 219.050 65.680 219.900 ;
        RECT 65.780 219.050 66.630 219.900 ;
        RECT 67.230 219.050 68.080 219.900 ;
        RECT 68.180 219.050 69.030 219.900 ;
        RECT 71.630 220.100 72.280 220.750 ;
        RECT 72.430 220.100 73.080 220.750 ;
        RECT 73.230 220.100 73.880 220.750 ;
        RECT 75.580 220.100 76.230 220.750 ;
        RECT 76.380 220.100 77.030 220.750 ;
        RECT 77.180 220.100 77.830 220.750 ;
        RECT 71.630 219.250 72.280 219.900 ;
        RECT 72.430 219.250 73.080 219.900 ;
        RECT 73.230 219.250 73.880 219.900 ;
        RECT 75.580 219.250 76.230 219.900 ;
        RECT 76.380 219.250 77.030 219.900 ;
        RECT 77.180 219.250 77.830 219.900 ;
        RECT 80.430 220.100 81.280 220.950 ;
        RECT 81.380 220.100 82.230 220.950 ;
        RECT 82.830 220.100 83.680 220.950 ;
        RECT 83.780 220.100 84.630 220.950 ;
        RECT 84.830 220.100 85.680 220.950 ;
        RECT 85.780 220.100 86.630 220.950 ;
        RECT 87.230 220.100 88.080 220.950 ;
        RECT 88.180 220.100 89.030 220.950 ;
        RECT 103.780 221.050 104.630 221.900 ;
        RECT 104.830 221.050 105.680 221.900 ;
        RECT 63.780 218.100 64.630 218.950 ;
        RECT 64.830 218.100 65.680 218.950 ;
        RECT 80.430 219.050 81.280 219.900 ;
        RECT 81.380 219.050 82.230 219.900 ;
        RECT 82.830 219.050 83.680 219.900 ;
        RECT 83.780 219.050 84.630 219.900 ;
        RECT 84.830 219.050 85.680 219.900 ;
        RECT 85.780 219.050 86.630 219.900 ;
        RECT 87.230 219.050 88.080 219.900 ;
        RECT 88.180 219.050 89.030 219.900 ;
        RECT 91.630 220.100 92.280 220.750 ;
        RECT 92.430 220.100 93.080 220.750 ;
        RECT 93.230 220.100 93.880 220.750 ;
        RECT 95.580 220.100 96.230 220.750 ;
        RECT 96.380 220.100 97.030 220.750 ;
        RECT 97.180 220.100 97.830 220.750 ;
        RECT 91.630 219.250 92.280 219.900 ;
        RECT 92.430 219.250 93.080 219.900 ;
        RECT 93.230 219.250 93.880 219.900 ;
        RECT 95.580 219.250 96.230 219.900 ;
        RECT 96.380 219.250 97.030 219.900 ;
        RECT 97.180 219.250 97.830 219.900 ;
        RECT 100.430 220.100 101.280 220.950 ;
        RECT 101.380 220.100 102.230 220.950 ;
        RECT 102.830 220.100 103.680 220.950 ;
        RECT 103.780 220.100 104.630 220.950 ;
        RECT 104.830 220.100 105.680 220.950 ;
        RECT 105.780 220.100 106.630 220.950 ;
        RECT 107.230 220.100 108.080 220.950 ;
        RECT 108.180 220.100 109.030 220.950 ;
        RECT 123.780 221.050 124.630 221.900 ;
        RECT 83.780 218.100 84.630 218.950 ;
        RECT 84.830 218.100 85.680 218.950 ;
        RECT 100.430 219.050 101.280 219.900 ;
        RECT 101.380 219.050 102.230 219.900 ;
        RECT 102.830 219.050 103.680 219.900 ;
        RECT 103.780 219.050 104.630 219.900 ;
        RECT 104.830 219.050 105.680 219.900 ;
        RECT 105.780 219.050 106.630 219.900 ;
        RECT 107.230 219.050 108.080 219.900 ;
        RECT 108.180 219.050 109.030 219.900 ;
        RECT 111.630 220.100 112.280 220.750 ;
        RECT 112.430 220.100 113.080 220.750 ;
        RECT 113.230 220.100 113.880 220.750 ;
        RECT 115.580 220.100 116.230 220.750 ;
        RECT 116.380 220.100 117.030 220.750 ;
        RECT 117.180 220.100 117.830 220.750 ;
        RECT 111.630 219.250 112.280 219.900 ;
        RECT 112.430 219.250 113.080 219.900 ;
        RECT 113.230 219.250 113.880 219.900 ;
        RECT 115.580 219.250 116.230 219.900 ;
        RECT 116.380 219.250 117.030 219.900 ;
        RECT 117.180 219.250 117.830 219.900 ;
        RECT 120.430 220.100 121.280 220.950 ;
        RECT 121.380 220.100 122.230 220.950 ;
        RECT 122.830 220.100 123.680 220.950 ;
        RECT 123.780 220.100 124.630 220.950 ;
        RECT 103.780 218.100 104.630 218.950 ;
        RECT 104.830 218.100 105.680 218.950 ;
        RECT 120.430 219.050 121.280 219.900 ;
        RECT 121.380 219.050 122.230 219.900 ;
        RECT 122.830 219.050 123.680 219.900 ;
        RECT 123.780 219.050 124.630 219.900 ;
        RECT 123.780 218.100 124.630 218.950 ;
        RECT 4.830 216.650 5.680 217.500 ;
        RECT 23.780 216.650 24.630 217.500 ;
        RECT 24.830 216.650 25.680 217.500 ;
        RECT 43.780 216.650 44.630 217.500 ;
        RECT 44.830 216.650 45.680 217.500 ;
        RECT 63.780 216.650 64.630 217.500 ;
        RECT 64.830 216.650 65.680 217.500 ;
        RECT 83.780 216.650 84.630 217.500 ;
        RECT 84.830 216.650 85.680 217.500 ;
        RECT 103.780 216.650 104.630 217.500 ;
        RECT 104.830 216.650 105.680 217.500 ;
        RECT 123.780 216.650 124.630 217.500 ;
        RECT 4.830 215.700 5.680 216.550 ;
        RECT 23.780 215.700 24.630 216.550 ;
        RECT 24.830 215.700 25.680 216.550 ;
        RECT 43.780 215.700 44.630 216.550 ;
        RECT 44.830 215.700 45.680 216.550 ;
        RECT 63.780 215.700 64.630 216.550 ;
        RECT 64.830 215.700 65.680 216.550 ;
        RECT 83.780 215.700 84.630 216.550 ;
        RECT 84.830 215.700 85.680 216.550 ;
        RECT 103.780 215.700 104.630 216.550 ;
        RECT 104.830 215.700 105.680 216.550 ;
        RECT 123.780 215.700 124.630 216.550 ;
        RECT 4.830 212.450 5.480 213.100 ;
        RECT 4.830 211.650 5.480 212.300 ;
        RECT 4.830 210.850 5.480 211.500 ;
        RECT 4.830 208.500 5.480 209.150 ;
        RECT 4.830 207.700 5.480 208.350 ;
        RECT 4.830 206.900 5.480 207.550 ;
        RECT 23.980 212.450 24.630 213.100 ;
        RECT 24.830 212.450 25.480 213.100 ;
        RECT 23.980 211.650 24.630 212.300 ;
        RECT 24.830 211.650 25.480 212.300 ;
        RECT 23.980 210.850 24.630 211.500 ;
        RECT 24.830 210.850 25.480 211.500 ;
        RECT 23.980 208.500 24.630 209.150 ;
        RECT 24.830 208.500 25.480 209.150 ;
        RECT 23.980 207.700 24.630 208.350 ;
        RECT 24.830 207.700 25.480 208.350 ;
        RECT 23.980 206.900 24.630 207.550 ;
        RECT 24.830 206.900 25.480 207.550 ;
        RECT 43.980 212.450 44.630 213.100 ;
        RECT 44.830 212.450 45.480 213.100 ;
        RECT 43.980 211.650 44.630 212.300 ;
        RECT 44.830 211.650 45.480 212.300 ;
        RECT 43.980 210.850 44.630 211.500 ;
        RECT 44.830 210.850 45.480 211.500 ;
        RECT 43.980 208.500 44.630 209.150 ;
        RECT 44.830 208.500 45.480 209.150 ;
        RECT 43.980 207.700 44.630 208.350 ;
        RECT 44.830 207.700 45.480 208.350 ;
        RECT 43.980 206.900 44.630 207.550 ;
        RECT 44.830 206.900 45.480 207.550 ;
        RECT 63.980 212.450 64.630 213.100 ;
        RECT 64.830 212.450 65.480 213.100 ;
        RECT 63.980 211.650 64.630 212.300 ;
        RECT 64.830 211.650 65.480 212.300 ;
        RECT 63.980 210.850 64.630 211.500 ;
        RECT 64.830 210.850 65.480 211.500 ;
        RECT 63.980 208.500 64.630 209.150 ;
        RECT 64.830 208.500 65.480 209.150 ;
        RECT 63.980 207.700 64.630 208.350 ;
        RECT 64.830 207.700 65.480 208.350 ;
        RECT 63.980 206.900 64.630 207.550 ;
        RECT 64.830 206.900 65.480 207.550 ;
        RECT 83.980 212.450 84.630 213.100 ;
        RECT 84.830 212.450 85.480 213.100 ;
        RECT 83.980 211.650 84.630 212.300 ;
        RECT 84.830 211.650 85.480 212.300 ;
        RECT 83.980 210.850 84.630 211.500 ;
        RECT 84.830 210.850 85.480 211.500 ;
        RECT 83.980 208.500 84.630 209.150 ;
        RECT 84.830 208.500 85.480 209.150 ;
        RECT 83.980 207.700 84.630 208.350 ;
        RECT 84.830 207.700 85.480 208.350 ;
        RECT 83.980 206.900 84.630 207.550 ;
        RECT 84.830 206.900 85.480 207.550 ;
        RECT 103.980 212.450 104.630 213.100 ;
        RECT 104.830 212.450 105.480 213.100 ;
        RECT 103.980 211.650 104.630 212.300 ;
        RECT 104.830 211.650 105.480 212.300 ;
        RECT 103.980 210.850 104.630 211.500 ;
        RECT 104.830 210.850 105.480 211.500 ;
        RECT 103.980 208.500 104.630 209.150 ;
        RECT 104.830 208.500 105.480 209.150 ;
        RECT 103.980 207.700 104.630 208.350 ;
        RECT 104.830 207.700 105.480 208.350 ;
        RECT 103.980 206.900 104.630 207.550 ;
        RECT 104.830 206.900 105.480 207.550 ;
        RECT 123.980 212.450 124.630 213.100 ;
        RECT 123.980 211.650 124.630 212.300 ;
        RECT 123.980 210.850 124.630 211.500 ;
        RECT 123.980 208.500 124.630 209.150 ;
        RECT 123.980 207.700 124.630 208.350 ;
        RECT 123.980 206.900 124.630 207.550 ;
        RECT 4.830 203.450 5.680 204.300 ;
        RECT 23.780 203.450 24.630 204.300 ;
        RECT 24.830 203.450 25.680 204.300 ;
        RECT 43.780 203.450 44.630 204.300 ;
        RECT 44.830 203.450 45.680 204.300 ;
        RECT 63.780 203.450 64.630 204.300 ;
        RECT 64.830 203.450 65.680 204.300 ;
        RECT 83.780 203.450 84.630 204.300 ;
        RECT 84.830 203.450 85.680 204.300 ;
        RECT 103.780 203.450 104.630 204.300 ;
        RECT 104.830 203.450 105.680 204.300 ;
        RECT 123.780 203.450 124.630 204.300 ;
        RECT 4.830 202.500 5.680 203.350 ;
        RECT 23.780 202.500 24.630 203.350 ;
        RECT 24.830 202.500 25.680 203.350 ;
        RECT 43.780 202.500 44.630 203.350 ;
        RECT 44.830 202.500 45.680 203.350 ;
        RECT 63.780 202.500 64.630 203.350 ;
        RECT 64.830 202.500 65.680 203.350 ;
        RECT 83.780 202.500 84.630 203.350 ;
        RECT 84.830 202.500 85.680 203.350 ;
        RECT 103.780 202.500 104.630 203.350 ;
        RECT 104.830 202.500 105.680 203.350 ;
        RECT 123.780 202.500 124.630 203.350 ;
        RECT 4.830 201.050 5.680 201.900 ;
        RECT 4.830 200.100 5.680 200.950 ;
        RECT 5.780 200.100 6.630 200.950 ;
        RECT 7.230 200.100 8.080 200.950 ;
        RECT 8.180 200.100 9.030 200.950 ;
        RECT 23.780 201.050 24.630 201.900 ;
        RECT 24.830 201.050 25.680 201.900 ;
        RECT 11.630 200.100 12.280 200.750 ;
        RECT 12.430 200.100 13.080 200.750 ;
        RECT 13.230 200.100 13.880 200.750 ;
        RECT 15.580 200.100 16.230 200.750 ;
        RECT 16.380 200.100 17.030 200.750 ;
        RECT 17.180 200.100 17.830 200.750 ;
        RECT 20.430 200.100 21.280 200.950 ;
        RECT 21.380 200.100 22.230 200.950 ;
        RECT 22.830 200.100 23.680 200.950 ;
        RECT 23.780 200.100 24.630 200.950 ;
        RECT 24.830 200.100 25.680 200.950 ;
        RECT 25.780 200.100 26.630 200.950 ;
        RECT 27.230 200.100 28.080 200.950 ;
        RECT 28.180 200.100 29.030 200.950 ;
        RECT 43.780 201.050 44.630 201.900 ;
        RECT 44.830 201.050 45.680 201.900 ;
        RECT 31.630 200.100 32.280 200.750 ;
        RECT 32.430 200.100 33.080 200.750 ;
        RECT 33.230 200.100 33.880 200.750 ;
        RECT 35.580 200.100 36.230 200.750 ;
        RECT 36.380 200.100 37.030 200.750 ;
        RECT 37.180 200.100 37.830 200.750 ;
        RECT 40.430 200.100 41.280 200.950 ;
        RECT 41.380 200.100 42.230 200.950 ;
        RECT 42.830 200.100 43.680 200.950 ;
        RECT 43.780 200.100 44.630 200.950 ;
        RECT 44.830 200.100 45.680 200.950 ;
        RECT 45.780 200.100 46.630 200.950 ;
        RECT 47.230 200.100 48.080 200.950 ;
        RECT 48.180 200.100 49.030 200.950 ;
        RECT 63.780 201.050 64.630 201.900 ;
        RECT 64.830 201.050 65.680 201.900 ;
        RECT 51.630 200.100 52.280 200.750 ;
        RECT 52.430 200.100 53.080 200.750 ;
        RECT 53.230 200.100 53.880 200.750 ;
        RECT 55.580 200.100 56.230 200.750 ;
        RECT 56.380 200.100 57.030 200.750 ;
        RECT 57.180 200.100 57.830 200.750 ;
        RECT 60.430 200.100 61.280 200.950 ;
        RECT 61.380 200.100 62.230 200.950 ;
        RECT 62.830 200.100 63.680 200.950 ;
        RECT 63.780 200.100 64.630 200.950 ;
        RECT 64.830 200.100 65.680 200.950 ;
        RECT 65.780 200.100 66.630 200.950 ;
        RECT 67.230 200.100 68.080 200.950 ;
        RECT 68.180 200.100 69.030 200.950 ;
        RECT 83.780 201.050 84.630 201.900 ;
        RECT 84.830 201.050 85.680 201.900 ;
        RECT 71.630 200.100 72.280 200.750 ;
        RECT 72.430 200.100 73.080 200.750 ;
        RECT 73.230 200.100 73.880 200.750 ;
        RECT 75.580 200.100 76.230 200.750 ;
        RECT 76.380 200.100 77.030 200.750 ;
        RECT 77.180 200.100 77.830 200.750 ;
        RECT 80.430 200.100 81.280 200.950 ;
        RECT 81.380 200.100 82.230 200.950 ;
        RECT 82.830 200.100 83.680 200.950 ;
        RECT 83.780 200.100 84.630 200.950 ;
        RECT 84.830 200.100 85.680 200.950 ;
        RECT 85.780 200.100 86.630 200.950 ;
        RECT 87.230 200.100 88.080 200.950 ;
        RECT 88.180 200.100 89.030 200.950 ;
        RECT 103.780 201.050 104.630 201.900 ;
        RECT 104.830 201.050 105.680 201.900 ;
        RECT 91.630 200.100 92.280 200.750 ;
        RECT 92.430 200.100 93.080 200.750 ;
        RECT 93.230 200.100 93.880 200.750 ;
        RECT 95.580 200.100 96.230 200.750 ;
        RECT 96.380 200.100 97.030 200.750 ;
        RECT 97.180 200.100 97.830 200.750 ;
        RECT 100.430 200.100 101.280 200.950 ;
        RECT 101.380 200.100 102.230 200.950 ;
        RECT 102.830 200.100 103.680 200.950 ;
        RECT 103.780 200.100 104.630 200.950 ;
        RECT 104.830 200.100 105.680 200.950 ;
        RECT 105.780 200.100 106.630 200.950 ;
        RECT 107.230 200.100 108.080 200.950 ;
        RECT 108.180 200.100 109.030 200.950 ;
        RECT 123.780 201.050 124.630 201.900 ;
        RECT 111.630 200.100 112.280 200.750 ;
        RECT 112.430 200.100 113.080 200.750 ;
        RECT 113.230 200.100 113.880 200.750 ;
        RECT 115.580 200.100 116.230 200.750 ;
        RECT 116.380 200.100 117.030 200.750 ;
        RECT 117.180 200.100 117.830 200.750 ;
        RECT 120.430 200.100 121.280 200.950 ;
        RECT 121.380 200.100 122.230 200.950 ;
        RECT 122.830 200.100 123.680 200.950 ;
        RECT 123.780 200.100 124.630 200.950 ;
        RECT 11.245 179.305 11.565 179.625 ;
        RECT 11.685 179.305 12.005 179.625 ;
        RECT 11.245 178.905 11.565 179.225 ;
        RECT 11.685 178.905 12.005 179.225 ;
        RECT 20.960 179.205 21.280 179.525 ;
        RECT 21.400 179.205 21.720 179.525 ;
        RECT 20.960 178.805 21.280 179.125 ;
        RECT 21.400 178.805 21.720 179.125 ;
        RECT 12.680 161.995 13.000 162.315 ;
        RECT 13.120 161.995 13.440 162.315 ;
        RECT 11.630 139.250 12.280 139.900 ;
        RECT 12.430 139.250 13.080 139.900 ;
        RECT 13.230 139.250 13.880 139.900 ;
        RECT 15.580 139.250 16.230 139.900 ;
        RECT 16.380 139.250 17.030 139.900 ;
        RECT 17.180 139.250 17.830 139.900 ;
        RECT 31.630 139.250 32.280 139.900 ;
        RECT 32.430 139.250 33.080 139.900 ;
        RECT 33.230 139.250 33.880 139.900 ;
        RECT 35.580 139.250 36.230 139.900 ;
        RECT 36.380 139.250 37.030 139.900 ;
        RECT 37.180 139.250 37.830 139.900 ;
        RECT 51.630 139.250 52.280 139.900 ;
        RECT 52.430 139.250 53.080 139.900 ;
        RECT 53.230 139.250 53.880 139.900 ;
        RECT 55.580 139.250 56.230 139.900 ;
        RECT 56.380 139.250 57.030 139.900 ;
        RECT 57.180 139.250 57.830 139.900 ;
        RECT 71.630 139.250 72.280 139.900 ;
        RECT 72.430 139.250 73.080 139.900 ;
        RECT 73.230 139.250 73.880 139.900 ;
        RECT 75.580 139.250 76.230 139.900 ;
        RECT 76.380 139.250 77.030 139.900 ;
        RECT 77.180 139.250 77.830 139.900 ;
        RECT 91.630 139.250 92.280 139.900 ;
        RECT 92.430 139.250 93.080 139.900 ;
        RECT 93.230 139.250 93.880 139.900 ;
        RECT 95.580 139.250 96.230 139.900 ;
        RECT 96.380 139.250 97.030 139.900 ;
        RECT 97.180 139.250 97.830 139.900 ;
        RECT 111.630 139.250 112.280 139.900 ;
        RECT 112.430 139.250 113.080 139.900 ;
        RECT 113.230 139.250 113.880 139.900 ;
        RECT 115.580 139.250 116.230 139.900 ;
        RECT 116.380 139.250 117.030 139.900 ;
        RECT 117.180 139.250 117.830 139.900 ;
        RECT 4.830 132.450 5.480 133.100 ;
        RECT 4.830 131.650 5.480 132.300 ;
        RECT 4.830 130.850 5.480 131.500 ;
        RECT 4.830 128.500 5.480 129.150 ;
        RECT 4.830 127.700 5.480 128.350 ;
        RECT 4.830 126.900 5.480 127.550 ;
        RECT 23.980 132.450 24.630 133.100 ;
        RECT 24.830 132.450 25.480 133.100 ;
        RECT 23.980 131.650 24.630 132.300 ;
        RECT 24.830 131.650 25.480 132.300 ;
        RECT 23.980 130.850 24.630 131.500 ;
        RECT 24.830 130.850 25.480 131.500 ;
        RECT 23.980 128.500 24.630 129.150 ;
        RECT 24.830 128.500 25.480 129.150 ;
        RECT 23.980 127.700 24.630 128.350 ;
        RECT 24.830 127.700 25.480 128.350 ;
        RECT 23.980 126.900 24.630 127.550 ;
        RECT 24.830 126.900 25.480 127.550 ;
        RECT 43.980 132.450 44.630 133.100 ;
        RECT 44.830 132.450 45.480 133.100 ;
        RECT 43.980 131.650 44.630 132.300 ;
        RECT 44.830 131.650 45.480 132.300 ;
        RECT 43.980 130.850 44.630 131.500 ;
        RECT 44.830 130.850 45.480 131.500 ;
        RECT 43.980 128.500 44.630 129.150 ;
        RECT 44.830 128.500 45.480 129.150 ;
        RECT 43.980 127.700 44.630 128.350 ;
        RECT 44.830 127.700 45.480 128.350 ;
        RECT 43.980 126.900 44.630 127.550 ;
        RECT 44.830 126.900 45.480 127.550 ;
        RECT 63.980 132.450 64.630 133.100 ;
        RECT 64.830 132.450 65.480 133.100 ;
        RECT 63.980 131.650 64.630 132.300 ;
        RECT 64.830 131.650 65.480 132.300 ;
        RECT 63.980 130.850 64.630 131.500 ;
        RECT 64.830 130.850 65.480 131.500 ;
        RECT 63.980 128.500 64.630 129.150 ;
        RECT 64.830 128.500 65.480 129.150 ;
        RECT 63.980 127.700 64.630 128.350 ;
        RECT 64.830 127.700 65.480 128.350 ;
        RECT 63.980 126.900 64.630 127.550 ;
        RECT 64.830 126.900 65.480 127.550 ;
        RECT 83.980 132.450 84.630 133.100 ;
        RECT 84.830 132.450 85.480 133.100 ;
        RECT 83.980 131.650 84.630 132.300 ;
        RECT 84.830 131.650 85.480 132.300 ;
        RECT 83.980 130.850 84.630 131.500 ;
        RECT 84.830 130.850 85.480 131.500 ;
        RECT 83.980 128.500 84.630 129.150 ;
        RECT 84.830 128.500 85.480 129.150 ;
        RECT 83.980 127.700 84.630 128.350 ;
        RECT 84.830 127.700 85.480 128.350 ;
        RECT 83.980 126.900 84.630 127.550 ;
        RECT 84.830 126.900 85.480 127.550 ;
        RECT 103.980 132.450 104.630 133.100 ;
        RECT 104.830 132.450 105.480 133.100 ;
        RECT 103.980 131.650 104.630 132.300 ;
        RECT 104.830 131.650 105.480 132.300 ;
        RECT 103.980 130.850 104.630 131.500 ;
        RECT 104.830 130.850 105.480 131.500 ;
        RECT 103.980 128.500 104.630 129.150 ;
        RECT 104.830 128.500 105.480 129.150 ;
        RECT 103.980 127.700 104.630 128.350 ;
        RECT 104.830 127.700 105.480 128.350 ;
        RECT 103.980 126.900 104.630 127.550 ;
        RECT 104.830 126.900 105.480 127.550 ;
        RECT 123.980 132.450 124.630 133.100 ;
        RECT 123.980 131.650 124.630 132.300 ;
        RECT 123.980 130.850 124.630 131.500 ;
        RECT 123.980 128.500 124.630 129.150 ;
        RECT 123.980 127.700 124.630 128.350 ;
        RECT 123.980 126.900 124.630 127.550 ;
        RECT 11.630 120.100 12.280 120.750 ;
        RECT 12.430 120.100 13.080 120.750 ;
        RECT 13.230 120.100 13.880 120.750 ;
        RECT 15.580 120.100 16.230 120.750 ;
        RECT 16.380 120.100 17.030 120.750 ;
        RECT 17.180 120.100 17.830 120.750 ;
        RECT 11.630 119.250 12.280 119.900 ;
        RECT 12.430 119.250 13.080 119.900 ;
        RECT 13.230 119.250 13.880 119.900 ;
        RECT 15.580 119.250 16.230 119.900 ;
        RECT 16.380 119.250 17.030 119.900 ;
        RECT 17.180 119.250 17.830 119.900 ;
        RECT 31.630 120.100 32.280 120.750 ;
        RECT 32.430 120.100 33.080 120.750 ;
        RECT 33.230 120.100 33.880 120.750 ;
        RECT 35.580 120.100 36.230 120.750 ;
        RECT 36.380 120.100 37.030 120.750 ;
        RECT 37.180 120.100 37.830 120.750 ;
        RECT 31.630 119.250 32.280 119.900 ;
        RECT 32.430 119.250 33.080 119.900 ;
        RECT 33.230 119.250 33.880 119.900 ;
        RECT 35.580 119.250 36.230 119.900 ;
        RECT 36.380 119.250 37.030 119.900 ;
        RECT 37.180 119.250 37.830 119.900 ;
        RECT 51.630 120.100 52.280 120.750 ;
        RECT 52.430 120.100 53.080 120.750 ;
        RECT 53.230 120.100 53.880 120.750 ;
        RECT 55.580 120.100 56.230 120.750 ;
        RECT 56.380 120.100 57.030 120.750 ;
        RECT 57.180 120.100 57.830 120.750 ;
        RECT 51.630 119.250 52.280 119.900 ;
        RECT 52.430 119.250 53.080 119.900 ;
        RECT 53.230 119.250 53.880 119.900 ;
        RECT 55.580 119.250 56.230 119.900 ;
        RECT 56.380 119.250 57.030 119.900 ;
        RECT 57.180 119.250 57.830 119.900 ;
        RECT 71.630 120.100 72.280 120.750 ;
        RECT 72.430 120.100 73.080 120.750 ;
        RECT 73.230 120.100 73.880 120.750 ;
        RECT 75.580 120.100 76.230 120.750 ;
        RECT 76.380 120.100 77.030 120.750 ;
        RECT 77.180 120.100 77.830 120.750 ;
        RECT 71.630 119.250 72.280 119.900 ;
        RECT 72.430 119.250 73.080 119.900 ;
        RECT 73.230 119.250 73.880 119.900 ;
        RECT 75.580 119.250 76.230 119.900 ;
        RECT 76.380 119.250 77.030 119.900 ;
        RECT 77.180 119.250 77.830 119.900 ;
        RECT 91.630 120.100 92.280 120.750 ;
        RECT 92.430 120.100 93.080 120.750 ;
        RECT 93.230 120.100 93.880 120.750 ;
        RECT 95.580 120.100 96.230 120.750 ;
        RECT 96.380 120.100 97.030 120.750 ;
        RECT 97.180 120.100 97.830 120.750 ;
        RECT 91.630 119.250 92.280 119.900 ;
        RECT 92.430 119.250 93.080 119.900 ;
        RECT 93.230 119.250 93.880 119.900 ;
        RECT 95.580 119.250 96.230 119.900 ;
        RECT 96.380 119.250 97.030 119.900 ;
        RECT 97.180 119.250 97.830 119.900 ;
        RECT 111.630 120.100 112.280 120.750 ;
        RECT 112.430 120.100 113.080 120.750 ;
        RECT 113.230 120.100 113.880 120.750 ;
        RECT 115.580 120.100 116.230 120.750 ;
        RECT 116.380 120.100 117.030 120.750 ;
        RECT 117.180 120.100 117.830 120.750 ;
        RECT 111.630 119.250 112.280 119.900 ;
        RECT 112.430 119.250 113.080 119.900 ;
        RECT 113.230 119.250 113.880 119.900 ;
        RECT 115.580 119.250 116.230 119.900 ;
        RECT 116.380 119.250 117.030 119.900 ;
        RECT 117.180 119.250 117.830 119.900 ;
        RECT 4.830 112.450 5.480 113.100 ;
        RECT 4.830 111.650 5.480 112.300 ;
        RECT 4.830 110.850 5.480 111.500 ;
        RECT 4.830 108.500 5.480 109.150 ;
        RECT 4.830 107.700 5.480 108.350 ;
        RECT 4.830 106.900 5.480 107.550 ;
        RECT 23.980 112.450 24.630 113.100 ;
        RECT 24.830 112.450 25.480 113.100 ;
        RECT 23.980 111.650 24.630 112.300 ;
        RECT 24.830 111.650 25.480 112.300 ;
        RECT 23.980 110.850 24.630 111.500 ;
        RECT 24.830 110.850 25.480 111.500 ;
        RECT 23.980 108.500 24.630 109.150 ;
        RECT 24.830 108.500 25.480 109.150 ;
        RECT 23.980 107.700 24.630 108.350 ;
        RECT 24.830 107.700 25.480 108.350 ;
        RECT 23.980 106.900 24.630 107.550 ;
        RECT 24.830 106.900 25.480 107.550 ;
        RECT 43.980 112.450 44.630 113.100 ;
        RECT 44.830 112.450 45.480 113.100 ;
        RECT 43.980 111.650 44.630 112.300 ;
        RECT 44.830 111.650 45.480 112.300 ;
        RECT 43.980 110.850 44.630 111.500 ;
        RECT 44.830 110.850 45.480 111.500 ;
        RECT 43.980 108.500 44.630 109.150 ;
        RECT 44.830 108.500 45.480 109.150 ;
        RECT 43.980 107.700 44.630 108.350 ;
        RECT 44.830 107.700 45.480 108.350 ;
        RECT 43.980 106.900 44.630 107.550 ;
        RECT 44.830 106.900 45.480 107.550 ;
        RECT 63.980 112.450 64.630 113.100 ;
        RECT 64.830 112.450 65.480 113.100 ;
        RECT 63.980 111.650 64.630 112.300 ;
        RECT 64.830 111.650 65.480 112.300 ;
        RECT 63.980 110.850 64.630 111.500 ;
        RECT 64.830 110.850 65.480 111.500 ;
        RECT 63.980 108.500 64.630 109.150 ;
        RECT 64.830 108.500 65.480 109.150 ;
        RECT 63.980 107.700 64.630 108.350 ;
        RECT 64.830 107.700 65.480 108.350 ;
        RECT 63.980 106.900 64.630 107.550 ;
        RECT 64.830 106.900 65.480 107.550 ;
        RECT 83.980 112.450 84.630 113.100 ;
        RECT 84.830 112.450 85.480 113.100 ;
        RECT 83.980 111.650 84.630 112.300 ;
        RECT 84.830 111.650 85.480 112.300 ;
        RECT 83.980 110.850 84.630 111.500 ;
        RECT 84.830 110.850 85.480 111.500 ;
        RECT 83.980 108.500 84.630 109.150 ;
        RECT 84.830 108.500 85.480 109.150 ;
        RECT 83.980 107.700 84.630 108.350 ;
        RECT 84.830 107.700 85.480 108.350 ;
        RECT 83.980 106.900 84.630 107.550 ;
        RECT 84.830 106.900 85.480 107.550 ;
        RECT 103.980 112.450 104.630 113.100 ;
        RECT 104.830 112.450 105.480 113.100 ;
        RECT 103.980 111.650 104.630 112.300 ;
        RECT 104.830 111.650 105.480 112.300 ;
        RECT 103.980 110.850 104.630 111.500 ;
        RECT 104.830 110.850 105.480 111.500 ;
        RECT 103.980 108.500 104.630 109.150 ;
        RECT 104.830 108.500 105.480 109.150 ;
        RECT 103.980 107.700 104.630 108.350 ;
        RECT 104.830 107.700 105.480 108.350 ;
        RECT 103.980 106.900 104.630 107.550 ;
        RECT 104.830 106.900 105.480 107.550 ;
        RECT 123.980 112.450 124.630 113.100 ;
        RECT 123.980 111.650 124.630 112.300 ;
        RECT 123.980 110.850 124.630 111.500 ;
        RECT 123.980 108.500 124.630 109.150 ;
        RECT 123.980 107.700 124.630 108.350 ;
        RECT 123.980 106.900 124.630 107.550 ;
        RECT 11.630 100.100 12.280 100.750 ;
        RECT 12.430 100.100 13.080 100.750 ;
        RECT 13.230 100.100 13.880 100.750 ;
        RECT 15.580 100.100 16.230 100.750 ;
        RECT 16.380 100.100 17.030 100.750 ;
        RECT 17.180 100.100 17.830 100.750 ;
        RECT 11.630 99.250 12.280 99.900 ;
        RECT 12.430 99.250 13.080 99.900 ;
        RECT 13.230 99.250 13.880 99.900 ;
        RECT 15.580 99.250 16.230 99.900 ;
        RECT 16.380 99.250 17.030 99.900 ;
        RECT 17.180 99.250 17.830 99.900 ;
        RECT 31.630 100.100 32.280 100.750 ;
        RECT 32.430 100.100 33.080 100.750 ;
        RECT 33.230 100.100 33.880 100.750 ;
        RECT 35.580 100.100 36.230 100.750 ;
        RECT 36.380 100.100 37.030 100.750 ;
        RECT 37.180 100.100 37.830 100.750 ;
        RECT 31.630 99.250 32.280 99.900 ;
        RECT 32.430 99.250 33.080 99.900 ;
        RECT 33.230 99.250 33.880 99.900 ;
        RECT 35.580 99.250 36.230 99.900 ;
        RECT 36.380 99.250 37.030 99.900 ;
        RECT 37.180 99.250 37.830 99.900 ;
        RECT 51.630 100.100 52.280 100.750 ;
        RECT 52.430 100.100 53.080 100.750 ;
        RECT 53.230 100.100 53.880 100.750 ;
        RECT 55.580 100.100 56.230 100.750 ;
        RECT 56.380 100.100 57.030 100.750 ;
        RECT 57.180 100.100 57.830 100.750 ;
        RECT 51.630 99.250 52.280 99.900 ;
        RECT 52.430 99.250 53.080 99.900 ;
        RECT 53.230 99.250 53.880 99.900 ;
        RECT 55.580 99.250 56.230 99.900 ;
        RECT 56.380 99.250 57.030 99.900 ;
        RECT 57.180 99.250 57.830 99.900 ;
        RECT 71.630 100.100 72.280 100.750 ;
        RECT 72.430 100.100 73.080 100.750 ;
        RECT 73.230 100.100 73.880 100.750 ;
        RECT 75.580 100.100 76.230 100.750 ;
        RECT 76.380 100.100 77.030 100.750 ;
        RECT 77.180 100.100 77.830 100.750 ;
        RECT 71.630 99.250 72.280 99.900 ;
        RECT 72.430 99.250 73.080 99.900 ;
        RECT 73.230 99.250 73.880 99.900 ;
        RECT 75.580 99.250 76.230 99.900 ;
        RECT 76.380 99.250 77.030 99.900 ;
        RECT 77.180 99.250 77.830 99.900 ;
        RECT 91.630 100.100 92.280 100.750 ;
        RECT 92.430 100.100 93.080 100.750 ;
        RECT 93.230 100.100 93.880 100.750 ;
        RECT 95.580 100.100 96.230 100.750 ;
        RECT 96.380 100.100 97.030 100.750 ;
        RECT 97.180 100.100 97.830 100.750 ;
        RECT 91.630 99.250 92.280 99.900 ;
        RECT 92.430 99.250 93.080 99.900 ;
        RECT 93.230 99.250 93.880 99.900 ;
        RECT 95.580 99.250 96.230 99.900 ;
        RECT 96.380 99.250 97.030 99.900 ;
        RECT 97.180 99.250 97.830 99.900 ;
        RECT 111.630 100.100 112.280 100.750 ;
        RECT 112.430 100.100 113.080 100.750 ;
        RECT 113.230 100.100 113.880 100.750 ;
        RECT 115.580 100.100 116.230 100.750 ;
        RECT 116.380 100.100 117.030 100.750 ;
        RECT 117.180 100.100 117.830 100.750 ;
        RECT 111.630 99.250 112.280 99.900 ;
        RECT 112.430 99.250 113.080 99.900 ;
        RECT 113.230 99.250 113.880 99.900 ;
        RECT 115.580 99.250 116.230 99.900 ;
        RECT 116.380 99.250 117.030 99.900 ;
        RECT 117.180 99.250 117.830 99.900 ;
        RECT 4.830 92.450 5.480 93.100 ;
        RECT 4.830 91.650 5.480 92.300 ;
        RECT 4.830 90.850 5.480 91.500 ;
        RECT 4.830 88.500 5.480 89.150 ;
        RECT 4.830 87.700 5.480 88.350 ;
        RECT 4.830 86.900 5.480 87.550 ;
        RECT 23.980 92.450 24.630 93.100 ;
        RECT 24.830 92.450 25.480 93.100 ;
        RECT 23.980 91.650 24.630 92.300 ;
        RECT 24.830 91.650 25.480 92.300 ;
        RECT 23.980 90.850 24.630 91.500 ;
        RECT 24.830 90.850 25.480 91.500 ;
        RECT 23.980 88.500 24.630 89.150 ;
        RECT 24.830 88.500 25.480 89.150 ;
        RECT 23.980 87.700 24.630 88.350 ;
        RECT 24.830 87.700 25.480 88.350 ;
        RECT 23.980 86.900 24.630 87.550 ;
        RECT 24.830 86.900 25.480 87.550 ;
        RECT 43.980 92.450 44.630 93.100 ;
        RECT 44.830 92.450 45.480 93.100 ;
        RECT 43.980 91.650 44.630 92.300 ;
        RECT 44.830 91.650 45.480 92.300 ;
        RECT 43.980 90.850 44.630 91.500 ;
        RECT 44.830 90.850 45.480 91.500 ;
        RECT 43.980 88.500 44.630 89.150 ;
        RECT 44.830 88.500 45.480 89.150 ;
        RECT 43.980 87.700 44.630 88.350 ;
        RECT 44.830 87.700 45.480 88.350 ;
        RECT 43.980 86.900 44.630 87.550 ;
        RECT 44.830 86.900 45.480 87.550 ;
        RECT 63.980 92.450 64.630 93.100 ;
        RECT 64.830 92.450 65.480 93.100 ;
        RECT 63.980 91.650 64.630 92.300 ;
        RECT 64.830 91.650 65.480 92.300 ;
        RECT 63.980 90.850 64.630 91.500 ;
        RECT 64.830 90.850 65.480 91.500 ;
        RECT 63.980 88.500 64.630 89.150 ;
        RECT 64.830 88.500 65.480 89.150 ;
        RECT 63.980 87.700 64.630 88.350 ;
        RECT 64.830 87.700 65.480 88.350 ;
        RECT 63.980 86.900 64.630 87.550 ;
        RECT 64.830 86.900 65.480 87.550 ;
        RECT 83.980 92.450 84.630 93.100 ;
        RECT 84.830 92.450 85.480 93.100 ;
        RECT 83.980 91.650 84.630 92.300 ;
        RECT 84.830 91.650 85.480 92.300 ;
        RECT 83.980 90.850 84.630 91.500 ;
        RECT 84.830 90.850 85.480 91.500 ;
        RECT 83.980 88.500 84.630 89.150 ;
        RECT 84.830 88.500 85.480 89.150 ;
        RECT 83.980 87.700 84.630 88.350 ;
        RECT 84.830 87.700 85.480 88.350 ;
        RECT 83.980 86.900 84.630 87.550 ;
        RECT 84.830 86.900 85.480 87.550 ;
        RECT 103.980 92.450 104.630 93.100 ;
        RECT 104.830 92.450 105.480 93.100 ;
        RECT 103.980 91.650 104.630 92.300 ;
        RECT 104.830 91.650 105.480 92.300 ;
        RECT 103.980 90.850 104.630 91.500 ;
        RECT 104.830 90.850 105.480 91.500 ;
        RECT 103.980 88.500 104.630 89.150 ;
        RECT 104.830 88.500 105.480 89.150 ;
        RECT 103.980 87.700 104.630 88.350 ;
        RECT 104.830 87.700 105.480 88.350 ;
        RECT 103.980 86.900 104.630 87.550 ;
        RECT 104.830 86.900 105.480 87.550 ;
        RECT 123.980 92.450 124.630 93.100 ;
        RECT 123.980 91.650 124.630 92.300 ;
        RECT 123.980 90.850 124.630 91.500 ;
        RECT 123.980 88.500 124.630 89.150 ;
        RECT 123.980 87.700 124.630 88.350 ;
        RECT 123.980 86.900 124.630 87.550 ;
        RECT 11.630 80.100 12.280 80.750 ;
        RECT 12.430 80.100 13.080 80.750 ;
        RECT 13.230 80.100 13.880 80.750 ;
        RECT 15.580 80.100 16.230 80.750 ;
        RECT 16.380 80.100 17.030 80.750 ;
        RECT 17.180 80.100 17.830 80.750 ;
        RECT 11.630 79.250 12.280 79.900 ;
        RECT 12.430 79.250 13.080 79.900 ;
        RECT 13.230 79.250 13.880 79.900 ;
        RECT 15.580 79.250 16.230 79.900 ;
        RECT 16.380 79.250 17.030 79.900 ;
        RECT 17.180 79.250 17.830 79.900 ;
        RECT 31.630 80.100 32.280 80.750 ;
        RECT 32.430 80.100 33.080 80.750 ;
        RECT 33.230 80.100 33.880 80.750 ;
        RECT 35.580 80.100 36.230 80.750 ;
        RECT 36.380 80.100 37.030 80.750 ;
        RECT 37.180 80.100 37.830 80.750 ;
        RECT 31.630 79.250 32.280 79.900 ;
        RECT 32.430 79.250 33.080 79.900 ;
        RECT 33.230 79.250 33.880 79.900 ;
        RECT 35.580 79.250 36.230 79.900 ;
        RECT 36.380 79.250 37.030 79.900 ;
        RECT 37.180 79.250 37.830 79.900 ;
        RECT 51.630 80.100 52.280 80.750 ;
        RECT 52.430 80.100 53.080 80.750 ;
        RECT 53.230 80.100 53.880 80.750 ;
        RECT 55.580 80.100 56.230 80.750 ;
        RECT 56.380 80.100 57.030 80.750 ;
        RECT 57.180 80.100 57.830 80.750 ;
        RECT 51.630 79.250 52.280 79.900 ;
        RECT 52.430 79.250 53.080 79.900 ;
        RECT 53.230 79.250 53.880 79.900 ;
        RECT 55.580 79.250 56.230 79.900 ;
        RECT 56.380 79.250 57.030 79.900 ;
        RECT 57.180 79.250 57.830 79.900 ;
        RECT 71.630 80.100 72.280 80.750 ;
        RECT 72.430 80.100 73.080 80.750 ;
        RECT 73.230 80.100 73.880 80.750 ;
        RECT 75.580 80.100 76.230 80.750 ;
        RECT 76.380 80.100 77.030 80.750 ;
        RECT 77.180 80.100 77.830 80.750 ;
        RECT 71.630 79.250 72.280 79.900 ;
        RECT 72.430 79.250 73.080 79.900 ;
        RECT 73.230 79.250 73.880 79.900 ;
        RECT 75.580 79.250 76.230 79.900 ;
        RECT 76.380 79.250 77.030 79.900 ;
        RECT 77.180 79.250 77.830 79.900 ;
        RECT 91.630 80.100 92.280 80.750 ;
        RECT 92.430 80.100 93.080 80.750 ;
        RECT 93.230 80.100 93.880 80.750 ;
        RECT 95.580 80.100 96.230 80.750 ;
        RECT 96.380 80.100 97.030 80.750 ;
        RECT 97.180 80.100 97.830 80.750 ;
        RECT 91.630 79.250 92.280 79.900 ;
        RECT 92.430 79.250 93.080 79.900 ;
        RECT 93.230 79.250 93.880 79.900 ;
        RECT 95.580 79.250 96.230 79.900 ;
        RECT 96.380 79.250 97.030 79.900 ;
        RECT 97.180 79.250 97.830 79.900 ;
        RECT 111.630 80.100 112.280 80.750 ;
        RECT 112.430 80.100 113.080 80.750 ;
        RECT 113.230 80.100 113.880 80.750 ;
        RECT 115.580 80.100 116.230 80.750 ;
        RECT 116.380 80.100 117.030 80.750 ;
        RECT 117.180 80.100 117.830 80.750 ;
        RECT 111.630 79.250 112.280 79.900 ;
        RECT 112.430 79.250 113.080 79.900 ;
        RECT 113.230 79.250 113.880 79.900 ;
        RECT 115.580 79.250 116.230 79.900 ;
        RECT 116.380 79.250 117.030 79.900 ;
        RECT 117.180 79.250 117.830 79.900 ;
        RECT 4.830 72.450 5.480 73.100 ;
        RECT 4.830 71.650 5.480 72.300 ;
        RECT 4.830 70.850 5.480 71.500 ;
        RECT 4.830 68.500 5.480 69.150 ;
        RECT 4.830 67.700 5.480 68.350 ;
        RECT 4.830 66.900 5.480 67.550 ;
        RECT 23.980 72.450 24.630 73.100 ;
        RECT 24.830 72.450 25.480 73.100 ;
        RECT 23.980 71.650 24.630 72.300 ;
        RECT 24.830 71.650 25.480 72.300 ;
        RECT 23.980 70.850 24.630 71.500 ;
        RECT 24.830 70.850 25.480 71.500 ;
        RECT 23.980 68.500 24.630 69.150 ;
        RECT 24.830 68.500 25.480 69.150 ;
        RECT 23.980 67.700 24.630 68.350 ;
        RECT 24.830 67.700 25.480 68.350 ;
        RECT 23.980 66.900 24.630 67.550 ;
        RECT 24.830 66.900 25.480 67.550 ;
        RECT 43.980 72.450 44.630 73.100 ;
        RECT 44.830 72.450 45.480 73.100 ;
        RECT 43.980 71.650 44.630 72.300 ;
        RECT 44.830 71.650 45.480 72.300 ;
        RECT 43.980 70.850 44.630 71.500 ;
        RECT 44.830 70.850 45.480 71.500 ;
        RECT 43.980 68.500 44.630 69.150 ;
        RECT 44.830 68.500 45.480 69.150 ;
        RECT 43.980 67.700 44.630 68.350 ;
        RECT 44.830 67.700 45.480 68.350 ;
        RECT 43.980 66.900 44.630 67.550 ;
        RECT 44.830 66.900 45.480 67.550 ;
        RECT 63.980 72.450 64.630 73.100 ;
        RECT 64.830 72.450 65.480 73.100 ;
        RECT 63.980 71.650 64.630 72.300 ;
        RECT 64.830 71.650 65.480 72.300 ;
        RECT 63.980 70.850 64.630 71.500 ;
        RECT 64.830 70.850 65.480 71.500 ;
        RECT 63.980 68.500 64.630 69.150 ;
        RECT 64.830 68.500 65.480 69.150 ;
        RECT 63.980 67.700 64.630 68.350 ;
        RECT 64.830 67.700 65.480 68.350 ;
        RECT 63.980 66.900 64.630 67.550 ;
        RECT 64.830 66.900 65.480 67.550 ;
        RECT 83.980 72.450 84.630 73.100 ;
        RECT 84.830 72.450 85.480 73.100 ;
        RECT 83.980 71.650 84.630 72.300 ;
        RECT 84.830 71.650 85.480 72.300 ;
        RECT 83.980 70.850 84.630 71.500 ;
        RECT 84.830 70.850 85.480 71.500 ;
        RECT 83.980 68.500 84.630 69.150 ;
        RECT 84.830 68.500 85.480 69.150 ;
        RECT 83.980 67.700 84.630 68.350 ;
        RECT 84.830 67.700 85.480 68.350 ;
        RECT 83.980 66.900 84.630 67.550 ;
        RECT 84.830 66.900 85.480 67.550 ;
        RECT 103.980 72.450 104.630 73.100 ;
        RECT 104.830 72.450 105.480 73.100 ;
        RECT 103.980 71.650 104.630 72.300 ;
        RECT 104.830 71.650 105.480 72.300 ;
        RECT 103.980 70.850 104.630 71.500 ;
        RECT 104.830 70.850 105.480 71.500 ;
        RECT 103.980 68.500 104.630 69.150 ;
        RECT 104.830 68.500 105.480 69.150 ;
        RECT 103.980 67.700 104.630 68.350 ;
        RECT 104.830 67.700 105.480 68.350 ;
        RECT 103.980 66.900 104.630 67.550 ;
        RECT 104.830 66.900 105.480 67.550 ;
        RECT 123.980 72.450 124.630 73.100 ;
        RECT 123.980 71.650 124.630 72.300 ;
        RECT 123.980 70.850 124.630 71.500 ;
        RECT 123.980 68.500 124.630 69.150 ;
        RECT 123.980 67.700 124.630 68.350 ;
        RECT 123.980 66.900 124.630 67.550 ;
        RECT 11.630 60.100 12.280 60.750 ;
        RECT 12.430 60.100 13.080 60.750 ;
        RECT 13.230 60.100 13.880 60.750 ;
        RECT 15.580 60.100 16.230 60.750 ;
        RECT 16.380 60.100 17.030 60.750 ;
        RECT 17.180 60.100 17.830 60.750 ;
        RECT 11.630 59.250 12.280 59.900 ;
        RECT 12.430 59.250 13.080 59.900 ;
        RECT 13.230 59.250 13.880 59.900 ;
        RECT 15.580 59.250 16.230 59.900 ;
        RECT 16.380 59.250 17.030 59.900 ;
        RECT 17.180 59.250 17.830 59.900 ;
        RECT 31.630 60.100 32.280 60.750 ;
        RECT 32.430 60.100 33.080 60.750 ;
        RECT 33.230 60.100 33.880 60.750 ;
        RECT 35.580 60.100 36.230 60.750 ;
        RECT 36.380 60.100 37.030 60.750 ;
        RECT 37.180 60.100 37.830 60.750 ;
        RECT 31.630 59.250 32.280 59.900 ;
        RECT 32.430 59.250 33.080 59.900 ;
        RECT 33.230 59.250 33.880 59.900 ;
        RECT 35.580 59.250 36.230 59.900 ;
        RECT 36.380 59.250 37.030 59.900 ;
        RECT 37.180 59.250 37.830 59.900 ;
        RECT 51.630 60.100 52.280 60.750 ;
        RECT 52.430 60.100 53.080 60.750 ;
        RECT 53.230 60.100 53.880 60.750 ;
        RECT 55.580 60.100 56.230 60.750 ;
        RECT 56.380 60.100 57.030 60.750 ;
        RECT 57.180 60.100 57.830 60.750 ;
        RECT 51.630 59.250 52.280 59.900 ;
        RECT 52.430 59.250 53.080 59.900 ;
        RECT 53.230 59.250 53.880 59.900 ;
        RECT 55.580 59.250 56.230 59.900 ;
        RECT 56.380 59.250 57.030 59.900 ;
        RECT 57.180 59.250 57.830 59.900 ;
        RECT 71.630 60.100 72.280 60.750 ;
        RECT 72.430 60.100 73.080 60.750 ;
        RECT 73.230 60.100 73.880 60.750 ;
        RECT 75.580 60.100 76.230 60.750 ;
        RECT 76.380 60.100 77.030 60.750 ;
        RECT 77.180 60.100 77.830 60.750 ;
        RECT 71.630 59.250 72.280 59.900 ;
        RECT 72.430 59.250 73.080 59.900 ;
        RECT 73.230 59.250 73.880 59.900 ;
        RECT 75.580 59.250 76.230 59.900 ;
        RECT 76.380 59.250 77.030 59.900 ;
        RECT 77.180 59.250 77.830 59.900 ;
        RECT 91.630 60.100 92.280 60.750 ;
        RECT 92.430 60.100 93.080 60.750 ;
        RECT 93.230 60.100 93.880 60.750 ;
        RECT 95.580 60.100 96.230 60.750 ;
        RECT 96.380 60.100 97.030 60.750 ;
        RECT 97.180 60.100 97.830 60.750 ;
        RECT 91.630 59.250 92.280 59.900 ;
        RECT 92.430 59.250 93.080 59.900 ;
        RECT 93.230 59.250 93.880 59.900 ;
        RECT 95.580 59.250 96.230 59.900 ;
        RECT 96.380 59.250 97.030 59.900 ;
        RECT 97.180 59.250 97.830 59.900 ;
        RECT 111.630 60.100 112.280 60.750 ;
        RECT 112.430 60.100 113.080 60.750 ;
        RECT 113.230 60.100 113.880 60.750 ;
        RECT 115.580 60.100 116.230 60.750 ;
        RECT 116.380 60.100 117.030 60.750 ;
        RECT 117.180 60.100 117.830 60.750 ;
        RECT 111.630 59.250 112.280 59.900 ;
        RECT 112.430 59.250 113.080 59.900 ;
        RECT 113.230 59.250 113.880 59.900 ;
        RECT 115.580 59.250 116.230 59.900 ;
        RECT 116.380 59.250 117.030 59.900 ;
        RECT 117.180 59.250 117.830 59.900 ;
        RECT 4.830 52.450 5.480 53.100 ;
        RECT 4.830 51.650 5.480 52.300 ;
        RECT 4.830 50.850 5.480 51.500 ;
        RECT 4.830 48.500 5.480 49.150 ;
        RECT 4.830 47.700 5.480 48.350 ;
        RECT 4.830 46.900 5.480 47.550 ;
        RECT 23.980 52.450 24.630 53.100 ;
        RECT 24.830 52.450 25.480 53.100 ;
        RECT 23.980 51.650 24.630 52.300 ;
        RECT 24.830 51.650 25.480 52.300 ;
        RECT 23.980 50.850 24.630 51.500 ;
        RECT 24.830 50.850 25.480 51.500 ;
        RECT 23.980 48.500 24.630 49.150 ;
        RECT 24.830 48.500 25.480 49.150 ;
        RECT 23.980 47.700 24.630 48.350 ;
        RECT 24.830 47.700 25.480 48.350 ;
        RECT 23.980 46.900 24.630 47.550 ;
        RECT 24.830 46.900 25.480 47.550 ;
        RECT 43.980 52.450 44.630 53.100 ;
        RECT 44.830 52.450 45.480 53.100 ;
        RECT 43.980 51.650 44.630 52.300 ;
        RECT 44.830 51.650 45.480 52.300 ;
        RECT 43.980 50.850 44.630 51.500 ;
        RECT 44.830 50.850 45.480 51.500 ;
        RECT 43.980 48.500 44.630 49.150 ;
        RECT 44.830 48.500 45.480 49.150 ;
        RECT 43.980 47.700 44.630 48.350 ;
        RECT 44.830 47.700 45.480 48.350 ;
        RECT 43.980 46.900 44.630 47.550 ;
        RECT 44.830 46.900 45.480 47.550 ;
        RECT 63.980 52.450 64.630 53.100 ;
        RECT 64.830 52.450 65.480 53.100 ;
        RECT 63.980 51.650 64.630 52.300 ;
        RECT 64.830 51.650 65.480 52.300 ;
        RECT 63.980 50.850 64.630 51.500 ;
        RECT 64.830 50.850 65.480 51.500 ;
        RECT 63.980 48.500 64.630 49.150 ;
        RECT 64.830 48.500 65.480 49.150 ;
        RECT 63.980 47.700 64.630 48.350 ;
        RECT 64.830 47.700 65.480 48.350 ;
        RECT 63.980 46.900 64.630 47.550 ;
        RECT 64.830 46.900 65.480 47.550 ;
        RECT 83.980 52.450 84.630 53.100 ;
        RECT 84.830 52.450 85.480 53.100 ;
        RECT 83.980 51.650 84.630 52.300 ;
        RECT 84.830 51.650 85.480 52.300 ;
        RECT 83.980 50.850 84.630 51.500 ;
        RECT 84.830 50.850 85.480 51.500 ;
        RECT 83.980 48.500 84.630 49.150 ;
        RECT 84.830 48.500 85.480 49.150 ;
        RECT 83.980 47.700 84.630 48.350 ;
        RECT 84.830 47.700 85.480 48.350 ;
        RECT 83.980 46.900 84.630 47.550 ;
        RECT 84.830 46.900 85.480 47.550 ;
        RECT 103.980 52.450 104.630 53.100 ;
        RECT 104.830 52.450 105.480 53.100 ;
        RECT 103.980 51.650 104.630 52.300 ;
        RECT 104.830 51.650 105.480 52.300 ;
        RECT 103.980 50.850 104.630 51.500 ;
        RECT 104.830 50.850 105.480 51.500 ;
        RECT 103.980 48.500 104.630 49.150 ;
        RECT 104.830 48.500 105.480 49.150 ;
        RECT 103.980 47.700 104.630 48.350 ;
        RECT 104.830 47.700 105.480 48.350 ;
        RECT 103.980 46.900 104.630 47.550 ;
        RECT 104.830 46.900 105.480 47.550 ;
        RECT 123.980 52.450 124.630 53.100 ;
        RECT 123.980 51.650 124.630 52.300 ;
        RECT 123.980 50.850 124.630 51.500 ;
        RECT 123.980 48.500 124.630 49.150 ;
        RECT 123.980 47.700 124.630 48.350 ;
        RECT 123.980 46.900 124.630 47.550 ;
        RECT 11.630 40.100 12.280 40.750 ;
        RECT 12.430 40.100 13.080 40.750 ;
        RECT 13.230 40.100 13.880 40.750 ;
        RECT 15.580 40.100 16.230 40.750 ;
        RECT 16.380 40.100 17.030 40.750 ;
        RECT 17.180 40.100 17.830 40.750 ;
        RECT 11.630 39.250 12.280 39.900 ;
        RECT 12.430 39.250 13.080 39.900 ;
        RECT 13.230 39.250 13.880 39.900 ;
        RECT 15.580 39.250 16.230 39.900 ;
        RECT 16.380 39.250 17.030 39.900 ;
        RECT 17.180 39.250 17.830 39.900 ;
        RECT 31.630 40.100 32.280 40.750 ;
        RECT 32.430 40.100 33.080 40.750 ;
        RECT 33.230 40.100 33.880 40.750 ;
        RECT 35.580 40.100 36.230 40.750 ;
        RECT 36.380 40.100 37.030 40.750 ;
        RECT 37.180 40.100 37.830 40.750 ;
        RECT 31.630 39.250 32.280 39.900 ;
        RECT 32.430 39.250 33.080 39.900 ;
        RECT 33.230 39.250 33.880 39.900 ;
        RECT 35.580 39.250 36.230 39.900 ;
        RECT 36.380 39.250 37.030 39.900 ;
        RECT 37.180 39.250 37.830 39.900 ;
        RECT 51.630 40.100 52.280 40.750 ;
        RECT 52.430 40.100 53.080 40.750 ;
        RECT 53.230 40.100 53.880 40.750 ;
        RECT 55.580 40.100 56.230 40.750 ;
        RECT 56.380 40.100 57.030 40.750 ;
        RECT 57.180 40.100 57.830 40.750 ;
        RECT 51.630 39.250 52.280 39.900 ;
        RECT 52.430 39.250 53.080 39.900 ;
        RECT 53.230 39.250 53.880 39.900 ;
        RECT 55.580 39.250 56.230 39.900 ;
        RECT 56.380 39.250 57.030 39.900 ;
        RECT 57.180 39.250 57.830 39.900 ;
        RECT 71.630 40.100 72.280 40.750 ;
        RECT 72.430 40.100 73.080 40.750 ;
        RECT 73.230 40.100 73.880 40.750 ;
        RECT 75.580 40.100 76.230 40.750 ;
        RECT 76.380 40.100 77.030 40.750 ;
        RECT 77.180 40.100 77.830 40.750 ;
        RECT 71.630 39.250 72.280 39.900 ;
        RECT 72.430 39.250 73.080 39.900 ;
        RECT 73.230 39.250 73.880 39.900 ;
        RECT 75.580 39.250 76.230 39.900 ;
        RECT 76.380 39.250 77.030 39.900 ;
        RECT 77.180 39.250 77.830 39.900 ;
        RECT 91.630 40.100 92.280 40.750 ;
        RECT 92.430 40.100 93.080 40.750 ;
        RECT 93.230 40.100 93.880 40.750 ;
        RECT 95.580 40.100 96.230 40.750 ;
        RECT 96.380 40.100 97.030 40.750 ;
        RECT 97.180 40.100 97.830 40.750 ;
        RECT 91.630 39.250 92.280 39.900 ;
        RECT 92.430 39.250 93.080 39.900 ;
        RECT 93.230 39.250 93.880 39.900 ;
        RECT 95.580 39.250 96.230 39.900 ;
        RECT 96.380 39.250 97.030 39.900 ;
        RECT 97.180 39.250 97.830 39.900 ;
        RECT 111.630 40.100 112.280 40.750 ;
        RECT 112.430 40.100 113.080 40.750 ;
        RECT 113.230 40.100 113.880 40.750 ;
        RECT 115.580 40.100 116.230 40.750 ;
        RECT 116.380 40.100 117.030 40.750 ;
        RECT 117.180 40.100 117.830 40.750 ;
        RECT 111.630 39.250 112.280 39.900 ;
        RECT 112.430 39.250 113.080 39.900 ;
        RECT 113.230 39.250 113.880 39.900 ;
        RECT 115.580 39.250 116.230 39.900 ;
        RECT 116.380 39.250 117.030 39.900 ;
        RECT 117.180 39.250 117.830 39.900 ;
        RECT 4.830 32.450 5.480 33.100 ;
        RECT 4.830 31.650 5.480 32.300 ;
        RECT 4.830 30.850 5.480 31.500 ;
        RECT 4.830 28.500 5.480 29.150 ;
        RECT 4.830 27.700 5.480 28.350 ;
        RECT 4.830 26.900 5.480 27.550 ;
        RECT 23.980 32.450 24.630 33.100 ;
        RECT 24.830 32.450 25.480 33.100 ;
        RECT 23.980 31.650 24.630 32.300 ;
        RECT 24.830 31.650 25.480 32.300 ;
        RECT 23.980 30.850 24.630 31.500 ;
        RECT 24.830 30.850 25.480 31.500 ;
        RECT 23.980 28.500 24.630 29.150 ;
        RECT 24.830 28.500 25.480 29.150 ;
        RECT 23.980 27.700 24.630 28.350 ;
        RECT 24.830 27.700 25.480 28.350 ;
        RECT 23.980 26.900 24.630 27.550 ;
        RECT 24.830 26.900 25.480 27.550 ;
        RECT 43.980 32.450 44.630 33.100 ;
        RECT 44.830 32.450 45.480 33.100 ;
        RECT 43.980 31.650 44.630 32.300 ;
        RECT 44.830 31.650 45.480 32.300 ;
        RECT 43.980 30.850 44.630 31.500 ;
        RECT 44.830 30.850 45.480 31.500 ;
        RECT 43.980 28.500 44.630 29.150 ;
        RECT 44.830 28.500 45.480 29.150 ;
        RECT 43.980 27.700 44.630 28.350 ;
        RECT 44.830 27.700 45.480 28.350 ;
        RECT 43.980 26.900 44.630 27.550 ;
        RECT 44.830 26.900 45.480 27.550 ;
        RECT 63.980 32.450 64.630 33.100 ;
        RECT 64.830 32.450 65.480 33.100 ;
        RECT 63.980 31.650 64.630 32.300 ;
        RECT 64.830 31.650 65.480 32.300 ;
        RECT 63.980 30.850 64.630 31.500 ;
        RECT 64.830 30.850 65.480 31.500 ;
        RECT 63.980 28.500 64.630 29.150 ;
        RECT 64.830 28.500 65.480 29.150 ;
        RECT 63.980 27.700 64.630 28.350 ;
        RECT 64.830 27.700 65.480 28.350 ;
        RECT 63.980 26.900 64.630 27.550 ;
        RECT 64.830 26.900 65.480 27.550 ;
        RECT 83.980 32.450 84.630 33.100 ;
        RECT 84.830 32.450 85.480 33.100 ;
        RECT 83.980 31.650 84.630 32.300 ;
        RECT 84.830 31.650 85.480 32.300 ;
        RECT 83.980 30.850 84.630 31.500 ;
        RECT 84.830 30.850 85.480 31.500 ;
        RECT 83.980 28.500 84.630 29.150 ;
        RECT 84.830 28.500 85.480 29.150 ;
        RECT 83.980 27.700 84.630 28.350 ;
        RECT 84.830 27.700 85.480 28.350 ;
        RECT 83.980 26.900 84.630 27.550 ;
        RECT 84.830 26.900 85.480 27.550 ;
        RECT 103.980 32.450 104.630 33.100 ;
        RECT 104.830 32.450 105.480 33.100 ;
        RECT 103.980 31.650 104.630 32.300 ;
        RECT 104.830 31.650 105.480 32.300 ;
        RECT 103.980 30.850 104.630 31.500 ;
        RECT 104.830 30.850 105.480 31.500 ;
        RECT 103.980 28.500 104.630 29.150 ;
        RECT 104.830 28.500 105.480 29.150 ;
        RECT 103.980 27.700 104.630 28.350 ;
        RECT 104.830 27.700 105.480 28.350 ;
        RECT 103.980 26.900 104.630 27.550 ;
        RECT 104.830 26.900 105.480 27.550 ;
        RECT 123.980 32.450 124.630 33.100 ;
        RECT 123.980 31.650 124.630 32.300 ;
        RECT 123.980 30.850 124.630 31.500 ;
        RECT 123.980 28.500 124.630 29.150 ;
        RECT 123.980 27.700 124.630 28.350 ;
        RECT 123.980 26.900 124.630 27.550 ;
        RECT 11.630 20.100 12.280 20.750 ;
        RECT 12.430 20.100 13.080 20.750 ;
        RECT 13.230 20.100 13.880 20.750 ;
        RECT 15.580 20.100 16.230 20.750 ;
        RECT 16.380 20.100 17.030 20.750 ;
        RECT 17.180 20.100 17.830 20.750 ;
        RECT 11.630 19.250 12.280 19.900 ;
        RECT 12.430 19.250 13.080 19.900 ;
        RECT 13.230 19.250 13.880 19.900 ;
        RECT 15.580 19.250 16.230 19.900 ;
        RECT 16.380 19.250 17.030 19.900 ;
        RECT 17.180 19.250 17.830 19.900 ;
        RECT 31.630 20.100 32.280 20.750 ;
        RECT 32.430 20.100 33.080 20.750 ;
        RECT 33.230 20.100 33.880 20.750 ;
        RECT 35.580 20.100 36.230 20.750 ;
        RECT 36.380 20.100 37.030 20.750 ;
        RECT 37.180 20.100 37.830 20.750 ;
        RECT 31.630 19.250 32.280 19.900 ;
        RECT 32.430 19.250 33.080 19.900 ;
        RECT 33.230 19.250 33.880 19.900 ;
        RECT 35.580 19.250 36.230 19.900 ;
        RECT 36.380 19.250 37.030 19.900 ;
        RECT 37.180 19.250 37.830 19.900 ;
        RECT 51.630 20.100 52.280 20.750 ;
        RECT 52.430 20.100 53.080 20.750 ;
        RECT 53.230 20.100 53.880 20.750 ;
        RECT 55.580 20.100 56.230 20.750 ;
        RECT 56.380 20.100 57.030 20.750 ;
        RECT 57.180 20.100 57.830 20.750 ;
        RECT 51.630 19.250 52.280 19.900 ;
        RECT 52.430 19.250 53.080 19.900 ;
        RECT 53.230 19.250 53.880 19.900 ;
        RECT 55.580 19.250 56.230 19.900 ;
        RECT 56.380 19.250 57.030 19.900 ;
        RECT 57.180 19.250 57.830 19.900 ;
        RECT 71.630 20.100 72.280 20.750 ;
        RECT 72.430 20.100 73.080 20.750 ;
        RECT 73.230 20.100 73.880 20.750 ;
        RECT 75.580 20.100 76.230 20.750 ;
        RECT 76.380 20.100 77.030 20.750 ;
        RECT 77.180 20.100 77.830 20.750 ;
        RECT 71.630 19.250 72.280 19.900 ;
        RECT 72.430 19.250 73.080 19.900 ;
        RECT 73.230 19.250 73.880 19.900 ;
        RECT 75.580 19.250 76.230 19.900 ;
        RECT 76.380 19.250 77.030 19.900 ;
        RECT 77.180 19.250 77.830 19.900 ;
        RECT 91.630 20.100 92.280 20.750 ;
        RECT 92.430 20.100 93.080 20.750 ;
        RECT 93.230 20.100 93.880 20.750 ;
        RECT 95.580 20.100 96.230 20.750 ;
        RECT 96.380 20.100 97.030 20.750 ;
        RECT 97.180 20.100 97.830 20.750 ;
        RECT 91.630 19.250 92.280 19.900 ;
        RECT 92.430 19.250 93.080 19.900 ;
        RECT 93.230 19.250 93.880 19.900 ;
        RECT 95.580 19.250 96.230 19.900 ;
        RECT 96.380 19.250 97.030 19.900 ;
        RECT 97.180 19.250 97.830 19.900 ;
        RECT 111.630 20.100 112.280 20.750 ;
        RECT 112.430 20.100 113.080 20.750 ;
        RECT 113.230 20.100 113.880 20.750 ;
        RECT 115.580 20.100 116.230 20.750 ;
        RECT 116.380 20.100 117.030 20.750 ;
        RECT 117.180 20.100 117.830 20.750 ;
        RECT 111.630 19.250 112.280 19.900 ;
        RECT 112.430 19.250 113.080 19.900 ;
        RECT 113.230 19.250 113.880 19.900 ;
        RECT 115.580 19.250 116.230 19.900 ;
        RECT 116.380 19.250 117.030 19.900 ;
        RECT 117.180 19.250 117.830 19.900 ;
        RECT 4.830 12.450 5.480 13.100 ;
        RECT 4.830 11.650 5.480 12.300 ;
        RECT 4.830 10.850 5.480 11.500 ;
        RECT 4.830 8.500 5.480 9.150 ;
        RECT 4.830 7.700 5.480 8.350 ;
        RECT 4.830 6.900 5.480 7.550 ;
        RECT 23.980 12.450 24.630 13.100 ;
        RECT 24.830 12.450 25.480 13.100 ;
        RECT 23.980 11.650 24.630 12.300 ;
        RECT 24.830 11.650 25.480 12.300 ;
        RECT 23.980 10.850 24.630 11.500 ;
        RECT 24.830 10.850 25.480 11.500 ;
        RECT 23.980 8.500 24.630 9.150 ;
        RECT 24.830 8.500 25.480 9.150 ;
        RECT 23.980 7.700 24.630 8.350 ;
        RECT 24.830 7.700 25.480 8.350 ;
        RECT 23.980 6.900 24.630 7.550 ;
        RECT 24.830 6.900 25.480 7.550 ;
        RECT 43.980 12.450 44.630 13.100 ;
        RECT 44.830 12.450 45.480 13.100 ;
        RECT 43.980 11.650 44.630 12.300 ;
        RECT 44.830 11.650 45.480 12.300 ;
        RECT 43.980 10.850 44.630 11.500 ;
        RECT 44.830 10.850 45.480 11.500 ;
        RECT 43.980 8.500 44.630 9.150 ;
        RECT 44.830 8.500 45.480 9.150 ;
        RECT 43.980 7.700 44.630 8.350 ;
        RECT 44.830 7.700 45.480 8.350 ;
        RECT 43.980 6.900 44.630 7.550 ;
        RECT 44.830 6.900 45.480 7.550 ;
        RECT 63.980 12.450 64.630 13.100 ;
        RECT 64.830 12.450 65.480 13.100 ;
        RECT 63.980 11.650 64.630 12.300 ;
        RECT 64.830 11.650 65.480 12.300 ;
        RECT 63.980 10.850 64.630 11.500 ;
        RECT 64.830 10.850 65.480 11.500 ;
        RECT 63.980 8.500 64.630 9.150 ;
        RECT 64.830 8.500 65.480 9.150 ;
        RECT 63.980 7.700 64.630 8.350 ;
        RECT 64.830 7.700 65.480 8.350 ;
        RECT 63.980 6.900 64.630 7.550 ;
        RECT 64.830 6.900 65.480 7.550 ;
        RECT 83.980 12.450 84.630 13.100 ;
        RECT 84.830 12.450 85.480 13.100 ;
        RECT 83.980 11.650 84.630 12.300 ;
        RECT 84.830 11.650 85.480 12.300 ;
        RECT 83.980 10.850 84.630 11.500 ;
        RECT 84.830 10.850 85.480 11.500 ;
        RECT 83.980 8.500 84.630 9.150 ;
        RECT 84.830 8.500 85.480 9.150 ;
        RECT 83.980 7.700 84.630 8.350 ;
        RECT 84.830 7.700 85.480 8.350 ;
        RECT 83.980 6.900 84.630 7.550 ;
        RECT 84.830 6.900 85.480 7.550 ;
        RECT 103.980 12.450 104.630 13.100 ;
        RECT 104.830 12.450 105.480 13.100 ;
        RECT 103.980 11.650 104.630 12.300 ;
        RECT 104.830 11.650 105.480 12.300 ;
        RECT 103.980 10.850 104.630 11.500 ;
        RECT 104.830 10.850 105.480 11.500 ;
        RECT 103.980 8.500 104.630 9.150 ;
        RECT 104.830 8.500 105.480 9.150 ;
        RECT 103.980 7.700 104.630 8.350 ;
        RECT 104.830 7.700 105.480 8.350 ;
        RECT 103.980 6.900 104.630 7.550 ;
        RECT 104.830 6.900 105.480 7.550 ;
        RECT 123.980 12.450 124.630 13.100 ;
        RECT 123.980 11.650 124.630 12.300 ;
        RECT 123.980 10.850 124.630 11.500 ;
        RECT 123.980 8.500 124.630 9.150 ;
        RECT 123.980 7.700 124.630 8.350 ;
        RECT 123.980 6.900 124.630 7.550 ;
        RECT 11.630 0.100 12.280 0.750 ;
        RECT 12.430 0.100 13.080 0.750 ;
        RECT 13.230 0.100 13.880 0.750 ;
        RECT 15.580 0.100 16.230 0.750 ;
        RECT 16.380 0.100 17.030 0.750 ;
        RECT 17.180 0.100 17.830 0.750 ;
        RECT 31.630 0.100 32.280 0.750 ;
        RECT 32.430 0.100 33.080 0.750 ;
        RECT 33.230 0.100 33.880 0.750 ;
        RECT 35.580 0.100 36.230 0.750 ;
        RECT 36.380 0.100 37.030 0.750 ;
        RECT 37.180 0.100 37.830 0.750 ;
        RECT 51.630 0.100 52.280 0.750 ;
        RECT 52.430 0.100 53.080 0.750 ;
        RECT 53.230 0.100 53.880 0.750 ;
        RECT 55.580 0.100 56.230 0.750 ;
        RECT 56.380 0.100 57.030 0.750 ;
        RECT 57.180 0.100 57.830 0.750 ;
        RECT 71.630 0.100 72.280 0.750 ;
        RECT 72.430 0.100 73.080 0.750 ;
        RECT 73.230 0.100 73.880 0.750 ;
        RECT 75.580 0.100 76.230 0.750 ;
        RECT 76.380 0.100 77.030 0.750 ;
        RECT 77.180 0.100 77.830 0.750 ;
        RECT 91.630 0.100 92.280 0.750 ;
        RECT 92.430 0.100 93.080 0.750 ;
        RECT 93.230 0.100 93.880 0.750 ;
        RECT 95.580 0.100 96.230 0.750 ;
        RECT 96.380 0.100 97.030 0.750 ;
        RECT 97.180 0.100 97.830 0.750 ;
        RECT 111.630 0.100 112.280 0.750 ;
        RECT 112.430 0.100 113.080 0.750 ;
        RECT 113.230 0.100 113.880 0.750 ;
        RECT 115.580 0.100 116.230 0.750 ;
        RECT 116.380 0.100 117.030 0.750 ;
        RECT 117.180 0.100 117.830 0.750 ;
      LAYER met4 ;
        RECT 4.730 338.950 9.130 340.000 ;
        RECT 4.730 335.600 5.780 338.950 ;
        RECT 11.530 338.550 17.930 340.000 ;
        RECT 20.330 338.950 29.130 340.000 ;
        RECT 6.180 333.200 23.280 338.550 ;
        RECT 23.680 335.600 25.780 338.950 ;
        RECT 31.530 338.550 37.930 340.000 ;
        RECT 40.330 338.950 49.130 340.000 ;
        RECT 26.180 333.200 43.280 338.550 ;
        RECT 43.680 335.600 45.780 338.950 ;
        RECT 51.530 338.550 57.930 340.000 ;
        RECT 60.330 338.950 69.130 340.000 ;
        RECT 46.180 333.200 63.280 338.550 ;
        RECT 63.680 335.600 65.780 338.950 ;
        RECT 71.530 338.550 77.930 340.000 ;
        RECT 80.330 338.950 89.130 340.000 ;
        RECT 66.180 333.200 83.280 338.550 ;
        RECT 83.680 335.600 85.780 338.950 ;
        RECT 91.530 338.550 97.930 340.000 ;
        RECT 100.330 338.950 109.130 340.000 ;
        RECT 86.180 333.200 103.280 338.550 ;
        RECT 103.680 335.600 105.780 338.950 ;
        RECT 111.530 338.550 117.930 340.000 ;
        RECT 120.330 338.950 124.730 340.000 ;
        RECT 106.180 333.200 123.280 338.550 ;
        RECT 123.680 335.600 124.730 338.950 ;
        RECT 4.730 326.800 124.730 333.200 ;
        RECT 4.730 321.050 5.780 324.400 ;
        RECT 6.180 321.450 23.280 326.800 ;
        RECT 4.730 318.950 9.130 321.050 ;
        RECT 4.730 315.600 5.780 318.950 ;
        RECT 11.530 318.550 17.930 321.450 ;
        RECT 23.680 321.050 25.780 324.400 ;
        RECT 26.180 321.450 43.280 326.800 ;
        RECT 20.330 318.950 29.130 321.050 ;
        RECT 6.180 313.200 23.280 318.550 ;
        RECT 23.680 315.600 25.780 318.950 ;
        RECT 31.530 318.550 37.930 321.450 ;
        RECT 43.680 321.050 45.780 324.400 ;
        RECT 46.180 321.450 63.280 326.800 ;
        RECT 40.330 318.950 49.130 321.050 ;
        RECT 26.180 313.200 43.280 318.550 ;
        RECT 43.680 315.600 45.780 318.950 ;
        RECT 51.530 318.550 57.930 321.450 ;
        RECT 63.680 321.050 65.780 324.400 ;
        RECT 66.180 321.450 83.280 326.800 ;
        RECT 60.330 318.950 69.130 321.050 ;
        RECT 46.180 313.200 63.280 318.550 ;
        RECT 63.680 315.600 65.780 318.950 ;
        RECT 71.530 318.550 77.930 321.450 ;
        RECT 83.680 321.050 85.780 324.400 ;
        RECT 86.180 321.450 103.280 326.800 ;
        RECT 80.330 318.950 89.130 321.050 ;
        RECT 66.180 313.200 83.280 318.550 ;
        RECT 83.680 315.600 85.780 318.950 ;
        RECT 91.530 318.550 97.930 321.450 ;
        RECT 103.680 321.050 105.780 324.400 ;
        RECT 106.180 321.450 123.280 326.800 ;
        RECT 100.330 318.950 109.130 321.050 ;
        RECT 86.180 313.200 103.280 318.550 ;
        RECT 103.680 315.600 105.780 318.950 ;
        RECT 111.530 318.550 117.930 321.450 ;
        RECT 123.680 321.050 124.730 324.400 ;
        RECT 120.330 318.950 124.730 321.050 ;
        RECT 106.180 313.200 123.280 318.550 ;
        RECT 123.680 315.600 124.730 318.950 ;
        RECT 4.730 306.800 124.730 313.200 ;
        RECT 4.730 301.050 5.780 304.400 ;
        RECT 6.180 301.450 23.280 306.800 ;
        RECT 4.730 298.950 9.130 301.050 ;
        RECT 4.730 295.600 5.780 298.950 ;
        RECT 11.530 298.550 17.930 301.450 ;
        RECT 23.680 301.050 25.780 304.400 ;
        RECT 26.180 301.450 43.280 306.800 ;
        RECT 20.330 298.950 29.130 301.050 ;
        RECT 6.180 293.200 23.280 298.550 ;
        RECT 23.680 295.600 25.780 298.950 ;
        RECT 31.530 298.550 37.930 301.450 ;
        RECT 43.680 301.050 45.780 304.400 ;
        RECT 46.180 301.450 63.280 306.800 ;
        RECT 40.330 298.950 49.130 301.050 ;
        RECT 26.180 293.200 43.280 298.550 ;
        RECT 43.680 295.600 45.780 298.950 ;
        RECT 51.530 298.550 57.930 301.450 ;
        RECT 63.680 301.050 65.780 304.400 ;
        RECT 66.180 301.450 83.280 306.800 ;
        RECT 60.330 298.950 69.130 301.050 ;
        RECT 46.180 293.200 63.280 298.550 ;
        RECT 63.680 295.600 65.780 298.950 ;
        RECT 71.530 298.550 77.930 301.450 ;
        RECT 83.680 301.050 85.780 304.400 ;
        RECT 86.180 301.450 103.280 306.800 ;
        RECT 80.330 298.950 89.130 301.050 ;
        RECT 66.180 293.200 83.280 298.550 ;
        RECT 83.680 295.600 85.780 298.950 ;
        RECT 91.530 298.550 97.930 301.450 ;
        RECT 103.680 301.050 105.780 304.400 ;
        RECT 106.180 301.450 123.280 306.800 ;
        RECT 100.330 298.950 109.130 301.050 ;
        RECT 86.180 293.200 103.280 298.550 ;
        RECT 103.680 295.600 105.780 298.950 ;
        RECT 111.530 298.550 117.930 301.450 ;
        RECT 123.680 301.050 124.730 304.400 ;
        RECT 120.330 298.950 124.730 301.050 ;
        RECT 106.180 293.200 123.280 298.550 ;
        RECT 123.680 295.600 124.730 298.950 ;
        RECT 4.730 286.800 124.730 293.200 ;
        RECT 4.730 281.050 5.780 284.400 ;
        RECT 6.180 281.450 23.280 286.800 ;
        RECT 4.730 278.950 9.130 281.050 ;
        RECT 4.730 275.600 5.780 278.950 ;
        RECT 11.530 278.550 17.930 281.450 ;
        RECT 23.680 281.050 25.780 284.400 ;
        RECT 26.180 281.450 43.280 286.800 ;
        RECT 20.330 278.950 29.130 281.050 ;
        RECT 6.180 273.200 23.280 278.550 ;
        RECT 23.680 275.600 25.780 278.950 ;
        RECT 31.530 278.550 37.930 281.450 ;
        RECT 43.680 281.050 45.780 284.400 ;
        RECT 46.180 281.450 63.280 286.800 ;
        RECT 40.330 278.950 49.130 281.050 ;
        RECT 26.180 273.200 43.280 278.550 ;
        RECT 43.680 275.600 45.780 278.950 ;
        RECT 51.530 278.550 57.930 281.450 ;
        RECT 63.680 281.050 65.780 284.400 ;
        RECT 66.180 281.450 83.280 286.800 ;
        RECT 60.330 278.950 69.130 281.050 ;
        RECT 46.180 273.200 63.280 278.550 ;
        RECT 63.680 275.600 65.780 278.950 ;
        RECT 71.530 278.550 77.930 281.450 ;
        RECT 83.680 281.050 85.780 284.400 ;
        RECT 86.180 281.450 103.280 286.800 ;
        RECT 80.330 278.950 89.130 281.050 ;
        RECT 66.180 273.200 83.280 278.550 ;
        RECT 83.680 275.600 85.780 278.950 ;
        RECT 91.530 278.550 97.930 281.450 ;
        RECT 103.680 281.050 105.780 284.400 ;
        RECT 106.180 281.450 123.280 286.800 ;
        RECT 100.330 278.950 109.130 281.050 ;
        RECT 86.180 273.200 103.280 278.550 ;
        RECT 103.680 275.600 105.780 278.950 ;
        RECT 111.530 278.550 117.930 281.450 ;
        RECT 123.680 281.050 124.730 284.400 ;
        RECT 120.330 278.950 124.730 281.050 ;
        RECT 106.180 273.200 123.280 278.550 ;
        RECT 123.680 275.600 124.730 278.950 ;
        RECT 4.730 266.800 124.730 273.200 ;
        RECT 4.730 261.050 5.780 264.400 ;
        RECT 6.180 261.450 23.280 266.800 ;
        RECT 4.730 258.950 9.130 261.050 ;
        RECT 4.730 255.600 5.780 258.950 ;
        RECT 11.530 258.550 17.930 261.450 ;
        RECT 23.680 261.050 25.780 264.400 ;
        RECT 26.180 261.450 43.280 266.800 ;
        RECT 20.330 258.950 29.130 261.050 ;
        RECT 6.180 253.200 23.280 258.550 ;
        RECT 23.680 255.600 25.780 258.950 ;
        RECT 31.530 258.550 37.930 261.450 ;
        RECT 43.680 261.050 45.780 264.400 ;
        RECT 46.180 261.450 63.280 266.800 ;
        RECT 40.330 258.950 49.130 261.050 ;
        RECT 26.180 253.200 43.280 258.550 ;
        RECT 43.680 255.600 45.780 258.950 ;
        RECT 51.530 258.550 57.930 261.450 ;
        RECT 63.680 261.050 65.780 264.400 ;
        RECT 66.180 261.450 83.280 266.800 ;
        RECT 60.330 258.950 69.130 261.050 ;
        RECT 46.180 253.200 63.280 258.550 ;
        RECT 63.680 255.600 65.780 258.950 ;
        RECT 71.530 258.550 77.930 261.450 ;
        RECT 83.680 261.050 85.780 264.400 ;
        RECT 86.180 261.450 103.280 266.800 ;
        RECT 80.330 258.950 89.130 261.050 ;
        RECT 66.180 253.200 83.280 258.550 ;
        RECT 83.680 255.600 85.780 258.950 ;
        RECT 91.530 258.550 97.930 261.450 ;
        RECT 103.680 261.050 105.780 264.400 ;
        RECT 106.180 261.450 123.280 266.800 ;
        RECT 100.330 258.950 109.130 261.050 ;
        RECT 86.180 253.200 103.280 258.550 ;
        RECT 103.680 255.600 105.780 258.950 ;
        RECT 111.530 258.550 117.930 261.450 ;
        RECT 123.680 261.050 124.730 264.400 ;
        RECT 120.330 258.950 124.730 261.050 ;
        RECT 106.180 253.200 123.280 258.550 ;
        RECT 123.680 255.600 124.730 258.950 ;
        RECT 4.730 246.800 124.730 253.200 ;
        RECT 4.730 241.050 5.780 244.400 ;
        RECT 6.180 241.450 23.280 246.800 ;
        RECT 4.730 238.950 9.130 241.050 ;
        RECT 4.730 235.600 5.780 238.950 ;
        RECT 11.530 238.550 17.930 241.450 ;
        RECT 23.680 241.050 25.780 244.400 ;
        RECT 26.180 241.450 43.280 246.800 ;
        RECT 20.330 238.950 29.130 241.050 ;
        RECT 6.180 233.200 23.280 238.550 ;
        RECT 23.680 235.600 25.780 238.950 ;
        RECT 31.530 238.550 37.930 241.450 ;
        RECT 43.680 241.050 45.780 244.400 ;
        RECT 46.180 241.450 63.280 246.800 ;
        RECT 40.330 238.950 49.130 241.050 ;
        RECT 26.180 233.200 43.280 238.550 ;
        RECT 43.680 235.600 45.780 238.950 ;
        RECT 51.530 238.550 57.930 241.450 ;
        RECT 63.680 241.050 65.780 244.400 ;
        RECT 66.180 241.450 83.280 246.800 ;
        RECT 60.330 238.950 69.130 241.050 ;
        RECT 46.180 233.200 63.280 238.550 ;
        RECT 63.680 235.600 65.780 238.950 ;
        RECT 71.530 238.550 77.930 241.450 ;
        RECT 83.680 241.050 85.780 244.400 ;
        RECT 86.180 241.450 103.280 246.800 ;
        RECT 80.330 238.950 89.130 241.050 ;
        RECT 66.180 233.200 83.280 238.550 ;
        RECT 83.680 235.600 85.780 238.950 ;
        RECT 91.530 238.550 97.930 241.450 ;
        RECT 103.680 241.050 105.780 244.400 ;
        RECT 106.180 241.450 123.280 246.800 ;
        RECT 100.330 238.950 109.130 241.050 ;
        RECT 86.180 233.200 103.280 238.550 ;
        RECT 103.680 235.600 105.780 238.950 ;
        RECT 111.530 238.550 117.930 241.450 ;
        RECT 123.680 241.050 124.730 244.400 ;
        RECT 120.330 238.950 124.730 241.050 ;
        RECT 106.180 233.200 123.280 238.550 ;
        RECT 123.680 235.600 124.730 238.950 ;
        RECT 4.730 226.800 124.730 233.200 ;
        RECT 4.730 221.050 5.780 224.400 ;
        RECT 6.180 221.450 23.280 226.800 ;
        RECT 4.730 218.950 9.130 221.050 ;
        RECT 4.730 215.600 5.780 218.950 ;
        RECT 11.530 218.550 17.930 221.450 ;
        RECT 23.680 221.050 25.780 224.400 ;
        RECT 26.180 221.450 43.280 226.800 ;
        RECT 20.330 218.950 29.130 221.050 ;
        RECT 6.180 213.200 23.280 218.550 ;
        RECT 23.680 215.600 25.780 218.950 ;
        RECT 31.530 218.550 37.930 221.450 ;
        RECT 43.680 221.050 45.780 224.400 ;
        RECT 46.180 221.450 63.280 226.800 ;
        RECT 40.330 218.950 49.130 221.050 ;
        RECT 26.180 213.200 43.280 218.550 ;
        RECT 43.680 215.600 45.780 218.950 ;
        RECT 51.530 218.550 57.930 221.450 ;
        RECT 63.680 221.050 65.780 224.400 ;
        RECT 66.180 221.450 83.280 226.800 ;
        RECT 60.330 218.950 69.130 221.050 ;
        RECT 46.180 213.200 63.280 218.550 ;
        RECT 63.680 215.600 65.780 218.950 ;
        RECT 71.530 218.550 77.930 221.450 ;
        RECT 83.680 221.050 85.780 224.400 ;
        RECT 86.180 221.450 103.280 226.800 ;
        RECT 80.330 218.950 89.130 221.050 ;
        RECT 66.180 213.200 83.280 218.550 ;
        RECT 83.680 215.600 85.780 218.950 ;
        RECT 91.530 218.550 97.930 221.450 ;
        RECT 103.680 221.050 105.780 224.400 ;
        RECT 106.180 221.450 123.280 226.800 ;
        RECT 100.330 218.950 109.130 221.050 ;
        RECT 86.180 213.200 103.280 218.550 ;
        RECT 103.680 215.600 105.780 218.950 ;
        RECT 111.530 218.550 117.930 221.450 ;
        RECT 123.680 221.050 124.730 224.400 ;
        RECT 120.330 218.950 124.730 221.050 ;
        RECT 106.180 213.200 123.280 218.550 ;
        RECT 123.680 215.600 124.730 218.950 ;
        RECT 4.730 206.800 124.730 213.200 ;
        RECT 4.730 201.050 5.780 204.400 ;
        RECT 6.180 201.450 23.280 206.800 ;
        RECT 4.730 200.000 9.130 201.050 ;
        RECT 11.530 200.000 17.930 201.450 ;
        RECT 23.680 201.050 25.780 204.400 ;
        RECT 26.180 201.450 43.280 206.800 ;
        RECT 20.330 200.000 29.130 201.050 ;
        RECT 31.530 200.000 37.930 201.450 ;
        RECT 43.680 201.050 45.780 204.400 ;
        RECT 46.180 201.450 63.280 206.800 ;
        RECT 40.330 200.000 49.130 201.050 ;
        RECT 51.530 200.000 57.930 201.450 ;
        RECT 63.680 201.050 65.780 204.400 ;
        RECT 66.180 201.450 83.280 206.800 ;
        RECT 60.330 200.000 69.130 201.050 ;
        RECT 71.530 200.000 77.930 201.450 ;
        RECT 83.680 201.050 85.780 204.400 ;
        RECT 86.180 201.450 103.280 206.800 ;
        RECT 80.330 200.000 89.130 201.050 ;
        RECT 91.530 200.000 97.930 201.450 ;
        RECT 103.680 201.050 105.780 204.400 ;
        RECT 106.180 201.450 123.280 206.800 ;
        RECT 100.330 200.000 109.130 201.050 ;
        RECT 111.530 200.000 117.930 201.450 ;
        RECT 123.680 201.050 124.730 204.400 ;
        RECT 120.330 200.000 124.730 201.050 ;
        RECT 11.530 179.710 14.340 200.000 ;
        RECT 11.230 178.875 14.340 179.710 ;
        RECT 11.530 178.870 14.340 178.875 ;
        RECT 20.595 178.770 22.450 200.000 ;
        RECT 11.530 140.000 13.690 162.380 ;
        RECT 11.530 138.550 17.930 140.000 ;
        RECT 31.530 138.550 37.930 140.000 ;
        RECT 51.530 138.550 57.930 140.000 ;
        RECT 71.530 138.550 77.930 140.000 ;
        RECT 91.530 138.550 97.930 140.000 ;
        RECT 111.530 138.550 117.930 140.000 ;
        RECT 6.180 133.200 23.280 138.550 ;
        RECT 26.180 133.200 43.280 138.550 ;
        RECT 46.180 133.200 63.280 138.550 ;
        RECT 66.180 133.200 83.280 138.550 ;
        RECT 86.180 133.200 103.280 138.550 ;
        RECT 106.180 133.200 123.280 138.550 ;
        RECT 4.730 126.800 124.730 133.200 ;
        RECT 6.180 121.450 23.280 126.800 ;
        RECT 26.180 121.450 43.280 126.800 ;
        RECT 46.180 121.450 63.280 126.800 ;
        RECT 66.180 121.450 83.280 126.800 ;
        RECT 86.180 121.450 103.280 126.800 ;
        RECT 106.180 121.450 123.280 126.800 ;
        RECT 11.530 118.550 17.930 121.450 ;
        RECT 31.530 118.550 37.930 121.450 ;
        RECT 51.530 118.550 57.930 121.450 ;
        RECT 71.530 118.550 77.930 121.450 ;
        RECT 91.530 118.550 97.930 121.450 ;
        RECT 111.530 118.550 117.930 121.450 ;
        RECT 6.180 113.200 23.280 118.550 ;
        RECT 26.180 113.200 43.280 118.550 ;
        RECT 46.180 113.200 63.280 118.550 ;
        RECT 66.180 113.200 83.280 118.550 ;
        RECT 86.180 113.200 103.280 118.550 ;
        RECT 106.180 113.200 123.280 118.550 ;
        RECT 4.730 106.800 124.730 113.200 ;
        RECT 6.180 101.450 23.280 106.800 ;
        RECT 26.180 101.450 43.280 106.800 ;
        RECT 46.180 101.450 63.280 106.800 ;
        RECT 66.180 101.450 83.280 106.800 ;
        RECT 86.180 101.450 103.280 106.800 ;
        RECT 106.180 101.450 123.280 106.800 ;
        RECT 11.530 98.550 17.930 101.450 ;
        RECT 31.530 98.550 37.930 101.450 ;
        RECT 51.530 98.550 57.930 101.450 ;
        RECT 71.530 98.550 77.930 101.450 ;
        RECT 91.530 98.550 97.930 101.450 ;
        RECT 111.530 98.550 117.930 101.450 ;
        RECT 6.180 93.200 23.280 98.550 ;
        RECT 26.180 93.200 43.280 98.550 ;
        RECT 46.180 93.200 63.280 98.550 ;
        RECT 66.180 93.200 83.280 98.550 ;
        RECT 86.180 93.200 103.280 98.550 ;
        RECT 106.180 93.200 123.280 98.550 ;
        RECT 4.730 86.800 124.730 93.200 ;
        RECT 6.180 81.450 23.280 86.800 ;
        RECT 26.180 81.450 43.280 86.800 ;
        RECT 46.180 81.450 63.280 86.800 ;
        RECT 66.180 81.450 83.280 86.800 ;
        RECT 86.180 81.450 103.280 86.800 ;
        RECT 106.180 81.450 123.280 86.800 ;
        RECT 11.530 78.550 17.930 81.450 ;
        RECT 31.530 78.550 37.930 81.450 ;
        RECT 51.530 78.550 57.930 81.450 ;
        RECT 71.530 78.550 77.930 81.450 ;
        RECT 91.530 78.550 97.930 81.450 ;
        RECT 111.530 78.550 117.930 81.450 ;
        RECT 6.180 73.200 23.280 78.550 ;
        RECT 26.180 73.200 43.280 78.550 ;
        RECT 46.180 73.200 63.280 78.550 ;
        RECT 66.180 73.200 83.280 78.550 ;
        RECT 86.180 73.200 103.280 78.550 ;
        RECT 106.180 73.200 123.280 78.550 ;
        RECT 4.730 66.800 124.730 73.200 ;
        RECT 6.180 61.450 23.280 66.800 ;
        RECT 26.180 61.450 43.280 66.800 ;
        RECT 46.180 61.450 63.280 66.800 ;
        RECT 66.180 61.450 83.280 66.800 ;
        RECT 86.180 61.450 103.280 66.800 ;
        RECT 106.180 61.450 123.280 66.800 ;
        RECT 11.530 58.550 17.930 61.450 ;
        RECT 31.530 58.550 37.930 61.450 ;
        RECT 51.530 58.550 57.930 61.450 ;
        RECT 71.530 58.550 77.930 61.450 ;
        RECT 91.530 58.550 97.930 61.450 ;
        RECT 111.530 58.550 117.930 61.450 ;
        RECT 6.180 53.200 23.280 58.550 ;
        RECT 26.180 53.200 43.280 58.550 ;
        RECT 46.180 53.200 63.280 58.550 ;
        RECT 66.180 53.200 83.280 58.550 ;
        RECT 86.180 53.200 103.280 58.550 ;
        RECT 106.180 53.200 123.280 58.550 ;
        RECT 4.730 46.800 124.730 53.200 ;
        RECT 6.180 41.450 23.280 46.800 ;
        RECT 26.180 41.450 43.280 46.800 ;
        RECT 46.180 41.450 63.280 46.800 ;
        RECT 66.180 41.450 83.280 46.800 ;
        RECT 86.180 41.450 103.280 46.800 ;
        RECT 106.180 41.450 123.280 46.800 ;
        RECT 11.530 38.550 17.930 41.450 ;
        RECT 31.530 38.550 37.930 41.450 ;
        RECT 51.530 38.550 57.930 41.450 ;
        RECT 71.530 38.550 77.930 41.450 ;
        RECT 91.530 38.550 97.930 41.450 ;
        RECT 111.530 38.550 117.930 41.450 ;
        RECT 6.180 33.200 23.280 38.550 ;
        RECT 26.180 33.200 43.280 38.550 ;
        RECT 46.180 33.200 63.280 38.550 ;
        RECT 66.180 33.200 83.280 38.550 ;
        RECT 86.180 33.200 103.280 38.550 ;
        RECT 106.180 33.200 123.280 38.550 ;
        RECT 4.730 26.800 124.730 33.200 ;
        RECT 6.180 21.450 23.280 26.800 ;
        RECT 26.180 21.450 43.280 26.800 ;
        RECT 46.180 21.450 63.280 26.800 ;
        RECT 66.180 21.450 83.280 26.800 ;
        RECT 86.180 21.450 103.280 26.800 ;
        RECT 106.180 21.450 123.280 26.800 ;
        RECT 11.530 18.550 17.930 21.450 ;
        RECT 31.530 18.550 37.930 21.450 ;
        RECT 51.530 18.550 57.930 21.450 ;
        RECT 71.530 18.550 77.930 21.450 ;
        RECT 91.530 18.550 97.930 21.450 ;
        RECT 111.530 18.550 117.930 21.450 ;
        RECT 6.180 13.200 23.280 18.550 ;
        RECT 26.180 13.200 43.280 18.550 ;
        RECT 46.180 13.200 63.280 18.550 ;
        RECT 66.180 13.200 83.280 18.550 ;
        RECT 86.180 13.200 103.280 18.550 ;
        RECT 106.180 13.200 123.280 18.550 ;
        RECT 4.730 6.800 124.730 13.200 ;
        RECT 6.180 1.450 23.280 6.800 ;
        RECT 26.180 1.450 43.280 6.800 ;
        RECT 46.180 1.450 63.280 6.800 ;
        RECT 66.180 1.450 83.280 6.800 ;
        RECT 86.180 1.450 103.280 6.800 ;
        RECT 106.180 1.450 123.280 6.800 ;
        RECT 11.530 0.000 17.930 1.450 ;
        RECT 31.530 0.000 37.930 1.450 ;
        RECT 51.530 0.000 57.930 1.450 ;
        RECT 71.530 0.000 77.930 1.450 ;
        RECT 91.530 0.000 97.930 1.450 ;
        RECT 111.530 0.000 117.930 1.450 ;
  END
END adc_vcm_generator
END LIBRARY

