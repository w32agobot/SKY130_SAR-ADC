** sch_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_array_matrix/adc_array_matrix_8Cap_12Bit.sch
.subckt adc_array_matrix_8Cap_12Bit VDD VSS sample sample_n col_n[15] col_n[14] col_n[13] col_n[12]
+ col_n[11] col_n[10] col_n[9] col_n[8] col_n[7] col_n[6] col_n[5] col_n[4] col_n[3] col_n[2] col_n[1] col_n[0]
+ colon_n[15] colon_n[14] colon_n[13] colon_n[12] colon_n[11] colon_n[10] colon_n[9] colon_n[8] colon_n[7]
+ colon_n[6] colon_n[5] colon_n[4] colon_n[3] colon_n[2] colon_n[1] colon_n[0] row_n[31] row_n[30] row_n[29]
+ row_n[28] row_n[27] row_n[26] row_n[25] row_n[24] row_n[23] row_n[22] row_n[21] row_n[20] row_n[19] row_n[18]
+ row_n[17] row_n[16] row_n[15] row_n[14] row_n[13] row_n[12] row_n[11] row_n[10] row_n[9] row_n[8] row_n[7]
+ row_n[6] row_n[5] row_n[4] row_n[3] row_n[2] row_n[1] row_n[0] vcom en_n_bit[2] en_n_bit[1] en_n_bit[0]
+ analog_in sw sw_n ctop
*.PININFO VDD:B VSS:B sample:I sample_n:I col_n[15:0]:I colon_n[15:0]:I row_n[31:0]:I vcom:B
*+ en_n_bit[2:0]:I analog_in:I sw:I sw_n:I ctop:B
x1 VDD ctop vcom col_n[0] colon_n[0] net2 net1 VSS row_n[0] adc_array_wafflecap_8_8
x2 VDD ctop vcom col_n[0] colon_n[0] net2 net1 VSS row_n[1] adc_array_wafflecap_8_8
x3 VDD ctop vcom col_n[0] colon_n[0] net2 net1 VSS row_n[2] adc_array_wafflecap_8_8
x4 VDD ctop vcom col_n[0] colon_n[0] net2 net1 VSS row_n[3] adc_array_wafflecap_8_8
x5 VDD ctop vcom col_n[0] colon_n[0] net2 net1 VSS row_n[4] adc_array_wafflecap_8_8
x6 VDD ctop vcom col_n[0] colon_n[0] net2 net1 VSS row_n[5] adc_array_wafflecap_8_8
x7 VDD ctop vcom col_n[0] colon_n[0] net2 net1 VSS row_n[6] adc_array_wafflecap_8_8
x8 VDD ctop vcom col_n[0] colon_n[0] net2 net1 VSS row_n[7] adc_array_wafflecap_8_8
x9 VDD ctop vcom col_n[0] colon_n[0] net2 net1 VSS row_n[8] adc_array_wafflecap_8_8
x10 VDD ctop vcom col_n[0] colon_n[0] net2 net1 VSS row_n[9] adc_array_wafflecap_8_8
x11 VDD ctop vcom col_n[0] colon_n[0] net2 net1 VSS row_n[10] adc_array_wafflecap_8_8
x12 VDD ctop vcom col_n[0] colon_n[0] net2 net1 VSS row_n[11] adc_array_wafflecap_8_8
x13 VDD ctop vcom col_n[0] colon_n[0] net2 net1 VSS row_n[12] adc_array_wafflecap_8_8
x14 VDD ctop vcom col_n[0] colon_n[0] net2 net1 VSS row_n[13] adc_array_wafflecap_8_8
x15 VDD ctop vcom col_n[0] colon_n[0] net2 net1 VSS row_n[14] adc_array_wafflecap_8_8
x16 VDD ctop vcom col_n[0] colon_n[0] net2 net1 VSS row_n[15] adc_array_wafflecap_8_8
x17 VDD ctop vcom col_n[0] colon_n[0] net2 net1 VSS row_n[16] adc_array_wafflecap_8_8
x18 VDD ctop vcom col_n[0] colon_n[0] net2 net1 VSS row_n[17] adc_array_wafflecap_8_8
x19 VDD ctop vcom col_n[0] colon_n[0] net2 net1 VSS row_n[18] adc_array_wafflecap_8_8
x20 VDD ctop vcom col_n[0] colon_n[0] net2 net1 VSS row_n[19] adc_array_wafflecap_8_8
x21 VDD ctop vcom col_n[0] colon_n[0] net2 net1 VSS row_n[20] adc_array_wafflecap_8_8
x22 VDD ctop vcom col_n[0] colon_n[0] net2 net1 VSS row_n[21] adc_array_wafflecap_8_8
x23 VDD ctop vcom col_n[0] colon_n[0] net2 net1 VSS row_n[22] adc_array_wafflecap_8_8
x24 VDD ctop vcom col_n[0] colon_n[0] net2 net1 VSS row_n[23] adc_array_wafflecap_8_8
x25 VDD ctop vcom col_n[0] colon_n[0] net2 net1 VSS row_n[24] adc_array_wafflecap_8_8
x26 VDD ctop vcom col_n[0] colon_n[0] net2 net1 VSS row_n[25] adc_array_wafflecap_8_8
x27 VDD ctop vcom col_n[0] colon_n[0] net2 net1 VSS row_n[26] adc_array_wafflecap_8_8
x28 VDD ctop vcom col_n[0] colon_n[0] net2 net1 VSS row_n[27] adc_array_wafflecap_8_8
x29 VDD ctop vcom col_n[0] colon_n[0] net2 net1 VSS row_n[28] adc_array_wafflecap_8_8
x30 VDD ctop vcom col_n[0] colon_n[0] net2 net1 VSS row_n[29] adc_array_wafflecap_8_8
x31 VDD ctop vcom col_n[0] colon_n[0] net2 net1 VSS row_n[30] adc_array_wafflecap_8_8
x32 VDD ctop vcom col_n[0] colon_n[0] net2 net1 VSS row_n[31] adc_array_wafflecap_8_8
x33 VDD ctop vcom col_n[1] colon_n[1] net4 net3 VSS row_n[0] adc_array_wafflecap_8_8
x34 VDD ctop vcom col_n[1] colon_n[1] net4 net3 VSS row_n[1] adc_array_wafflecap_8_8
x35 VDD ctop vcom col_n[1] colon_n[1] net4 net3 VSS row_n[2] adc_array_wafflecap_8_8
x36 VDD ctop vcom col_n[1] colon_n[1] net4 net3 VSS row_n[3] adc_array_wafflecap_8_8
x37 VDD ctop vcom col_n[1] colon_n[1] net4 net3 VSS row_n[4] adc_array_wafflecap_8_8
x38 VDD ctop vcom col_n[1] colon_n[1] net4 net3 VSS row_n[5] adc_array_wafflecap_8_8
x39 VDD ctop vcom col_n[1] colon_n[1] net4 net3 VSS row_n[6] adc_array_wafflecap_8_8
x40 VDD ctop vcom col_n[1] colon_n[1] net4 net3 VSS row_n[7] adc_array_wafflecap_8_8
x41 VDD ctop vcom col_n[1] colon_n[1] net4 net3 VSS row_n[8] adc_array_wafflecap_8_8
x42 VDD ctop vcom col_n[1] colon_n[1] net4 net3 VSS row_n[9] adc_array_wafflecap_8_8
x43 VDD ctop vcom col_n[1] colon_n[1] net4 net3 VSS row_n[10] adc_array_wafflecap_8_8
x44 VDD ctop vcom col_n[1] colon_n[1] net4 net3 VSS row_n[11] adc_array_wafflecap_8_8
x45 VDD ctop vcom col_n[1] colon_n[1] net4 net3 VSS row_n[12] adc_array_wafflecap_8_8
x46 VDD ctop vcom col_n[1] colon_n[1] net4 net3 VSS row_n[13] adc_array_wafflecap_8_8
x47 VDD ctop vcom col_n[1] colon_n[1] net4 net3 VSS row_n[14] adc_array_wafflecap_8_8
x48 VDD ctop vcom col_n[1] colon_n[1] net4 net3 VSS row_n[15] adc_array_wafflecap_8_8
x49 VDD ctop vcom col_n[1] colon_n[1] net4 net3 VSS row_n[16] adc_array_wafflecap_8_8
x50 VDD ctop vcom col_n[1] colon_n[1] net4 net3 VSS row_n[17] adc_array_wafflecap_8_8
x51 VDD ctop vcom col_n[1] colon_n[1] net4 net3 VSS row_n[18] adc_array_wafflecap_8_8
x52 VDD ctop vcom col_n[1] colon_n[1] net4 net3 VSS row_n[19] adc_array_wafflecap_8_8
x53 VDD ctop vcom col_n[1] colon_n[1] net4 net3 VSS row_n[20] adc_array_wafflecap_8_8
x54 VDD ctop vcom col_n[1] colon_n[1] net4 net3 VSS row_n[21] adc_array_wafflecap_8_8
x55 VDD ctop vcom col_n[1] colon_n[1] net4 net3 VSS row_n[22] adc_array_wafflecap_8_8
x56 VDD ctop vcom col_n[1] colon_n[1] net4 net3 VSS row_n[23] adc_array_wafflecap_8_8
x57 VDD ctop vcom col_n[1] colon_n[1] net4 net3 VSS row_n[24] adc_array_wafflecap_8_8
x58 VDD ctop vcom col_n[1] colon_n[1] net4 net3 VSS row_n[25] adc_array_wafflecap_8_8
x59 VDD ctop vcom col_n[1] colon_n[1] net4 net3 VSS row_n[26] adc_array_wafflecap_8_8
x60 VDD ctop vcom col_n[1] colon_n[1] net4 net3 VSS row_n[27] adc_array_wafflecap_8_8
x61 VDD ctop vcom col_n[1] colon_n[1] net4 net3 VSS row_n[28] adc_array_wafflecap_8_8
x62 VDD ctop vcom col_n[1] colon_n[1] net4 net3 VSS row_n[29] adc_array_wafflecap_8_8
x63 VDD ctop vcom col_n[1] colon_n[1] net4 net3 VSS row_n[30] adc_array_wafflecap_8_8
x64 VDD ctop vcom col_n[1] colon_n[1] net4 net3 VSS row_n[31] adc_array_wafflecap_8_8
x65 VDD ctop vcom col_n[2] colon_n[2] net6 net5 VSS row_n[0] adc_array_wafflecap_8_8
x66 VDD ctop vcom col_n[2] colon_n[2] net6 net5 VSS row_n[1] adc_array_wafflecap_8_8
x67 VDD ctop vcom col_n[2] colon_n[2] net6 net5 VSS row_n[2] adc_array_wafflecap_8_8
x68 VDD ctop vcom col_n[2] colon_n[2] net6 net5 VSS row_n[3] adc_array_wafflecap_8_8
x69 VDD ctop vcom col_n[2] colon_n[2] net6 net5 VSS row_n[4] adc_array_wafflecap_8_8
x70 VDD ctop vcom col_n[2] colon_n[2] net6 net5 VSS row_n[5] adc_array_wafflecap_8_8
x71 VDD ctop vcom col_n[2] colon_n[2] net6 net5 VSS row_n[6] adc_array_wafflecap_8_8
x72 VDD ctop vcom col_n[2] colon_n[2] net6 net5 VSS row_n[7] adc_array_wafflecap_8_8
x73 VDD ctop vcom col_n[2] colon_n[2] net6 net5 VSS row_n[8] adc_array_wafflecap_8_8
x74 VDD ctop vcom col_n[2] colon_n[2] net6 net5 VSS row_n[9] adc_array_wafflecap_8_8
x75 VDD ctop vcom col_n[2] colon_n[2] net6 net5 VSS row_n[10] adc_array_wafflecap_8_8
x76 VDD ctop vcom col_n[2] colon_n[2] net6 net5 VSS row_n[11] adc_array_wafflecap_8_8
x77 VDD ctop vcom col_n[2] colon_n[2] net6 net5 VSS row_n[12] adc_array_wafflecap_8_8
x78 VDD ctop vcom col_n[2] colon_n[2] net6 net5 VSS row_n[13] adc_array_wafflecap_8_8
x79 VDD ctop vcom col_n[2] colon_n[2] net6 net5 VSS row_n[14] adc_array_wafflecap_8_8
x80 VDD ctop vcom col_n[2] colon_n[2] net6 net5 VSS row_n[15] adc_array_wafflecap_8_8
x81 VDD ctop vcom col_n[2] colon_n[2] net6 net5 VSS row_n[16] adc_array_wafflecap_8_8
x82 VDD ctop vcom col_n[2] colon_n[2] net6 net5 VSS row_n[17] adc_array_wafflecap_8_8
x83 VDD ctop vcom col_n[2] colon_n[2] net6 net5 VSS row_n[18] adc_array_wafflecap_8_8
x84 VDD ctop vcom col_n[2] colon_n[2] net6 net5 VSS row_n[19] adc_array_wafflecap_8_8
x85 VDD ctop vcom col_n[2] colon_n[2] net6 net5 VSS row_n[20] adc_array_wafflecap_8_8
x86 VDD ctop vcom col_n[2] colon_n[2] net6 net5 VSS row_n[21] adc_array_wafflecap_8_8
x87 VDD ctop vcom col_n[2] colon_n[2] net6 net5 VSS row_n[22] adc_array_wafflecap_8_8
x88 VDD ctop vcom col_n[2] colon_n[2] net6 net5 VSS row_n[23] adc_array_wafflecap_8_8
x89 VDD ctop vcom col_n[2] colon_n[2] net6 net5 VSS row_n[24] adc_array_wafflecap_8_8
x90 VDD ctop vcom col_n[2] colon_n[2] net6 net5 VSS row_n[25] adc_array_wafflecap_8_8
x91 VDD ctop vcom col_n[2] colon_n[2] net6 net5 VSS row_n[26] adc_array_wafflecap_8_8
x92 VDD ctop vcom col_n[2] colon_n[2] net6 net5 VSS row_n[27] adc_array_wafflecap_8_8
x93 VDD ctop vcom col_n[2] colon_n[2] net6 net5 VSS row_n[28] adc_array_wafflecap_8_8
x94 VDD ctop vcom col_n[2] colon_n[2] net6 net5 VSS row_n[29] adc_array_wafflecap_8_8
x95 VDD ctop vcom col_n[2] colon_n[2] net6 net5 VSS row_n[30] adc_array_wafflecap_8_8
x96 VDD ctop vcom col_n[2] colon_n[2] net6 net5 VSS row_n[31] adc_array_wafflecap_8_8
x97 VDD ctop vcom col_n[3] colon_n[3] net8 net7 VSS row_n[0] adc_array_wafflecap_8_8
x98 VDD ctop vcom col_n[3] colon_n[3] net8 net7 VSS row_n[1] adc_array_wafflecap_8_8
x99 VDD ctop vcom col_n[3] colon_n[3] net8 net7 VSS row_n[2] adc_array_wafflecap_8_8
x100 VDD ctop vcom col_n[3] colon_n[3] net8 net7 VSS row_n[3] adc_array_wafflecap_8_8
x101 VDD ctop vcom col_n[3] colon_n[3] net8 net7 VSS row_n[4] adc_array_wafflecap_8_8
x102 VDD ctop vcom col_n[3] colon_n[3] net8 net7 VSS row_n[5] adc_array_wafflecap_8_8
x103 VDD ctop vcom col_n[3] colon_n[3] net8 net7 VSS row_n[6] adc_array_wafflecap_8_8
x104 VDD ctop vcom col_n[3] colon_n[3] net8 net7 VSS row_n[7] adc_array_wafflecap_8_8
x105 VDD ctop vcom col_n[3] colon_n[3] net8 net7 VSS row_n[8] adc_array_wafflecap_8_8
x106 VDD ctop vcom col_n[3] colon_n[3] net8 net7 VSS row_n[9] adc_array_wafflecap_8_8
x107 VDD ctop vcom col_n[3] colon_n[3] net8 net7 VSS row_n[10] adc_array_wafflecap_8_8
x108 VDD ctop vcom col_n[3] colon_n[3] net8 net7 VSS row_n[11] adc_array_wafflecap_8_8
x109 VDD ctop vcom col_n[3] colon_n[3] net8 net7 VSS row_n[12] adc_array_wafflecap_8_8
x110 VDD ctop vcom col_n[3] colon_n[3] net8 net7 VSS row_n[13] adc_array_wafflecap_8_8
x111 VDD ctop vcom col_n[3] colon_n[3] net8 net7 VSS row_n[14] adc_array_wafflecap_8_8
x112 VDD ctop vcom col_n[3] colon_n[3] net8 net7 VSS row_n[15] adc_array_wafflecap_8_8
x113 VDD ctop vcom col_n[3] colon_n[3] net8 net7 VSS row_n[16] adc_array_wafflecap_8_8
x114 VDD ctop vcom col_n[3] colon_n[3] net8 net7 VSS row_n[17] adc_array_wafflecap_8_8
x115 VDD ctop vcom col_n[3] colon_n[3] net8 net7 VSS row_n[18] adc_array_wafflecap_8_8
x116 VDD ctop vcom col_n[3] colon_n[3] net8 net7 VSS row_n[19] adc_array_wafflecap_8_8
x117 VDD ctop vcom col_n[3] colon_n[3] net8 net7 VSS row_n[20] adc_array_wafflecap_8_8
x118 VDD ctop vcom col_n[3] colon_n[3] net8 net7 VSS row_n[21] adc_array_wafflecap_8_8
x119 VDD ctop vcom col_n[3] colon_n[3] net8 net7 VSS row_n[22] adc_array_wafflecap_8_8
x120 VDD ctop vcom col_n[3] colon_n[3] net8 net7 VSS row_n[23] adc_array_wafflecap_8_8
x121 VDD ctop vcom col_n[3] colon_n[3] net8 net7 VSS row_n[24] adc_array_wafflecap_8_8
x122 VDD ctop vcom col_n[3] colon_n[3] net8 net7 VSS row_n[25] adc_array_wafflecap_8_8
x123 VDD ctop vcom col_n[3] colon_n[3] net8 net7 VSS row_n[26] adc_array_wafflecap_8_8
x124 VDD ctop vcom col_n[3] colon_n[3] net8 net7 VSS row_n[27] adc_array_wafflecap_8_8
x125 VDD ctop vcom col_n[3] colon_n[3] net8 net7 VSS row_n[28] adc_array_wafflecap_8_8
x126 VDD ctop vcom col_n[3] colon_n[3] net8 net7 VSS row_n[29] adc_array_wafflecap_8_8
x127 VDD ctop vcom col_n[3] colon_n[3] net8 net7 VSS row_n[30] adc_array_wafflecap_8_8
x128 VDD ctop vcom col_n[3] colon_n[3] net8 net7 VSS row_n[31] adc_array_wafflecap_8_8
x129 VDD ctop vcom col_n[4] colon_n[4] net10 net9 VSS row_n[0] adc_array_wafflecap_8_8
x130 VDD ctop vcom col_n[4] colon_n[4] net10 net9 VSS row_n[1] adc_array_wafflecap_8_8
x131 VDD ctop vcom col_n[4] colon_n[4] net10 net9 VSS row_n[2] adc_array_wafflecap_8_8
x132 VDD ctop vcom col_n[4] colon_n[4] net10 net9 VSS row_n[3] adc_array_wafflecap_8_8
x133 VDD ctop vcom col_n[4] colon_n[4] net10 net9 VSS row_n[4] adc_array_wafflecap_8_8
x134 VDD ctop vcom col_n[4] colon_n[4] net10 net9 VSS row_n[5] adc_array_wafflecap_8_8
x135 VDD ctop vcom col_n[4] colon_n[4] net10 net9 VSS row_n[6] adc_array_wafflecap_8_8
x136 VDD ctop vcom col_n[4] colon_n[4] net10 net9 VSS row_n[7] adc_array_wafflecap_8_8
x137 VDD ctop vcom col_n[4] colon_n[4] net10 net9 VSS row_n[8] adc_array_wafflecap_8_8
x138 VDD ctop vcom col_n[4] colon_n[4] net10 net9 VSS row_n[9] adc_array_wafflecap_8_8
x139 VDD ctop vcom col_n[4] colon_n[4] net10 net9 VSS row_n[10] adc_array_wafflecap_8_8
x140 VDD ctop vcom col_n[4] colon_n[4] net10 net9 VSS row_n[11] adc_array_wafflecap_8_8
x141 VDD ctop vcom col_n[4] colon_n[4] net10 net9 VSS row_n[12] adc_array_wafflecap_8_8
x142 VDD ctop vcom col_n[4] colon_n[4] net10 net9 VSS row_n[13] adc_array_wafflecap_8_8
x143 VDD ctop vcom col_n[4] colon_n[4] net10 net9 VSS row_n[14] adc_array_wafflecap_8_8
x144 VDD ctop vcom col_n[4] colon_n[4] net10 net9 VSS row_n[15] adc_array_wafflecap_8_8
x145 VDD ctop vcom col_n[4] colon_n[4] net10 net9 VSS row_n[16] adc_array_wafflecap_8_8
x146 VDD ctop vcom col_n[4] colon_n[4] net10 net9 VSS row_n[17] adc_array_wafflecap_8_8
x147 VDD ctop vcom col_n[4] colon_n[4] net10 net9 VSS row_n[18] adc_array_wafflecap_8_8
x148 VDD ctop vcom col_n[4] colon_n[4] net10 net9 VSS row_n[19] adc_array_wafflecap_8_8
x149 VDD ctop vcom col_n[4] colon_n[4] net10 net9 VSS row_n[20] adc_array_wafflecap_8_8
x150 VDD ctop vcom col_n[4] colon_n[4] net10 net9 VSS row_n[21] adc_array_wafflecap_8_8
x151 VDD ctop vcom col_n[4] colon_n[4] net10 net9 VSS row_n[22] adc_array_wafflecap_8_8
x152 VDD ctop vcom col_n[4] colon_n[4] net10 net9 VSS row_n[23] adc_array_wafflecap_8_8
x153 VDD ctop vcom col_n[4] colon_n[4] net10 net9 VSS row_n[24] adc_array_wafflecap_8_8
x154 VDD ctop vcom col_n[4] colon_n[4] net10 net9 VSS row_n[25] adc_array_wafflecap_8_8
x155 VDD ctop vcom col_n[4] colon_n[4] net10 net9 VSS row_n[26] adc_array_wafflecap_8_8
x156 VDD ctop vcom col_n[4] colon_n[4] net10 net9 VSS row_n[27] adc_array_wafflecap_8_8
x157 VDD ctop vcom col_n[4] colon_n[4] net10 net9 VSS row_n[28] adc_array_wafflecap_8_8
x158 VDD ctop vcom col_n[4] colon_n[4] net10 net9 VSS row_n[29] adc_array_wafflecap_8_8
x159 VDD ctop vcom col_n[4] colon_n[4] net10 net9 VSS row_n[30] adc_array_wafflecap_8_8
x160 VDD ctop vcom col_n[4] colon_n[4] net10 net9 VSS row_n[31] adc_array_wafflecap_8_8
x161 VDD ctop vcom col_n[5] colon_n[5] net12 net11 VSS row_n[0] adc_array_wafflecap_8_8
x162 VDD ctop vcom col_n[5] colon_n[5] net12 net11 VSS row_n[1] adc_array_wafflecap_8_8
x163 VDD ctop vcom col_n[5] colon_n[5] net12 net11 VSS row_n[2] adc_array_wafflecap_8_8
x164 VDD ctop vcom col_n[5] colon_n[5] net12 net11 VSS row_n[3] adc_array_wafflecap_8_8
x165 VDD ctop vcom col_n[5] colon_n[5] net12 net11 VSS row_n[4] adc_array_wafflecap_8_8
x166 VDD ctop vcom col_n[5] colon_n[5] net12 net11 VSS row_n[5] adc_array_wafflecap_8_8
x167 VDD ctop vcom col_n[5] colon_n[5] net12 net11 VSS row_n[6] adc_array_wafflecap_8_8
x168 VDD ctop vcom col_n[5] colon_n[5] net12 net11 VSS row_n[7] adc_array_wafflecap_8_8
x169 VDD ctop vcom col_n[5] colon_n[5] net12 net11 VSS row_n[8] adc_array_wafflecap_8_8
x170 VDD ctop vcom col_n[5] colon_n[5] net12 net11 VSS row_n[9] adc_array_wafflecap_8_8
x171 VDD ctop vcom col_n[5] colon_n[5] net12 net11 VSS row_n[10] adc_array_wafflecap_8_8
x172 VDD ctop vcom col_n[5] colon_n[5] net12 net11 VSS row_n[11] adc_array_wafflecap_8_8
x173 VDD ctop vcom col_n[5] colon_n[5] net12 net11 VSS row_n[12] adc_array_wafflecap_8_8
x174 VDD ctop vcom col_n[5] colon_n[5] net12 net11 VSS row_n[13] adc_array_wafflecap_8_8
x175 VDD ctop vcom col_n[5] colon_n[5] net12 net11 VSS row_n[14] adc_array_wafflecap_8_8
x176 VDD ctop vcom col_n[5] colon_n[5] net12 net11 VSS row_n[15] adc_array_wafflecap_8_8
x177 VDD ctop vcom col_n[5] colon_n[5] net12 net11 VSS row_n[16] adc_array_wafflecap_8_8
x178 VDD ctop vcom col_n[5] colon_n[5] net12 net11 VSS row_n[17] adc_array_wafflecap_8_8
x179 VDD ctop vcom col_n[5] colon_n[5] net12 net11 VSS row_n[18] adc_array_wafflecap_8_8
x180 VDD ctop vcom col_n[5] colon_n[5] net12 net11 VSS row_n[19] adc_array_wafflecap_8_8
x181 VDD ctop vcom col_n[5] colon_n[5] net12 net11 VSS row_n[20] adc_array_wafflecap_8_8
x182 VDD ctop vcom col_n[5] colon_n[5] net12 net11 VSS row_n[21] adc_array_wafflecap_8_8
x183 VDD ctop vcom col_n[5] colon_n[5] net12 net11 VSS row_n[22] adc_array_wafflecap_8_8
x184 VDD ctop vcom col_n[5] colon_n[5] net12 net11 VSS row_n[23] adc_array_wafflecap_8_8
x185 VDD ctop vcom col_n[5] colon_n[5] net12 net11 VSS row_n[24] adc_array_wafflecap_8_8
x186 VDD ctop vcom col_n[5] colon_n[5] net12 net11 VSS row_n[25] adc_array_wafflecap_8_8
x187 VDD ctop vcom col_n[5] colon_n[5] net12 net11 VSS row_n[26] adc_array_wafflecap_8_8
x188 VDD ctop vcom col_n[5] colon_n[5] net12 net11 VSS row_n[27] adc_array_wafflecap_8_8
x189 VDD ctop vcom col_n[5] colon_n[5] net12 net11 VSS row_n[28] adc_array_wafflecap_8_8
x190 VDD ctop vcom col_n[5] colon_n[5] net12 net11 VSS row_n[29] adc_array_wafflecap_8_8
x191 VDD ctop vcom col_n[5] colon_n[5] net12 net11 VSS row_n[30] adc_array_wafflecap_8_8
x192 VDD ctop vcom col_n[5] colon_n[5] net12 net11 VSS row_n[31] adc_array_wafflecap_8_8
x193 VDD ctop vcom col_n[6] colon_n[6] net14 net13 VSS row_n[0] adc_array_wafflecap_8_8
x194 VDD ctop vcom col_n[6] colon_n[6] net14 net13 VSS row_n[1] adc_array_wafflecap_8_8
x195 VDD ctop vcom col_n[6] colon_n[6] net14 net13 VSS row_n[2] adc_array_wafflecap_8_8
x196 VDD ctop vcom col_n[6] colon_n[6] net14 net13 VSS row_n[3] adc_array_wafflecap_8_8
x197 VDD ctop vcom col_n[6] colon_n[6] net14 net13 VSS row_n[4] adc_array_wafflecap_8_8
x198 VDD ctop vcom col_n[6] colon_n[6] net14 net13 VSS row_n[5] adc_array_wafflecap_8_8
x199 VDD ctop vcom col_n[6] colon_n[6] net14 net13 VSS row_n[6] adc_array_wafflecap_8_8
x200 VDD ctop vcom col_n[6] colon_n[6] net14 net13 VSS row_n[7] adc_array_wafflecap_8_8
x201 VDD ctop vcom col_n[6] colon_n[6] net14 net13 VSS row_n[8] adc_array_wafflecap_8_8
x202 VDD ctop vcom col_n[6] colon_n[6] net14 net13 VSS row_n[9] adc_array_wafflecap_8_8
x203 VDD ctop vcom col_n[6] colon_n[6] net14 net13 VSS row_n[10] adc_array_wafflecap_8_8
x204 VDD ctop vcom col_n[6] colon_n[6] net14 net13 VSS row_n[11] adc_array_wafflecap_8_8
x205 VDD ctop vcom col_n[6] colon_n[6] net14 net13 VSS row_n[12] adc_array_wafflecap_8_8
x206 VDD ctop vcom col_n[6] colon_n[6] net14 net13 VSS row_n[13] adc_array_wafflecap_8_8
x207 VDD ctop vcom col_n[6] colon_n[6] net14 net13 VSS row_n[14] adc_array_wafflecap_8_8
x208 VDD ctop vcom col_n[6] colon_n[6] net14 net13 VSS row_n[15] adc_array_wafflecap_8_8
x209 VDD ctop vcom col_n[6] colon_n[6] net14 net13 VSS row_n[16] adc_array_wafflecap_8_8
x210 VDD ctop vcom col_n[6] colon_n[6] net14 net13 VSS row_n[17] adc_array_wafflecap_8_8
x211 VDD ctop vcom col_n[6] colon_n[6] net14 net13 VSS row_n[18] adc_array_wafflecap_8_8
x212 VDD ctop vcom col_n[6] colon_n[6] net14 net13 VSS row_n[19] adc_array_wafflecap_8_8
x213 VDD ctop vcom col_n[6] colon_n[6] net14 net13 VSS row_n[20] adc_array_wafflecap_8_8
x214 VDD ctop vcom col_n[6] colon_n[6] net14 net13 VSS row_n[21] adc_array_wafflecap_8_8
x215 VDD ctop vcom col_n[6] colon_n[6] net14 net13 VSS row_n[22] adc_array_wafflecap_8_8
x216 VDD ctop vcom col_n[6] colon_n[6] net14 net13 VSS row_n[23] adc_array_wafflecap_8_8
x217 VDD ctop vcom col_n[6] colon_n[6] net14 net13 VSS row_n[24] adc_array_wafflecap_8_8
x218 VDD ctop vcom col_n[6] colon_n[6] net14 net13 VSS row_n[25] adc_array_wafflecap_8_8
x219 VDD ctop vcom col_n[6] colon_n[6] net14 net13 VSS row_n[26] adc_array_wafflecap_8_8
x220 VDD ctop vcom col_n[6] colon_n[6] net14 net13 VSS row_n[27] adc_array_wafflecap_8_8
x221 VDD ctop vcom col_n[6] colon_n[6] net14 net13 VSS row_n[28] adc_array_wafflecap_8_8
x222 VDD ctop vcom col_n[6] colon_n[6] net14 net13 VSS row_n[29] adc_array_wafflecap_8_8
x223 VDD ctop vcom col_n[6] colon_n[6] net14 net13 VSS row_n[30] adc_array_wafflecap_8_8
x224 VDD ctop vcom col_n[6] colon_n[6] net14 net13 VSS row_n[31] adc_array_wafflecap_8_8
x225 VDD ctop vcom col_n[7] colon_n[7] net16 net15 VSS row_n[0] adc_array_wafflecap_8_8
x226 VDD ctop vcom col_n[7] colon_n[7] net16 net15 VSS row_n[1] adc_array_wafflecap_8_8
x227 VDD ctop vcom col_n[7] colon_n[7] net16 net15 VSS row_n[2] adc_array_wafflecap_8_8
x228 VDD ctop vcom col_n[7] colon_n[7] net16 net15 VSS row_n[3] adc_array_wafflecap_8_8
x229 VDD ctop vcom col_n[7] colon_n[7] net16 net15 VSS row_n[4] adc_array_wafflecap_8_8
x230 VDD ctop vcom col_n[7] colon_n[7] net16 net15 VSS row_n[5] adc_array_wafflecap_8_8
x231 VDD ctop vcom col_n[7] colon_n[7] net16 net15 VSS row_n[6] adc_array_wafflecap_8_8
x232 VDD ctop vcom col_n[7] colon_n[7] net16 net15 VSS row_n[7] adc_array_wafflecap_8_8
x233 VDD ctop vcom col_n[7] colon_n[7] net16 net15 VSS row_n[8] adc_array_wafflecap_8_8
x234 VDD ctop vcom col_n[7] colon_n[7] net16 net15 VSS row_n[9] adc_array_wafflecap_8_8
x235 VDD ctop vcom col_n[7] colon_n[7] net16 net15 VSS row_n[10] adc_array_wafflecap_8_8
x236 VDD ctop vcom col_n[7] colon_n[7] net16 net15 VSS row_n[11] adc_array_wafflecap_8_8
x237 VDD ctop vcom col_n[7] colon_n[7] net16 net15 VSS row_n[12] adc_array_wafflecap_8_8
x238 VDD ctop vcom col_n[7] colon_n[7] net16 net15 VSS row_n[13] adc_array_wafflecap_8_8
x239 VDD ctop vcom col_n[7] colon_n[7] net16 net15 VSS row_n[14] adc_array_wafflecap_8_8
x240 VDD ctop vcom col_n[7] colon_n[7] net16 net15 VSS row_n[15] adc_array_wafflecap_8_8
x241 VDD ctop vcom col_n[7] colon_n[7] net16 net15 VSS row_n[16] adc_array_wafflecap_8_8
x242 VDD ctop vcom col_n[7] colon_n[7] net16 net15 VSS row_n[17] adc_array_wafflecap_8_8
x243 VDD ctop vcom col_n[7] colon_n[7] net16 net15 VSS row_n[18] adc_array_wafflecap_8_8
x244 VDD ctop vcom col_n[7] colon_n[7] net16 net15 VSS row_n[19] adc_array_wafflecap_8_8
x245 VDD ctop vcom col_n[7] colon_n[7] net16 net15 VSS row_n[20] adc_array_wafflecap_8_8
x246 VDD ctop vcom col_n[7] colon_n[7] net16 net15 VSS row_n[21] adc_array_wafflecap_8_8
x247 VDD ctop vcom col_n[7] colon_n[7] net16 net15 VSS row_n[22] adc_array_wafflecap_8_8
x248 VDD ctop vcom col_n[7] colon_n[7] net16 net15 VSS row_n[23] adc_array_wafflecap_8_8
x249 VDD ctop vcom col_n[7] colon_n[7] net16 net15 VSS row_n[24] adc_array_wafflecap_8_8
x250 VDD ctop vcom col_n[7] colon_n[7] net16 net15 VSS row_n[25] adc_array_wafflecap_8_8
x251 VDD ctop vcom col_n[7] colon_n[7] net16 net15 VSS row_n[26] adc_array_wafflecap_8_8
x252 VDD ctop vcom col_n[7] colon_n[7] net16 net15 VSS row_n[27] adc_array_wafflecap_8_8
x253 VDD ctop vcom col_n[7] colon_n[7] net16 net15 VSS row_n[28] adc_array_wafflecap_8_8
x254 VDD ctop vcom col_n[7] colon_n[7] net16 net15 VSS row_n[29] adc_array_wafflecap_8_8
x255 VDD ctop vcom col_n[7] colon_n[7] net16 net15 VSS row_n[30] adc_array_wafflecap_8_8
x256 VDD ctop vcom col_n[7] colon_n[7] net16 net15 VSS row_n[31] adc_array_wafflecap_8_8
x257 VDD ctop vcom col_n[8] colon_n[8] net18 net17 VSS row_n[0] adc_array_wafflecap_8_8
x258 VDD ctop vcom col_n[8] colon_n[8] net18 net17 VSS row_n[1] adc_array_wafflecap_8_8
x259 VDD ctop vcom col_n[8] colon_n[8] net18 net17 VSS row_n[2] adc_array_wafflecap_8_8
x260 VDD ctop vcom col_n[8] colon_n[8] net18 net17 VSS row_n[3] adc_array_wafflecap_8_8
x261 VDD ctop vcom col_n[8] colon_n[8] net18 net17 VSS row_n[4] adc_array_wafflecap_8_8
x262 VDD ctop vcom col_n[8] colon_n[8] net18 net17 VSS row_n[5] adc_array_wafflecap_8_8
x263 VDD ctop vcom col_n[8] colon_n[8] net18 net17 VSS row_n[6] adc_array_wafflecap_8_8
x264 VDD ctop vcom col_n[8] colon_n[8] net18 net17 VSS row_n[7] adc_array_wafflecap_8_8
x265 VDD ctop vcom col_n[8] colon_n[8] net18 net17 VSS row_n[8] adc_array_wafflecap_8_8
x266 VDD ctop vcom col_n[8] colon_n[8] net18 net17 VSS row_n[9] adc_array_wafflecap_8_8
x267 VDD ctop vcom col_n[8] colon_n[8] net18 net17 VSS row_n[10] adc_array_wafflecap_8_8
x268 VDD ctop vcom col_n[8] colon_n[8] net18 net17 VSS row_n[11] adc_array_wafflecap_8_8
x269 VDD ctop vcom col_n[8] colon_n[8] net18 net17 VSS row_n[12] adc_array_wafflecap_8_8
x270 VDD ctop vcom col_n[8] colon_n[8] net18 net17 VSS row_n[13] adc_array_wafflecap_8_8
x271 VDD ctop vcom col_n[8] colon_n[8] net18 net17 VSS row_n[14] adc_array_wafflecap_8_8
x272 VDD ctop vcom col_n[8] colon_n[8] net18 net17 VSS row_n[15] adc_array_wafflecap_8_8
x273 VDD ctop vcom col_n[8] colon_n[8] net18 net17 VSS row_n[16] adc_array_wafflecap_8_8
x274 VDD ctop vcom col_n[8] colon_n[8] net18 net17 VSS row_n[17] adc_array_wafflecap_8_8
x275 VDD ctop vcom col_n[8] colon_n[8] net18 net17 VSS row_n[18] adc_array_wafflecap_8_8
x276 VDD ctop vcom col_n[8] colon_n[8] net18 net17 VSS row_n[19] adc_array_wafflecap_8_8
x277 VDD ctop vcom col_n[8] colon_n[8] net18 net17 VSS row_n[20] adc_array_wafflecap_8_8
x278 VDD ctop vcom col_n[8] colon_n[8] net18 net17 VSS row_n[21] adc_array_wafflecap_8_8
x279 VDD ctop vcom col_n[8] colon_n[8] net18 net17 VSS row_n[22] adc_array_wafflecap_8_8
x280 VDD ctop vcom col_n[8] colon_n[8] net18 net17 VSS row_n[23] adc_array_wafflecap_8_8
x281 VDD ctop vcom col_n[8] colon_n[8] net18 net17 VSS row_n[24] adc_array_wafflecap_8_8
x282 VDD ctop vcom col_n[8] colon_n[8] net18 net17 VSS row_n[25] adc_array_wafflecap_8_8
x283 VDD ctop vcom col_n[8] colon_n[8] net18 net17 VSS row_n[26] adc_array_wafflecap_8_8
x284 VDD ctop vcom col_n[8] colon_n[8] net18 net17 VSS row_n[27] adc_array_wafflecap_8_8
x285 VDD ctop vcom col_n[8] colon_n[8] net18 net17 VSS row_n[28] adc_array_wafflecap_8_8
x286 VDD ctop vcom col_n[8] colon_n[8] net18 net17 VSS row_n[29] adc_array_wafflecap_8_8
x287 VDD ctop vcom col_n[8] colon_n[8] net18 net17 VSS row_n[30] adc_array_wafflecap_8_8
x288 VDD ctop vcom col_n[8] colon_n[8] net18 net17 VSS row_n[31] adc_array_wafflecap_8_8
x289 VDD ctop vcom col_n[9] colon_n[9] net20 net19 VSS row_n[0] adc_array_wafflecap_8_8
x290 VDD ctop vcom col_n[9] colon_n[9] net20 net19 VSS row_n[1] adc_array_wafflecap_8_8
x291 VDD ctop vcom col_n[9] colon_n[9] net20 net19 VSS row_n[2] adc_array_wafflecap_8_8
x292 VDD ctop vcom col_n[9] colon_n[9] net20 net19 VSS row_n[3] adc_array_wafflecap_8_8
x293 VDD ctop vcom col_n[9] colon_n[9] net20 net19 VSS row_n[4] adc_array_wafflecap_8_8
x294 VDD ctop vcom col_n[9] colon_n[9] net20 net19 VSS row_n[5] adc_array_wafflecap_8_8
x295 VDD ctop vcom col_n[9] colon_n[9] net20 net19 VSS row_n[6] adc_array_wafflecap_8_8
x296 VDD ctop vcom col_n[9] colon_n[9] net20 net19 VSS row_n[7] adc_array_wafflecap_8_8
x297 VDD ctop vcom col_n[9] colon_n[9] net20 net19 VSS row_n[8] adc_array_wafflecap_8_8
x298 VDD ctop vcom col_n[9] colon_n[9] net20 net19 VSS row_n[9] adc_array_wafflecap_8_8
x299 VDD ctop vcom col_n[9] colon_n[9] net20 net19 VSS row_n[10] adc_array_wafflecap_8_8
x300 VDD ctop vcom col_n[9] colon_n[9] net20 net19 VSS row_n[11] adc_array_wafflecap_8_8
x301 VDD ctop vcom col_n[9] colon_n[9] net20 net19 VSS row_n[12] adc_array_wafflecap_8_8
x302 VDD ctop vcom col_n[9] colon_n[9] net20 net19 VSS row_n[13] adc_array_wafflecap_8_8
x303 VDD ctop vcom col_n[9] colon_n[9] net20 net19 VSS row_n[14] adc_array_wafflecap_8_8
x304 VDD ctop vcom col_n[9] colon_n[9] net20 net19 VSS row_n[15] adc_array_wafflecap_8_8
x305 VDD ctop vcom col_n[9] colon_n[9] net20 net19 VSS row_n[16] adc_array_wafflecap_8_8
x306 VDD ctop vcom col_n[9] colon_n[9] net20 net19 VSS row_n[17] adc_array_wafflecap_8_8
x307 VDD ctop vcom col_n[9] colon_n[9] net20 net19 VSS row_n[18] adc_array_wafflecap_8_8
x308 VDD ctop vcom col_n[9] colon_n[9] net20 net19 VSS row_n[19] adc_array_wafflecap_8_8
x309 VDD ctop vcom col_n[9] colon_n[9] net20 net19 VSS row_n[20] adc_array_wafflecap_8_8
x310 VDD ctop vcom col_n[9] colon_n[9] net20 net19 VSS row_n[21] adc_array_wafflecap_8_8
x311 VDD ctop vcom col_n[9] colon_n[9] net20 net19 VSS row_n[22] adc_array_wafflecap_8_8
x312 VDD ctop vcom col_n[9] colon_n[9] net20 net19 VSS row_n[23] adc_array_wafflecap_8_8
x313 VDD ctop vcom col_n[9] colon_n[9] net20 net19 VSS row_n[24] adc_array_wafflecap_8_8
x314 VDD ctop vcom col_n[9] colon_n[9] net20 net19 VSS row_n[25] adc_array_wafflecap_8_8
x315 VDD ctop vcom col_n[9] colon_n[9] net20 net19 VSS row_n[26] adc_array_wafflecap_8_8
x316 VDD ctop vcom col_n[9] colon_n[9] net20 net19 VSS row_n[27] adc_array_wafflecap_8_8
x317 VDD ctop vcom col_n[9] colon_n[9] net20 net19 VSS row_n[28] adc_array_wafflecap_8_8
x318 VDD ctop vcom col_n[9] colon_n[9] net20 net19 VSS row_n[29] adc_array_wafflecap_8_8
x319 VDD ctop vcom col_n[9] colon_n[9] net20 net19 VSS row_n[30] adc_array_wafflecap_8_8
x320 VDD ctop vcom col_n[9] colon_n[9] net20 net19 VSS row_n[31] adc_array_wafflecap_8_8
x321 VDD ctop vcom col_n[10] colon_n[10] net22 net21 VSS row_n[0] adc_array_wafflecap_8_8
x322 VDD ctop vcom col_n[10] colon_n[10] net22 net21 VSS row_n[1] adc_array_wafflecap_8_8
x323 VDD ctop vcom col_n[10] colon_n[10] net22 net21 VSS row_n[2] adc_array_wafflecap_8_8
x324 VDD ctop vcom col_n[10] colon_n[10] net22 net21 VSS row_n[3] adc_array_wafflecap_8_8
x325 VDD ctop vcom col_n[10] colon_n[10] net22 net21 VSS row_n[4] adc_array_wafflecap_8_8
x326 VDD ctop vcom col_n[10] colon_n[10] net22 net21 VSS row_n[5] adc_array_wafflecap_8_8
x327 VDD ctop vcom col_n[10] colon_n[10] net22 net21 VSS row_n[6] adc_array_wafflecap_8_8
x328 VDD ctop vcom col_n[10] colon_n[10] net22 net21 VSS row_n[7] adc_array_wafflecap_8_8
x329 VDD ctop vcom col_n[10] colon_n[10] net22 net21 VSS row_n[8] adc_array_wafflecap_8_8
x330 VDD ctop vcom col_n[10] colon_n[10] net22 net21 VSS row_n[9] adc_array_wafflecap_8_8
x331 VDD ctop vcom col_n[10] colon_n[10] net22 net21 VSS row_n[10] adc_array_wafflecap_8_8
x332 VDD ctop vcom col_n[10] colon_n[10] net22 net21 VSS row_n[11] adc_array_wafflecap_8_8
x333 VDD ctop vcom col_n[10] colon_n[10] net22 net21 VSS row_n[12] adc_array_wafflecap_8_8
x334 VDD ctop vcom col_n[10] colon_n[10] net22 net21 VSS row_n[13] adc_array_wafflecap_8_8
x335 VDD ctop vcom col_n[10] colon_n[10] net22 net21 VSS row_n[14] adc_array_wafflecap_8_8
x336 VDD ctop vcom col_n[10] colon_n[10] net22 net21 VSS row_n[15] adc_array_wafflecap_8_8
x337 VDD ctop vcom col_n[10] colon_n[10] net22 net21 VSS row_n[16] adc_array_wafflecap_8_8
x338 VDD ctop vcom col_n[10] colon_n[10] net22 net21 VSS row_n[17] adc_array_wafflecap_8_8
x339 VDD ctop vcom col_n[10] colon_n[10] net22 net21 VSS row_n[18] adc_array_wafflecap_8_8
x340 VDD ctop vcom col_n[10] colon_n[10] net22 net21 VSS row_n[19] adc_array_wafflecap_8_8
x341 VDD ctop vcom col_n[10] colon_n[10] net22 net21 VSS row_n[20] adc_array_wafflecap_8_8
x342 VDD ctop vcom col_n[10] colon_n[10] net22 net21 VSS row_n[21] adc_array_wafflecap_8_8
x343 VDD ctop vcom col_n[10] colon_n[10] net22 net21 VSS row_n[22] adc_array_wafflecap_8_8
x344 VDD ctop vcom col_n[10] colon_n[10] net22 net21 VSS row_n[23] adc_array_wafflecap_8_8
x345 VDD ctop vcom col_n[10] colon_n[10] net22 net21 VSS row_n[24] adc_array_wafflecap_8_8
x346 VDD ctop vcom col_n[10] colon_n[10] net22 net21 VSS row_n[25] adc_array_wafflecap_8_8
x347 VDD ctop vcom col_n[10] colon_n[10] net22 net21 VSS row_n[26] adc_array_wafflecap_8_8
x348 VDD ctop vcom col_n[10] colon_n[10] net22 net21 VSS row_n[27] adc_array_wafflecap_8_8
x349 VDD ctop vcom col_n[10] colon_n[10] net22 net21 VSS row_n[28] adc_array_wafflecap_8_8
x350 VDD ctop vcom col_n[10] colon_n[10] net22 net21 VSS row_n[29] adc_array_wafflecap_8_8
x351 VDD ctop vcom col_n[10] colon_n[10] net22 net21 VSS row_n[30] adc_array_wafflecap_8_8
x352 VDD ctop vcom col_n[10] colon_n[10] net22 net21 VSS row_n[31] adc_array_wafflecap_8_8
x353 VDD ctop vcom col_n[11] colon_n[11] net24 net23 VSS row_n[0] adc_array_wafflecap_8_8
x354 VDD ctop vcom col_n[11] colon_n[11] net24 net23 VSS row_n[1] adc_array_wafflecap_8_8
x355 VDD ctop vcom col_n[11] colon_n[11] net24 net23 VSS row_n[2] adc_array_wafflecap_8_8
x356 VDD ctop vcom col_n[11] colon_n[11] net24 net23 VSS row_n[3] adc_array_wafflecap_8_8
x357 VDD ctop vcom col_n[11] colon_n[11] net24 net23 VSS row_n[4] adc_array_wafflecap_8_8
x358 VDD ctop vcom col_n[11] colon_n[11] net24 net23 VSS row_n[5] adc_array_wafflecap_8_8
x359 VDD ctop vcom col_n[11] colon_n[11] net24 net23 VSS row_n[6] adc_array_wafflecap_8_8
x360 VDD ctop vcom col_n[11] colon_n[11] net24 net23 VSS row_n[7] adc_array_wafflecap_8_8
x361 VDD ctop vcom col_n[11] colon_n[11] net24 net23 VSS row_n[8] adc_array_wafflecap_8_8
x362 VDD ctop vcom col_n[11] colon_n[11] net24 net23 VSS row_n[9] adc_array_wafflecap_8_8
x363 VDD ctop vcom col_n[11] colon_n[11] net24 net23 VSS row_n[10] adc_array_wafflecap_8_8
x364 VDD ctop vcom col_n[11] colon_n[11] net24 net23 VSS row_n[11] adc_array_wafflecap_8_8
x365 VDD ctop vcom col_n[11] colon_n[11] net24 net23 VSS row_n[12] adc_array_wafflecap_8_8
x366 VDD ctop vcom col_n[11] colon_n[11] net24 net23 VSS row_n[13] adc_array_wafflecap_8_8
x367 VDD ctop vcom col_n[11] colon_n[11] net24 net23 VSS row_n[14] adc_array_wafflecap_8_8
x368 VDD ctop vcom col_n[11] colon_n[11] net24 net23 VSS row_n[15] adc_array_wafflecap_8_8
x369 VDD ctop vcom col_n[11] colon_n[11] net24 net23 VSS row_n[16] adc_array_wafflecap_8_8
x370 VDD ctop vcom col_n[11] colon_n[11] net24 net23 VSS row_n[17] adc_array_wafflecap_8_8
x371 VDD ctop vcom col_n[11] colon_n[11] net24 net23 VSS row_n[18] adc_array_wafflecap_8_8
x372 VDD ctop vcom col_n[11] colon_n[11] net24 net23 VSS row_n[19] adc_array_wafflecap_8_8
x373 VDD ctop vcom col_n[11] colon_n[11] net24 net23 VSS row_n[20] adc_array_wafflecap_8_8
x374 VDD ctop vcom col_n[11] colon_n[11] net24 net23 VSS row_n[21] adc_array_wafflecap_8_8
x375 VDD ctop vcom col_n[11] colon_n[11] net24 net23 VSS row_n[22] adc_array_wafflecap_8_8
x376 VDD ctop vcom col_n[11] colon_n[11] net24 net23 VSS row_n[23] adc_array_wafflecap_8_8
x377 VDD ctop vcom col_n[11] colon_n[11] net24 net23 VSS row_n[24] adc_array_wafflecap_8_8
x378 VDD ctop vcom col_n[11] colon_n[11] net24 net23 VSS row_n[25] adc_array_wafflecap_8_8
x379 VDD ctop vcom col_n[11] colon_n[11] net24 net23 VSS row_n[26] adc_array_wafflecap_8_8
x380 VDD ctop vcom col_n[11] colon_n[11] net24 net23 VSS row_n[27] adc_array_wafflecap_8_8
x381 VDD ctop vcom col_n[11] colon_n[11] net24 net23 VSS row_n[28] adc_array_wafflecap_8_8
x382 VDD ctop vcom col_n[11] colon_n[11] net24 net23 VSS row_n[29] adc_array_wafflecap_8_8
x383 VDD ctop vcom col_n[11] colon_n[11] net24 net23 VSS row_n[30] adc_array_wafflecap_8_8
x384 VDD ctop vcom col_n[11] colon_n[11] net24 net23 VSS row_n[31] adc_array_wafflecap_8_8
x385 VDD ctop vcom col_n[12] colon_n[12] net26 net25 VSS row_n[0] adc_array_wafflecap_8_8
x386 VDD ctop vcom col_n[12] colon_n[12] net26 net25 VSS row_n[1] adc_array_wafflecap_8_8
x387 VDD ctop vcom col_n[12] colon_n[12] net26 net25 VSS row_n[2] adc_array_wafflecap_8_8
x388 VDD ctop vcom col_n[12] colon_n[12] net26 net25 VSS row_n[3] adc_array_wafflecap_8_8
x389 VDD ctop vcom col_n[12] colon_n[12] net26 net25 VSS row_n[4] adc_array_wafflecap_8_8
x390 VDD ctop vcom col_n[12] colon_n[12] net26 net25 VSS row_n[5] adc_array_wafflecap_8_8
x391 VDD ctop vcom col_n[12] colon_n[12] net26 net25 VSS row_n[6] adc_array_wafflecap_8_8
x392 VDD ctop vcom col_n[12] colon_n[12] net26 net25 VSS row_n[7] adc_array_wafflecap_8_8
x393 VDD ctop vcom col_n[12] colon_n[12] net26 net25 VSS row_n[8] adc_array_wafflecap_8_8
x394 VDD ctop vcom col_n[12] colon_n[12] net26 net25 VSS row_n[9] adc_array_wafflecap_8_8
x395 VDD ctop vcom col_n[12] colon_n[12] net26 net25 VSS row_n[10] adc_array_wafflecap_8_8
x396 VDD ctop vcom col_n[12] colon_n[12] net26 net25 VSS row_n[11] adc_array_wafflecap_8_8
x397 VDD ctop vcom col_n[12] colon_n[12] net26 net25 VSS row_n[12] adc_array_wafflecap_8_8
x398 VDD ctop vcom col_n[12] colon_n[12] net26 net25 VSS row_n[13] adc_array_wafflecap_8_8
x399 VDD ctop vcom col_n[12] colon_n[12] net26 net25 VSS row_n[14] adc_array_wafflecap_8_8
x400 VDD ctop vcom col_n[12] colon_n[12] net26 net25 VSS row_n[15] adc_array_wafflecap_8_8
x401 VDD ctop vcom col_n[12] colon_n[12] net26 net25 VSS row_n[16] adc_array_wafflecap_8_8
x402 VDD ctop vcom col_n[12] colon_n[12] net26 net25 VSS row_n[17] adc_array_wafflecap_8_8
x403 VDD ctop vcom col_n[12] colon_n[12] net26 net25 VSS row_n[18] adc_array_wafflecap_8_8
x404 VDD ctop vcom col_n[12] colon_n[12] net26 net25 VSS row_n[19] adc_array_wafflecap_8_8
x405 VDD ctop vcom col_n[12] colon_n[12] net26 net25 VSS row_n[20] adc_array_wafflecap_8_8
x406 VDD ctop vcom col_n[12] colon_n[12] net26 net25 VSS row_n[21] adc_array_wafflecap_8_8
x407 VDD ctop vcom col_n[12] colon_n[12] net26 net25 VSS row_n[22] adc_array_wafflecap_8_8
x408 VDD ctop vcom col_n[12] colon_n[12] net26 net25 VSS row_n[23] adc_array_wafflecap_8_8
x409 VDD ctop vcom col_n[12] colon_n[12] net26 net25 VSS row_n[24] adc_array_wafflecap_8_8
x410 VDD ctop vcom col_n[12] colon_n[12] net26 net25 VSS row_n[25] adc_array_wafflecap_8_8
x411 VDD ctop vcom col_n[12] colon_n[12] net26 net25 VSS row_n[26] adc_array_wafflecap_8_8
x412 VDD ctop vcom col_n[12] colon_n[12] net26 net25 VSS row_n[27] adc_array_wafflecap_8_8
x413 VDD ctop vcom col_n[12] colon_n[12] net26 net25 VSS row_n[28] adc_array_wafflecap_8_8
x414 VDD ctop vcom col_n[12] colon_n[12] net26 net25 VSS row_n[29] adc_array_wafflecap_8_8
x415 VDD ctop vcom col_n[12] colon_n[12] net26 net25 VSS row_n[30] adc_array_wafflecap_8_8
x416 VDD ctop vcom col_n[12] colon_n[12] net26 net25 VSS row_n[31] adc_array_wafflecap_8_8
x417 VDD ctop vcom col_n[13] colon_n[13] net28 net27 VSS row_n[0] adc_array_wafflecap_8_8
x418 VDD ctop vcom col_n[13] colon_n[13] net28 net27 VSS row_n[1] adc_array_wafflecap_8_8
x419 VDD ctop vcom col_n[13] colon_n[13] net28 net27 VSS row_n[2] adc_array_wafflecap_8_8
x420 VDD ctop vcom col_n[13] colon_n[13] net28 net27 VSS row_n[3] adc_array_wafflecap_8_8
x421 VDD ctop vcom col_n[13] colon_n[13] net28 net27 VSS row_n[4] adc_array_wafflecap_8_8
x422 VDD ctop vcom col_n[13] colon_n[13] net28 net27 VSS row_n[5] adc_array_wafflecap_8_8
x423 VDD ctop vcom col_n[13] colon_n[13] net28 net27 VSS row_n[6] adc_array_wafflecap_8_8
x424 VDD ctop vcom col_n[13] colon_n[13] net28 net27 VSS row_n[7] adc_array_wafflecap_8_8
x425 VDD ctop vcom col_n[13] colon_n[13] net28 net27 VSS row_n[8] adc_array_wafflecap_8_8
x426 VDD ctop vcom col_n[13] colon_n[13] net28 net27 VSS row_n[9] adc_array_wafflecap_8_8
x427 VDD ctop vcom col_n[13] colon_n[13] net28 net27 VSS row_n[10] adc_array_wafflecap_8_8
x428 VDD ctop vcom col_n[13] colon_n[13] net28 net27 VSS row_n[11] adc_array_wafflecap_8_8
x429 VDD ctop vcom col_n[13] colon_n[13] net28 net27 VSS row_n[12] adc_array_wafflecap_8_8
x430 VDD ctop vcom col_n[13] colon_n[13] net28 net27 VSS row_n[13] adc_array_wafflecap_8_8
x431 VDD ctop vcom col_n[13] colon_n[13] net28 net27 VSS row_n[14] adc_array_wafflecap_8_8
x432 VDD ctop vcom col_n[13] colon_n[13] net28 net27 VSS row_n[15] adc_array_wafflecap_8_8
x433 VDD ctop vcom col_n[13] colon_n[13] net28 net27 VSS row_n[16] adc_array_wafflecap_8_8
x434 VDD ctop vcom col_n[13] colon_n[13] net28 net27 VSS row_n[17] adc_array_wafflecap_8_8
x435 VDD ctop vcom col_n[13] colon_n[13] net28 net27 VSS row_n[18] adc_array_wafflecap_8_8
x436 VDD ctop vcom col_n[13] colon_n[13] net28 net27 VSS row_n[19] adc_array_wafflecap_8_8
x437 VDD ctop vcom col_n[13] colon_n[13] net28 net27 VSS row_n[20] adc_array_wafflecap_8_8
x438 VDD ctop vcom col_n[13] colon_n[13] net28 net27 VSS row_n[21] adc_array_wafflecap_8_8
x439 VDD ctop vcom col_n[13] colon_n[13] net28 net27 VSS row_n[22] adc_array_wafflecap_8_8
x440 VDD ctop vcom col_n[13] colon_n[13] net28 net27 VSS row_n[23] adc_array_wafflecap_8_8
x441 VDD ctop vcom col_n[13] colon_n[13] net28 net27 VSS row_n[24] adc_array_wafflecap_8_8
x442 VDD ctop vcom col_n[13] colon_n[13] net28 net27 VSS row_n[25] adc_array_wafflecap_8_8
x443 VDD ctop vcom col_n[13] colon_n[13] net28 net27 VSS row_n[26] adc_array_wafflecap_8_8
x444 VDD ctop vcom col_n[13] colon_n[13] net28 net27 VSS row_n[27] adc_array_wafflecap_8_8
x445 VDD ctop vcom col_n[13] colon_n[13] net28 net27 VSS row_n[28] adc_array_wafflecap_8_8
x446 VDD ctop vcom col_n[13] colon_n[13] net28 net27 VSS row_n[29] adc_array_wafflecap_8_8
x447 VDD ctop vcom col_n[13] colon_n[13] net28 net27 VSS row_n[30] adc_array_wafflecap_8_8
x448 VDD ctop vcom col_n[13] colon_n[13] net28 net27 VSS row_n[31] adc_array_wafflecap_8_8
x449 VDD ctop vcom col_n[14] colon_n[14] net30 net29 VSS row_n[0] adc_array_wafflecap_8_8
x450 VDD ctop vcom col_n[14] colon_n[14] net30 net29 VSS row_n[1] adc_array_wafflecap_8_8
x451 VDD ctop vcom col_n[14] colon_n[14] net30 net29 VSS row_n[2] adc_array_wafflecap_8_8
x452 VDD ctop vcom col_n[14] colon_n[14] net30 net29 VSS row_n[3] adc_array_wafflecap_8_8
x453 VDD ctop vcom col_n[14] colon_n[14] net30 net29 VSS row_n[4] adc_array_wafflecap_8_8
x454 VDD ctop vcom col_n[14] colon_n[14] net30 net29 VSS row_n[5] adc_array_wafflecap_8_8
x455 VDD ctop vcom col_n[14] colon_n[14] net30 net29 VSS row_n[6] adc_array_wafflecap_8_8
x456 VDD ctop vcom col_n[14] colon_n[14] net30 net29 VSS row_n[7] adc_array_wafflecap_8_8
x457 VDD ctop vcom col_n[14] colon_n[14] net30 net29 VSS row_n[8] adc_array_wafflecap_8_8
x458 VDD ctop vcom col_n[14] colon_n[14] net30 net29 VSS row_n[9] adc_array_wafflecap_8_8
x459 VDD ctop vcom col_n[14] colon_n[14] net30 net29 VSS row_n[10] adc_array_wafflecap_8_8
x460 VDD ctop vcom col_n[14] colon_n[14] net30 net29 VSS row_n[11] adc_array_wafflecap_8_8
x461 VDD ctop vcom col_n[14] colon_n[14] net30 net29 VSS row_n[12] adc_array_wafflecap_8_8
x462 VDD ctop vcom col_n[14] colon_n[14] net30 net29 VSS row_n[13] adc_array_wafflecap_8_8
x463 VDD ctop vcom col_n[14] colon_n[14] net30 net29 VSS row_n[14] adc_array_wafflecap_8_8
x464 VDD ctop vcom col_n[14] colon_n[14] net30 net29 VSS row_n[15] adc_array_wafflecap_8_8
x465 VDD ctop vcom col_n[14] colon_n[14] net30 net29 VSS row_n[16] adc_array_wafflecap_8_8
x466 VDD ctop vcom col_n[14] colon_n[14] net30 net29 VSS row_n[17] adc_array_wafflecap_8_8
x467 VDD ctop vcom col_n[14] colon_n[14] net30 net29 VSS row_n[18] adc_array_wafflecap_8_8
x468 VDD ctop vcom col_n[14] colon_n[14] net30 net29 VSS row_n[19] adc_array_wafflecap_8_8
x469 VDD ctop vcom col_n[14] colon_n[14] net30 net29 VSS row_n[20] adc_array_wafflecap_8_8
x470 VDD ctop vcom col_n[14] colon_n[14] net30 net29 VSS row_n[21] adc_array_wafflecap_8_8
x471 VDD ctop vcom col_n[14] colon_n[14] net30 net29 VSS row_n[22] adc_array_wafflecap_8_8
x472 VDD ctop vcom col_n[14] colon_n[14] net30 net29 VSS row_n[23] adc_array_wafflecap_8_8
x473 VDD ctop vcom col_n[14] colon_n[14] net30 net29 VSS row_n[24] adc_array_wafflecap_8_8
x474 VDD ctop vcom col_n[14] colon_n[14] net30 net29 VSS row_n[25] adc_array_wafflecap_8_8
x475 VDD ctop vcom col_n[14] colon_n[14] net30 net29 VSS row_n[26] adc_array_wafflecap_8_8
x476 VDD ctop vcom col_n[14] colon_n[14] net30 net29 VSS row_n[27] adc_array_wafflecap_8_8
x477 VDD ctop vcom col_n[14] colon_n[14] net30 net29 VSS row_n[28] adc_array_wafflecap_8_8
x478 VDD ctop vcom col_n[14] colon_n[14] net30 net29 VSS row_n[29] adc_array_wafflecap_8_8
x479 VDD ctop vcom col_n[14] colon_n[14] net30 net29 VSS row_n[30] adc_array_wafflecap_8_8
x480 VDD ctop vcom col_n[14] colon_n[14] net30 net29 VSS row_n[31] adc_array_wafflecap_8_8
x481 VDD ctop vcom col_n[15] colon_n[15] net32 net31 VSS row_n[0] adc_array_wafflecap_8_8
x482 VDD ctop vcom col_n[15] colon_n[15] net32 net31 VSS row_n[1] adc_array_wafflecap_8_8
x483 VDD ctop vcom col_n[15] colon_n[15] net32 net31 VSS row_n[2] adc_array_wafflecap_8_8
x484 VDD ctop vcom col_n[15] colon_n[15] net32 net31 VSS row_n[3] adc_array_wafflecap_8_8
x485 VDD ctop vcom col_n[15] colon_n[15] net32 net31 VSS row_n[4] adc_array_wafflecap_8_8
x486 VDD ctop vcom col_n[15] colon_n[15] net32 net31 VSS row_n[5] adc_array_wafflecap_8_8
x487 VDD ctop vcom col_n[15] colon_n[15] net32 net31 VSS row_n[6] adc_array_wafflecap_8_8
x488 VDD ctop vcom col_n[15] colon_n[15] net32 net31 VSS row_n[7] adc_array_wafflecap_8_8
x489 VDD ctop vcom col_n[15] colon_n[15] net32 net31 VSS row_n[8] adc_array_wafflecap_8_8
x490 VDD ctop vcom col_n[15] colon_n[15] net32 net31 VSS row_n[9] adc_array_wafflecap_8_8
x491 VDD ctop vcom col_n[15] colon_n[15] net32 net31 VSS row_n[10] adc_array_wafflecap_8_8
x492 VDD ctop vcom col_n[15] colon_n[15] net32 net31 VSS row_n[11] adc_array_wafflecap_8_8
x493 VDD ctop vcom col_n[15] colon_n[15] net32 net31 VSS row_n[12] adc_array_wafflecap_8_8
x494 VDD ctop vcom col_n[15] colon_n[15] net32 net31 VSS row_n[13] adc_array_wafflecap_8_8
x495 VDD ctop vcom col_n[15] colon_n[15] net32 net31 VSS row_n[14] adc_array_wafflecap_8_8
x496 VDD ctop vcom col_n[15] colon_n[15] net32 net31 VSS row_n[15] adc_array_wafflecap_8_8
x497 VDD ctop vcom col_n[15] colon_n[15] net32 net31 VSS row_n[16] adc_array_wafflecap_8_8
x498 VDD ctop vcom col_n[15] colon_n[15] net32 net31 VSS row_n[17] adc_array_wafflecap_8_8
x499 VDD ctop vcom col_n[15] colon_n[15] net32 net31 VSS row_n[18] adc_array_wafflecap_8_8
x500 VDD ctop vcom col_n[15] colon_n[15] net32 net31 VSS row_n[19] adc_array_wafflecap_8_8
x501 VDD ctop vcom col_n[15] colon_n[15] net32 net31 VSS row_n[20] adc_array_wafflecap_8_8
x502 VDD ctop vcom col_n[15] colon_n[15] net32 net31 VSS row_n[21] adc_array_wafflecap_8_8
x503 VDD ctop vcom col_n[15] colon_n[15] net32 net31 VSS row_n[22] adc_array_wafflecap_8_8
x504 VDD ctop vcom col_n[15] colon_n[15] net32 net31 VSS row_n[23] adc_array_wafflecap_8_8
x505 VDD ctop vcom col_n[15] colon_n[15] net32 net31 VSS row_n[24] adc_array_wafflecap_8_8
x506 VDD ctop vcom col_n[15] colon_n[15] net32 net31 VSS row_n[25] adc_array_wafflecap_8_8
x507 VDD ctop vcom col_n[15] colon_n[15] net32 net31 VSS row_n[26] adc_array_wafflecap_8_8
x508 VDD ctop vcom col_n[15] colon_n[15] net32 net31 VSS row_n[27] adc_array_wafflecap_8_8
x509 VDD ctop vcom col_n[15] colon_n[15] net32 net31 VSS row_n[28] adc_array_wafflecap_8_8
x510 VDD ctop vcom col_n[15] colon_n[15] net32 net31 VSS row_n[29] adc_array_wafflecap_8_8
x511 VDD ctop vcom col_n[15] colon_n[15] net32 net31 VSS row_n[30] adc_array_wafflecap_8_8
x512 VDD ctop vcom col_n[15] colon_n[15] net32 net31 VSS row_n[31] adc_array_wafflecap_8_8
x1025 VDD ctop vcom col_n[0] colon_n[0] sample_n sample VSS VDD net2 net1 adc_array_wafflecap_8_Drv
x1026 VDD ctop vcom col_n[1] colon_n[1] sample_n sample VSS VDD net4 net3 adc_array_wafflecap_8_Drv
x1027 VDD ctop vcom col_n[2] colon_n[2] sample_n sample VSS VDD net6 net5 adc_array_wafflecap_8_Drv
x1028 VDD ctop vcom col_n[3] colon_n[3] sample_n sample VSS VDD net8 net7 adc_array_wafflecap_8_Drv
x1029 VDD ctop vcom col_n[4] colon_n[4] sample_n sample VSS VDD net10 net9 adc_array_wafflecap_8_Drv
x1030 VDD ctop vcom col_n[5] colon_n[5] sample_n sample VSS VDD net12 net11
+ adc_array_wafflecap_8_Drv
x1031 VDD ctop vcom col_n[6] colon_n[6] sample_n sample VSS VDD net14 net13
+ adc_array_wafflecap_8_Drv
x1032 VDD ctop vcom col_n[7] colon_n[7] sample_n sample VSS VDD net16 net15
+ adc_array_wafflecap_8_Drv
x1033 VDD ctop vcom col_n[8] colon_n[8] sample_n sample VSS VDD net18 net17
+ adc_array_wafflecap_8_Drv
x1034 VDD ctop vcom col_n[9] colon_n[9] sample_n sample VSS VDD net20 net19
+ adc_array_wafflecap_8_Drv
x1035 VDD ctop vcom col_n[10] colon_n[10] sample_n sample VSS VDD net22 net21
+ adc_array_wafflecap_8_Drv
x1036 VDD ctop vcom col_n[11] colon_n[11] sample_n sample VSS VDD net24 net23
+ adc_array_wafflecap_8_Drv
x1037 VDD ctop vcom col_n[12] colon_n[12] sample_n sample VSS VDD net26 net25
+ adc_array_wafflecap_8_Drv
x1038 VDD ctop vcom col_n[13] colon_n[13] sample_n sample VSS VDD net28 net27
+ adc_array_wafflecap_8_Drv
x1039 VDD ctop vcom col_n[14] colon_n[14] sample_n sample VSS VDD net30 net29
+ adc_array_wafflecap_8_Drv
x1040 VDD ctop vcom col_n[15] colon_n[15] sample_n sample VSS VDD net32 net31
+ adc_array_wafflecap_8_Drv
x1057 VDD ctop vcom VSS VSS VDD VSS VSS VDD adc_array_wafflecap_8_Dummy
x1058 VDD ctop vcom VSS VSS VDD VSS VSS row_n[0] adc_array_wafflecap_8_Dummy
x1059 VDD ctop vcom VSS VSS VDD VSS VSS row_n[1] adc_array_wafflecap_8_Dummy
x1061 VDD ctop vcom VSS VSS VDD VSS VSS row_n[3] adc_array_wafflecap_8_Dummy
x1062 VDD ctop vcom VSS VSS VDD VSS VSS row_n[4] adc_array_wafflecap_8_Dummy
x1063 VDD ctop vcom VSS VSS VDD VSS VSS row_n[5] adc_array_wafflecap_8_Dummy
x1064 VDD ctop vcom VSS VSS VDD VSS VSS row_n[6] adc_array_wafflecap_8_Dummy
x1065 VDD ctop vcom VSS VSS VDD VSS VSS row_n[7] adc_array_wafflecap_8_Dummy
x1067 VDD ctop vcom VSS VSS VDD VSS VSS row_n[9] adc_array_wafflecap_8_Dummy
x1069 VDD ctop vcom VSS VSS VDD VSS VSS row_n[11] adc_array_wafflecap_8_Dummy
x1071 VDD ctop vcom VSS VSS VDD VSS VSS row_n[13] adc_array_wafflecap_8_Dummy
x1072 VDD ctop vcom VSS VSS VDD VSS VSS row_n[14] adc_array_wafflecap_8_Dummy
x1073 VDD ctop vcom VSS VSS VDD VSS VSS row_n[15] adc_array_wafflecap_8_Dummy
x1075 VDD ctop vcom VSS VSS VDD VSS VSS row_n[17] adc_array_wafflecap_8_Dummy
x1077 VDD ctop vcom VSS VSS VDD VSS VSS row_n[19] adc_array_wafflecap_8_Dummy
x1078 VDD ctop vcom VSS VSS VDD VSS VSS row_n[20] adc_array_wafflecap_8_Dummy
x1079 VDD ctop vcom VSS VSS VDD VSS VSS row_n[21] adc_array_wafflecap_8_Dummy
x1080 VDD ctop vcom VSS VSS VDD VSS VSS row_n[22] adc_array_wafflecap_8_Dummy
x1081 VDD ctop vcom VSS VSS VDD VSS VSS row_n[23] adc_array_wafflecap_8_Dummy
x1083 VDD ctop vcom VSS VSS VDD VSS VSS row_n[25] adc_array_wafflecap_8_Dummy
x1085 VDD ctop vcom VSS VSS VDD VSS VSS row_n[12] adc_array_wafflecap_8_Dummy
x1086 VDD ctop vcom VSS VSS VDD VSS VSS row_n[28] adc_array_wafflecap_8_Dummy
x1087 VDD ctop vcom VSS VSS VDD VSS VSS row_n[29] adc_array_wafflecap_8_Dummy
x1088 VDD ctop vcom VSS VSS VDD VSS VSS row_n[30] adc_array_wafflecap_8_Dummy
x1089 VDD ctop vcom VSS VSS VDD VSS VSS row_n[27] adc_array_wafflecap_8_Dummy
x1090 VDD ctop vcom VSS VSS VDD VSS VSS VDD adc_array_wafflecap_8_Dummy
x1091 VDD ctop vcom VDD VDD VDD VSS VSS VDD adc_array_wafflecap_8_Dummy
x1092 VDD ctop vcom VDD VDD VDD VSS VSS row_n[0] adc_array_wafflecap_8_Dummy
x1093 VDD ctop vcom VDD VDD VDD VSS VSS row_n[1] adc_array_wafflecap_8_Dummy
x1094 VDD ctop vcom VDD VDD VDD VSS VSS row_n[2] adc_array_wafflecap_8_Dummy
x1095 VDD ctop vcom VDD VDD VDD VSS VSS row_n[3] adc_array_wafflecap_8_Dummy
x1096 VDD ctop vcom VDD VDD VDD VSS VSS row_n[4] adc_array_wafflecap_8_Dummy
x1097 VDD ctop vcom VDD VDD VDD VSS VSS row_n[5] adc_array_wafflecap_8_Dummy
x1098 VDD ctop vcom VDD VDD VDD VSS VSS row_n[6] adc_array_wafflecap_8_Dummy
x1099 VDD ctop vcom VDD VDD VDD VSS VSS row_n[7] adc_array_wafflecap_8_Dummy
x1100 VDD ctop vcom VDD VDD VDD VSS VSS row_n[8] adc_array_wafflecap_8_Dummy
x1101 VDD ctop vcom VDD VDD VDD VSS VSS row_n[9] adc_array_wafflecap_8_Dummy
x1102 VDD ctop vcom VDD VDD VDD VSS VSS row_n[10] adc_array_wafflecap_8_Dummy
x1103 VDD ctop vcom VDD VDD VDD VSS VSS row_n[11] adc_array_wafflecap_8_Dummy
x1104 VDD ctop vcom VDD VDD VDD VSS VSS row_n[12] adc_array_wafflecap_8_Dummy
x1105 VDD ctop vcom VDD VDD VDD VSS VSS row_n[13] adc_array_wafflecap_8_Dummy
x1106 VDD ctop vcom VDD VDD VDD VSS VSS row_n[14] adc_array_wafflecap_8_Dummy
x1107 VDD ctop vcom VDD VDD VDD VSS VSS row_n[15] adc_array_wafflecap_8_Dummy
x1108 VDD ctop vcom VDD VDD VDD VSS VSS row_n[16] adc_array_wafflecap_8_Dummy
x1109 VDD ctop vcom VDD VDD VDD VSS VSS row_n[17] adc_array_wafflecap_8_Dummy
x1110 VDD ctop vcom VDD VDD VDD VSS VSS row_n[18] adc_array_wafflecap_8_Dummy
x1111 VDD ctop vcom VDD VDD VDD VSS VSS row_n[19] adc_array_wafflecap_8_Dummy
x1112 VDD ctop vcom VDD VDD VDD VSS VSS row_n[20] adc_array_wafflecap_8_Dummy
x1113 VDD ctop vcom VDD VDD VDD VSS VSS row_n[21] adc_array_wafflecap_8_Dummy
x1114 VDD ctop vcom VDD VDD VDD VSS VSS row_n[22] adc_array_wafflecap_8_Dummy
x1115 VDD ctop vcom VDD VDD VDD VSS VSS row_n[23] adc_array_wafflecap_8_Dummy
x1116 VDD ctop vcom VDD VDD VDD VSS VSS row_n[24] adc_array_wafflecap_8_Dummy
x1117 VDD ctop vcom VDD VDD VDD VSS VSS row_n[25] adc_array_wafflecap_8_Dummy
x1118 VDD ctop vcom VDD VDD VDD VSS VSS row_n[26] adc_array_wafflecap_8_Dummy
x1119 VDD ctop vcom VDD VDD VDD VSS VSS row_n[27] adc_array_wafflecap_8_Dummy
x1120 VDD ctop vcom VDD VDD VDD VSS VSS row_n[28] adc_array_wafflecap_8_Dummy
x1121 VDD ctop vcom VDD VDD VDD VSS VSS row_n[29] adc_array_wafflecap_8_Dummy
x1122 VDD ctop vcom VDD VDD VDD VSS VSS row_n[30] adc_array_wafflecap_8_Dummy
x1123 VDD ctop vcom VDD VDD VDD VSS VSS row_n[31] adc_array_wafflecap_8_Dummy
x1124 VDD ctop vcom VDD VDD VDD VSS VSS VDD adc_array_wafflecap_8_Dummy
x1125 VDD ctop vcom col_n[0] colon_n[0] net2 net1 VSS VDD adc_array_wafflecap_8_Dummy
x1126 VDD ctop vcom col_n[1] colon_n[1] net4 net3 VSS VDD adc_array_wafflecap_8_Dummy
x1127 VDD ctop vcom col_n[2] colon_n[2] net6 net5 VSS VDD adc_array_wafflecap_8_Dummy
x1128 VDD ctop vcom col_n[3] colon_n[3] net8 net7 VSS VDD adc_array_wafflecap_8_Dummy
x1129 VDD ctop vcom col_n[4] colon_n[4] net10 net9 VSS VDD adc_array_wafflecap_8_Dummy
x1130 VDD ctop vcom col_n[5] colon_n[5] net12 net11 VSS VDD adc_array_wafflecap_8_Dummy
x1131 VDD ctop vcom col_n[6] colon_n[6] net14 net13 VSS VDD adc_array_wafflecap_8_Dummy
x1132 VDD ctop vcom col_n[7] colon_n[7] net16 net15 VSS VDD adc_array_wafflecap_8_Dummy
x1133 VDD ctop vcom col_n[8] colon_n[8] net18 net17 VSS VDD adc_array_wafflecap_8_Dummy
x1134 VDD ctop vcom col_n[9] colon_n[9] net20 net19 VSS VDD adc_array_wafflecap_8_Dummy
x1135 VDD ctop vcom col_n[10] colon_n[10] net22 net21 VSS VDD adc_array_wafflecap_8_Dummy
x1136 VDD ctop vcom col_n[11] colon_n[11] net24 net23 VSS VDD adc_array_wafflecap_8_Dummy
x1137 VDD ctop vcom col_n[12] colon_n[12] net26 net25 VSS VDD adc_array_wafflecap_8_Dummy
x1138 VDD ctop vcom col_n[13] colon_n[13] net28 net27 VSS VDD adc_array_wafflecap_8_Dummy
x1139 VDD ctop vcom col_n[14] colon_n[14] net30 net29 VSS VDD adc_array_wafflecap_8_Dummy
x1140 VDD ctop vcom col_n[15] colon_n[15] net32 net31 VSS VDD adc_array_wafflecap_8_Dummy
x513 VDD ctop vcom VSS VSS VDD VSS VSS row_n[2] adc_array_wafflecap_8_Dummy
x514 VDD ctop vcom VSS VSS VDD VSS VSS row_n[10] adc_array_wafflecap_8_Dummy
x515 VDD ctop vcom VSS VSS VDD VSS VSS row_n[18] adc_array_wafflecap_8_Dummy
x516 VDD ctop vcom VSS VSS VDD VSS VSS row_n[26] adc_array_wafflecap_8_Dummy
x517 VDD ctop vcom VSS VSS VDD VSS VSS row_n[8] en_n_bit[2] adc_array_wafflecap_8_4
x518 VDD ctop vcom VSS VSS VDD VSS VSS row_n[16] en_n_bit[1] adc_array_wafflecap_8_2
x519 VDD ctop vcom VSS VSS VDD VSS VSS row_n[24] en_n_bit[0] adc_array_wafflecap_8_1
x520 VDD ctop vcom VSS VSS VDD VSS VSS row_n[31] sw analog_in sw_n adc_array_wafflecap_8_Gate
.ends

* expanding   symbol:  /foss/designs/SKY130_SAR-ADC/xschem/adc_array_cap/adc_array_wafflecap_8_8.sym
*+ # of pins=9
** sym_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_array_cap/adc_array_wafflecap_8_8.sym
** sch_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_array_cap/adc_array_wafflecap_8_8.sch
.subckt adc_array_wafflecap_8_8  VDD ctop vcom col_n colon_n sample_n sample VSS row_n
*.PININFO vcom:B VDD:B ctop:B VSS:B row_n:I col_n:I colon_n:I sample_n:I sample:I
x1 VDD row_n cbot col_n colon_n sample_n vcom sample VSS adc_array_circuit_150n_8
.ends


* expanding   symbol:
*+  /foss/designs/SKY130_SAR-ADC/xschem/adc_array_cap/adc_array_wafflecap_8_Drv.sym # of pins=11
** sym_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_array_cap/adc_array_wafflecap_8_Drv.sym
** sch_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_array_cap/adc_array_wafflecap_8_Drv.sch
.subckt adc_array_wafflecap_8_Drv  VDD ctop vcom col_n colon_n sample_n_i sample_i VSS row_n
+ sample_n_o sample_o
*.PININFO sample_n_i:I sample_i:I vcom:B VDD:B ctop:B VSS:B sample_n_o:O sample_o:O row_n:I col_n:I
*+ colon_n:I
x1 VDD row_n col_n colon_n sample_n_i vcom sample_i VSS sample_n_o sample_o
+ adc_array_circuit_150n_Drv
.ends


* expanding   symbol:
*+  /foss/designs/SKY130_SAR-ADC/xschem/adc_array_cap/adc_array_wafflecap_8_Dummy.sym # of pins=9
** sym_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_array_cap/adc_array_wafflecap_8_Dummy.sym
** sch_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_array_cap/adc_array_wafflecap_8_Dummy.sch
.subckt adc_array_wafflecap_8_Dummy  VDD ctop vcom col_n colon_n sample_n sample VSS row_n
*.PININFO vcom:B VDD:B ctop:B VSS:B row_n:I col_n:I colon_n:I sample_n:I sample:I
x1 VDD row_n cbot col_n colon_n sample_n vcom sample VSS adc_array_circuit_150n_8
.ends


* expanding   symbol:  /foss/designs/SKY130_SAR-ADC/xschem/adc_array_cap/adc_array_wafflecap_8_4.sym
*+ # of pins=10
** sym_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_array_cap/adc_array_wafflecap_8_4.sym
** sch_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_array_cap/adc_array_wafflecap_8_4.sch
.subckt adc_array_wafflecap_8_4  VDD ctop vcom col_n colon_n sample_n sample VSS row_n en_n
*.PININFO vcom:B VDD:B ctop:B VSS:B en_n:I row_n:I col_n:I colon_n:I sample_n:I sample:I
x1 VDD row_n cbot col_n colon_n sample_n vcom sample VSS en_n adc_array_circuit_150n_4
.ends


* expanding   symbol:  /foss/designs/SKY130_SAR-ADC/xschem/adc_array_cap/adc_array_wafflecap_8_2.sym
*+ # of pins=10
** sym_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_array_cap/adc_array_wafflecap_8_2.sym
** sch_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_array_cap/adc_array_wafflecap_8_2.sch
.subckt adc_array_wafflecap_8_2  VDD ctop vcom col_n colon_n sample_n sample VSS row_n en_n
*.PININFO vcom:B VDD:B ctop:B VSS:B en_n:I row_n:I col_n:I colon_n:I sample_n:I sample:I
x1 VDD row_n cbot col_n colon_n sample_n vcom sample VSS en_n adc_array_circuit_150n_2
.ends


* expanding   symbol:  /foss/designs/SKY130_SAR-ADC/xschem/adc_array_cap/adc_array_wafflecap_8_1.sym
*+ # of pins=10
** sym_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_array_cap/adc_array_wafflecap_8_1.sym
** sch_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_array_cap/adc_array_wafflecap_8_1.sch
.subckt adc_array_wafflecap_8_1  VDD ctop vcom col_n colon_n sample_n sample VSS row_n en_n
*.PININFO vcom:B VDD:B ctop:B VSS:B en_n:I row_n:I col_n:I colon_n:I sample_n:I sample:I
x1 VDD row_n cbot col_n colon_n sample_n vcom sample VSS en_n adc_array_circuit_150n_1
.ends


* expanding   symbol:
*+  /foss/designs/SKY130_SAR-ADC/xschem/adc_array_cap/adc_array_wafflecap_8_Gate.sym # of pins=12
** sym_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_array_cap/adc_array_wafflecap_8_Gate.sym
** sch_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_array_cap/adc_array_wafflecap_8_Gate.sch
.subckt adc_array_wafflecap_8_Gate  VDD ctop vcom col_n colon_n sample_n sample VSS row_n sw in sw_n
*.PININFO vcom:B VDD:B ctop:B VSS:B row_n:I col_n:I colon_n:I sample_n:I sample:I in:B sw:I sw_n:I
x1 VDD row_n col_n colon_n sample_n vcom sample VSS ctop in sw_n sw adc_array_circuit_150n_gate
.ends


* expanding   symbol:
*+  /foss/designs/SKY130_SAR-ADC/xschem/adc_array_circuit/adc_array_circuit_150n_8.sym # of pins=9
** sym_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_array_circuit/adc_array_circuit_150n_8.sym
** sch_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_array_circuit/adc_array_circuit_150n_8.sch
.subckt adc_array_circuit_150n_8  VDD row_n Cbot col_n colon_n sample_n vcom sample VSS
*.PININFO sample_n:I sample:I vcom:B row_n:I col_n:I colon_n:I VDD:B VSS:B Cbot:B
XM1 vcom sample Cbot VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 vcom sample_n Cbot VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 vdrv sample_n Cbot VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 vdrv sample Cbot VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 vint1 col_n vdrv VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM6 VDD row_n vint1 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM7 VDD colon_n vdrv VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM8 vint2 colon_n vdrv VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM9 VSS row_n vint2 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM10 VSS col_n vint2 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:
*+  /foss/designs/SKY130_SAR-ADC/xschem/adc_array_circuit/adc_array_circuit_150n_Drv.sym # of pins=10
** sym_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_array_circuit/adc_array_circuit_150n_Drv.sym
** sch_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_array_circuit/adc_array_circuit_150n_Drv.sch
.subckt adc_array_circuit_150n_Drv  VDD row_n col_n colon_n sample_n_i vcom sample_i VSS sample_n_o
+ sample_o
*.PININFO sample_n_i:I sample_i:I vcom:B row_n:I col_n:I colon_n:I VDD:B VSS:B sample_o:O
*+ sample_n_o:O
XM6 VDD sample_n_i sample_o VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1.6 nf=2 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM7 VDD sample_i sample_n_o VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1.6 nf=2 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM9 VSS sample_i sample_n_o VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.84 nf=2 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM10 VSS sample_n_i sample_o VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.84 nf=2 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:
*+  /foss/designs/SKY130_SAR-ADC/xschem/adc_array_circuit/adc_array_circuit_150n_4.sym # of pins=10
** sym_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_array_circuit/adc_array_circuit_150n_4.sym
** sch_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_array_circuit/adc_array_circuit_150n_4.sch
.subckt adc_array_circuit_150n_4  VDD row_n Cbot col_n colon_n sample_n vcom sample VSS en_n
*.PININFO sample_n:I sample:I vcom:B row_n:I col_n:I colon_n:I VDD:B VSS:B Cbot:B en_n:I
XM1 vcom sample Cbot VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 vcom sample_n Cbot VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 vdrv sample_n Cbot VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 vdrv sample Cbot VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 vint1 en_n vdrv VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM6 VDD en_n vint1 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM7 VDD en_n vdrv VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM8 vint2 en_n vdrv VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM9 VSS en_n vint2 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM10 VSS en_n vint2 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:
*+  /foss/designs/SKY130_SAR-ADC/xschem/adc_array_circuit/adc_array_circuit_150n_2.sym # of pins=10
** sym_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_array_circuit/adc_array_circuit_150n_2.sym
** sch_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_array_circuit/adc_array_circuit_150n_2.sch
.subckt adc_array_circuit_150n_2  VDD row_n Cbot col_n colon_n sample_n vcom sample VSS en_n
*.PININFO sample_n:I sample:I vcom:B row_n:I col_n:I colon_n:I VDD:B VSS:B Cbot:B en_n:I
XM1 vcom sample Cbot VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 vcom sample_n Cbot VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 vdrv sample_n Cbot VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 vdrv sample Cbot VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 vint1 en_n vdrv VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM6 VDD en_n vint1 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM7 VDD en_n vdrv VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM8 vint2 en_n vdrv VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM9 VSS en_n vint2 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM10 VSS en_n vint2 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:
*+  /foss/designs/SKY130_SAR-ADC/xschem/adc_array_circuit/adc_array_circuit_150n_1.sym # of pins=10
** sym_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_array_circuit/adc_array_circuit_150n_1.sym
** sch_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_array_circuit/adc_array_circuit_150n_1.sch
.subckt adc_array_circuit_150n_1  VDD row_n Cbot col_n colon_n sample_n vcom sample VSS en_n
*.PININFO sample_n:I sample:I vcom:B row_n:I col_n:I colon_n:I VDD:B VSS:B Cbot:B en_n:I
XM1 vcom sample Cbot VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 vcom sample_n Cbot VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 vdrv sample_n Cbot VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 vdrv sample Cbot VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 vint1 en_n vdrv VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM6 VDD en_n vint1 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM7 VDD en_n vdrv VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM8 vint2 en_n vdrv VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM9 VSS en_n vint2 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM10 VSS en_n vint2 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:
*+  /foss/designs/SKY130_SAR-ADC/xschem/adc_array_circuit/adc_array_circuit_150n_gate.sym # of pins=12
** sym_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_array_circuit/adc_array_circuit_150n_gate.sym
** sch_path: /foss/designs/SKY130_SAR-ADC/xschem/adc_array_circuit/adc_array_circuit_150n_gate.sch
.subckt adc_array_circuit_150n_gate  VDD row_n col_n colon_n sample_n vcom sample VSS out in sw_n sw
*.PININFO sw:I sw_n:I vcom:B row_n:I col_n:I colon_n:I VDD:B VSS:B sample:I sample_n:I in:B out:B
XM1 in sw_n out VDD sky130_fd_pr__pfet_01v8 L=1 W=2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 in sw out VSS sky130_fd_pr__nfet_01v8 L=0.5 W=1 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.end
