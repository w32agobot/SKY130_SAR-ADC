magic
tech sky130A
magscale 1 2
timestamp 1662392255
<< nwell >>
rect -38 244 1862 582
<< pwell >>
rect -38 -18 1862 174
<< nmos >>
rect 56 80 856 164
rect 1030 80 1060 164
rect 1126 80 1156 164
rect 1222 80 1252 164
rect 1318 80 1348 164
rect 1532 80 1562 164
<< pmos >>
rect 56 308 856 468
rect 1030 308 1060 468
rect 1126 308 1156 468
rect 1222 308 1252 468
rect 1318 308 1348 468
rect 1600 308 1630 468
<< ndiff >>
rect -2 152 56 164
rect -2 92 10 152
rect 44 92 56 152
rect -2 80 56 92
rect 856 152 914 164
rect 856 92 868 152
rect 902 92 914 152
rect 856 80 914 92
rect 968 152 1030 164
rect 968 92 980 152
rect 1014 92 1030 152
rect 968 80 1030 92
rect 1060 152 1126 164
rect 1060 92 1076 152
rect 1110 92 1126 152
rect 1060 80 1126 92
rect 1156 152 1222 164
rect 1156 92 1172 152
rect 1206 92 1222 152
rect 1156 80 1222 92
rect 1252 152 1318 164
rect 1252 92 1268 152
rect 1302 92 1318 152
rect 1252 80 1318 92
rect 1348 152 1410 164
rect 1348 92 1364 152
rect 1398 92 1410 152
rect 1348 80 1410 92
rect 1470 152 1532 164
rect 1470 92 1482 152
rect 1516 92 1532 152
rect 1470 80 1532 92
rect 1562 152 1624 164
rect 1562 92 1578 152
rect 1612 92 1624 152
rect 1562 80 1624 92
<< pdiff >>
rect -2 456 56 468
rect -2 320 10 456
rect 44 320 56 456
rect -2 308 56 320
rect 856 456 914 468
rect 856 320 868 456
rect 902 320 914 456
rect 856 308 914 320
rect 968 456 1030 468
rect 968 320 980 456
rect 1014 320 1030 456
rect 968 308 1030 320
rect 1060 456 1126 468
rect 1060 320 1076 456
rect 1110 320 1126 456
rect 1060 308 1126 320
rect 1156 456 1222 468
rect 1156 320 1172 456
rect 1206 320 1222 456
rect 1156 308 1222 320
rect 1252 456 1318 468
rect 1252 320 1268 456
rect 1302 320 1318 456
rect 1252 308 1318 320
rect 1348 456 1410 468
rect 1348 320 1364 456
rect 1398 320 1410 456
rect 1348 308 1410 320
rect 1538 456 1600 468
rect 1538 320 1550 456
rect 1584 320 1600 456
rect 1538 308 1600 320
rect 1630 456 1718 468
rect 1630 320 1646 456
rect 1680 320 1718 456
rect 1630 308 1718 320
<< ndiffc >>
rect 10 92 44 152
rect 868 92 902 152
rect 980 92 1014 152
rect 1076 92 1110 152
rect 1172 92 1206 152
rect 1268 92 1302 152
rect 1364 92 1398 152
rect 1482 92 1516 152
rect 1578 92 1612 152
<< pdiffc >>
rect 10 320 44 456
rect 868 320 902 456
rect 980 320 1014 456
rect 1076 320 1110 456
rect 1172 320 1206 456
rect 1268 320 1302 456
rect 1364 320 1398 456
rect 1550 320 1584 456
rect 1646 320 1680 456
<< psubdiff >>
rect 94 -18 1730 26
<< poly >>
rect 56 468 856 494
rect 1030 468 1060 494
rect 1126 468 1156 494
rect 1222 468 1252 494
rect 1318 468 1348 494
rect 1600 468 1630 494
rect 56 282 856 308
rect 1030 282 1060 308
rect 1126 282 1156 308
rect 1222 282 1252 308
rect 1318 282 1348 308
rect 1600 282 1630 308
rect 56 266 182 282
rect -32 256 182 266
rect -32 210 -16 256
rect 32 210 182 256
rect -32 200 182 210
rect 898 248 988 258
rect 1030 252 1348 282
rect 1030 248 1060 252
rect 898 246 1060 248
rect 898 212 938 246
rect 972 212 1060 246
rect 898 206 1060 212
rect 898 202 988 206
rect 56 190 182 200
rect 56 164 856 190
rect 1030 164 1060 206
rect 1126 164 1156 252
rect 1222 164 1252 252
rect 1318 164 1348 252
rect 1392 252 1458 262
rect 1392 218 1408 252
rect 1442 220 1458 252
rect 1532 252 1630 282
rect 1532 220 1562 252
rect 1442 218 1562 220
rect 1392 190 1562 218
rect 1532 164 1562 190
rect 56 54 856 80
rect 1030 54 1060 80
rect 1126 54 1156 80
rect 1222 54 1252 80
rect 1318 54 1348 80
rect 1532 54 1562 80
<< polycont >>
rect -16 210 32 256
rect 938 212 972 246
rect 1408 218 1442 252
<< locali >>
rect 0 561 1824 562
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1824 561
rect 0 526 1824 527
rect 10 456 44 472
rect 10 304 44 320
rect 868 456 902 472
rect -32 256 48 260
rect -32 210 -16 256
rect 32 210 48 256
rect -32 206 48 210
rect 868 258 902 320
rect 980 456 1014 472
rect 980 304 1014 320
rect 1076 456 1110 526
rect 1076 304 1110 320
rect 1172 456 1206 472
rect 1172 304 1206 320
rect 1268 456 1302 472
rect 1268 304 1302 320
rect 1364 456 1398 472
rect 1364 304 1398 320
rect 1476 270 1510 526
rect 1544 456 1584 472
rect 1544 320 1550 456
rect 1544 304 1584 320
rect 1646 456 1680 472
rect 1646 270 1680 320
rect 868 246 988 258
rect 868 212 916 246
rect 972 212 988 246
rect 868 202 988 212
rect 1408 252 1442 268
rect 1476 236 1612 270
rect 1646 236 1694 270
rect 1408 202 1442 218
rect 10 152 44 168
rect 10 76 44 92
rect 868 152 902 202
rect 868 76 902 92
rect 980 152 1014 168
rect 980 76 1014 92
rect 1076 152 1110 168
rect 1076 18 1110 92
rect 1172 152 1206 168
rect 1172 76 1206 92
rect 1268 76 1302 92
rect 1364 152 1398 168
rect 1364 76 1398 92
rect 1482 152 1516 168
rect 1482 76 1516 92
rect 1578 152 1612 236
rect 1578 76 1612 92
rect 1660 18 1694 236
rect 0 -18 28 18
rect 64 17 1824 18
rect 64 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1824 17
rect 64 -18 1824 -17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 10 320 44 456
rect 868 320 902 456
rect 980 320 1014 456
rect 1172 320 1206 456
rect 1268 320 1302 376
rect 1364 320 1398 456
rect 1550 340 1584 456
rect 916 212 938 246
rect 938 212 972 246
rect 1408 218 1442 252
rect 10 92 44 152
rect 868 92 902 152
rect 980 92 1014 152
rect 1172 92 1206 152
rect 1268 152 1302 178
rect 1268 144 1302 152
rect 1364 92 1398 152
rect 1482 92 1516 132
rect 28 -18 64 18
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
<< metal1 >>
rect 0 561 1824 594
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1824 561
rect 0 496 1824 527
rect 4 456 50 496
rect 4 320 10 456
rect 44 320 50 456
rect 4 308 50 320
rect 862 456 908 468
rect 862 320 868 456
rect 902 320 908 456
rect 862 258 908 320
rect 974 456 1020 468
rect 974 320 980 456
rect 1014 400 1020 456
rect 1166 456 1590 468
rect 1166 400 1172 456
rect 1014 362 1172 400
rect 1014 320 1020 362
rect 974 308 1020 320
rect 1166 320 1172 362
rect 1206 434 1364 456
rect 1206 320 1212 434
rect 1166 308 1212 320
rect 1262 376 1308 406
rect 1262 320 1268 376
rect 1302 320 1308 376
rect 862 256 988 258
rect 862 204 916 256
rect 972 204 988 256
rect 862 202 988 204
rect 1262 248 1308 320
rect 1358 320 1364 434
rect 1398 434 1550 456
rect 1398 320 1404 434
rect 1544 340 1550 434
rect 1584 340 1590 456
rect 1544 328 1590 340
rect 1358 308 1404 320
rect 1396 252 1454 258
rect 1396 248 1408 252
rect 1262 220 1408 248
rect 4 152 50 164
rect 4 92 10 152
rect 44 92 50 152
rect 4 48 50 92
rect 862 152 908 202
rect 1262 178 1308 220
rect 1396 218 1408 220
rect 1442 248 1454 252
rect 1442 220 1824 248
rect 1442 218 1454 220
rect 1396 212 1454 218
rect 862 92 868 152
rect 902 92 908 152
rect 862 80 908 92
rect 974 152 1020 164
rect 974 92 980 152
rect 1014 138 1020 152
rect 1166 152 1212 164
rect 1166 138 1172 152
rect 1014 104 1172 138
rect 1014 92 1020 104
rect 974 80 1020 92
rect 1166 92 1172 104
rect 1206 104 1212 152
rect 1262 144 1268 178
rect 1302 144 1308 178
rect 1262 132 1308 144
rect 1358 152 1404 164
rect 1358 104 1364 152
rect 1206 92 1364 104
rect 1398 108 1404 152
rect 1476 132 1522 144
rect 1476 108 1482 132
rect 1398 92 1482 108
rect 1516 92 1522 132
rect 1166 80 1522 92
rect 1166 76 1496 80
rect 0 44 1824 48
rect 0 40 1472 44
rect 0 18 246 40
rect 0 -18 28 18
rect 64 17 246 18
rect 304 17 1472 40
rect 1530 17 1824 44
rect 64 -17 121 17
rect 155 -17 213 17
rect 304 -12 305 17
rect 247 -17 305 -12
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -12 1472 17
rect 1443 -17 1501 -12
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1824 17
rect 64 -18 1824 -17
rect 0 -48 1824 -18
<< via1 >>
rect 916 246 972 256
rect 916 212 972 246
rect 916 204 972 212
rect 246 17 304 40
rect 1472 17 1530 44
rect 246 -12 247 17
rect 247 -12 304 17
rect 1472 -12 1501 17
rect 1501 -12 1530 17
<< metal2 >>
rect 912 260 992 290
rect 912 258 922 260
rect 898 256 922 258
rect 898 204 916 256
rect 898 202 922 204
rect 978 202 992 260
rect 912 168 992 202
rect 212 44 340 48
rect 212 -12 246 44
rect 304 -12 340 44
rect 212 -18 340 -12
rect 1436 44 1564 48
rect 1436 -12 1472 44
rect 1530 -12 1564 44
rect 1436 -18 1564 -12
<< via2 >>
rect 922 256 978 260
rect 922 204 972 256
rect 972 204 978 256
rect 922 202 978 204
rect 246 40 304 44
rect 246 -12 304 40
rect 1472 -12 1530 44
<< metal3 >>
rect 54 54 850 496
rect 912 264 992 290
rect 912 200 918 264
rect 982 200 992 264
rect 912 168 992 200
rect 1056 54 1788 496
rect 212 44 340 54
rect 212 -12 246 44
rect 304 -12 340 44
rect 212 -18 340 -12
rect 1436 44 1564 54
rect 1436 -12 1472 44
rect 1530 -12 1564 44
rect 1436 -18 1564 -12
<< via3 >>
rect 918 260 982 264
rect 918 202 922 260
rect 922 202 978 260
rect 978 202 982 260
rect 918 200 982 202
<< mimcap >>
rect 86 264 822 468
rect 86 200 736 264
rect 800 200 822 264
rect 86 82 822 200
rect 1084 264 1736 468
rect 1084 200 1100 264
rect 1164 200 1736 264
rect 1084 82 1736 200
<< mimcapcontact >>
rect 736 200 800 264
rect 1100 200 1164 264
<< metal4 >>
rect 912 268 992 290
rect 732 264 1170 268
rect 732 200 736 264
rect 800 200 918 264
rect 982 200 1100 264
rect 1164 200 1170 264
rect 732 194 1170 200
rect 912 168 992 194
<< labels >>
rlabel locali -16 210 32 256 7 in
port 2 w
rlabel metal1 0 496 1824 594 7 VPWR
port 1 w
rlabel nwell 28 526 64 562 7 VPB
port 6 w
rlabel metal1 1794 220 1824 248 3 out
port 3 e
rlabel metal1 0 -48 0 48 7 VGND
port 4 w
rlabel metal1 1824 -48 1824 48 3 VGND
port 4 e
rlabel locali 868 76 902 76 5 cap_top
rlabel psubdiff 120 -14 156 22 7 VNB
port 5 w
<< end >>
