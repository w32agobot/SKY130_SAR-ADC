magic
tech sky130A
timestamp 1661513809
<< nwell >>
rect -4 2 253 230
<< nmos >>
rect 45 -74 60 -32
rect 93 -74 108 -32
<< pmos >>
rect 45 53 60 133
rect 93 53 108 133
rect 141 53 156 133
rect 189 53 204 133
<< ndiff >>
rect 14 -38 45 -32
rect 14 -68 20 -38
rect 37 -68 45 -38
rect 14 -74 45 -68
rect 60 -38 93 -32
rect 60 -68 68 -38
rect 85 -68 93 -38
rect 60 -74 93 -68
rect 108 -38 139 -32
rect 108 -68 116 -38
rect 133 -68 139 -38
rect 108 -74 139 -68
<< pdiff >>
rect 14 127 45 133
rect 14 59 20 127
rect 37 59 45 127
rect 14 53 45 59
rect 60 127 93 133
rect 60 59 68 127
rect 85 59 93 127
rect 60 53 93 59
rect 108 127 141 133
rect 108 59 116 127
rect 133 59 141 127
rect 108 53 141 59
rect 156 127 189 133
rect 156 59 164 127
rect 181 59 189 127
rect 156 53 189 59
rect 204 127 235 133
rect 204 59 212 127
rect 229 59 235 127
rect 204 53 235 59
<< ndiffc >>
rect 20 -68 37 -38
rect 68 -68 85 -38
rect 116 -68 133 -38
<< pdiffc >>
rect 20 59 37 127
rect 68 59 85 127
rect 116 59 133 127
rect 164 59 181 127
rect 212 59 229 127
<< psubdiff >>
rect 56 -118 68 -101
rect 85 -118 99 -101
<< nsubdiff >>
rect 33 195 48 212
rect 65 195 82 212
rect 99 195 116 212
rect 133 195 150 212
rect 167 195 184 212
rect 201 195 222 212
<< psubdiffcont >>
rect 68 -118 85 -101
<< nsubdiffcont >>
rect 48 195 65 212
rect 82 195 99 212
rect 116 195 133 212
rect 150 195 167 212
rect 184 195 201 212
<< poly >>
rect 23 174 156 182
rect 23 157 28 174
rect 45 167 156 174
rect 45 157 60 167
rect 23 149 60 157
rect 45 133 60 149
rect 93 133 108 146
rect 141 133 156 167
rect 189 133 204 146
rect 45 -32 60 53
rect 93 37 108 53
rect 141 40 156 53
rect 81 29 108 37
rect 81 12 86 29
rect 103 19 108 29
rect 189 19 204 53
rect 103 12 204 19
rect 81 4 204 12
rect 93 -32 108 4
rect 45 -87 60 -74
rect 93 -87 108 -74
<< polycont >>
rect 28 157 45 174
rect 86 12 103 29
<< locali >>
rect 40 195 48 212
rect 65 195 82 212
rect 99 195 116 212
rect 133 195 150 212
rect 167 195 184 212
rect 201 195 215 212
rect 20 174 53 178
rect 20 157 28 174
rect 45 157 53 174
rect 20 152 53 157
rect 20 127 37 135
rect 20 -38 37 59
rect 68 127 85 135
rect 68 51 85 59
rect 116 127 133 195
rect 116 51 133 59
rect 164 127 181 135
rect 164 51 181 59
rect 212 127 229 135
rect 78 29 111 33
rect 78 12 86 29
rect 103 12 111 29
rect 78 7 111 12
rect 212 -1 229 59
rect 126 -20 229 -1
rect 126 -30 143 -20
rect 20 -76 37 -68
rect 68 -38 85 -30
rect 68 -101 85 -68
rect 116 -38 143 -30
rect 133 -68 143 -38
rect 116 -76 143 -68
rect 56 -118 68 -101
rect 85 -118 99 -101
<< viali >>
rect 86 12 103 29
rect 20 -68 37 -38
rect 116 -68 133 -38
<< metal1 >>
rect 78 31 111 33
rect 12 29 111 31
rect 12 13 86 29
rect 78 12 86 13
rect 103 12 111 29
rect 78 7 111 12
rect 17 -38 40 -32
rect 17 -68 20 -38
rect 37 -46 40 -38
rect 113 -38 136 -32
rect 113 -46 116 -38
rect 37 -60 116 -46
rect 37 -68 40 -60
rect 17 -74 40 -68
rect 113 -68 116 -60
rect 133 -68 136 -38
rect 113 -74 136 -68
<< comment >>
rect 61 58 71 132
rect 115 58 134 126
rect 178 55 188 129
rect 69 -65 83 -41
<< labels >>
rlabel locali 40 195 40 212 7 VDD
port 1 w
rlabel locali 229 -20 229 -1 3 Q
port 7 e
rlabel metal1 12 13 12 31 7 B
port 6 w
rlabel locali 20 152 20 178 7 A
port 8 w
rlabel locali 56 -118 56 -101 7 VSS
port 4 w
<< end >>
