* SPICE3 file created from adc_array_wafflecap_9_5ux5u_4870aF.ext - technology: sky130A

.subckt adc_array_wafflecap_9_5ux5u_4870aF ctop cbot
C0 cbot ctop 4.87fF
.ends
