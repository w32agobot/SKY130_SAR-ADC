magic
tech sky130A
timestamp 1661515501
<< nwell >>
rect 0 120 505 348
<< nmos >>
rect 49 44 64 86
rect 97 44 112 86
rect 297 44 312 86
rect 345 44 360 86
<< pmos >>
rect 49 171 64 251
rect 97 171 112 251
rect 145 171 160 251
rect 193 171 208 251
rect 297 171 312 251
rect 345 171 360 251
rect 393 171 408 251
rect 441 171 456 251
<< ndiff >>
rect 18 80 49 86
rect 18 50 24 80
rect 41 50 49 80
rect 18 44 49 50
rect 64 80 97 86
rect 64 50 72 80
rect 89 50 97 80
rect 64 44 97 50
rect 112 80 143 86
rect 112 50 120 80
rect 137 50 143 80
rect 112 44 143 50
rect 266 80 297 86
rect 266 50 272 80
rect 289 50 297 80
rect 266 44 297 50
rect 312 80 345 86
rect 312 50 320 80
rect 337 50 345 80
rect 312 44 345 50
rect 360 80 391 86
rect 360 50 368 80
rect 385 50 391 80
rect 360 44 391 50
<< pdiff >>
rect 18 245 49 251
rect 18 177 24 245
rect 41 177 49 245
rect 18 171 49 177
rect 64 245 97 251
rect 64 177 72 245
rect 89 177 97 245
rect 64 171 97 177
rect 112 245 145 251
rect 112 177 120 245
rect 137 177 145 245
rect 112 171 145 177
rect 160 245 193 251
rect 160 177 168 245
rect 185 177 193 245
rect 160 171 193 177
rect 208 245 239 251
rect 208 177 216 245
rect 233 177 239 245
rect 208 171 239 177
rect 266 245 297 251
rect 266 177 272 245
rect 289 177 297 245
rect 266 171 297 177
rect 312 245 345 251
rect 312 177 320 245
rect 337 177 345 245
rect 312 171 345 177
rect 360 245 393 251
rect 360 177 368 245
rect 385 177 393 245
rect 360 171 393 177
rect 408 245 441 251
rect 408 177 416 245
rect 433 177 441 245
rect 408 171 441 177
rect 456 245 487 251
rect 456 177 464 245
rect 481 177 487 245
rect 456 171 487 177
<< ndiffc >>
rect 24 50 41 80
rect 72 50 89 80
rect 120 50 137 80
rect 272 50 289 80
rect 320 50 337 80
rect 368 50 385 80
<< pdiffc >>
rect 24 177 41 245
rect 72 177 89 245
rect 120 177 137 245
rect 168 177 185 245
rect 216 177 233 245
rect 272 177 289 245
rect 320 177 337 245
rect 368 177 385 245
rect 416 177 433 245
rect 464 177 481 245
<< psubdiff >>
rect 60 0 72 17
rect 89 0 103 17
rect 308 0 320 17
rect 337 0 351 17
<< nsubdiff >>
rect 37 313 52 330
rect 69 313 86 330
rect 103 313 120 330
rect 137 313 154 330
rect 171 313 188 330
rect 205 313 226 330
rect 285 313 300 330
rect 317 313 334 330
rect 351 313 368 330
rect 385 313 402 330
rect 419 313 436 330
rect 453 313 474 330
<< psubdiffcont >>
rect 72 0 89 17
rect 320 0 337 17
<< nsubdiffcont >>
rect 52 313 69 330
rect 86 313 103 330
rect 120 313 137 330
rect 154 313 171 330
rect 188 313 205 330
rect 300 313 317 330
rect 334 313 351 330
rect 368 313 385 330
rect 402 313 419 330
rect 436 313 453 330
<< poly >>
rect 27 292 160 300
rect 27 275 32 292
rect 49 285 160 292
rect 49 275 64 285
rect 27 267 64 275
rect 49 251 64 267
rect 97 251 112 264
rect 145 251 160 285
rect 275 292 408 300
rect 275 275 280 292
rect 297 285 408 292
rect 297 275 312 285
rect 275 267 312 275
rect 193 251 208 264
rect 297 251 312 267
rect 345 251 360 264
rect 393 251 408 285
rect 441 251 456 264
rect 49 114 64 171
rect 97 155 112 171
rect 145 158 160 171
rect 85 147 112 155
rect 85 130 90 147
rect 107 137 112 147
rect 193 137 208 171
rect 107 130 208 137
rect 85 122 208 130
rect 0 98 64 114
rect 49 86 64 98
rect 97 86 112 122
rect 297 86 312 171
rect 345 155 360 171
rect 393 158 408 171
rect 333 147 360 155
rect 333 130 338 147
rect 355 137 360 147
rect 441 137 456 171
rect 355 130 456 137
rect 333 122 456 130
rect 345 86 360 122
rect 49 31 64 44
rect 97 31 112 44
rect 297 31 312 44
rect 345 31 360 44
<< polycont >>
rect 32 275 49 292
rect 280 275 297 292
rect 90 130 107 147
rect 338 130 355 147
<< locali >>
rect 44 313 52 330
rect 69 313 86 330
rect 103 313 120 330
rect 137 313 154 330
rect 171 313 188 330
rect 205 313 300 330
rect 317 313 334 330
rect 351 313 368 330
rect 385 313 402 330
rect 419 313 436 330
rect 453 313 467 330
rect 24 292 57 296
rect 24 275 32 292
rect 49 275 57 292
rect 24 270 57 275
rect 24 245 41 253
rect 24 80 41 177
rect 72 245 89 253
rect 72 169 89 177
rect 120 245 137 313
rect 272 293 305 296
rect 272 275 280 293
rect 297 275 305 293
rect 272 270 305 275
rect 120 169 137 177
rect 168 245 185 253
rect 168 169 185 177
rect 216 245 233 253
rect 82 147 115 151
rect 82 130 90 147
rect 107 130 115 147
rect 82 125 115 130
rect 216 122 233 177
rect 272 245 289 253
rect 216 119 240 122
rect 216 117 220 119
rect 130 102 220 117
rect 237 102 240 119
rect 130 98 240 102
rect 130 88 147 98
rect 24 42 41 50
rect 72 80 89 88
rect 72 17 89 50
rect 120 80 147 88
rect 137 50 147 80
rect 120 42 147 50
rect 272 80 289 177
rect 320 245 337 253
rect 320 169 337 177
rect 368 245 385 313
rect 368 169 385 177
rect 416 245 433 253
rect 416 169 433 177
rect 464 245 481 253
rect 330 147 363 151
rect 330 130 338 147
rect 355 130 363 147
rect 330 125 363 130
rect 464 117 481 177
rect 378 98 481 117
rect 378 88 395 98
rect 272 42 289 50
rect 320 80 337 88
rect 320 17 337 50
rect 368 80 395 88
rect 385 50 395 80
rect 368 42 395 50
rect 59 0 72 17
rect 89 0 320 17
rect 337 0 352 17
<< viali >>
rect 280 292 297 293
rect 280 276 297 292
rect 90 130 107 147
rect 220 102 237 119
rect 24 50 41 80
rect 120 50 137 80
rect 338 130 355 147
rect 272 50 289 80
rect 368 50 385 80
<< metal1 >>
rect -3 296 58 299
rect -3 293 303 296
rect -3 282 280 293
rect 272 276 280 282
rect 297 276 303 293
rect 272 273 303 276
rect 82 149 115 151
rect 330 150 363 151
rect 324 149 483 150
rect 16 147 195 149
rect 16 131 90 147
rect 82 130 90 131
rect 107 131 195 147
rect 107 130 115 131
rect 82 125 115 130
rect 21 80 44 86
rect 21 50 24 80
rect 41 72 44 80
rect 117 80 140 86
rect 117 72 120 80
rect 41 58 120 72
rect 41 50 44 58
rect 21 44 44 50
rect 117 50 120 58
rect 137 50 140 80
rect 177 75 195 131
rect 222 147 483 149
rect 222 131 338 147
rect 222 125 240 131
rect 330 130 338 131
rect 355 132 483 147
rect 355 130 363 132
rect 330 125 363 130
rect 216 119 240 125
rect 216 102 220 119
rect 237 102 240 119
rect 216 96 240 102
rect 269 80 292 86
rect 269 75 272 80
rect 177 57 272 75
rect 117 44 140 50
rect 269 50 272 57
rect 289 72 292 80
rect 365 80 388 86
rect 365 72 368 80
rect 289 58 368 72
rect 289 50 292 58
rect 269 44 292 50
rect 365 50 368 58
rect 385 50 388 80
rect 365 44 388 50
<< comment >>
rect 65 176 75 250
rect 119 176 138 244
rect 182 173 192 247
rect 313 176 323 250
rect 367 176 386 244
rect 430 173 440 247
rect 73 53 87 77
rect 321 53 335 77
<< labels >>
rlabel poly 0 98 0 114 7 R
port 1 w
rlabel metal1 -3 283 -3 299 7 S
port 7 w
rlabel locali 44 313 44 330 7 VDD
port 4 w
rlabel locali 481 98 481 118 3 QN
port 2 e
rlabel metal1 483 132 483 150 3 Q
port 6 e
rlabel locali 59 0 59 17 7 VSS
port 5 w
rlabel locali 292 313 292 330 7 NOR_1/VDD
rlabel locali 481 98 481 117 3 NOR_1/Q
rlabel metal1 264 131 264 149 7 NOR_1/B
rlabel locali 272 270 272 296 7 NOR_1/A
rlabel locali 308 0 308 17 7 NOR_1/VSS
rlabel locali 44 313 44 330 7 NOR_0/VDD
rlabel locali 233 98 233 117 3 NOR_0/Q
rlabel metal1 16 131 16 149 7 NOR_0/B
rlabel locali 24 270 24 296 7 NOR_0/A
rlabel locali 60 0 60 17 7 NOR_0/VSS
<< end >>
