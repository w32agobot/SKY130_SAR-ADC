magic
tech sky130A
magscale 1 2
timestamp 1662821229
<< nwell >>
rect -38 414 2338 582
rect -38 247 946 414
rect 1648 247 2338 414
<< pwell >>
rect 946 214 1648 414
rect 1 -17 2299 214
<< nmos >>
rect 85 95 851 179
rect 1072 71 1522 346
rect 1694 71 1724 155
rect 1790 71 1820 155
rect 1999 71 2029 155
rect 2095 71 2125 155
<< pmos >>
rect 1753 329 1783 489
rect 1849 329 1879 489
rect 2087 329 2117 489
rect 2183 329 2213 489
<< pmoslvt >>
rect 85 283 851 443
<< ndiff >>
rect 1014 334 1072 346
rect 27 142 85 179
rect 27 107 39 142
rect 73 107 85 142
rect 27 95 85 107
rect 851 159 909 179
rect 851 107 863 159
rect 897 107 909 159
rect 851 95 909 107
rect 1014 79 1026 334
rect 1060 79 1072 334
rect 1014 71 1072 79
rect 1522 334 1580 346
rect 1522 79 1534 334
rect 1568 79 1580 334
rect 1522 71 1580 79
rect 1634 143 1694 155
rect 1634 83 1644 143
rect 1678 83 1694 143
rect 1634 71 1694 83
rect 1724 143 1790 155
rect 1724 85 1740 143
rect 1774 85 1790 143
rect 1724 71 1790 85
rect 1820 143 1878 155
rect 1820 85 1836 143
rect 1870 85 1878 143
rect 1820 71 1878 85
rect 1937 124 1999 155
rect 1937 85 1949 124
rect 1983 85 1999 124
rect 1937 71 1999 85
rect 2029 143 2095 155
rect 2029 85 2045 143
rect 2079 85 2095 143
rect 2029 71 2095 85
rect 2125 143 2187 155
rect 2125 85 2141 143
rect 2175 85 2187 143
rect 2125 71 2187 85
<< pdiff >>
rect 1693 477 1753 489
rect 27 431 85 443
rect 27 379 39 431
rect 73 379 85 431
rect 27 283 85 379
rect 851 431 909 443
rect 851 305 863 431
rect 897 305 909 431
rect 851 283 909 305
rect 1693 341 1703 477
rect 1737 341 1753 477
rect 1693 329 1753 341
rect 1783 475 1849 489
rect 1783 354 1799 475
rect 1833 354 1849 475
rect 1783 329 1849 354
rect 1879 475 1939 489
rect 1879 341 1895 475
rect 1929 341 1939 475
rect 1879 329 1939 341
rect 2025 475 2087 489
rect 2025 400 2037 475
rect 2071 400 2087 475
rect 2025 329 2087 400
rect 2117 475 2183 489
rect 2117 341 2133 475
rect 2167 341 2183 475
rect 2117 329 2183 341
rect 2213 475 2273 489
rect 2213 341 2229 475
rect 2263 341 2273 475
rect 2213 329 2273 341
<< ndiffc >>
rect 39 107 73 142
rect 863 107 897 159
rect 1026 79 1060 334
rect 1534 79 1568 334
rect 1644 83 1678 143
rect 1740 85 1774 143
rect 1836 85 1870 143
rect 1949 85 1983 124
rect 2045 85 2079 143
rect 2141 85 2175 143
<< pdiffc >>
rect 39 379 73 431
rect 863 305 897 431
rect 1703 341 1737 477
rect 1799 354 1833 475
rect 1895 341 1929 475
rect 2037 400 2071 475
rect 2133 341 2167 475
rect 2229 341 2263 475
<< poly >>
rect 1753 489 1783 515
rect 1849 489 1879 515
rect 2087 489 2117 515
rect 2183 489 2213 515
rect 85 443 851 479
rect 1072 418 1522 438
rect 1072 384 1121 418
rect 1475 384 1522 418
rect 1072 346 1522 384
rect 85 243 851 283
rect 924 243 980 259
rect 85 209 934 243
rect 968 209 980 243
rect 85 179 851 209
rect 924 193 980 209
rect 85 69 851 95
rect 1753 314 1783 329
rect 1849 314 1879 329
rect 1753 284 1879 314
rect 2087 305 2117 329
rect 2183 305 2213 329
rect 1753 248 1783 284
rect 1694 236 1783 248
rect 2087 275 2213 305
rect 2087 265 2180 275
rect 1694 202 1733 236
rect 1767 214 1783 236
rect 1916 227 1982 238
rect 1767 202 1820 214
rect 1694 184 1820 202
rect 1694 155 1724 184
rect 1790 155 1820 184
rect 1916 193 1932 227
rect 1966 219 1982 227
rect 2087 231 2130 265
rect 2164 231 2180 265
rect 2087 219 2180 231
rect 1966 193 2125 219
rect 1916 189 2125 193
rect 1916 182 2029 189
rect 1999 155 2029 182
rect 2095 155 2125 189
rect 1072 32 1522 71
rect 1694 44 1724 71
rect 1790 44 1820 71
rect 1999 44 2029 71
rect 2095 44 2125 71
<< polycont >>
rect 1121 384 1475 418
rect 934 209 968 243
rect 1733 202 1767 236
rect 1932 193 1966 227
rect 2130 231 2164 265
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2300 561
rect 1703 477 1737 527
rect 39 431 73 447
rect 38 379 39 400
rect 38 361 73 379
rect 863 431 897 447
rect 1095 418 1499 425
rect 1095 384 1121 418
rect 1475 384 1499 418
rect 1095 374 1499 384
rect 1026 336 1060 350
rect 1534 336 1568 351
rect 863 289 897 305
rect 1024 334 1568 336
rect 21 243 75 264
rect 21 209 934 243
rect 968 209 985 243
rect 21 198 75 209
rect 863 159 897 175
rect 39 142 73 158
rect 39 91 73 107
rect 863 73 897 107
rect 1024 79 1026 334
rect 1060 79 1534 334
rect 1703 325 1737 341
rect 1799 475 1833 491
rect 1799 325 1833 354
rect 1895 475 1929 491
rect 1634 268 1668 279
rect 1634 235 1678 268
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 1024 17 1568 79
rect 1644 143 1678 235
rect 1712 202 1723 236
rect 1767 202 1783 236
rect 1895 228 1929 341
rect 1963 296 1997 527
rect 2031 475 2071 491
rect 2031 400 2037 475
rect 2031 383 2071 400
rect 2133 475 2167 491
rect 2133 309 2167 341
rect 2229 475 2269 491
rect 2263 341 2269 475
rect 2229 325 2269 341
rect 1963 262 2079 296
rect 1895 227 1982 228
rect 1895 210 1932 227
rect 1836 193 1932 210
rect 1966 193 1982 227
rect 1836 176 1929 193
rect 1644 17 1678 83
rect 1740 143 1774 159
rect 1740 69 1774 85
rect 1836 143 1870 176
rect 2045 143 2079 262
rect 2114 231 2130 265
rect 2164 231 2181 265
rect 2135 193 2181 231
rect 1836 69 1870 85
rect 1949 133 1983 143
rect 1949 69 1983 85
rect 2045 69 2079 85
rect 2141 143 2175 159
rect 2141 69 2175 85
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2300 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 39 379 73 431
rect 863 305 897 417
rect 1228 384 1264 418
rect 1326 384 1362 418
rect 39 107 73 142
rect 863 107 897 143
rect 1799 354 1833 445
rect 1634 279 1668 313
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 18
rect 1723 202 1733 236
rect 1733 202 1767 236
rect 2037 412 2071 451
rect 2133 341 2167 389
rect 2229 361 2263 443
rect 1740 105 1774 143
rect 1949 124 1983 133
rect 1949 99 1983 124
rect 2141 105 2175 139
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
<< metal1 >>
rect 0 561 2300 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2300 561
rect 0 496 2300 527
rect 33 431 79 496
rect 1793 451 2269 458
rect 1793 445 2037 451
rect 33 379 39 431
rect 73 379 79 431
rect 33 362 79 379
rect 857 417 903 439
rect 38 361 73 362
rect 857 305 863 417
rect 897 316 903 417
rect 1216 418 1374 424
rect 1216 384 1228 418
rect 1264 384 1326 418
rect 1362 384 1374 418
rect 1216 378 1374 384
rect 1273 336 1318 378
rect 1793 354 1799 445
rect 1833 430 2037 445
rect 1833 354 1839 430
rect 2031 412 2037 430
rect 2071 443 2269 451
rect 2071 430 2229 443
rect 2071 412 2077 430
rect 2031 400 2077 412
rect 1793 342 1839 354
rect 2127 389 2173 402
rect 2127 341 2133 389
rect 2167 341 2173 389
rect 2223 361 2229 430
rect 2263 361 2269 443
rect 2223 349 2269 361
rect 1010 316 1588 336
rect 897 305 1588 316
rect 857 285 1588 305
rect 982 223 1588 285
rect 1622 314 1674 320
rect 2127 314 2173 341
rect 1622 313 2173 314
rect 1622 279 1634 313
rect 1668 279 2173 313
rect 1622 275 2173 279
rect 1622 273 1674 275
rect 1693 236 1783 242
rect 1693 223 1723 236
rect 982 202 1723 223
rect 1767 202 1783 236
rect 982 184 1783 202
rect 982 157 1588 184
rect 33 142 79 155
rect 33 107 39 142
rect 73 107 79 142
rect 33 48 79 107
rect 856 143 1588 157
rect 856 107 863 143
rect 897 107 1588 143
rect 856 95 1588 107
rect 1010 93 1588 95
rect 1734 143 1780 155
rect 1734 105 1740 143
rect 1774 121 1780 143
rect 2129 139 2187 147
rect 1937 133 1995 139
rect 1937 121 1949 133
rect 1774 105 1949 121
rect 1734 99 1949 105
rect 1983 121 1995 133
rect 2129 121 2141 139
rect 1983 105 2141 121
rect 2175 113 2187 139
rect 2175 105 2181 113
rect 1983 99 2181 105
rect 1734 93 2181 99
rect 0 18 2300 48
rect 0 17 949 18
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 17 2300 18
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2300 17
rect 0 -48 2300 -17
<< labels >>
flabel metal1 s 0 496 2300 592 0 FreeSans 160 0 0 0 VPWR
port 1 nsew power bidirectional abutment
flabel metal1 s 0 -48 2300 48 0 FreeSans 160 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 673 527 707 561 0 FreeSans 160 0 0 0 VPWR
port 1 nsew power bidirectional abutment
flabel metal1 s 673 -17 707 17 0 FreeSans 160 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel nwell s 673 527 707 561 0 FreeSans 160 0 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 673 -17 707 17 0 FreeSans 160 0 0 0 VNB
port 6 nsew ground bidirectional
flabel locali s 40 221 74 255 7 FreeSans 160 0 0 0 in
port 2 nsew signal input
rlabel locali 863 161 897 161 1 cap_top
flabel locali s 2141 207 2175 241 0 FreeSans 160 0 0 0 out
port 3 nsew signal output
flabel metal1 s 1317 -17 1351 17 0 FreeSans 160 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel pwell s 1317 -17 1351 17 0 FreeSans 160 0 0 0 VNB
port 6 nsew ground bidirectional
flabel metal1 s 949 -16 983 18 0 FreeSans 160 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 121 -17 155 17 0 FreeSans 160 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 121 527 155 561 0 FreeSans 160 0 0 0 VPWR
port 1 nsew power bidirectional abutment
flabel nwell s 121 527 155 561 0 FreeSans 160 0 0 0 VPB
port 5 nsew power bidirectional
flabel metal1 s 2145 527 2179 561 0 FreeSans 160 0 0 0 VPWR
port 1 nsew power bidirectional abutment
flabel nwell s 2145 527 2179 561 0 FreeSans 160 0 0 0 VPB
port 5 nsew power bidirectional
flabel metal1 s 1961 527 1995 561 0 FreeSans 160 0 0 0 VPWR
port 1 nsew power bidirectional abutment
flabel nwell s 1961 527 1995 561 0 FreeSans 160 0 0 0 VPB
port 5 nsew power bidirectional
flabel metal1 s 1501 527 1535 561 0 FreeSans 160 0 0 0 VPWR
port 1 nsew power bidirectional abutment
flabel nwell s 1501 527 1535 561 0 FreeSans 160 0 0 0 VPB
port 5 nsew power bidirectional
flabel metal1 s 1869 -17 1903 17 0 FreeSans 160 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel pwell s 1869 -17 1903 17 0 FreeSans 160 0 0 0 VNB
port 6 nsew ground bidirectional
flabel pwell s 121 -17 155 17 0 FreeSans 160 0 0 0 VNB
port 6 nsew ground bidirectional
flabel pwell s 949 -16 983 18 0 FreeSans 160 0 0 0 VNB
port 6 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 2300 544
string LEFclass CORE
string LEForigin 0 0
string LEFsite unithd
string LEFsource USER
<< end >>
