magic
tech sky130A
timestamp 1663932020
<< nwell >>
rect 0 253 47 440
rect 451 253 502 440
<< locali >>
rect 57 443 74 502
rect 427 443 444 502
rect 57 0 74 64
rect 427 0 444 64
<< metal1 >>
rect 0 399 47 427
rect 451 399 502 427
rect 0 370 47 385
rect 451 370 502 385
rect 0 256 47 270
rect 451 256 502 270
rect 0 215 47 229
rect 451 215 502 229
rect 0 187 47 201
rect 451 187 502 201
rect 0 110 47 124
rect 451 110 502 124
rect 0 68 47 96
rect 451 68 502 96
<< metal2 >>
rect 209 484 258 486
<< metal4 >>
rect 92 454 122 467
<< comment >>
rect 69 375 154 399
rect 215 378 281 402
rect 69 130 97 375
rect 156 345 184 375
rect 150 130 178 159
rect 179 157 203 344
rect 215 281 239 378
rect 282 358 303 381
rect 299 302 316 358
rect 279 301 316 302
rect 279 281 300 301
rect 215 279 300 281
rect 215 257 279 279
rect 69 129 178 130
rect 69 106 153 129
rect 215 103 239 257
rect 280 239 301 261
rect 280 238 318 239
rect 301 99 318 238
rect 335 99 358 401
use adc_array_circuit_drv  adc_array_circuit_drv_0
timestamp 1663066618
transform 1 0 -70 0 1 -221
box 117 285 521 664
use adc_array_top_drv adc_array_top_drv_0
timestamp 1659615172
transform 1 0 0 0 1 0
box 0 0 502 502
<< labels >>
rlabel metal1 0 399 0 427 7 vdd
port 2 w
rlabel metal1 0 256 0 270 7 colon_n
port 3 w
rlabel metal1 0 215 0 229 7 col_n
port 4 w
rlabel metal1 0 110 0 124 7 vcom
port 5 w
rlabel metal1 0 68 0 96 7 VSS
port 6 w
rlabel locali 427 0 444 0 5 row_n
port 7 s
rlabel metal4 92 467 122 467 1 ctop
port 1 n
rlabel metal2 209 486 258 486 1 cbot
rlabel metal1 0 187 0 201 7 sample_i
port 12 w
rlabel metal1 0 370 0 385 7 sample_n_i
port 13 w
rlabel metal1 502 370 502 385 3 sample_n_o
port 14 e
rlabel metal1 502 187 502 201 3 sample_o
port 15 e
<< end >>
