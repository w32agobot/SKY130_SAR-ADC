magic
tech sky130A
magscale 1 2
timestamp 1661178173
<< error_p >>
rect -70 50 -10 2250
rect 10 50 70 2250
rect -70 -2250 -10 -50
rect 10 -2250 70 -50
<< metal3 >>
rect -1509 2222 -10 2250
rect -1509 78 -94 2222
rect -30 78 -10 2222
rect -1509 50 -10 78
rect 10 2222 1509 2250
rect 10 78 1425 2222
rect 1489 78 1509 2222
rect 10 50 1509 78
rect -1509 -78 -10 -50
rect -1509 -2222 -94 -78
rect -30 -2222 -10 -78
rect -1509 -2250 -10 -2222
rect 10 -78 1509 -50
rect 10 -2222 1425 -78
rect 1489 -2222 1509 -78
rect 10 -2250 1509 -2222
<< via3 >>
rect -94 78 -30 2222
rect 1425 78 1489 2222
rect -94 -2222 -30 -78
rect 1425 -2222 1489 -78
<< mimcap >>
rect -1409 2110 -209 2150
rect -1409 190 -1369 2110
rect -249 190 -209 2110
rect -1409 150 -209 190
rect 110 2110 1310 2150
rect 110 190 150 2110
rect 1270 190 1310 2110
rect 110 150 1310 190
rect -1409 -190 -209 -150
rect -1409 -2110 -1369 -190
rect -249 -2110 -209 -190
rect -1409 -2150 -209 -2110
rect 110 -190 1310 -150
rect 110 -2110 150 -190
rect 1270 -2110 1310 -190
rect 110 -2150 1310 -2110
<< mimcapcontact >>
rect -1369 190 -249 2110
rect 150 190 1270 2110
rect -1369 -2110 -249 -190
rect 150 -2110 1270 -190
<< metal4 >>
rect -861 2111 -757 2300
rect -141 2238 -37 2300
rect -141 2222 -14 2238
rect -1370 2110 -248 2111
rect -1370 190 -1369 2110
rect -249 190 -248 2110
rect -1370 189 -248 190
rect -861 -189 -757 189
rect -141 78 -94 2222
rect -30 78 -14 2222
rect 658 2111 762 2300
rect 1378 2238 1482 2300
rect 1378 2222 1505 2238
rect 149 2110 1271 2111
rect 149 190 150 2110
rect 1270 190 1271 2110
rect 149 189 1271 190
rect -141 62 -14 78
rect -141 -62 -37 62
rect -141 -78 -14 -62
rect -1370 -190 -248 -189
rect -1370 -2110 -1369 -190
rect -249 -2110 -248 -190
rect -1370 -2111 -248 -2110
rect -861 -2300 -757 -2111
rect -141 -2222 -94 -78
rect -30 -2222 -14 -78
rect 658 -189 762 189
rect 1378 78 1425 2222
rect 1489 78 1505 2222
rect 1378 62 1505 78
rect 1378 -62 1482 62
rect 1378 -78 1505 -62
rect 149 -190 1271 -189
rect 149 -2110 150 -190
rect 1270 -2110 1271 -190
rect 149 -2111 1271 -2110
rect -141 -2238 -14 -2222
rect -141 -2300 -37 -2238
rect 658 -2300 762 -2111
rect 1378 -2222 1425 -78
rect 1489 -2222 1505 -78
rect 1378 -2238 1505 -2222
rect 1378 -2300 1482 -2238
<< properties >>
string FIXED_BBOX 10 50 1410 2250
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 6 l 10 val 126.08 carea 2.00 cperi 0.19 nx 2 ny 2 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
