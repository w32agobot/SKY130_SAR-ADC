magic
tech sky130A
timestamp 1666978453
<< metal1 >>
rect 0 0 4500 4500
<< properties >>
string FIXED_BBOX 0 0 4500 4500
string LEFclass BLOCK
string LEForigin 0 0
string LEFsource USER
<< end >>
