magic
tech sky130A
magscale 1 2
timestamp 1679612785
<< nwell >>
rect 0 464 1004 880
<< nmos >>
rect 227 236 257 356
rect 431 236 461 356
rect 632 236 662 356
rect 745 236 775 356
<< pmos >>
rect 227 502 257 742
rect 431 502 461 742
rect 632 502 662 742
rect 745 502 775 742
<< ndiff >>
rect 170 348 227 356
rect 170 244 182 348
rect 216 244 227 348
rect 170 236 227 244
rect 257 348 314 356
rect 257 244 268 348
rect 302 244 314 348
rect 257 236 314 244
rect 374 279 431 356
rect 374 244 386 279
rect 420 244 431 279
rect 374 236 431 244
rect 461 334 518 356
rect 461 244 472 334
rect 506 244 518 334
rect 461 236 518 244
rect 575 336 632 356
rect 575 244 587 336
rect 621 244 632 336
rect 575 236 632 244
rect 662 278 745 356
rect 662 244 673 278
rect 734 244 745 278
rect 662 236 745 244
rect 775 334 832 356
rect 775 244 786 334
rect 820 244 832 334
rect 775 236 832 244
<< pdiff >>
rect 170 734 227 742
rect 170 518 182 734
rect 216 518 227 734
rect 170 502 227 518
rect 257 734 314 742
rect 257 518 268 734
rect 302 518 314 734
rect 257 502 314 518
rect 374 734 431 742
rect 374 586 386 734
rect 420 586 431 734
rect 374 502 431 586
rect 461 734 518 742
rect 461 518 472 734
rect 506 518 518 734
rect 461 502 518 518
rect 575 734 632 742
rect 575 518 587 734
rect 621 518 632 734
rect 575 502 632 518
rect 662 734 745 742
rect 662 586 673 734
rect 734 586 745 734
rect 662 502 745 586
rect 775 734 832 742
rect 775 518 786 734
rect 820 518 832 734
rect 775 502 832 518
<< ndiffc >>
rect 182 244 216 348
rect 268 244 302 348
rect 386 244 420 279
rect 472 244 506 334
rect 587 244 621 336
rect 673 244 734 278
rect 786 244 820 334
<< pdiffc >>
rect 182 518 216 734
rect 268 518 302 734
rect 386 586 420 734
rect 472 518 506 734
rect 587 518 621 734
rect 673 586 734 734
rect 786 518 820 734
<< psubdiff >>
rect 279 148 326 182
rect 360 148 430 182
rect 464 148 534 182
rect 568 148 628 182
rect 662 148 726 182
rect 760 148 792 182
<< nsubdiff >>
rect 198 838 302 844
rect 198 804 222 838
rect 256 804 302 838
rect 198 798 302 804
rect 414 838 806 844
rect 414 804 441 838
rect 475 804 534 838
rect 568 804 630 838
rect 664 804 724 838
rect 758 804 806 838
rect 414 798 806 804
<< psubdiffcont >>
rect 326 148 360 182
rect 430 148 464 182
rect 534 148 568 182
rect 628 148 662 182
rect 726 148 760 182
<< nsubdiffcont >>
rect 222 804 256 838
rect 441 804 475 838
rect 534 804 568 838
rect 630 804 664 838
rect 724 804 758 838
<< poly >>
rect 324 838 390 848
rect 324 804 340 838
rect 374 804 390 838
rect 324 794 390 804
rect 227 742 257 770
rect 227 486 257 502
rect 125 456 257 486
rect 125 168 155 456
rect 329 414 359 794
rect 431 742 461 770
rect 632 742 662 770
rect 745 742 775 770
rect 431 463 461 502
rect 632 487 662 502
rect 227 384 359 414
rect 401 434 461 463
rect 556 457 662 487
rect 745 474 775 502
rect 556 452 587 457
rect 401 400 415 434
rect 449 400 461 434
rect 401 384 461 400
rect 503 441 587 452
rect 503 407 519 441
rect 553 407 587 441
rect 503 401 587 407
rect 704 436 775 474
rect 704 402 714 436
rect 748 402 775 436
rect 503 396 662 401
rect 227 356 257 384
rect 431 356 461 384
rect 556 371 662 396
rect 704 371 775 402
rect 632 356 662 371
rect 745 356 775 371
rect 227 210 257 236
rect 431 210 461 236
rect 632 210 662 236
rect 745 210 775 236
rect 125 158 256 168
rect 125 124 198 158
rect 232 124 256 158
rect 125 112 256 124
<< polycont >>
rect 340 804 374 838
rect 415 400 449 434
rect 519 407 553 441
rect 714 402 748 436
rect 198 124 232 158
<< locali >>
rect 34 922 182 1004
rect 34 888 48 922
rect 136 888 182 922
rect 34 882 182 888
rect 910 922 970 1004
rect 910 888 922 922
rect 956 888 970 922
rect 910 882 970 888
rect 34 706 148 882
rect 182 838 820 844
rect 182 804 222 838
rect 256 804 340 838
rect 374 804 441 838
rect 475 804 534 838
rect 568 804 630 838
rect 664 804 724 838
rect 758 804 820 838
rect 182 798 820 804
rect 34 630 48 706
rect 130 630 148 706
rect 34 340 148 630
rect 34 292 48 340
rect 132 292 148 340
rect 34 102 148 292
rect 182 734 216 750
rect 182 390 216 518
rect 182 228 216 244
rect 268 734 302 750
rect 386 734 420 798
rect 386 570 420 586
rect 472 734 506 750
rect 268 348 302 518
rect 471 518 472 536
rect 587 734 621 750
rect 506 518 517 530
rect 471 502 517 518
rect 483 457 517 502
rect 673 734 734 798
rect 673 570 734 586
rect 786 734 820 750
rect 415 434 449 450
rect 445 387 449 400
rect 415 384 449 387
rect 483 441 553 457
rect 483 407 519 441
rect 483 391 553 407
rect 483 350 517 391
rect 472 334 517 350
rect 370 244 386 279
rect 420 244 436 279
rect 506 319 517 334
rect 587 336 621 518
rect 692 436 752 474
rect 692 417 714 436
rect 692 383 702 417
rect 748 402 752 436
rect 736 383 752 402
rect 692 371 752 383
rect 268 227 302 244
rect 386 182 420 244
rect 472 228 506 244
rect 786 334 820 518
rect 587 228 621 244
rect 655 244 673 278
rect 734 244 752 278
rect 655 236 752 244
rect 673 182 734 236
rect 786 228 820 244
rect 182 124 198 182
rect 232 148 326 182
rect 360 148 430 182
rect 464 148 534 182
rect 568 148 628 182
rect 662 148 726 182
rect 760 148 814 182
rect 232 124 248 148
rect 854 108 970 882
rect 34 68 46 102
rect 136 90 148 102
rect 910 102 970 108
rect 136 68 182 90
rect 34 0 182 68
rect 910 68 922 102
rect 958 68 970 102
rect 910 0 970 68
<< viali >>
rect 48 888 136 922
rect 922 888 956 922
rect 222 804 256 838
rect 340 804 374 838
rect 441 804 475 838
rect 534 804 568 838
rect 630 804 664 838
rect 724 804 758 838
rect 48 630 130 706
rect 48 292 132 340
rect 182 348 216 390
rect 182 340 216 348
rect 786 663 820 701
rect 411 400 415 421
rect 415 400 445 421
rect 411 387 445 400
rect 268 298 302 337
rect 702 402 714 417
rect 714 402 736 417
rect 702 383 736 402
rect 587 293 621 327
rect 198 158 232 182
rect 198 148 232 158
rect 326 148 360 182
rect 430 148 464 182
rect 534 148 568 182
rect 628 148 662 182
rect 726 148 760 182
rect 46 68 136 102
rect 922 68 958 102
<< metal1 >>
rect 34 922 182 1004
rect 34 888 48 922
rect 136 888 182 922
rect 34 882 182 888
rect 910 922 970 1004
rect 910 888 922 922
rect 956 888 970 922
rect 910 882 970 888
rect 0 838 1004 854
rect 0 804 222 838
rect 256 804 340 838
rect 374 804 441 838
rect 475 804 534 838
rect 568 804 630 838
rect 664 804 724 838
rect 758 804 1004 838
rect 0 798 1004 804
rect 0 740 158 770
rect 780 740 1004 770
rect 34 706 142 712
rect 34 630 48 706
rect 130 630 142 706
rect 780 701 826 740
rect 780 663 786 701
rect 820 663 826 701
rect 780 651 826 663
rect 34 624 142 630
rect 0 568 1004 596
rect 0 512 1004 540
rect 121 458 865 483
rect 0 455 1004 458
rect 0 430 158 455
rect 837 430 1004 455
rect 187 421 457 427
rect 187 402 411 421
rect 0 399 411 402
rect 0 390 222 399
rect 0 374 182 390
rect 34 340 144 346
rect 34 292 48 340
rect 132 292 144 340
rect 176 340 182 374
rect 216 340 222 390
rect 399 387 411 399
rect 445 387 457 421
rect 399 381 457 387
rect 485 417 751 427
rect 485 399 702 417
rect 485 351 513 399
rect 690 383 702 399
rect 736 383 751 417
rect 690 371 751 383
rect 799 374 1004 402
rect 176 328 222 340
rect 260 337 513 351
rect 34 286 144 292
rect 260 298 268 337
rect 302 313 513 337
rect 799 333 827 374
rect 575 327 827 333
rect 302 298 308 313
rect 260 286 308 298
rect 575 293 587 327
rect 621 305 827 327
rect 621 293 635 305
rect 575 286 635 293
rect 0 220 1004 258
rect 0 182 1004 192
rect 0 148 198 182
rect 232 148 326 182
rect 360 148 430 182
rect 464 148 534 182
rect 568 148 628 182
rect 662 148 726 182
rect 760 148 1004 182
rect 0 136 1004 148
rect 34 102 182 108
rect 34 68 46 102
rect 136 68 182 102
rect 34 0 182 68
rect 910 102 970 108
rect 910 68 922 102
rect 958 68 970 102
rect 910 0 970 68
<< metal2 >>
rect 32 962 972 972
rect 32 906 42 962
rect 98 906 138 962
rect 194 906 234 962
rect 290 906 330 962
rect 386 906 426 962
rect 482 906 522 962
rect 578 906 618 962
rect 674 906 714 962
rect 770 906 810 962
rect 866 906 906 962
rect 962 906 972 962
rect 32 866 972 906
rect 32 810 42 866
rect 98 810 330 866
rect 386 810 618 866
rect 674 810 906 866
rect 962 810 972 866
rect 32 770 972 810
rect 32 714 42 770
rect 98 714 330 770
rect 386 714 618 770
rect 674 714 906 770
rect 962 714 972 770
rect 32 674 972 714
rect 32 618 42 674
rect 98 618 138 674
rect 194 618 234 674
rect 290 618 330 674
rect 386 618 426 674
rect 482 618 522 674
rect 578 618 618 674
rect 674 618 714 674
rect 770 618 810 674
rect 866 618 906 674
rect 962 618 972 674
rect 32 608 972 618
rect 32 578 396 608
rect 32 522 42 578
rect 98 522 330 578
rect 386 522 396 578
rect 608 578 972 608
rect 32 482 396 522
rect 32 426 42 482
rect 98 426 330 482
rect 386 426 396 482
rect 460 460 544 544
rect 608 522 618 578
rect 674 522 906 578
rect 962 522 972 578
rect 608 482 972 522
rect 32 396 396 426
rect 608 426 618 482
rect 674 426 906 482
rect 962 426 972 482
rect 608 396 972 426
rect 32 386 972 396
rect 32 330 42 386
rect 98 330 138 386
rect 194 330 234 386
rect 290 330 330 386
rect 386 330 426 386
rect 482 330 522 386
rect 578 330 618 386
rect 674 330 714 386
rect 770 330 810 386
rect 866 330 906 386
rect 962 330 972 386
rect 32 290 972 330
rect 32 234 42 290
rect 98 234 330 290
rect 386 234 618 290
rect 674 234 906 290
rect 962 234 972 290
rect 32 194 972 234
rect 32 138 42 194
rect 98 138 330 194
rect 386 138 618 194
rect 674 138 906 194
rect 962 138 972 194
rect 32 98 972 138
rect 32 42 42 98
rect 98 42 138 98
rect 194 42 234 98
rect 290 42 330 98
rect 386 42 426 98
rect 482 42 522 98
rect 578 42 618 98
rect 674 42 714 98
rect 770 42 810 98
rect 866 42 906 98
rect 962 42 972 98
rect 32 32 972 42
<< via2 >>
rect 42 906 98 962
rect 138 906 194 962
rect 234 906 290 962
rect 330 906 386 962
rect 426 906 482 962
rect 522 906 578 962
rect 618 906 674 962
rect 714 906 770 962
rect 810 906 866 962
rect 906 906 962 962
rect 42 810 98 866
rect 330 810 386 866
rect 618 810 674 866
rect 906 810 962 866
rect 42 714 98 770
rect 330 714 386 770
rect 618 714 674 770
rect 906 714 962 770
rect 42 618 98 674
rect 138 618 194 674
rect 234 618 290 674
rect 330 618 386 674
rect 426 618 482 674
rect 522 618 578 674
rect 618 618 674 674
rect 714 618 770 674
rect 810 618 866 674
rect 906 618 962 674
rect 42 522 98 578
rect 330 522 386 578
rect 42 426 98 482
rect 330 426 386 482
rect 618 522 674 578
rect 906 522 962 578
rect 618 426 674 482
rect 906 426 962 482
rect 42 330 98 386
rect 138 330 194 386
rect 234 330 290 386
rect 330 330 386 386
rect 426 330 482 386
rect 522 330 578 386
rect 618 330 674 386
rect 714 330 770 386
rect 810 330 866 386
rect 906 330 962 386
rect 42 234 98 290
rect 330 234 386 290
rect 618 234 674 290
rect 906 234 962 290
rect 42 138 98 194
rect 330 138 386 194
rect 618 138 674 194
rect 906 138 962 194
rect 42 42 98 98
rect 138 42 194 98
rect 234 42 290 98
rect 330 42 386 98
rect 426 42 482 98
rect 522 42 578 98
rect 618 42 674 98
rect 714 42 770 98
rect 810 42 866 98
rect 906 42 962 98
<< metal3 >>
rect 36 962 968 968
rect 36 906 42 962
rect 98 906 138 962
rect 194 906 234 962
rect 290 906 330 962
rect 386 906 426 962
rect 482 906 522 962
rect 578 906 618 962
rect 674 906 714 962
rect 770 906 810 962
rect 866 906 906 962
rect 962 906 968 962
rect 36 900 968 906
rect 36 866 104 900
rect 36 810 42 866
rect 98 810 104 866
rect 324 866 392 900
rect 36 770 104 810
rect 36 714 42 770
rect 98 714 104 770
rect 164 824 264 840
rect 164 756 180 824
rect 248 756 264 824
rect 164 740 264 756
rect 324 810 330 866
rect 386 810 392 866
rect 612 866 680 900
rect 324 770 392 810
rect 36 680 104 714
rect 324 714 330 770
rect 386 714 392 770
rect 452 824 552 840
rect 452 756 468 824
rect 536 756 552 824
rect 452 740 552 756
rect 612 810 618 866
rect 674 810 680 866
rect 900 866 968 900
rect 612 770 680 810
rect 324 680 392 714
rect 612 714 618 770
rect 674 714 680 770
rect 740 824 840 840
rect 740 756 756 824
rect 824 756 840 824
rect 740 740 840 756
rect 900 810 906 866
rect 962 810 968 866
rect 900 770 968 810
rect 612 680 680 714
rect 900 714 906 770
rect 962 714 968 770
rect 900 680 968 714
rect 36 674 968 680
rect 36 618 42 674
rect 98 618 138 674
rect 194 618 234 674
rect 290 618 330 674
rect 386 618 426 674
rect 482 618 522 674
rect 578 618 618 674
rect 674 618 714 674
rect 770 618 810 674
rect 866 618 906 674
rect 962 618 968 674
rect 36 612 968 618
rect 36 578 104 612
rect 36 522 42 578
rect 98 522 104 578
rect 324 578 392 612
rect 36 482 104 522
rect 36 426 42 482
rect 98 426 104 482
rect 164 536 264 552
rect 164 468 180 536
rect 248 468 264 536
rect 164 452 264 468
rect 324 522 330 578
rect 386 522 392 578
rect 324 482 392 522
rect 36 392 104 426
rect 324 426 330 482
rect 386 426 392 482
rect 324 392 392 426
rect 612 578 680 612
rect 612 522 618 578
rect 674 522 680 578
rect 900 578 968 612
rect 612 482 680 522
rect 612 426 618 482
rect 674 426 680 482
rect 740 536 840 552
rect 740 468 756 536
rect 824 468 840 536
rect 740 452 840 468
rect 900 522 906 578
rect 962 522 968 578
rect 900 482 968 522
rect 612 392 680 426
rect 900 426 906 482
rect 962 426 968 482
rect 900 392 968 426
rect 36 386 968 392
rect 36 330 42 386
rect 98 330 138 386
rect 194 330 234 386
rect 290 330 330 386
rect 386 330 426 386
rect 482 330 522 386
rect 578 330 618 386
rect 674 330 714 386
rect 770 330 810 386
rect 866 330 906 386
rect 962 330 968 386
rect 36 324 968 330
rect 36 290 104 324
rect 36 234 42 290
rect 98 234 104 290
rect 324 290 392 324
rect 36 194 104 234
rect 36 138 42 194
rect 98 138 104 194
rect 164 248 264 264
rect 164 180 180 248
rect 248 180 264 248
rect 164 164 264 180
rect 324 234 330 290
rect 386 234 392 290
rect 612 290 680 324
rect 324 194 392 234
rect 36 104 104 138
rect 324 138 330 194
rect 386 138 392 194
rect 452 248 552 264
rect 452 180 468 248
rect 536 180 552 248
rect 452 164 552 180
rect 612 234 618 290
rect 674 234 680 290
rect 900 290 968 324
rect 612 194 680 234
rect 324 104 392 138
rect 612 138 618 194
rect 674 138 680 194
rect 740 248 840 264
rect 740 180 756 248
rect 824 180 840 248
rect 740 164 840 180
rect 900 234 906 290
rect 962 234 968 290
rect 900 194 968 234
rect 612 104 680 138
rect 900 138 906 194
rect 962 138 968 194
rect 900 104 968 138
rect 36 98 968 104
rect 36 42 42 98
rect 98 42 138 98
rect 194 42 234 98
rect 290 42 330 98
rect 386 42 426 98
rect 482 42 522 98
rect 578 42 618 98
rect 674 42 714 98
rect 770 42 810 98
rect 866 42 906 98
rect 962 42 968 98
rect 36 36 968 42
<< via3 >>
rect 180 756 248 824
rect 468 756 536 824
rect 756 756 824 824
rect 180 468 248 536
rect 756 468 824 536
rect 180 180 248 248
rect 468 180 536 248
rect 756 180 824 248
<< metal4 >>
rect 184 840 244 934
rect 472 840 532 934
rect 760 840 820 934
rect 164 824 264 840
rect 164 820 180 824
rect 70 760 180 820
rect 164 756 180 760
rect 248 820 264 824
rect 452 824 552 840
rect 452 820 468 824
rect 248 760 468 820
rect 248 756 264 760
rect 164 740 264 756
rect 452 756 468 760
rect 536 820 552 824
rect 740 824 840 840
rect 740 820 756 824
rect 536 760 756 820
rect 536 756 552 760
rect 452 740 552 756
rect 740 756 756 760
rect 824 820 840 824
rect 824 760 934 820
rect 824 756 840 760
rect 740 740 840 756
rect 184 552 244 740
rect 472 646 532 740
rect 760 552 820 740
rect 164 536 264 552
rect 164 532 180 536
rect 70 472 180 532
rect 164 468 180 472
rect 248 532 264 536
rect 740 536 840 552
rect 740 532 756 536
rect 248 472 358 532
rect 646 472 756 532
rect 248 468 264 472
rect 164 452 264 468
rect 740 468 756 472
rect 824 532 840 536
rect 824 472 934 532
rect 824 468 840 472
rect 740 452 840 468
rect 184 264 244 452
rect 472 264 532 358
rect 760 264 820 452
rect 164 248 264 264
rect 164 244 180 248
rect 70 184 180 244
rect 164 180 180 184
rect 248 244 264 248
rect 452 248 552 264
rect 452 244 468 248
rect 248 184 468 244
rect 248 180 264 184
rect 164 164 264 180
rect 452 180 468 184
rect 536 244 552 248
rect 740 248 840 264
rect 740 244 756 248
rect 536 184 756 244
rect 536 180 552 184
rect 452 164 552 180
rect 740 180 756 184
rect 824 244 840 248
rect 824 184 934 244
rect 824 180 840 184
rect 740 164 840 180
rect 184 70 244 164
rect 472 70 532 164
rect 760 70 820 164
<< comment >>
rect 0 972 32 1004
rect 972 972 1004 1004
rect 138 750 308 798
rect 430 756 562 804
rect 138 260 194 750
rect 312 690 368 750
rect 358 428 406 688
rect 430 562 478 756
rect 564 716 606 762
rect 598 608 632 716
rect 576 604 632 608
rect 558 602 632 604
rect 558 576 608 602
rect 544 562 600 576
rect 430 558 600 562
rect 430 544 576 558
rect 430 514 558 544
rect 430 460 478 514
rect 560 478 602 522
rect 560 476 636 478
rect 428 428 478 460
rect 358 396 428 428
rect 300 260 356 318
rect 358 314 406 396
rect 138 258 356 260
rect 138 212 306 258
rect 430 206 478 428
rect 602 198 636 476
rect 670 198 716 802
rect 0 0 32 32
rect 972 0 1004 32
<< labels >>
flabel metal1 837 798 1004 854 0 FreeSans 160 0 0 0 VDD
port 1 e power bidirectional
flabel metal1 0 136 1004 192 0 FreeSans 320 0 0 0 VSS
port 2 nsew ground bidirectional
flabel metal4 472 874 532 934 1 FreeSans 160 0 0 0 ctop
port 4 n
flabel metal1 34 0 182 108 5 FreeSans 320 0 0 0 col
port 5 s
flabel metal1 34 882 182 1004 1 FreeSans 320 0 0 0 col
port 5 n
flabel metal1 910 882 970 1004 1 FreeSans 320 0 0 0 col_n
port 6 n
flabel metal1 846 430 1004 458 0 FreeSans 160 0 0 0 row_n
port 7 e
flabel metal1 0 512 155 540 0 FreeSans 160 0 0 0 rowon_n
port 8 w
flabel metal1 849 512 1004 540 0 FreeSans 160 0 0 0 rowon_n
port 8 e
flabel metal1 846 374 1004 402 0 FreeSans 160 0 0 0 sample_o
port 10 e
flabel metal1 846 740 1004 770 0 FreeSans 160 0 0 0 sample_n_o
port 12 nsew
flabel metal1 0 568 156 596 7 FreeSans 160 0 0 0 off_n
port 13 w
flabel metal1 848 568 1004 596 3 FreeSans 160 0 0 0 off_n
port 13 e
rlabel metal2 500 972 500 972 1 cbot
flabel metal1 910 0 970 108 1 FreeSans 320 0 0 0 col_n
port 6 s
flabel metal1 0 798 167 854 0 FreeSans 160 0 0 0 VDD
port 1 w power bidirectional
flabel metal1 0 740 158 770 0 FreeSans 160 0 0 0 sample_n_i
port 11 nsew
flabel metal1 0 374 158 402 0 FreeSans 160 0 0 0 sample_i
port 9 w
flabel metal1 0 430 158 458 0 FreeSans 160 0 0 0 row_n
port 7 w
flabel metal1 0 220 1004 258 0 FreeSans 320 0 0 0 vcom
port 3 nsew
<< end >>
