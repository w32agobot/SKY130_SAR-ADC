* SPICE3 file created from adc_array_fingercap_8(8)x392aF_23um2.ext - technology: sky130A

C0 ctop cbot 3.66fF
C1 ctop VSUBS 0.55fF
C2 cbot VSUBS 1.90fF
