* SPICE3 file created from extract.ext - technology: sky130A

C0 dummy_bot bot_2 14.82fF
C1 dummy_bot bot_8 12.90fF
C2 top_1 bot_1 30.59fF
C3 dummy_bot bot_1 14.82fF
C4 bot_4 dummy_bot 14.82fF
C5 bot_1 m4_11832_164# 3.62fF
C6 dummy_bot dummy_top 269.06fF
C7 top_8 bot_8 29.82fF
C8 bot_2 m4_8352_164# 3.55fF
C9 bot_4 top_4 32.51fF
C10 top_2 bot_2 31.19fF
C11 bot_4 m4_4872_164# 2.41fF
C12 dummy_top VSUBS 3.52fF
C13 bot_1 VSUBS 2.68fF
C14 bot_2 VSUBS 2.68fF
C15 bot_4 VSUBS 2.68fF
C16 bot_8 VSUBS 2.07fF
C17 dummy_bot VSUBS 33.21fF
