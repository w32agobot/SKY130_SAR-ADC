magic
tech sky130A
timestamp 1661762619
<< metal2 >>
rect 14 2245 334 2250
rect 14 2213 19 2245
rect 51 2213 297 2245
rect 329 2213 334 2245
rect 14 2121 334 2213
rect 14 2089 19 2121
rect 51 2089 297 2121
rect 329 2089 334 2121
rect 14 1997 334 2089
rect 14 1965 19 1997
rect 51 1965 297 1997
rect 329 1978 334 1997
rect 362 2245 682 2250
rect 362 2213 367 2245
rect 399 2213 645 2245
rect 677 2213 682 2245
rect 362 2121 682 2213
rect 362 2089 367 2121
rect 399 2089 645 2121
rect 677 2089 682 2121
rect 362 1997 682 2089
rect 362 1978 367 1997
rect 329 1965 367 1978
rect 399 1965 645 1997
rect 677 1978 682 1997
rect 710 2245 1030 2250
rect 710 2213 715 2245
rect 747 2213 993 2245
rect 1025 2213 1030 2245
rect 710 2121 1030 2213
rect 710 2089 715 2121
rect 747 2089 993 2121
rect 1025 2089 1030 2121
rect 710 1997 1030 2089
rect 710 1978 715 1997
rect 677 1965 715 1978
rect 747 1965 993 1997
rect 1025 1978 1030 1997
rect 1058 2245 1378 2250
rect 1058 2213 1063 2245
rect 1095 2213 1341 2245
rect 1373 2213 1378 2245
rect 1058 2121 1378 2213
rect 1058 2089 1063 2121
rect 1095 2089 1341 2121
rect 1373 2089 1378 2121
rect 1058 1997 1378 2089
rect 1058 1978 1063 1997
rect 1025 1965 1063 1978
rect 1095 1965 1341 1997
rect 1373 1978 1378 1997
rect 1406 2245 1726 2250
rect 1406 2213 1411 2245
rect 1443 2213 1689 2245
rect 1721 2213 1726 2245
rect 1406 2121 1726 2213
rect 1406 2089 1411 2121
rect 1443 2089 1689 2121
rect 1721 2089 1726 2121
rect 1406 1997 1726 2089
rect 1406 1978 1411 1997
rect 1373 1965 1411 1978
rect 1443 1965 1689 1997
rect 1721 1978 1726 1997
rect 1754 2245 2074 2250
rect 1754 2213 1759 2245
rect 1791 2213 2037 2245
rect 2069 2213 2074 2245
rect 1754 2121 2074 2213
rect 1754 2089 1759 2121
rect 1791 2089 2037 2121
rect 2069 2089 2074 2121
rect 1754 1997 2074 2089
rect 1754 1978 1759 1997
rect 1721 1965 1759 1978
rect 1791 1965 2037 1997
rect 2069 1978 2074 1997
rect 2102 2245 2422 2250
rect 2102 2213 2107 2245
rect 2139 2213 2385 2245
rect 2417 2213 2422 2245
rect 2102 2121 2422 2213
rect 2102 2089 2107 2121
rect 2139 2089 2385 2121
rect 2417 2089 2422 2121
rect 2102 1997 2422 2089
rect 2102 1978 2107 1997
rect 2069 1965 2107 1978
rect 2139 1965 2385 1997
rect 2417 1978 2422 1997
rect 2450 2245 2770 2250
rect 2450 2213 2455 2245
rect 2487 2213 2733 2245
rect 2765 2213 2770 2245
rect 2450 2121 2770 2213
rect 2450 2089 2455 2121
rect 2487 2089 2733 2121
rect 2765 2089 2770 2121
rect 2450 1997 2770 2089
rect 2450 1978 2455 1997
rect 2417 1965 2455 1978
rect 2487 1965 2733 1997
rect 2765 1978 2770 1997
rect 2798 2245 3118 2250
rect 2798 2213 2803 2245
rect 2835 2213 3081 2245
rect 3113 2213 3118 2245
rect 2798 2121 3118 2213
rect 2798 2089 2803 2121
rect 2835 2089 3081 2121
rect 3113 2089 3118 2121
rect 2798 1997 3118 2089
rect 2798 1978 2803 1997
rect 2765 1965 2803 1978
rect 2835 1965 3081 1997
rect 3113 1978 3118 1997
rect 3146 2245 3466 2250
rect 3146 2213 3151 2245
rect 3183 2213 3429 2245
rect 3461 2213 3466 2245
rect 3146 2121 3466 2213
rect 3146 2089 3151 2121
rect 3183 2089 3429 2121
rect 3461 2089 3466 2121
rect 3146 1997 3466 2089
rect 3146 1978 3151 1997
rect 3113 1965 3151 1978
rect 3183 1965 3429 1997
rect 3461 1978 3466 1997
rect 3494 2245 3814 2250
rect 3494 2213 3499 2245
rect 3531 2213 3777 2245
rect 3809 2213 3814 2245
rect 3494 2121 3814 2213
rect 3494 2089 3499 2121
rect 3531 2089 3777 2121
rect 3809 2089 3814 2121
rect 3494 1997 3814 2089
rect 3494 1978 3499 1997
rect 3461 1965 3499 1978
rect 3531 1965 3777 1997
rect 3809 1978 3814 1997
rect 3842 2245 4162 2250
rect 3842 2213 3847 2245
rect 3879 2213 4125 2245
rect 4157 2213 4162 2245
rect 3842 2121 4162 2213
rect 3842 2089 3847 2121
rect 3879 2089 4125 2121
rect 4157 2089 4162 2121
rect 3842 1997 4162 2089
rect 3842 1978 3847 1997
rect 3809 1965 3847 1978
rect 3879 1965 4125 1997
rect 4157 1978 4162 1997
rect 4190 2245 4510 2250
rect 4190 2213 4195 2245
rect 4227 2213 4473 2245
rect 4505 2213 4510 2245
rect 4190 2121 4510 2213
rect 4190 2089 4195 2121
rect 4227 2089 4473 2121
rect 4505 2089 4510 2121
rect 4190 1997 4510 2089
rect 4190 1978 4195 1997
rect 4157 1965 4195 1978
rect 4227 1965 4473 1997
rect 4505 1978 4510 1997
rect 4538 2245 4858 2250
rect 4538 2213 4543 2245
rect 4575 2213 4821 2245
rect 4853 2213 4858 2245
rect 4538 2121 4858 2213
rect 4538 2089 4543 2121
rect 4575 2089 4821 2121
rect 4853 2089 4858 2121
rect 4538 1997 4858 2089
rect 4538 1978 4543 1997
rect 4505 1965 4543 1978
rect 4575 1965 4821 1997
rect 4853 1978 4858 1997
rect 4886 2245 5206 2250
rect 4886 2213 4891 2245
rect 4923 2213 5169 2245
rect 5201 2213 5206 2245
rect 4886 2121 5206 2213
rect 4886 2089 4891 2121
rect 4923 2089 5169 2121
rect 5201 2089 5206 2121
rect 4886 1997 5206 2089
rect 4886 1978 4891 1997
rect 4853 1965 4891 1978
rect 4923 1965 5169 1997
rect 5201 1978 5206 1997
rect 5234 2245 5554 2250
rect 5234 2213 5239 2245
rect 5271 2213 5517 2245
rect 5549 2213 5554 2245
rect 5234 2121 5554 2213
rect 5234 2089 5239 2121
rect 5271 2089 5517 2121
rect 5549 2089 5554 2121
rect 5234 1997 5554 2089
rect 5234 1978 5239 1997
rect 5201 1965 5239 1978
rect 5271 1965 5517 1997
rect 5549 1978 5554 1997
rect 5582 2245 5902 2250
rect 5582 2213 5587 2245
rect 5619 2213 5865 2245
rect 5897 2213 5902 2245
rect 5582 2121 5902 2213
rect 5582 2089 5587 2121
rect 5619 2089 5865 2121
rect 5897 2089 5902 2121
rect 5582 1997 5902 2089
rect 5582 1978 5587 1997
rect 5549 1965 5587 1978
rect 5619 1965 5865 1997
rect 5897 1978 5902 1997
rect 5930 2245 6250 2250
rect 5930 2213 5935 2245
rect 5967 2213 6213 2245
rect 6245 2213 6250 2245
rect 5930 2121 6250 2213
rect 5930 2089 5935 2121
rect 5967 2089 6213 2121
rect 6245 2089 6250 2121
rect 5930 1997 6250 2089
rect 5930 1978 5935 1997
rect 5897 1965 5935 1978
rect 5967 1965 6213 1997
rect 6245 1978 6250 1997
rect 6278 2245 6598 2250
rect 6278 2213 6283 2245
rect 6315 2213 6561 2245
rect 6593 2213 6598 2245
rect 6278 2121 6598 2213
rect 6278 2089 6283 2121
rect 6315 2089 6561 2121
rect 6593 2089 6598 2121
rect 6278 1997 6598 2089
rect 6278 1978 6283 1997
rect 6245 1965 6283 1978
rect 6315 1965 6561 1997
rect 6593 1978 6598 1997
rect 6626 2245 6946 2250
rect 6626 2213 6631 2245
rect 6663 2213 6909 2245
rect 6941 2213 6946 2245
rect 6626 2121 6946 2213
rect 6626 2089 6631 2121
rect 6663 2089 6909 2121
rect 6941 2089 6946 2121
rect 6626 1997 6946 2089
rect 6626 1978 6631 1997
rect 6593 1965 6631 1978
rect 6663 1965 6909 1997
rect 6941 1965 6946 1997
rect 14 1964 6946 1965
rect 14 1873 334 1964
rect 14 1841 19 1873
rect 51 1841 297 1873
rect 329 1841 334 1873
rect 14 1749 334 1841
rect 14 1717 19 1749
rect 51 1717 297 1749
rect 329 1717 334 1749
rect 14 1712 334 1717
rect 362 1873 682 1964
rect 362 1841 367 1873
rect 399 1841 645 1873
rect 677 1841 682 1873
rect 362 1749 682 1841
rect 362 1717 367 1749
rect 399 1717 645 1749
rect 677 1717 682 1749
rect 362 1712 682 1717
rect 710 1873 1030 1964
rect 710 1841 715 1873
rect 747 1841 993 1873
rect 1025 1841 1030 1873
rect 710 1749 1030 1841
rect 710 1717 715 1749
rect 747 1717 993 1749
rect 1025 1717 1030 1749
rect 710 1712 1030 1717
rect 1058 1873 1378 1964
rect 1058 1841 1063 1873
rect 1095 1841 1341 1873
rect 1373 1841 1378 1873
rect 1058 1749 1378 1841
rect 1058 1717 1063 1749
rect 1095 1717 1341 1749
rect 1373 1717 1378 1749
rect 1058 1712 1378 1717
rect 1406 1873 1726 1964
rect 1406 1841 1411 1873
rect 1443 1841 1689 1873
rect 1721 1841 1726 1873
rect 1406 1749 1726 1841
rect 1406 1717 1411 1749
rect 1443 1717 1689 1749
rect 1721 1717 1726 1749
rect 1406 1712 1726 1717
rect 1754 1873 2074 1964
rect 1754 1841 1759 1873
rect 1791 1841 2037 1873
rect 2069 1841 2074 1873
rect 1754 1749 2074 1841
rect 1754 1717 1759 1749
rect 1791 1717 2037 1749
rect 2069 1717 2074 1749
rect 1754 1712 2074 1717
rect 2102 1873 2422 1964
rect 2102 1841 2107 1873
rect 2139 1841 2385 1873
rect 2417 1841 2422 1873
rect 2102 1749 2422 1841
rect 2102 1717 2107 1749
rect 2139 1717 2385 1749
rect 2417 1717 2422 1749
rect 2102 1712 2422 1717
rect 2450 1873 2770 1964
rect 2450 1841 2455 1873
rect 2487 1841 2733 1873
rect 2765 1841 2770 1873
rect 2450 1749 2770 1841
rect 2450 1717 2455 1749
rect 2487 1717 2733 1749
rect 2765 1717 2770 1749
rect 2450 1712 2770 1717
rect 2798 1873 3118 1964
rect 2798 1841 2803 1873
rect 2835 1841 3081 1873
rect 3113 1841 3118 1873
rect 2798 1749 3118 1841
rect 2798 1717 2803 1749
rect 2835 1717 3081 1749
rect 3113 1717 3118 1749
rect 2798 1712 3118 1717
rect 3146 1873 3466 1964
rect 3146 1841 3151 1873
rect 3183 1841 3429 1873
rect 3461 1841 3466 1873
rect 3146 1749 3466 1841
rect 3146 1717 3151 1749
rect 3183 1717 3429 1749
rect 3461 1717 3466 1749
rect 3146 1712 3466 1717
rect 3494 1873 3814 1964
rect 3494 1841 3499 1873
rect 3531 1841 3777 1873
rect 3809 1841 3814 1873
rect 3494 1749 3814 1841
rect 3494 1717 3499 1749
rect 3531 1717 3777 1749
rect 3809 1717 3814 1749
rect 3494 1712 3814 1717
rect 3842 1873 4162 1964
rect 3842 1841 3847 1873
rect 3879 1841 4125 1873
rect 4157 1841 4162 1873
rect 3842 1749 4162 1841
rect 3842 1717 3847 1749
rect 3879 1717 4125 1749
rect 4157 1717 4162 1749
rect 3842 1712 4162 1717
rect 4190 1873 4510 1964
rect 4190 1841 4195 1873
rect 4227 1841 4473 1873
rect 4505 1841 4510 1873
rect 4190 1749 4510 1841
rect 4190 1717 4195 1749
rect 4227 1717 4473 1749
rect 4505 1717 4510 1749
rect 4190 1712 4510 1717
rect 4538 1873 4858 1964
rect 4538 1841 4543 1873
rect 4575 1841 4821 1873
rect 4853 1841 4858 1873
rect 4538 1749 4858 1841
rect 4538 1717 4543 1749
rect 4575 1717 4821 1749
rect 4853 1717 4858 1749
rect 4538 1712 4858 1717
rect 4886 1873 5206 1964
rect 4886 1841 4891 1873
rect 4923 1841 5169 1873
rect 5201 1841 5206 1873
rect 4886 1749 5206 1841
rect 4886 1717 4891 1749
rect 4923 1717 5169 1749
rect 5201 1717 5206 1749
rect 4886 1712 5206 1717
rect 5234 1873 5554 1964
rect 5234 1841 5239 1873
rect 5271 1841 5517 1873
rect 5549 1841 5554 1873
rect 5234 1749 5554 1841
rect 5234 1717 5239 1749
rect 5271 1717 5517 1749
rect 5549 1717 5554 1749
rect 5234 1712 5554 1717
rect 5582 1873 5902 1964
rect 5582 1841 5587 1873
rect 5619 1841 5865 1873
rect 5897 1841 5902 1873
rect 5582 1749 5902 1841
rect 5582 1717 5587 1749
rect 5619 1717 5865 1749
rect 5897 1717 5902 1749
rect 5582 1712 5902 1717
rect 5930 1873 6250 1964
rect 5930 1841 5935 1873
rect 5967 1841 6213 1873
rect 6245 1841 6250 1873
rect 5930 1749 6250 1841
rect 5930 1717 5935 1749
rect 5967 1717 6213 1749
rect 6245 1717 6250 1749
rect 5930 1712 6250 1717
rect 6278 1873 6598 1964
rect 6278 1841 6283 1873
rect 6315 1841 6561 1873
rect 6593 1841 6598 1873
rect 6278 1749 6598 1841
rect 6278 1717 6283 1749
rect 6315 1717 6561 1749
rect 6593 1717 6598 1749
rect 6278 1712 6598 1717
rect 6626 1873 6946 1964
rect 6626 1841 6631 1873
rect 6663 1841 6909 1873
rect 6941 1841 6946 1873
rect 6626 1749 6946 1841
rect 6626 1717 6631 1749
rect 6663 1717 6909 1749
rect 6941 1746 6946 1749
rect 6974 2245 7294 2250
rect 6974 2213 6979 2245
rect 7011 2213 7257 2245
rect 7289 2213 7294 2245
rect 6974 2121 7294 2213
rect 6974 2089 6979 2121
rect 7011 2089 7257 2121
rect 7289 2089 7294 2121
rect 6974 1997 7294 2089
rect 6974 1965 6979 1997
rect 7011 1965 7257 1997
rect 7289 1978 7294 1997
rect 7289 1965 7307 1978
rect 6974 1964 7307 1965
rect 6974 1873 7294 1964
rect 6974 1841 6979 1873
rect 7011 1841 7257 1873
rect 7289 1841 7294 1873
rect 6974 1749 7294 1841
rect 6974 1746 6979 1749
rect 6941 1728 6979 1746
rect 6941 1717 6946 1728
rect 6626 1712 6946 1717
rect 6974 1717 6979 1728
rect 7011 1717 7257 1749
rect 7289 1717 7294 1749
rect 6974 1712 7294 1717
rect 25 1684 45 1712
rect 1689 1684 1709 1712
rect 1768 1684 1788 1712
rect 3439 1684 3457 1712
rect 3785 1684 3805 1712
rect 5179 1684 5195 1712
rect 5524 1684 5540 1712
rect 6985 1684 7005 1712
rect 14 1679 334 1684
rect 14 1647 19 1679
rect 51 1647 297 1679
rect 329 1647 334 1679
rect 14 1555 334 1647
rect 14 1523 19 1555
rect 51 1523 297 1555
rect 329 1523 334 1555
rect 14 1431 334 1523
rect 14 1399 19 1431
rect 51 1399 297 1431
rect 329 1399 334 1431
rect 14 1307 334 1399
rect 14 1275 19 1307
rect 51 1275 297 1307
rect 329 1275 334 1307
rect 14 1183 334 1275
rect 14 1151 19 1183
rect 51 1151 297 1183
rect 329 1151 334 1183
rect 14 1146 334 1151
rect 362 1679 682 1684
rect 362 1647 367 1679
rect 399 1647 645 1679
rect 677 1647 682 1679
rect 362 1555 682 1647
rect 362 1523 367 1555
rect 399 1523 645 1555
rect 677 1523 682 1555
rect 362 1431 682 1523
rect 362 1399 367 1431
rect 399 1399 645 1431
rect 677 1399 682 1431
rect 362 1307 682 1399
rect 362 1275 367 1307
rect 399 1275 645 1307
rect 677 1302 682 1307
rect 710 1679 1030 1684
rect 710 1647 715 1679
rect 747 1647 993 1679
rect 1025 1647 1030 1679
rect 710 1555 1030 1647
rect 710 1523 715 1555
rect 747 1523 993 1555
rect 1025 1523 1030 1555
rect 710 1431 1030 1523
rect 710 1399 715 1431
rect 747 1399 993 1431
rect 1025 1399 1030 1431
rect 710 1307 1030 1399
rect 710 1302 715 1307
rect 677 1287 715 1302
rect 677 1275 682 1287
rect 362 1183 682 1275
rect 362 1151 367 1183
rect 399 1151 645 1183
rect 677 1151 682 1183
rect 362 1146 682 1151
rect 710 1275 715 1287
rect 747 1275 993 1307
rect 1025 1299 1030 1307
rect 1058 1679 1378 1684
rect 1058 1647 1063 1679
rect 1095 1647 1341 1679
rect 1373 1647 1378 1679
rect 1058 1555 1378 1647
rect 1058 1523 1063 1555
rect 1095 1523 1341 1555
rect 1373 1523 1378 1555
rect 1058 1431 1378 1523
rect 1058 1399 1063 1431
rect 1095 1399 1341 1431
rect 1373 1399 1378 1431
rect 1058 1307 1378 1399
rect 1058 1299 1063 1307
rect 1025 1284 1063 1299
rect 1025 1275 1030 1284
rect 710 1183 1030 1275
rect 710 1151 715 1183
rect 747 1151 993 1183
rect 1025 1151 1030 1183
rect 710 1146 1030 1151
rect 1058 1275 1063 1284
rect 1095 1275 1341 1307
rect 1373 1275 1378 1307
rect 1058 1183 1378 1275
rect 1058 1151 1063 1183
rect 1095 1151 1341 1183
rect 1373 1151 1378 1183
rect 1058 1146 1378 1151
rect 1406 1679 1726 1684
rect 1406 1647 1411 1679
rect 1443 1647 1689 1679
rect 1721 1647 1726 1679
rect 1406 1555 1726 1647
rect 1406 1523 1411 1555
rect 1443 1523 1689 1555
rect 1721 1523 1726 1555
rect 1406 1431 1726 1523
rect 1406 1399 1411 1431
rect 1443 1399 1689 1431
rect 1721 1399 1726 1431
rect 1406 1307 1726 1399
rect 1406 1275 1411 1307
rect 1443 1275 1689 1307
rect 1721 1275 1726 1307
rect 1406 1183 1726 1275
rect 1406 1151 1411 1183
rect 1443 1151 1689 1183
rect 1721 1151 1726 1183
rect 1406 1146 1726 1151
rect 1754 1679 2074 1684
rect 1754 1647 1759 1679
rect 1791 1647 2037 1679
rect 2069 1647 2074 1679
rect 1754 1555 2074 1647
rect 1754 1523 1759 1555
rect 1791 1523 2037 1555
rect 2069 1523 2074 1555
rect 1754 1431 2074 1523
rect 1754 1399 1759 1431
rect 1791 1399 2037 1431
rect 2069 1399 2074 1431
rect 1754 1307 2074 1399
rect 1754 1275 1759 1307
rect 1791 1275 2037 1307
rect 2069 1275 2074 1307
rect 1754 1183 2074 1275
rect 1754 1151 1759 1183
rect 1791 1151 2037 1183
rect 2069 1151 2074 1183
rect 1754 1146 2074 1151
rect 2102 1679 2422 1684
rect 2102 1647 2107 1679
rect 2139 1647 2385 1679
rect 2417 1647 2422 1679
rect 2102 1555 2422 1647
rect 2102 1523 2107 1555
rect 2139 1523 2385 1555
rect 2417 1523 2422 1555
rect 2102 1431 2422 1523
rect 2102 1399 2107 1431
rect 2139 1399 2385 1431
rect 2417 1399 2422 1431
rect 2102 1307 2422 1399
rect 2102 1275 2107 1307
rect 2139 1275 2385 1307
rect 2417 1275 2422 1307
rect 2102 1183 2422 1275
rect 2102 1151 2107 1183
rect 2139 1151 2385 1183
rect 2417 1177 2422 1183
rect 2450 1679 2770 1684
rect 2450 1647 2455 1679
rect 2487 1647 2733 1679
rect 2765 1647 2770 1679
rect 2450 1555 2770 1647
rect 2450 1523 2455 1555
rect 2487 1523 2733 1555
rect 2765 1523 2770 1555
rect 2450 1431 2770 1523
rect 2450 1399 2455 1431
rect 2487 1399 2733 1431
rect 2765 1399 2770 1431
rect 2450 1307 2770 1399
rect 2450 1275 2455 1307
rect 2487 1275 2733 1307
rect 2765 1275 2770 1307
rect 2450 1183 2770 1275
rect 2450 1177 2455 1183
rect 2417 1162 2455 1177
rect 2417 1151 2422 1162
rect 2102 1146 2422 1151
rect 2450 1151 2455 1162
rect 2487 1151 2733 1183
rect 2765 1174 2770 1183
rect 2798 1679 3118 1684
rect 2798 1647 2803 1679
rect 2835 1647 3081 1679
rect 3113 1647 3118 1679
rect 2798 1555 3118 1647
rect 2798 1523 2803 1555
rect 2835 1523 3081 1555
rect 3113 1523 3118 1555
rect 2798 1431 3118 1523
rect 2798 1399 2803 1431
rect 2835 1399 3081 1431
rect 3113 1399 3118 1431
rect 2798 1307 3118 1399
rect 2798 1275 2803 1307
rect 2835 1275 3081 1307
rect 3113 1275 3118 1307
rect 2798 1183 3118 1275
rect 2798 1174 2803 1183
rect 2765 1159 2803 1174
rect 2765 1151 2770 1159
rect 2450 1146 2770 1151
rect 2798 1151 2803 1159
rect 2835 1151 3081 1183
rect 3113 1151 3118 1183
rect 2798 1146 3118 1151
rect 3146 1679 3466 1684
rect 3146 1647 3151 1679
rect 3183 1647 3429 1679
rect 3461 1647 3466 1679
rect 3146 1555 3466 1647
rect 3146 1523 3151 1555
rect 3183 1523 3429 1555
rect 3461 1523 3466 1555
rect 3146 1431 3466 1523
rect 3146 1399 3151 1431
rect 3183 1399 3429 1431
rect 3461 1399 3466 1431
rect 3146 1307 3466 1399
rect 3146 1275 3151 1307
rect 3183 1275 3429 1307
rect 3461 1275 3466 1307
rect 3146 1183 3466 1275
rect 3146 1151 3151 1183
rect 3183 1151 3429 1183
rect 3461 1151 3466 1183
rect 3146 1146 3466 1151
rect 3494 1679 3814 1684
rect 3494 1647 3499 1679
rect 3531 1647 3777 1679
rect 3809 1647 3814 1679
rect 3494 1555 3814 1647
rect 3494 1523 3499 1555
rect 3531 1523 3777 1555
rect 3809 1523 3814 1555
rect 3494 1431 3814 1523
rect 3494 1399 3499 1431
rect 3531 1399 3777 1431
rect 3809 1399 3814 1431
rect 3494 1307 3814 1399
rect 3494 1275 3499 1307
rect 3531 1275 3777 1307
rect 3809 1275 3814 1307
rect 3494 1183 3814 1275
rect 3494 1151 3499 1183
rect 3531 1151 3777 1183
rect 3809 1151 3814 1183
rect 3494 1146 3814 1151
rect 3842 1679 4162 1684
rect 3842 1647 3847 1679
rect 3879 1647 4125 1679
rect 4157 1647 4162 1679
rect 3842 1555 4162 1647
rect 3842 1523 3847 1555
rect 3879 1523 4125 1555
rect 4157 1523 4162 1555
rect 3842 1431 4162 1523
rect 3842 1399 3847 1431
rect 3879 1399 4125 1431
rect 4157 1399 4162 1431
rect 3842 1307 4162 1399
rect 3842 1275 3847 1307
rect 3879 1275 4125 1307
rect 4157 1275 4162 1307
rect 3842 1183 4162 1275
rect 3842 1151 3847 1183
rect 3879 1151 4125 1183
rect 4157 1182 4162 1183
rect 4190 1679 4510 1684
rect 4190 1647 4195 1679
rect 4227 1647 4473 1679
rect 4505 1647 4510 1679
rect 4190 1555 4510 1647
rect 4190 1523 4195 1555
rect 4227 1523 4473 1555
rect 4505 1523 4510 1555
rect 4190 1431 4510 1523
rect 4190 1399 4195 1431
rect 4227 1399 4473 1431
rect 4505 1399 4510 1431
rect 4190 1307 4510 1399
rect 4190 1275 4195 1307
rect 4227 1275 4473 1307
rect 4505 1275 4510 1307
rect 4190 1183 4510 1275
rect 4190 1182 4195 1183
rect 4157 1167 4195 1182
rect 4157 1151 4162 1167
rect 3842 1146 4162 1151
rect 4190 1151 4195 1167
rect 4227 1151 4473 1183
rect 4505 1182 4510 1183
rect 4538 1679 4858 1684
rect 4538 1647 4543 1679
rect 4575 1647 4821 1679
rect 4853 1647 4858 1679
rect 4538 1555 4858 1647
rect 4538 1523 4543 1555
rect 4575 1523 4821 1555
rect 4853 1523 4858 1555
rect 4538 1431 4858 1523
rect 4538 1399 4543 1431
rect 4575 1399 4821 1431
rect 4853 1399 4858 1431
rect 4538 1307 4858 1399
rect 4538 1275 4543 1307
rect 4575 1275 4821 1307
rect 4853 1275 4858 1307
rect 4538 1183 4858 1275
rect 4538 1182 4543 1183
rect 4505 1167 4543 1182
rect 4505 1151 4510 1167
rect 4190 1146 4510 1151
rect 4538 1151 4543 1167
rect 4575 1151 4821 1183
rect 4853 1151 4858 1183
rect 4538 1146 4858 1151
rect 4886 1679 5206 1684
rect 4886 1647 4891 1679
rect 4923 1647 5169 1679
rect 5201 1647 5206 1679
rect 4886 1555 5206 1647
rect 4886 1523 4891 1555
rect 4923 1523 5169 1555
rect 5201 1523 5206 1555
rect 4886 1431 5206 1523
rect 4886 1399 4891 1431
rect 4923 1399 5169 1431
rect 5201 1399 5206 1431
rect 4886 1307 5206 1399
rect 4886 1275 4891 1307
rect 4923 1275 5169 1307
rect 5201 1275 5206 1307
rect 4886 1183 5206 1275
rect 4886 1151 4891 1183
rect 4923 1151 5169 1183
rect 5201 1151 5206 1183
rect 4886 1146 5206 1151
rect 5234 1679 5554 1684
rect 5234 1647 5239 1679
rect 5271 1647 5517 1679
rect 5549 1647 5554 1679
rect 5234 1555 5554 1647
rect 5234 1523 5239 1555
rect 5271 1523 5517 1555
rect 5549 1523 5554 1555
rect 5234 1431 5554 1523
rect 5234 1399 5239 1431
rect 5271 1399 5517 1431
rect 5549 1399 5554 1431
rect 5234 1307 5554 1399
rect 5234 1275 5239 1307
rect 5271 1275 5517 1307
rect 5549 1275 5554 1307
rect 5234 1183 5554 1275
rect 5234 1151 5239 1183
rect 5271 1151 5517 1183
rect 5549 1151 5554 1183
rect 5234 1146 5554 1151
rect 5582 1679 5902 1684
rect 5582 1647 5587 1679
rect 5619 1647 5865 1679
rect 5897 1647 5902 1679
rect 5582 1555 5902 1647
rect 5582 1523 5587 1555
rect 5619 1523 5865 1555
rect 5897 1523 5902 1555
rect 5582 1431 5902 1523
rect 5582 1399 5587 1431
rect 5619 1399 5865 1431
rect 5897 1399 5902 1431
rect 5582 1307 5902 1399
rect 5582 1275 5587 1307
rect 5619 1275 5865 1307
rect 5897 1275 5902 1307
rect 5582 1183 5902 1275
rect 5582 1151 5587 1183
rect 5619 1151 5865 1183
rect 5897 1177 5902 1183
rect 5930 1679 6250 1684
rect 5930 1647 5935 1679
rect 5967 1647 6213 1679
rect 6245 1647 6250 1679
rect 5930 1555 6250 1647
rect 5930 1523 5935 1555
rect 5967 1523 6213 1555
rect 6245 1523 6250 1555
rect 5930 1431 6250 1523
rect 5930 1399 5935 1431
rect 5967 1399 6213 1431
rect 6245 1399 6250 1431
rect 5930 1307 6250 1399
rect 5930 1275 5935 1307
rect 5967 1275 6213 1307
rect 6245 1275 6250 1307
rect 5930 1183 6250 1275
rect 5930 1177 5935 1183
rect 5897 1162 5935 1177
rect 5897 1151 5902 1162
rect 5582 1146 5902 1151
rect 5930 1151 5935 1162
rect 5967 1151 6213 1183
rect 6245 1182 6250 1183
rect 6278 1679 6598 1684
rect 6278 1647 6283 1679
rect 6315 1647 6561 1679
rect 6593 1647 6598 1679
rect 6278 1555 6598 1647
rect 6278 1523 6283 1555
rect 6315 1523 6561 1555
rect 6593 1523 6598 1555
rect 6278 1431 6598 1523
rect 6278 1399 6283 1431
rect 6315 1399 6561 1431
rect 6593 1399 6598 1431
rect 6278 1307 6598 1399
rect 6278 1275 6283 1307
rect 6315 1275 6561 1307
rect 6593 1275 6598 1307
rect 6278 1183 6598 1275
rect 6278 1182 6283 1183
rect 6245 1167 6283 1182
rect 6245 1151 6250 1167
rect 5930 1146 6250 1151
rect 6278 1151 6283 1167
rect 6315 1151 6561 1183
rect 6593 1151 6598 1183
rect 6278 1146 6598 1151
rect 6626 1679 6946 1684
rect 6626 1647 6631 1679
rect 6663 1647 6909 1679
rect 6941 1647 6946 1679
rect 6626 1555 6946 1647
rect 6626 1523 6631 1555
rect 6663 1523 6909 1555
rect 6941 1523 6946 1555
rect 6626 1431 6946 1523
rect 6626 1399 6631 1431
rect 6663 1399 6909 1431
rect 6941 1399 6946 1431
rect 6626 1307 6946 1399
rect 6626 1275 6631 1307
rect 6663 1275 6909 1307
rect 6941 1275 6946 1307
rect 6626 1183 6946 1275
rect 6626 1151 6631 1183
rect 6663 1151 6909 1183
rect 6941 1151 6946 1183
rect 6626 1146 6946 1151
rect 6974 1679 7294 1684
rect 6974 1647 6979 1679
rect 7011 1647 7257 1679
rect 7289 1647 7294 1679
rect 6974 1555 7294 1647
rect 6974 1523 6979 1555
rect 7011 1523 7257 1555
rect 7289 1523 7294 1555
rect 6974 1431 7294 1523
rect 6974 1399 6979 1431
rect 7011 1399 7257 1431
rect 7289 1399 7294 1431
rect 6974 1307 7294 1399
rect 6974 1275 6979 1307
rect 7011 1275 7257 1307
rect 7289 1275 7294 1307
rect 6974 1183 7294 1275
rect 6974 1151 6979 1183
rect 7011 1151 7257 1183
rect 7289 1151 7294 1183
rect 6974 1146 7294 1151
rect 25 1118 45 1146
rect 1000 1118 1015 1146
rect 1689 1118 1709 1146
rect 1768 1118 1788 1146
rect 2465 1118 2480 1146
rect 3292 1118 3322 1146
rect 3785 1118 3805 1146
rect 4484 1118 4499 1146
rect 4984 1118 4999 1146
rect 5524 1118 5540 1146
rect 6221 1118 6236 1146
rect 6715 1118 6734 1146
rect 6985 1118 7005 1146
rect 14 1113 334 1118
rect 14 1081 19 1113
rect 51 1081 297 1113
rect 329 1081 334 1113
rect 14 989 334 1081
rect 14 957 19 989
rect 51 957 297 989
rect 329 957 334 989
rect 14 865 334 957
rect 14 833 19 865
rect 51 833 297 865
rect 329 833 334 865
rect 14 741 334 833
rect 14 709 19 741
rect 51 709 297 741
rect 329 709 334 741
rect 14 617 334 709
rect 14 585 19 617
rect 51 585 297 617
rect 329 585 334 617
rect 14 580 334 585
rect 362 1113 682 1118
rect 362 1081 367 1113
rect 399 1081 645 1113
rect 677 1081 682 1113
rect 362 989 682 1081
rect 362 957 367 989
rect 399 957 645 989
rect 677 957 682 989
rect 362 865 682 957
rect 362 833 367 865
rect 399 833 645 865
rect 677 833 682 865
rect 362 741 682 833
rect 362 709 367 741
rect 399 709 645 741
rect 677 733 682 741
rect 710 1113 1030 1118
rect 710 1081 715 1113
rect 747 1081 993 1113
rect 1025 1081 1030 1113
rect 710 989 1030 1081
rect 710 957 715 989
rect 747 957 993 989
rect 1025 957 1030 989
rect 710 865 1030 957
rect 710 833 715 865
rect 747 833 993 865
rect 1025 833 1030 865
rect 710 741 1030 833
rect 710 733 715 741
rect 677 718 715 733
rect 677 709 682 718
rect 362 617 682 709
rect 362 585 367 617
rect 399 585 645 617
rect 677 585 682 617
rect 362 580 682 585
rect 710 709 715 718
rect 747 709 993 741
rect 1025 734 1030 741
rect 1058 1113 1378 1118
rect 1058 1081 1063 1113
rect 1095 1081 1341 1113
rect 1373 1081 1378 1113
rect 1058 989 1378 1081
rect 1058 957 1063 989
rect 1095 957 1341 989
rect 1373 957 1378 989
rect 1058 865 1378 957
rect 1058 833 1063 865
rect 1095 833 1341 865
rect 1373 833 1378 865
rect 1058 741 1378 833
rect 1058 734 1063 741
rect 1025 719 1063 734
rect 1025 709 1030 719
rect 710 617 1030 709
rect 710 585 715 617
rect 747 585 993 617
rect 1025 585 1030 617
rect 710 580 1030 585
rect 1058 709 1063 719
rect 1095 709 1341 741
rect 1373 709 1378 741
rect 1058 617 1378 709
rect 1058 585 1063 617
rect 1095 585 1341 617
rect 1373 585 1378 617
rect 1058 580 1378 585
rect 1406 1113 1726 1118
rect 1406 1081 1411 1113
rect 1443 1081 1689 1113
rect 1721 1081 1726 1113
rect 1406 989 1726 1081
rect 1406 957 1411 989
rect 1443 957 1689 989
rect 1721 957 1726 989
rect 1406 865 1726 957
rect 1406 833 1411 865
rect 1443 833 1689 865
rect 1721 833 1726 865
rect 1406 741 1726 833
rect 1406 709 1411 741
rect 1443 709 1689 741
rect 1721 709 1726 741
rect 1406 617 1726 709
rect 1406 585 1411 617
rect 1443 585 1689 617
rect 1721 585 1726 617
rect 1406 580 1726 585
rect 1754 1113 2074 1118
rect 1754 1081 1759 1113
rect 1791 1081 2037 1113
rect 2069 1081 2074 1113
rect 1754 989 2074 1081
rect 1754 957 1759 989
rect 1791 957 2037 989
rect 2069 957 2074 989
rect 1754 865 2074 957
rect 1754 833 1759 865
rect 1791 833 2037 865
rect 2069 833 2074 865
rect 1754 741 2074 833
rect 1754 709 1759 741
rect 1791 709 2037 741
rect 2069 709 2074 741
rect 1754 617 2074 709
rect 1754 585 1759 617
rect 1791 585 2037 617
rect 2069 585 2074 617
rect 1754 580 2074 585
rect 2102 1113 2422 1118
rect 2102 1081 2107 1113
rect 2139 1081 2385 1113
rect 2417 1081 2422 1113
rect 2102 989 2422 1081
rect 2102 957 2107 989
rect 2139 957 2385 989
rect 2417 957 2422 989
rect 2102 865 2422 957
rect 2102 833 2107 865
rect 2139 833 2385 865
rect 2417 833 2422 865
rect 2102 741 2422 833
rect 2102 709 2107 741
rect 2139 709 2385 741
rect 2417 709 2422 741
rect 2102 617 2422 709
rect 2102 585 2107 617
rect 2139 585 2385 617
rect 2417 610 2422 617
rect 2450 1113 2770 1118
rect 2450 1081 2455 1113
rect 2487 1081 2733 1113
rect 2765 1081 2770 1113
rect 2450 989 2770 1081
rect 2450 957 2455 989
rect 2487 957 2733 989
rect 2765 957 2770 989
rect 2450 865 2770 957
rect 2450 833 2455 865
rect 2487 833 2733 865
rect 2765 833 2770 865
rect 2450 741 2770 833
rect 2450 709 2455 741
rect 2487 709 2733 741
rect 2765 709 2770 741
rect 2450 617 2770 709
rect 2450 610 2455 617
rect 2417 595 2455 610
rect 2417 585 2422 595
rect 2102 580 2422 585
rect 2450 585 2455 595
rect 2487 585 2733 617
rect 2765 614 2770 617
rect 2798 1113 3118 1118
rect 2798 1081 2803 1113
rect 2835 1081 3081 1113
rect 3113 1081 3118 1113
rect 2798 989 3118 1081
rect 2798 957 2803 989
rect 2835 957 3081 989
rect 3113 957 3118 989
rect 2798 865 3118 957
rect 2798 833 2803 865
rect 2835 833 3081 865
rect 3113 833 3118 865
rect 2798 741 3118 833
rect 2798 709 2803 741
rect 2835 709 3081 741
rect 3113 709 3118 741
rect 2798 617 3118 709
rect 2798 614 2803 617
rect 2765 599 2803 614
rect 2765 585 2770 599
rect 2450 580 2770 585
rect 2798 585 2803 599
rect 2835 585 3081 617
rect 3113 585 3118 617
rect 2798 580 3118 585
rect 3146 1113 3466 1118
rect 3146 1081 3151 1113
rect 3183 1081 3429 1113
rect 3461 1081 3466 1113
rect 3146 989 3466 1081
rect 3146 957 3151 989
rect 3183 957 3429 989
rect 3461 957 3466 989
rect 3146 865 3466 957
rect 3146 833 3151 865
rect 3183 833 3429 865
rect 3461 833 3466 865
rect 3146 741 3466 833
rect 3146 709 3151 741
rect 3183 709 3429 741
rect 3461 709 3466 741
rect 3146 617 3466 709
rect 3146 585 3151 617
rect 3183 585 3429 617
rect 3461 585 3466 617
rect 3146 580 3466 585
rect 3494 1113 3814 1118
rect 3494 1081 3499 1113
rect 3531 1081 3777 1113
rect 3809 1081 3814 1113
rect 3494 989 3814 1081
rect 3494 957 3499 989
rect 3531 957 3777 989
rect 3809 957 3814 989
rect 3494 865 3814 957
rect 3494 833 3499 865
rect 3531 833 3777 865
rect 3809 833 3814 865
rect 3494 741 3814 833
rect 3494 709 3499 741
rect 3531 709 3777 741
rect 3809 709 3814 741
rect 3494 617 3814 709
rect 3494 585 3499 617
rect 3531 585 3777 617
rect 3809 585 3814 617
rect 3494 580 3814 585
rect 3842 1113 4162 1118
rect 3842 1081 3847 1113
rect 3879 1081 4125 1113
rect 4157 1081 4162 1113
rect 3842 989 4162 1081
rect 3842 957 3847 989
rect 3879 957 4125 989
rect 4157 957 4162 989
rect 3842 865 4162 957
rect 3842 833 3847 865
rect 3879 833 4125 865
rect 4157 833 4162 865
rect 3842 741 4162 833
rect 3842 709 3847 741
rect 3879 709 4125 741
rect 4157 709 4162 741
rect 3842 617 4162 709
rect 3842 585 3847 617
rect 3879 585 4125 617
rect 4157 614 4162 617
rect 4190 1113 4510 1118
rect 4190 1081 4195 1113
rect 4227 1081 4473 1113
rect 4505 1081 4510 1113
rect 4190 989 4510 1081
rect 4190 957 4195 989
rect 4227 957 4473 989
rect 4505 957 4510 989
rect 4190 865 4510 957
rect 4190 833 4195 865
rect 4227 833 4473 865
rect 4505 833 4510 865
rect 4190 741 4510 833
rect 4190 709 4195 741
rect 4227 709 4473 741
rect 4505 709 4510 741
rect 4190 617 4510 709
rect 4190 614 4195 617
rect 4157 599 4195 614
rect 4157 585 4162 599
rect 3842 580 4162 585
rect 4190 585 4195 599
rect 4227 585 4473 617
rect 4505 616 4510 617
rect 4538 1113 4858 1118
rect 4538 1081 4543 1113
rect 4575 1081 4821 1113
rect 4853 1081 4858 1113
rect 4538 989 4858 1081
rect 4538 957 4543 989
rect 4575 957 4821 989
rect 4853 957 4858 989
rect 4538 865 4858 957
rect 4538 833 4543 865
rect 4575 833 4821 865
rect 4853 833 4858 865
rect 4538 741 4858 833
rect 4538 709 4543 741
rect 4575 709 4821 741
rect 4853 709 4858 741
rect 4538 617 4858 709
rect 4538 616 4543 617
rect 4505 601 4543 616
rect 4505 585 4510 601
rect 4190 580 4510 585
rect 4538 585 4543 601
rect 4575 585 4821 617
rect 4853 585 4858 617
rect 4538 580 4858 585
rect 4886 1113 5206 1118
rect 4886 1081 4891 1113
rect 4923 1081 5169 1113
rect 5201 1081 5206 1113
rect 4886 989 5206 1081
rect 4886 957 4891 989
rect 4923 957 5169 989
rect 5201 957 5206 989
rect 4886 865 5206 957
rect 4886 833 4891 865
rect 4923 833 5169 865
rect 5201 833 5206 865
rect 4886 741 5206 833
rect 4886 709 4891 741
rect 4923 709 5169 741
rect 5201 709 5206 741
rect 4886 617 5206 709
rect 4886 585 4891 617
rect 4923 585 5169 617
rect 5201 585 5206 617
rect 4886 580 5206 585
rect 5234 1113 5554 1118
rect 5234 1081 5239 1113
rect 5271 1081 5517 1113
rect 5549 1081 5554 1113
rect 5234 989 5554 1081
rect 5234 957 5239 989
rect 5271 957 5517 989
rect 5549 957 5554 989
rect 5234 865 5554 957
rect 5234 833 5239 865
rect 5271 833 5517 865
rect 5549 833 5554 865
rect 5234 741 5554 833
rect 5234 709 5239 741
rect 5271 709 5517 741
rect 5549 709 5554 741
rect 5234 617 5554 709
rect 5234 585 5239 617
rect 5271 585 5517 617
rect 5549 585 5554 617
rect 5234 580 5554 585
rect 5582 1113 5902 1118
rect 5582 1081 5587 1113
rect 5619 1081 5865 1113
rect 5897 1081 5902 1113
rect 5582 989 5902 1081
rect 5582 957 5587 989
rect 5619 957 5865 989
rect 5897 957 5902 989
rect 5582 865 5902 957
rect 5582 833 5587 865
rect 5619 833 5865 865
rect 5897 833 5902 865
rect 5582 741 5902 833
rect 5582 709 5587 741
rect 5619 709 5865 741
rect 5897 709 5902 741
rect 5582 617 5902 709
rect 5930 1113 6250 1118
rect 5930 1081 5935 1113
rect 5967 1081 6213 1113
rect 6245 1081 6250 1113
rect 5930 989 6250 1081
rect 5930 957 5935 989
rect 5967 957 6213 989
rect 6245 957 6250 989
rect 5930 865 6250 957
rect 5930 833 5935 865
rect 5967 833 6213 865
rect 6245 833 6250 865
rect 5930 741 6250 833
rect 5930 709 5935 741
rect 5967 709 6213 741
rect 6245 709 6250 741
rect 5930 617 6250 709
rect 5582 585 5587 617
rect 5619 585 5865 617
rect 5897 602 5935 617
rect 5897 585 5902 602
rect 5582 580 5902 585
rect 5930 585 5935 602
rect 5967 585 6213 617
rect 6245 614 6250 617
rect 6278 1113 6598 1118
rect 6278 1081 6283 1113
rect 6315 1081 6561 1113
rect 6593 1081 6598 1113
rect 6278 989 6598 1081
rect 6278 957 6283 989
rect 6315 957 6561 989
rect 6593 957 6598 989
rect 6278 865 6598 957
rect 6278 833 6283 865
rect 6315 833 6561 865
rect 6593 833 6598 865
rect 6278 741 6598 833
rect 6278 709 6283 741
rect 6315 709 6561 741
rect 6593 709 6598 741
rect 6278 617 6598 709
rect 6278 614 6283 617
rect 6245 599 6283 614
rect 6245 585 6250 599
rect 5930 580 6250 585
rect 6278 585 6283 599
rect 6315 585 6561 617
rect 6593 585 6598 617
rect 6278 580 6598 585
rect 6626 1113 6946 1118
rect 6626 1081 6631 1113
rect 6663 1081 6909 1113
rect 6941 1081 6946 1113
rect 6626 989 6946 1081
rect 6626 957 6631 989
rect 6663 957 6909 989
rect 6941 957 6946 989
rect 6626 865 6946 957
rect 6626 833 6631 865
rect 6663 833 6909 865
rect 6941 833 6946 865
rect 6626 741 6946 833
rect 6626 709 6631 741
rect 6663 709 6909 741
rect 6941 709 6946 741
rect 6626 617 6946 709
rect 6626 585 6631 617
rect 6663 585 6909 617
rect 6941 585 6946 617
rect 6626 580 6946 585
rect 6974 1113 7294 1118
rect 6974 1081 6979 1113
rect 7011 1081 7257 1113
rect 7289 1081 7294 1113
rect 6974 989 7294 1081
rect 6974 957 6979 989
rect 7011 957 7257 989
rect 7289 957 7294 989
rect 6974 865 7294 957
rect 6974 833 6979 865
rect 7011 833 7257 865
rect 7289 833 7294 865
rect 6974 741 7294 833
rect 6974 709 6979 741
rect 7011 709 7257 741
rect 7289 709 7294 741
rect 6974 617 7294 709
rect 6974 585 6979 617
rect 7011 585 7257 617
rect 7289 585 7294 617
rect 6974 580 7294 585
rect 25 552 45 580
rect 1689 552 1709 580
rect 1768 552 1788 580
rect 2662 552 2676 580
rect 3292 552 3322 580
rect 3785 552 3805 580
rect 4418 552 4434 580
rect 4985 552 5000 580
rect 5524 552 5540 580
rect 6138 552 6152 580
rect 6713 552 6732 580
rect 6985 552 7005 580
rect 14 547 334 552
rect 14 515 19 547
rect 51 515 297 547
rect 329 515 334 547
rect 14 423 334 515
rect 14 391 19 423
rect 51 391 297 423
rect 329 391 334 423
rect 14 299 334 391
rect 14 267 19 299
rect 51 267 297 299
rect 329 267 334 299
rect 14 175 334 267
rect 14 143 19 175
rect 51 143 297 175
rect 329 163 334 175
rect 362 547 682 552
rect 362 515 367 547
rect 399 515 645 547
rect 677 515 682 547
rect 362 423 682 515
rect 362 391 367 423
rect 399 391 645 423
rect 677 391 682 423
rect 362 299 682 391
rect 362 267 367 299
rect 399 267 645 299
rect 677 267 682 299
rect 362 175 682 267
rect 362 163 367 175
rect 329 149 367 163
rect 329 143 334 149
rect 14 51 334 143
rect 14 19 19 51
rect 51 19 297 51
rect 329 19 334 51
rect 14 14 334 19
rect 362 143 367 149
rect 399 143 645 175
rect 677 163 682 175
rect 710 547 1030 552
rect 710 515 715 547
rect 747 515 993 547
rect 1025 515 1030 547
rect 710 423 1030 515
rect 710 391 715 423
rect 747 391 993 423
rect 1025 391 1030 423
rect 710 299 1030 391
rect 710 267 715 299
rect 747 267 993 299
rect 1025 267 1030 299
rect 710 175 1030 267
rect 710 163 715 175
rect 677 149 715 163
rect 677 143 682 149
rect 362 51 682 143
rect 362 19 367 51
rect 399 19 645 51
rect 677 19 682 51
rect 362 14 682 19
rect 710 143 715 149
rect 747 143 993 175
rect 1025 163 1030 175
rect 1058 547 1378 552
rect 1058 515 1063 547
rect 1095 515 1341 547
rect 1373 515 1378 547
rect 1058 423 1378 515
rect 1058 391 1063 423
rect 1095 391 1341 423
rect 1373 391 1378 423
rect 1058 299 1378 391
rect 1058 267 1063 299
rect 1095 267 1341 299
rect 1373 267 1378 299
rect 1058 175 1378 267
rect 1058 163 1063 175
rect 1025 149 1063 163
rect 1025 143 1030 149
rect 710 51 1030 143
rect 710 19 715 51
rect 747 19 993 51
rect 1025 19 1030 51
rect 710 14 1030 19
rect 1058 143 1063 149
rect 1095 143 1341 175
rect 1373 163 1378 175
rect 1406 547 1726 552
rect 1406 515 1411 547
rect 1443 515 1689 547
rect 1721 515 1726 547
rect 1406 423 1726 515
rect 1406 391 1411 423
rect 1443 391 1689 423
rect 1721 391 1726 423
rect 1406 299 1726 391
rect 1406 267 1411 299
rect 1443 267 1689 299
rect 1721 267 1726 299
rect 1406 175 1726 267
rect 1406 163 1411 175
rect 1373 149 1411 163
rect 1373 143 1378 149
rect 1058 51 1378 143
rect 1058 19 1063 51
rect 1095 19 1341 51
rect 1373 19 1378 51
rect 1058 14 1378 19
rect 1406 143 1411 149
rect 1443 143 1689 175
rect 1721 163 1726 175
rect 1754 547 2074 552
rect 1754 515 1759 547
rect 1791 515 2037 547
rect 2069 515 2074 547
rect 1754 423 2074 515
rect 1754 391 1759 423
rect 1791 391 2037 423
rect 2069 391 2074 423
rect 1754 299 2074 391
rect 1754 267 1759 299
rect 1791 267 2037 299
rect 2069 267 2074 299
rect 1754 175 2074 267
rect 1754 163 1759 175
rect 1721 149 1759 163
rect 1721 143 1726 149
rect 1406 51 1726 143
rect 1406 19 1411 51
rect 1443 19 1689 51
rect 1721 19 1726 51
rect 1406 14 1726 19
rect 1754 143 1759 149
rect 1791 143 2037 175
rect 2069 163 2074 175
rect 2102 547 2422 552
rect 2102 515 2107 547
rect 2139 515 2385 547
rect 2417 515 2422 547
rect 2102 423 2422 515
rect 2102 391 2107 423
rect 2139 391 2385 423
rect 2417 391 2422 423
rect 2102 299 2422 391
rect 2102 267 2107 299
rect 2139 267 2385 299
rect 2417 267 2422 299
rect 2102 175 2422 267
rect 2102 163 2107 175
rect 2069 149 2107 163
rect 2069 143 2074 149
rect 1754 51 2074 143
rect 1754 19 1759 51
rect 1791 19 2037 51
rect 2069 19 2074 51
rect 1754 14 2074 19
rect 2102 143 2107 149
rect 2139 143 2385 175
rect 2417 143 2422 175
rect 2102 51 2422 143
rect 2102 19 2107 51
rect 2139 19 2385 51
rect 2417 19 2422 51
rect 2102 14 2422 19
rect 2450 547 2770 552
rect 2450 515 2455 547
rect 2487 515 2733 547
rect 2765 515 2770 547
rect 2450 423 2770 515
rect 2450 391 2455 423
rect 2487 391 2733 423
rect 2765 391 2770 423
rect 2450 299 2770 391
rect 2450 267 2455 299
rect 2487 267 2733 299
rect 2765 267 2770 299
rect 2450 175 2770 267
rect 2450 143 2455 175
rect 2487 143 2733 175
rect 2765 143 2770 175
rect 2450 51 2770 143
rect 2450 19 2455 51
rect 2487 19 2733 51
rect 2765 19 2770 51
rect 2450 14 2770 19
rect 2798 547 3118 552
rect 2798 515 2803 547
rect 2835 515 3081 547
rect 3113 515 3118 547
rect 2798 423 3118 515
rect 2798 391 2803 423
rect 2835 391 3081 423
rect 3113 391 3118 423
rect 2798 299 3118 391
rect 2798 267 2803 299
rect 2835 267 3081 299
rect 3113 267 3118 299
rect 2798 175 3118 267
rect 2798 143 2803 175
rect 2835 143 3081 175
rect 3113 163 3118 175
rect 3146 547 3466 552
rect 3146 515 3151 547
rect 3183 515 3429 547
rect 3461 515 3466 547
rect 3146 423 3466 515
rect 3146 391 3151 423
rect 3183 391 3429 423
rect 3461 391 3466 423
rect 3146 299 3466 391
rect 3146 267 3151 299
rect 3183 267 3429 299
rect 3461 267 3466 299
rect 3146 175 3466 267
rect 3146 163 3151 175
rect 3113 149 3151 163
rect 3113 143 3118 149
rect 2798 51 3118 143
rect 2798 19 2803 51
rect 2835 19 3081 51
rect 3113 19 3118 51
rect 2798 14 3118 19
rect 3146 143 3151 149
rect 3183 143 3429 175
rect 3461 163 3466 175
rect 3494 547 3814 552
rect 3494 515 3499 547
rect 3531 515 3777 547
rect 3809 515 3814 547
rect 3494 423 3814 515
rect 3494 391 3499 423
rect 3531 391 3777 423
rect 3809 391 3814 423
rect 3494 299 3814 391
rect 3494 267 3499 299
rect 3531 267 3777 299
rect 3809 267 3814 299
rect 3494 175 3814 267
rect 3494 163 3499 175
rect 3461 149 3499 163
rect 3461 143 3466 149
rect 3146 51 3466 143
rect 3146 19 3151 51
rect 3183 19 3429 51
rect 3461 19 3466 51
rect 3146 14 3466 19
rect 3494 143 3499 149
rect 3531 143 3777 175
rect 3809 163 3814 175
rect 3842 547 4162 552
rect 3842 515 3847 547
rect 3879 515 4125 547
rect 4157 515 4162 547
rect 3842 423 4162 515
rect 3842 391 3847 423
rect 3879 391 4125 423
rect 4157 391 4162 423
rect 3842 299 4162 391
rect 3842 267 3847 299
rect 3879 267 4125 299
rect 4157 267 4162 299
rect 3842 175 4162 267
rect 3842 163 3847 175
rect 3809 149 3847 163
rect 3809 143 3814 149
rect 3494 51 3814 143
rect 3494 19 3499 51
rect 3531 19 3777 51
rect 3809 19 3814 51
rect 3494 14 3814 19
rect 3842 143 3847 149
rect 3879 143 4125 175
rect 4157 143 4162 175
rect 3842 51 4162 143
rect 3842 19 3847 51
rect 3879 19 4125 51
rect 4157 19 4162 51
rect 3842 14 4162 19
rect 4190 547 4510 552
rect 4190 515 4195 547
rect 4227 515 4473 547
rect 4505 515 4510 547
rect 4190 423 4510 515
rect 4190 391 4195 423
rect 4227 391 4473 423
rect 4505 391 4510 423
rect 4190 299 4510 391
rect 4190 267 4195 299
rect 4227 267 4473 299
rect 4505 267 4510 299
rect 4190 175 4510 267
rect 4190 143 4195 175
rect 4227 143 4473 175
rect 4505 143 4510 175
rect 4190 51 4510 143
rect 4190 19 4195 51
rect 4227 19 4473 51
rect 4505 19 4510 51
rect 4190 14 4510 19
rect 4538 547 4858 552
rect 4538 515 4543 547
rect 4575 515 4821 547
rect 4853 515 4858 547
rect 4538 423 4858 515
rect 4538 391 4543 423
rect 4575 391 4821 423
rect 4853 391 4858 423
rect 4538 299 4858 391
rect 4538 267 4543 299
rect 4575 267 4821 299
rect 4853 267 4858 299
rect 4538 175 4858 267
rect 4538 143 4543 175
rect 4575 143 4821 175
rect 4853 163 4858 175
rect 4886 547 5206 552
rect 4886 515 4891 547
rect 4923 515 5169 547
rect 5201 515 5206 547
rect 4886 423 5206 515
rect 4886 391 4891 423
rect 4923 391 5169 423
rect 5201 391 5206 423
rect 4886 299 5206 391
rect 4886 267 4891 299
rect 4923 267 5169 299
rect 5201 267 5206 299
rect 4886 175 5206 267
rect 4886 163 4891 175
rect 4853 149 4891 163
rect 4853 143 4858 149
rect 4538 51 4858 143
rect 4538 19 4543 51
rect 4575 19 4821 51
rect 4853 19 4858 51
rect 4538 14 4858 19
rect 4886 143 4891 149
rect 4923 143 5169 175
rect 5201 163 5206 175
rect 5234 547 5554 552
rect 5234 515 5239 547
rect 5271 515 5517 547
rect 5549 515 5554 547
rect 5234 423 5554 515
rect 5234 391 5239 423
rect 5271 391 5517 423
rect 5549 391 5554 423
rect 5234 299 5554 391
rect 5234 267 5239 299
rect 5271 267 5517 299
rect 5549 267 5554 299
rect 5234 175 5554 267
rect 5234 163 5239 175
rect 5201 149 5239 163
rect 5201 143 5206 149
rect 4886 51 5206 143
rect 4886 19 4891 51
rect 4923 19 5169 51
rect 5201 19 5206 51
rect 4886 14 5206 19
rect 5234 143 5239 149
rect 5271 143 5517 175
rect 5549 163 5554 175
rect 5582 547 5902 552
rect 5582 515 5587 547
rect 5619 515 5865 547
rect 5897 515 5902 547
rect 5582 423 5902 515
rect 5582 391 5587 423
rect 5619 391 5865 423
rect 5897 391 5902 423
rect 5582 299 5902 391
rect 5582 267 5587 299
rect 5619 267 5865 299
rect 5897 267 5902 299
rect 5582 175 5902 267
rect 5582 163 5587 175
rect 5549 149 5587 163
rect 5549 143 5554 149
rect 5234 51 5554 143
rect 5234 19 5239 51
rect 5271 19 5517 51
rect 5549 19 5554 51
rect 5234 14 5554 19
rect 5582 143 5587 149
rect 5619 143 5865 175
rect 5897 143 5902 175
rect 5582 51 5902 143
rect 5582 19 5587 51
rect 5619 19 5865 51
rect 5897 19 5902 51
rect 5582 14 5902 19
rect 5930 547 6250 552
rect 5930 515 5935 547
rect 5967 515 6213 547
rect 6245 515 6250 547
rect 5930 423 6250 515
rect 5930 391 5935 423
rect 5967 391 6213 423
rect 6245 391 6250 423
rect 5930 299 6250 391
rect 5930 267 5935 299
rect 5967 267 6213 299
rect 6245 267 6250 299
rect 5930 175 6250 267
rect 5930 143 5935 175
rect 5967 143 6213 175
rect 6245 143 6250 175
rect 5930 51 6250 143
rect 5930 19 5935 51
rect 5967 19 6213 51
rect 6245 19 6250 51
rect 5930 14 6250 19
rect 6278 547 6598 552
rect 6278 515 6283 547
rect 6315 515 6561 547
rect 6593 515 6598 547
rect 6278 423 6598 515
rect 6278 391 6283 423
rect 6315 391 6561 423
rect 6593 391 6598 423
rect 6278 299 6598 391
rect 6278 267 6283 299
rect 6315 267 6561 299
rect 6593 267 6598 299
rect 6278 175 6598 267
rect 6278 143 6283 175
rect 6315 143 6561 175
rect 6593 163 6598 175
rect 6626 547 6946 552
rect 6626 515 6631 547
rect 6663 515 6909 547
rect 6941 515 6946 547
rect 6626 423 6946 515
rect 6626 391 6631 423
rect 6663 391 6909 423
rect 6941 391 6946 423
rect 6626 299 6946 391
rect 6626 267 6631 299
rect 6663 267 6909 299
rect 6941 267 6946 299
rect 6626 175 6946 267
rect 6626 163 6631 175
rect 6593 149 6631 163
rect 6593 143 6598 149
rect 6278 51 6598 143
rect 6278 19 6283 51
rect 6315 19 6561 51
rect 6593 19 6598 51
rect 6278 14 6598 19
rect 6626 143 6631 149
rect 6663 143 6909 175
rect 6941 167 6946 175
rect 6974 547 7294 552
rect 6974 515 6979 547
rect 7011 515 7257 547
rect 7289 515 7294 547
rect 6974 423 7294 515
rect 6974 391 6979 423
rect 7011 391 7257 423
rect 7289 391 7294 423
rect 6974 299 7294 391
rect 6974 267 6979 299
rect 7011 267 7257 299
rect 7289 267 7294 299
rect 6974 175 7294 267
rect 6974 167 6979 175
rect 6941 149 6979 167
rect 6941 143 6946 149
rect 6626 51 6946 143
rect 6626 19 6631 51
rect 6663 19 6909 51
rect 6941 19 6946 51
rect 6626 14 6946 19
rect 6974 143 6979 149
rect 7011 143 7257 175
rect 7289 163 7294 175
rect 7289 149 7307 163
rect 7289 143 7294 149
rect 6974 51 7294 143
rect 6974 19 6979 51
rect 7011 19 7257 51
rect 7289 19 7294 51
rect 6974 14 7294 19
<< via2 >>
rect 19 2213 51 2245
rect 297 2213 329 2245
rect 19 2089 51 2121
rect 297 2089 329 2121
rect 19 1965 51 1997
rect 297 1965 329 1997
rect 367 2213 399 2245
rect 645 2213 677 2245
rect 367 2089 399 2121
rect 645 2089 677 2121
rect 367 1965 399 1997
rect 645 1965 677 1997
rect 715 2213 747 2245
rect 993 2213 1025 2245
rect 715 2089 747 2121
rect 993 2089 1025 2121
rect 715 1965 747 1997
rect 993 1965 1025 1997
rect 1063 2213 1095 2245
rect 1341 2213 1373 2245
rect 1063 2089 1095 2121
rect 1341 2089 1373 2121
rect 1063 1965 1095 1997
rect 1341 1965 1373 1997
rect 1411 2213 1443 2245
rect 1689 2213 1721 2245
rect 1411 2089 1443 2121
rect 1689 2089 1721 2121
rect 1411 1965 1443 1997
rect 1689 1965 1721 1997
rect 1759 2213 1791 2245
rect 2037 2213 2069 2245
rect 1759 2089 1791 2121
rect 2037 2089 2069 2121
rect 1759 1965 1791 1997
rect 2037 1965 2069 1997
rect 2107 2213 2139 2245
rect 2385 2213 2417 2245
rect 2107 2089 2139 2121
rect 2385 2089 2417 2121
rect 2107 1965 2139 1997
rect 2385 1965 2417 1997
rect 2455 2213 2487 2245
rect 2733 2213 2765 2245
rect 2455 2089 2487 2121
rect 2733 2089 2765 2121
rect 2455 1965 2487 1997
rect 2733 1965 2765 1997
rect 2803 2213 2835 2245
rect 3081 2213 3113 2245
rect 2803 2089 2835 2121
rect 3081 2089 3113 2121
rect 2803 1965 2835 1997
rect 3081 1965 3113 1997
rect 3151 2213 3183 2245
rect 3429 2213 3461 2245
rect 3151 2089 3183 2121
rect 3429 2089 3461 2121
rect 3151 1965 3183 1997
rect 3429 1965 3461 1997
rect 3499 2213 3531 2245
rect 3777 2213 3809 2245
rect 3499 2089 3531 2121
rect 3777 2089 3809 2121
rect 3499 1965 3531 1997
rect 3777 1965 3809 1997
rect 3847 2213 3879 2245
rect 4125 2213 4157 2245
rect 3847 2089 3879 2121
rect 4125 2089 4157 2121
rect 3847 1965 3879 1997
rect 4125 1965 4157 1997
rect 4195 2213 4227 2245
rect 4473 2213 4505 2245
rect 4195 2089 4227 2121
rect 4473 2089 4505 2121
rect 4195 1965 4227 1997
rect 4473 1965 4505 1997
rect 4543 2213 4575 2245
rect 4821 2213 4853 2245
rect 4543 2089 4575 2121
rect 4821 2089 4853 2121
rect 4543 1965 4575 1997
rect 4821 1965 4853 1997
rect 4891 2213 4923 2245
rect 5169 2213 5201 2245
rect 4891 2089 4923 2121
rect 5169 2089 5201 2121
rect 4891 1965 4923 1997
rect 5169 1965 5201 1997
rect 5239 2213 5271 2245
rect 5517 2213 5549 2245
rect 5239 2089 5271 2121
rect 5517 2089 5549 2121
rect 5239 1965 5271 1997
rect 5517 1965 5549 1997
rect 5587 2213 5619 2245
rect 5865 2213 5897 2245
rect 5587 2089 5619 2121
rect 5865 2089 5897 2121
rect 5587 1965 5619 1997
rect 5865 1965 5897 1997
rect 5935 2213 5967 2245
rect 6213 2213 6245 2245
rect 5935 2089 5967 2121
rect 6213 2089 6245 2121
rect 5935 1965 5967 1997
rect 6213 1965 6245 1997
rect 6283 2213 6315 2245
rect 6561 2213 6593 2245
rect 6283 2089 6315 2121
rect 6561 2089 6593 2121
rect 6283 1965 6315 1997
rect 6561 1965 6593 1997
rect 6631 2213 6663 2245
rect 6909 2213 6941 2245
rect 6631 2089 6663 2121
rect 6909 2089 6941 2121
rect 6631 1965 6663 1997
rect 6909 1965 6941 1997
rect 19 1841 51 1873
rect 297 1841 329 1873
rect 19 1717 51 1749
rect 297 1717 329 1749
rect 367 1841 399 1873
rect 645 1841 677 1873
rect 367 1717 399 1749
rect 645 1717 677 1749
rect 715 1841 747 1873
rect 993 1841 1025 1873
rect 715 1717 747 1749
rect 993 1717 1025 1749
rect 1063 1841 1095 1873
rect 1341 1841 1373 1873
rect 1063 1717 1095 1749
rect 1341 1717 1373 1749
rect 1411 1841 1443 1873
rect 1689 1841 1721 1873
rect 1411 1717 1443 1749
rect 1689 1717 1721 1749
rect 1759 1841 1791 1873
rect 2037 1841 2069 1873
rect 1759 1717 1791 1749
rect 2037 1717 2069 1749
rect 2107 1841 2139 1873
rect 2385 1841 2417 1873
rect 2107 1717 2139 1749
rect 2385 1717 2417 1749
rect 2455 1841 2487 1873
rect 2733 1841 2765 1873
rect 2455 1717 2487 1749
rect 2733 1717 2765 1749
rect 2803 1841 2835 1873
rect 3081 1841 3113 1873
rect 2803 1717 2835 1749
rect 3081 1717 3113 1749
rect 3151 1841 3183 1873
rect 3429 1841 3461 1873
rect 3151 1717 3183 1749
rect 3429 1717 3461 1749
rect 3499 1841 3531 1873
rect 3777 1841 3809 1873
rect 3499 1717 3531 1749
rect 3777 1717 3809 1749
rect 3847 1841 3879 1873
rect 4125 1841 4157 1873
rect 3847 1717 3879 1749
rect 4125 1717 4157 1749
rect 4195 1841 4227 1873
rect 4473 1841 4505 1873
rect 4195 1717 4227 1749
rect 4473 1717 4505 1749
rect 4543 1841 4575 1873
rect 4821 1841 4853 1873
rect 4543 1717 4575 1749
rect 4821 1717 4853 1749
rect 4891 1841 4923 1873
rect 5169 1841 5201 1873
rect 4891 1717 4923 1749
rect 5169 1717 5201 1749
rect 5239 1841 5271 1873
rect 5517 1841 5549 1873
rect 5239 1717 5271 1749
rect 5517 1717 5549 1749
rect 5587 1841 5619 1873
rect 5865 1841 5897 1873
rect 5587 1717 5619 1749
rect 5865 1717 5897 1749
rect 5935 1841 5967 1873
rect 6213 1841 6245 1873
rect 5935 1717 5967 1749
rect 6213 1717 6245 1749
rect 6283 1841 6315 1873
rect 6561 1841 6593 1873
rect 6283 1717 6315 1749
rect 6561 1717 6593 1749
rect 6631 1841 6663 1873
rect 6909 1841 6941 1873
rect 6631 1717 6663 1749
rect 6909 1717 6941 1749
rect 6979 2213 7011 2245
rect 7257 2213 7289 2245
rect 6979 2089 7011 2121
rect 7257 2089 7289 2121
rect 6979 1965 7011 1997
rect 7257 1965 7289 1997
rect 6979 1841 7011 1873
rect 7257 1841 7289 1873
rect 6979 1717 7011 1749
rect 7257 1717 7289 1749
rect 19 1647 51 1679
rect 297 1647 329 1679
rect 19 1523 51 1555
rect 297 1523 329 1555
rect 19 1399 51 1431
rect 297 1399 329 1431
rect 19 1275 51 1307
rect 297 1275 329 1307
rect 19 1151 51 1183
rect 297 1151 329 1183
rect 367 1647 399 1679
rect 645 1647 677 1679
rect 367 1523 399 1555
rect 645 1523 677 1555
rect 367 1399 399 1431
rect 645 1399 677 1431
rect 367 1275 399 1307
rect 645 1275 677 1307
rect 715 1647 747 1679
rect 993 1647 1025 1679
rect 715 1523 747 1555
rect 993 1523 1025 1555
rect 715 1399 747 1431
rect 993 1399 1025 1431
rect 367 1151 399 1183
rect 645 1151 677 1183
rect 715 1275 747 1307
rect 993 1275 1025 1307
rect 1063 1647 1095 1679
rect 1341 1647 1373 1679
rect 1063 1523 1095 1555
rect 1341 1523 1373 1555
rect 1063 1399 1095 1431
rect 1341 1399 1373 1431
rect 715 1151 747 1183
rect 993 1151 1025 1183
rect 1063 1275 1095 1307
rect 1341 1275 1373 1307
rect 1063 1151 1095 1183
rect 1341 1151 1373 1183
rect 1411 1647 1443 1679
rect 1689 1647 1721 1679
rect 1411 1523 1443 1555
rect 1689 1523 1721 1555
rect 1411 1399 1443 1431
rect 1689 1399 1721 1431
rect 1411 1275 1443 1307
rect 1689 1275 1721 1307
rect 1411 1151 1443 1183
rect 1689 1151 1721 1183
rect 1759 1647 1791 1679
rect 2037 1647 2069 1679
rect 1759 1523 1791 1555
rect 2037 1523 2069 1555
rect 1759 1399 1791 1431
rect 2037 1399 2069 1431
rect 1759 1275 1791 1307
rect 2037 1275 2069 1307
rect 1759 1151 1791 1183
rect 2037 1151 2069 1183
rect 2107 1647 2139 1679
rect 2385 1647 2417 1679
rect 2107 1523 2139 1555
rect 2385 1523 2417 1555
rect 2107 1399 2139 1431
rect 2385 1399 2417 1431
rect 2107 1275 2139 1307
rect 2385 1275 2417 1307
rect 2107 1151 2139 1183
rect 2385 1151 2417 1183
rect 2455 1647 2487 1679
rect 2733 1647 2765 1679
rect 2455 1523 2487 1555
rect 2733 1523 2765 1555
rect 2455 1399 2487 1431
rect 2733 1399 2765 1431
rect 2455 1275 2487 1307
rect 2733 1275 2765 1307
rect 2455 1151 2487 1183
rect 2733 1151 2765 1183
rect 2803 1647 2835 1679
rect 3081 1647 3113 1679
rect 2803 1523 2835 1555
rect 3081 1523 3113 1555
rect 2803 1399 2835 1431
rect 3081 1399 3113 1431
rect 2803 1275 2835 1307
rect 3081 1275 3113 1307
rect 2803 1151 2835 1183
rect 3081 1151 3113 1183
rect 3151 1647 3183 1679
rect 3429 1647 3461 1679
rect 3151 1523 3183 1555
rect 3429 1523 3461 1555
rect 3151 1399 3183 1431
rect 3429 1399 3461 1431
rect 3151 1275 3183 1307
rect 3429 1275 3461 1307
rect 3151 1151 3183 1183
rect 3429 1151 3461 1183
rect 3499 1647 3531 1679
rect 3777 1647 3809 1679
rect 3499 1523 3531 1555
rect 3777 1523 3809 1555
rect 3499 1399 3531 1431
rect 3777 1399 3809 1431
rect 3499 1275 3531 1307
rect 3777 1275 3809 1307
rect 3499 1151 3531 1183
rect 3777 1151 3809 1183
rect 3847 1647 3879 1679
rect 4125 1647 4157 1679
rect 3847 1523 3879 1555
rect 4125 1523 4157 1555
rect 3847 1399 3879 1431
rect 4125 1399 4157 1431
rect 3847 1275 3879 1307
rect 4125 1275 4157 1307
rect 3847 1151 3879 1183
rect 4125 1151 4157 1183
rect 4195 1647 4227 1679
rect 4473 1647 4505 1679
rect 4195 1523 4227 1555
rect 4473 1523 4505 1555
rect 4195 1399 4227 1431
rect 4473 1399 4505 1431
rect 4195 1275 4227 1307
rect 4473 1275 4505 1307
rect 4195 1151 4227 1183
rect 4473 1151 4505 1183
rect 4543 1647 4575 1679
rect 4821 1647 4853 1679
rect 4543 1523 4575 1555
rect 4821 1523 4853 1555
rect 4543 1399 4575 1431
rect 4821 1399 4853 1431
rect 4543 1275 4575 1307
rect 4821 1275 4853 1307
rect 4543 1151 4575 1183
rect 4821 1151 4853 1183
rect 4891 1647 4923 1679
rect 5169 1647 5201 1679
rect 4891 1523 4923 1555
rect 5169 1523 5201 1555
rect 4891 1399 4923 1431
rect 5169 1399 5201 1431
rect 4891 1275 4923 1307
rect 5169 1275 5201 1307
rect 4891 1151 4923 1183
rect 5169 1151 5201 1183
rect 5239 1647 5271 1679
rect 5517 1647 5549 1679
rect 5239 1523 5271 1555
rect 5517 1523 5549 1555
rect 5239 1399 5271 1431
rect 5517 1399 5549 1431
rect 5239 1275 5271 1307
rect 5517 1275 5549 1307
rect 5239 1151 5271 1183
rect 5517 1151 5549 1183
rect 5587 1647 5619 1679
rect 5865 1647 5897 1679
rect 5587 1523 5619 1555
rect 5865 1523 5897 1555
rect 5587 1399 5619 1431
rect 5865 1399 5897 1431
rect 5587 1275 5619 1307
rect 5865 1275 5897 1307
rect 5587 1151 5619 1183
rect 5865 1151 5897 1183
rect 5935 1647 5967 1679
rect 6213 1647 6245 1679
rect 5935 1523 5967 1555
rect 6213 1523 6245 1555
rect 5935 1399 5967 1431
rect 6213 1399 6245 1431
rect 5935 1275 5967 1307
rect 6213 1275 6245 1307
rect 5935 1151 5967 1183
rect 6213 1151 6245 1183
rect 6283 1647 6315 1679
rect 6561 1647 6593 1679
rect 6283 1523 6315 1555
rect 6561 1523 6593 1555
rect 6283 1399 6315 1431
rect 6561 1399 6593 1431
rect 6283 1275 6315 1307
rect 6561 1275 6593 1307
rect 6283 1151 6315 1183
rect 6561 1151 6593 1183
rect 6631 1647 6663 1679
rect 6909 1647 6941 1679
rect 6631 1523 6663 1555
rect 6909 1523 6941 1555
rect 6631 1399 6663 1431
rect 6909 1399 6941 1431
rect 6631 1275 6663 1307
rect 6909 1275 6941 1307
rect 6631 1151 6663 1183
rect 6909 1151 6941 1183
rect 6979 1647 7011 1679
rect 7257 1647 7289 1679
rect 6979 1523 7011 1555
rect 7257 1523 7289 1555
rect 6979 1399 7011 1431
rect 7257 1399 7289 1431
rect 6979 1275 7011 1307
rect 7257 1275 7289 1307
rect 6979 1151 7011 1183
rect 7257 1151 7289 1183
rect 19 1081 51 1113
rect 297 1081 329 1113
rect 19 957 51 989
rect 297 957 329 989
rect 19 833 51 865
rect 297 833 329 865
rect 19 709 51 741
rect 297 709 329 741
rect 19 585 51 617
rect 297 585 329 617
rect 367 1081 399 1113
rect 645 1081 677 1113
rect 367 957 399 989
rect 645 957 677 989
rect 367 833 399 865
rect 645 833 677 865
rect 367 709 399 741
rect 645 709 677 741
rect 715 1081 747 1113
rect 993 1081 1025 1113
rect 715 957 747 989
rect 993 957 1025 989
rect 715 833 747 865
rect 993 833 1025 865
rect 367 585 399 617
rect 645 585 677 617
rect 715 709 747 741
rect 993 709 1025 741
rect 1063 1081 1095 1113
rect 1341 1081 1373 1113
rect 1063 957 1095 989
rect 1341 957 1373 989
rect 1063 833 1095 865
rect 1341 833 1373 865
rect 715 585 747 617
rect 993 585 1025 617
rect 1063 709 1095 741
rect 1341 709 1373 741
rect 1063 585 1095 617
rect 1341 585 1373 617
rect 1411 1081 1443 1113
rect 1689 1081 1721 1113
rect 1411 957 1443 989
rect 1689 957 1721 989
rect 1411 833 1443 865
rect 1689 833 1721 865
rect 1411 709 1443 741
rect 1689 709 1721 741
rect 1411 585 1443 617
rect 1689 585 1721 617
rect 1759 1081 1791 1113
rect 2037 1081 2069 1113
rect 1759 957 1791 989
rect 2037 957 2069 989
rect 1759 833 1791 865
rect 2037 833 2069 865
rect 1759 709 1791 741
rect 2037 709 2069 741
rect 1759 585 1791 617
rect 2037 585 2069 617
rect 2107 1081 2139 1113
rect 2385 1081 2417 1113
rect 2107 957 2139 989
rect 2385 957 2417 989
rect 2107 833 2139 865
rect 2385 833 2417 865
rect 2107 709 2139 741
rect 2385 709 2417 741
rect 2107 585 2139 617
rect 2385 585 2417 617
rect 2455 1081 2487 1113
rect 2733 1081 2765 1113
rect 2455 957 2487 989
rect 2733 957 2765 989
rect 2455 833 2487 865
rect 2733 833 2765 865
rect 2455 709 2487 741
rect 2733 709 2765 741
rect 2455 585 2487 617
rect 2733 585 2765 617
rect 2803 1081 2835 1113
rect 3081 1081 3113 1113
rect 2803 957 2835 989
rect 3081 957 3113 989
rect 2803 833 2835 865
rect 3081 833 3113 865
rect 2803 709 2835 741
rect 3081 709 3113 741
rect 2803 585 2835 617
rect 3081 585 3113 617
rect 3151 1081 3183 1113
rect 3429 1081 3461 1113
rect 3151 957 3183 989
rect 3429 957 3461 989
rect 3151 833 3183 865
rect 3429 833 3461 865
rect 3151 709 3183 741
rect 3429 709 3461 741
rect 3151 585 3183 617
rect 3429 585 3461 617
rect 3499 1081 3531 1113
rect 3777 1081 3809 1113
rect 3499 957 3531 989
rect 3777 957 3809 989
rect 3499 833 3531 865
rect 3777 833 3809 865
rect 3499 709 3531 741
rect 3777 709 3809 741
rect 3499 585 3531 617
rect 3777 585 3809 617
rect 3847 1081 3879 1113
rect 4125 1081 4157 1113
rect 3847 957 3879 989
rect 4125 957 4157 989
rect 3847 833 3879 865
rect 4125 833 4157 865
rect 3847 709 3879 741
rect 4125 709 4157 741
rect 3847 585 3879 617
rect 4125 585 4157 617
rect 4195 1081 4227 1113
rect 4473 1081 4505 1113
rect 4195 957 4227 989
rect 4473 957 4505 989
rect 4195 833 4227 865
rect 4473 833 4505 865
rect 4195 709 4227 741
rect 4473 709 4505 741
rect 4195 585 4227 617
rect 4473 585 4505 617
rect 4543 1081 4575 1113
rect 4821 1081 4853 1113
rect 4543 957 4575 989
rect 4821 957 4853 989
rect 4543 833 4575 865
rect 4821 833 4853 865
rect 4543 709 4575 741
rect 4821 709 4853 741
rect 4543 585 4575 617
rect 4821 585 4853 617
rect 4891 1081 4923 1113
rect 5169 1081 5201 1113
rect 4891 957 4923 989
rect 5169 957 5201 989
rect 4891 833 4923 865
rect 5169 833 5201 865
rect 4891 709 4923 741
rect 5169 709 5201 741
rect 4891 585 4923 617
rect 5169 585 5201 617
rect 5239 1081 5271 1113
rect 5517 1081 5549 1113
rect 5239 957 5271 989
rect 5517 957 5549 989
rect 5239 833 5271 865
rect 5517 833 5549 865
rect 5239 709 5271 741
rect 5517 709 5549 741
rect 5239 585 5271 617
rect 5517 585 5549 617
rect 5587 1081 5619 1113
rect 5865 1081 5897 1113
rect 5587 957 5619 989
rect 5865 957 5897 989
rect 5587 833 5619 865
rect 5865 833 5897 865
rect 5587 709 5619 741
rect 5865 709 5897 741
rect 5935 1081 5967 1113
rect 6213 1081 6245 1113
rect 5935 957 5967 989
rect 6213 957 6245 989
rect 5935 833 5967 865
rect 6213 833 6245 865
rect 5935 709 5967 741
rect 6213 709 6245 741
rect 5587 585 5619 617
rect 5865 585 5897 617
rect 5935 585 5967 617
rect 6213 585 6245 617
rect 6283 1081 6315 1113
rect 6561 1081 6593 1113
rect 6283 957 6315 989
rect 6561 957 6593 989
rect 6283 833 6315 865
rect 6561 833 6593 865
rect 6283 709 6315 741
rect 6561 709 6593 741
rect 6283 585 6315 617
rect 6561 585 6593 617
rect 6631 1081 6663 1113
rect 6909 1081 6941 1113
rect 6631 957 6663 989
rect 6909 957 6941 989
rect 6631 833 6663 865
rect 6909 833 6941 865
rect 6631 709 6663 741
rect 6909 709 6941 741
rect 6631 585 6663 617
rect 6909 585 6941 617
rect 6979 1081 7011 1113
rect 7257 1081 7289 1113
rect 6979 957 7011 989
rect 7257 957 7289 989
rect 6979 833 7011 865
rect 7257 833 7289 865
rect 6979 709 7011 741
rect 7257 709 7289 741
rect 6979 585 7011 617
rect 7257 585 7289 617
rect 19 515 51 547
rect 297 515 329 547
rect 19 391 51 423
rect 297 391 329 423
rect 19 267 51 299
rect 297 267 329 299
rect 19 143 51 175
rect 297 143 329 175
rect 367 515 399 547
rect 645 515 677 547
rect 367 391 399 423
rect 645 391 677 423
rect 367 267 399 299
rect 645 267 677 299
rect 19 19 51 51
rect 297 19 329 51
rect 367 143 399 175
rect 645 143 677 175
rect 715 515 747 547
rect 993 515 1025 547
rect 715 391 747 423
rect 993 391 1025 423
rect 715 267 747 299
rect 993 267 1025 299
rect 367 19 399 51
rect 645 19 677 51
rect 715 143 747 175
rect 993 143 1025 175
rect 1063 515 1095 547
rect 1341 515 1373 547
rect 1063 391 1095 423
rect 1341 391 1373 423
rect 1063 267 1095 299
rect 1341 267 1373 299
rect 715 19 747 51
rect 993 19 1025 51
rect 1063 143 1095 175
rect 1341 143 1373 175
rect 1411 515 1443 547
rect 1689 515 1721 547
rect 1411 391 1443 423
rect 1689 391 1721 423
rect 1411 267 1443 299
rect 1689 267 1721 299
rect 1063 19 1095 51
rect 1341 19 1373 51
rect 1411 143 1443 175
rect 1689 143 1721 175
rect 1759 515 1791 547
rect 2037 515 2069 547
rect 1759 391 1791 423
rect 2037 391 2069 423
rect 1759 267 1791 299
rect 2037 267 2069 299
rect 1411 19 1443 51
rect 1689 19 1721 51
rect 1759 143 1791 175
rect 2037 143 2069 175
rect 2107 515 2139 547
rect 2385 515 2417 547
rect 2107 391 2139 423
rect 2385 391 2417 423
rect 2107 267 2139 299
rect 2385 267 2417 299
rect 1759 19 1791 51
rect 2037 19 2069 51
rect 2107 143 2139 175
rect 2385 143 2417 175
rect 2107 19 2139 51
rect 2385 19 2417 51
rect 2455 515 2487 547
rect 2733 515 2765 547
rect 2455 391 2487 423
rect 2733 391 2765 423
rect 2455 267 2487 299
rect 2733 267 2765 299
rect 2455 143 2487 175
rect 2733 143 2765 175
rect 2455 19 2487 51
rect 2733 19 2765 51
rect 2803 515 2835 547
rect 3081 515 3113 547
rect 2803 391 2835 423
rect 3081 391 3113 423
rect 2803 267 2835 299
rect 3081 267 3113 299
rect 2803 143 2835 175
rect 3081 143 3113 175
rect 3151 515 3183 547
rect 3429 515 3461 547
rect 3151 391 3183 423
rect 3429 391 3461 423
rect 3151 267 3183 299
rect 3429 267 3461 299
rect 2803 19 2835 51
rect 3081 19 3113 51
rect 3151 143 3183 175
rect 3429 143 3461 175
rect 3499 515 3531 547
rect 3777 515 3809 547
rect 3499 391 3531 423
rect 3777 391 3809 423
rect 3499 267 3531 299
rect 3777 267 3809 299
rect 3151 19 3183 51
rect 3429 19 3461 51
rect 3499 143 3531 175
rect 3777 143 3809 175
rect 3847 515 3879 547
rect 4125 515 4157 547
rect 3847 391 3879 423
rect 4125 391 4157 423
rect 3847 267 3879 299
rect 4125 267 4157 299
rect 3499 19 3531 51
rect 3777 19 3809 51
rect 3847 143 3879 175
rect 4125 143 4157 175
rect 3847 19 3879 51
rect 4125 19 4157 51
rect 4195 515 4227 547
rect 4473 515 4505 547
rect 4195 391 4227 423
rect 4473 391 4505 423
rect 4195 267 4227 299
rect 4473 267 4505 299
rect 4195 143 4227 175
rect 4473 143 4505 175
rect 4195 19 4227 51
rect 4473 19 4505 51
rect 4543 515 4575 547
rect 4821 515 4853 547
rect 4543 391 4575 423
rect 4821 391 4853 423
rect 4543 267 4575 299
rect 4821 267 4853 299
rect 4543 143 4575 175
rect 4821 143 4853 175
rect 4891 515 4923 547
rect 5169 515 5201 547
rect 4891 391 4923 423
rect 5169 391 5201 423
rect 4891 267 4923 299
rect 5169 267 5201 299
rect 4543 19 4575 51
rect 4821 19 4853 51
rect 4891 143 4923 175
rect 5169 143 5201 175
rect 5239 515 5271 547
rect 5517 515 5549 547
rect 5239 391 5271 423
rect 5517 391 5549 423
rect 5239 267 5271 299
rect 5517 267 5549 299
rect 4891 19 4923 51
rect 5169 19 5201 51
rect 5239 143 5271 175
rect 5517 143 5549 175
rect 5587 515 5619 547
rect 5865 515 5897 547
rect 5587 391 5619 423
rect 5865 391 5897 423
rect 5587 267 5619 299
rect 5865 267 5897 299
rect 5239 19 5271 51
rect 5517 19 5549 51
rect 5587 143 5619 175
rect 5865 143 5897 175
rect 5587 19 5619 51
rect 5865 19 5897 51
rect 5935 515 5967 547
rect 6213 515 6245 547
rect 5935 391 5967 423
rect 6213 391 6245 423
rect 5935 267 5967 299
rect 6213 267 6245 299
rect 5935 143 5967 175
rect 6213 143 6245 175
rect 5935 19 5967 51
rect 6213 19 6245 51
rect 6283 515 6315 547
rect 6561 515 6593 547
rect 6283 391 6315 423
rect 6561 391 6593 423
rect 6283 267 6315 299
rect 6561 267 6593 299
rect 6283 143 6315 175
rect 6561 143 6593 175
rect 6631 515 6663 547
rect 6909 515 6941 547
rect 6631 391 6663 423
rect 6909 391 6941 423
rect 6631 267 6663 299
rect 6909 267 6941 299
rect 6283 19 6315 51
rect 6561 19 6593 51
rect 6631 143 6663 175
rect 6909 143 6941 175
rect 6979 515 7011 547
rect 7257 515 7289 547
rect 6979 391 7011 423
rect 7257 391 7289 423
rect 6979 267 7011 299
rect 7257 267 7289 299
rect 6631 19 6663 51
rect 6909 19 6941 51
rect 6979 143 7011 175
rect 7257 143 7289 175
rect 6979 19 7011 51
rect 7257 19 7289 51
<< metal3 >>
rect 16 2246 54 2248
rect 294 2246 332 2248
rect 16 2245 83 2246
rect 16 2213 19 2245
rect 51 2213 83 2245
rect 16 2212 83 2213
rect 265 2245 332 2246
rect 265 2213 297 2245
rect 329 2213 332 2245
rect 265 2212 332 2213
rect 16 2210 54 2212
rect 294 2210 332 2212
rect 364 2246 402 2248
rect 642 2246 680 2248
rect 364 2245 431 2246
rect 364 2213 367 2245
rect 399 2213 431 2245
rect 364 2212 431 2213
rect 613 2245 680 2246
rect 613 2213 645 2245
rect 677 2213 680 2245
rect 613 2212 680 2213
rect 364 2210 402 2212
rect 642 2210 680 2212
rect 712 2246 750 2248
rect 990 2246 1028 2248
rect 712 2245 779 2246
rect 712 2213 715 2245
rect 747 2213 779 2245
rect 712 2212 779 2213
rect 961 2245 1028 2246
rect 961 2213 993 2245
rect 1025 2213 1028 2245
rect 961 2212 1028 2213
rect 712 2210 750 2212
rect 990 2210 1028 2212
rect 1060 2246 1098 2248
rect 1338 2246 1376 2248
rect 1060 2245 1127 2246
rect 1060 2213 1063 2245
rect 1095 2213 1127 2245
rect 1060 2212 1127 2213
rect 1309 2245 1376 2246
rect 1309 2213 1341 2245
rect 1373 2213 1376 2245
rect 1309 2212 1376 2213
rect 1060 2210 1098 2212
rect 1338 2210 1376 2212
rect 1408 2246 1446 2248
rect 1686 2246 1724 2248
rect 1408 2245 1475 2246
rect 1408 2213 1411 2245
rect 1443 2213 1475 2245
rect 1408 2212 1475 2213
rect 1657 2245 1724 2246
rect 1657 2213 1689 2245
rect 1721 2213 1724 2245
rect 1657 2212 1724 2213
rect 1408 2210 1446 2212
rect 1686 2210 1724 2212
rect 1756 2246 1794 2248
rect 2034 2246 2072 2248
rect 1756 2245 1823 2246
rect 1756 2213 1759 2245
rect 1791 2213 1823 2245
rect 1756 2212 1823 2213
rect 2005 2245 2072 2246
rect 2005 2213 2037 2245
rect 2069 2213 2072 2245
rect 2005 2212 2072 2213
rect 1756 2210 1794 2212
rect 2034 2210 2072 2212
rect 2104 2246 2142 2248
rect 2382 2246 2420 2248
rect 2104 2245 2171 2246
rect 2104 2213 2107 2245
rect 2139 2213 2171 2245
rect 2104 2212 2171 2213
rect 2353 2245 2420 2246
rect 2353 2213 2385 2245
rect 2417 2213 2420 2245
rect 2353 2212 2420 2213
rect 2104 2210 2142 2212
rect 2382 2210 2420 2212
rect 2452 2246 2490 2248
rect 2730 2246 2768 2248
rect 2452 2245 2519 2246
rect 2452 2213 2455 2245
rect 2487 2213 2519 2245
rect 2452 2212 2519 2213
rect 2701 2245 2768 2246
rect 2701 2213 2733 2245
rect 2765 2213 2768 2245
rect 2701 2212 2768 2213
rect 2452 2210 2490 2212
rect 2730 2210 2768 2212
rect 2800 2246 2838 2248
rect 3078 2246 3116 2248
rect 2800 2245 2867 2246
rect 2800 2213 2803 2245
rect 2835 2213 2867 2245
rect 2800 2212 2867 2213
rect 3049 2245 3116 2246
rect 3049 2213 3081 2245
rect 3113 2213 3116 2245
rect 3049 2212 3116 2213
rect 2800 2210 2838 2212
rect 3078 2210 3116 2212
rect 3148 2246 3186 2248
rect 3426 2246 3464 2248
rect 3148 2245 3215 2246
rect 3148 2213 3151 2245
rect 3183 2213 3215 2245
rect 3148 2212 3215 2213
rect 3397 2245 3464 2246
rect 3397 2213 3429 2245
rect 3461 2213 3464 2245
rect 3397 2212 3464 2213
rect 3148 2210 3186 2212
rect 3426 2210 3464 2212
rect 3496 2246 3534 2248
rect 3774 2246 3812 2248
rect 3496 2245 3563 2246
rect 3496 2213 3499 2245
rect 3531 2213 3563 2245
rect 3496 2212 3563 2213
rect 3745 2245 3812 2246
rect 3745 2213 3777 2245
rect 3809 2213 3812 2245
rect 3745 2212 3812 2213
rect 3496 2210 3534 2212
rect 3774 2210 3812 2212
rect 3844 2246 3882 2248
rect 4122 2246 4160 2248
rect 3844 2245 3911 2246
rect 3844 2213 3847 2245
rect 3879 2213 3911 2245
rect 3844 2212 3911 2213
rect 4093 2245 4160 2246
rect 4093 2213 4125 2245
rect 4157 2213 4160 2245
rect 4093 2212 4160 2213
rect 3844 2210 3882 2212
rect 4122 2210 4160 2212
rect 4192 2246 4230 2248
rect 4470 2246 4508 2248
rect 4192 2245 4259 2246
rect 4192 2213 4195 2245
rect 4227 2213 4259 2245
rect 4192 2212 4259 2213
rect 4441 2245 4508 2246
rect 4441 2213 4473 2245
rect 4505 2213 4508 2245
rect 4441 2212 4508 2213
rect 4192 2210 4230 2212
rect 4470 2210 4508 2212
rect 4540 2246 4578 2248
rect 4818 2246 4856 2248
rect 4540 2245 4607 2246
rect 4540 2213 4543 2245
rect 4575 2213 4607 2245
rect 4540 2212 4607 2213
rect 4789 2245 4856 2246
rect 4789 2213 4821 2245
rect 4853 2213 4856 2245
rect 4789 2212 4856 2213
rect 4540 2210 4578 2212
rect 4818 2210 4856 2212
rect 4888 2246 4926 2248
rect 5166 2246 5204 2248
rect 4888 2245 4955 2246
rect 4888 2213 4891 2245
rect 4923 2213 4955 2245
rect 4888 2212 4955 2213
rect 5137 2245 5204 2246
rect 5137 2213 5169 2245
rect 5201 2213 5204 2245
rect 5137 2212 5204 2213
rect 4888 2210 4926 2212
rect 5166 2210 5204 2212
rect 5236 2246 5274 2248
rect 5514 2246 5552 2248
rect 5236 2245 5303 2246
rect 5236 2213 5239 2245
rect 5271 2213 5303 2245
rect 5236 2212 5303 2213
rect 5485 2245 5552 2246
rect 5485 2213 5517 2245
rect 5549 2213 5552 2245
rect 5485 2212 5552 2213
rect 5236 2210 5274 2212
rect 5514 2210 5552 2212
rect 5584 2246 5622 2248
rect 5862 2246 5900 2248
rect 5584 2245 5651 2246
rect 5584 2213 5587 2245
rect 5619 2213 5651 2245
rect 5584 2212 5651 2213
rect 5833 2245 5900 2246
rect 5833 2213 5865 2245
rect 5897 2213 5900 2245
rect 5833 2212 5900 2213
rect 5584 2210 5622 2212
rect 5862 2210 5900 2212
rect 5932 2246 5970 2248
rect 6210 2246 6248 2248
rect 5932 2245 5999 2246
rect 5932 2213 5935 2245
rect 5967 2213 5999 2245
rect 5932 2212 5999 2213
rect 6181 2245 6248 2246
rect 6181 2213 6213 2245
rect 6245 2213 6248 2245
rect 6181 2212 6248 2213
rect 5932 2210 5970 2212
rect 6210 2210 6248 2212
rect 6280 2246 6318 2248
rect 6558 2246 6596 2248
rect 6280 2245 6347 2246
rect 6280 2213 6283 2245
rect 6315 2213 6347 2245
rect 6280 2212 6347 2213
rect 6529 2245 6596 2246
rect 6529 2213 6561 2245
rect 6593 2213 6596 2245
rect 6529 2212 6596 2213
rect 6280 2210 6318 2212
rect 6558 2210 6596 2212
rect 6628 2246 6666 2248
rect 6906 2246 6944 2248
rect 6628 2245 6695 2246
rect 6628 2213 6631 2245
rect 6663 2213 6695 2245
rect 6628 2212 6695 2213
rect 6877 2245 6944 2246
rect 6877 2213 6909 2245
rect 6941 2213 6944 2245
rect 6877 2212 6944 2213
rect 6628 2210 6666 2212
rect 6906 2210 6944 2212
rect 6976 2246 7014 2248
rect 7254 2246 7292 2248
rect 6976 2245 7043 2246
rect 6976 2213 6979 2245
rect 7011 2213 7043 2245
rect 6976 2212 7043 2213
rect 7225 2245 7292 2246
rect 7225 2213 7257 2245
rect 7289 2213 7292 2245
rect 7225 2212 7292 2213
rect 6976 2210 7014 2212
rect 7254 2210 7292 2212
rect 16 2122 54 2124
rect 294 2122 332 2124
rect 16 2121 83 2122
rect 16 2089 19 2121
rect 51 2089 83 2121
rect 16 2088 83 2089
rect 265 2121 332 2122
rect 265 2089 297 2121
rect 329 2089 332 2121
rect 265 2088 332 2089
rect 16 2086 54 2088
rect 294 2086 332 2088
rect 364 2122 402 2124
rect 642 2122 680 2124
rect 364 2121 431 2122
rect 364 2089 367 2121
rect 399 2089 431 2121
rect 364 2088 431 2089
rect 613 2121 680 2122
rect 613 2089 645 2121
rect 677 2089 680 2121
rect 613 2088 680 2089
rect 364 2086 402 2088
rect 642 2086 680 2088
rect 712 2122 750 2124
rect 990 2122 1028 2124
rect 712 2121 779 2122
rect 712 2089 715 2121
rect 747 2089 779 2121
rect 712 2088 779 2089
rect 961 2121 1028 2122
rect 961 2089 993 2121
rect 1025 2089 1028 2121
rect 961 2088 1028 2089
rect 712 2086 750 2088
rect 990 2086 1028 2088
rect 1060 2122 1098 2124
rect 1338 2122 1376 2124
rect 1060 2121 1127 2122
rect 1060 2089 1063 2121
rect 1095 2089 1127 2121
rect 1060 2088 1127 2089
rect 1309 2121 1376 2122
rect 1309 2089 1341 2121
rect 1373 2089 1376 2121
rect 1309 2088 1376 2089
rect 1060 2086 1098 2088
rect 1338 2086 1376 2088
rect 1408 2122 1446 2124
rect 1686 2122 1724 2124
rect 1408 2121 1475 2122
rect 1408 2089 1411 2121
rect 1443 2089 1475 2121
rect 1408 2088 1475 2089
rect 1657 2121 1724 2122
rect 1657 2089 1689 2121
rect 1721 2089 1724 2121
rect 1657 2088 1724 2089
rect 1408 2086 1446 2088
rect 1686 2086 1724 2088
rect 1756 2122 1794 2124
rect 2034 2122 2072 2124
rect 1756 2121 1823 2122
rect 1756 2089 1759 2121
rect 1791 2089 1823 2121
rect 1756 2088 1823 2089
rect 2005 2121 2072 2122
rect 2005 2089 2037 2121
rect 2069 2089 2072 2121
rect 2005 2088 2072 2089
rect 1756 2086 1794 2088
rect 2034 2086 2072 2088
rect 2104 2122 2142 2124
rect 2382 2122 2420 2124
rect 2104 2121 2171 2122
rect 2104 2089 2107 2121
rect 2139 2089 2171 2121
rect 2104 2088 2171 2089
rect 2353 2121 2420 2122
rect 2353 2089 2385 2121
rect 2417 2089 2420 2121
rect 2353 2088 2420 2089
rect 2104 2086 2142 2088
rect 2382 2086 2420 2088
rect 2452 2122 2490 2124
rect 2730 2122 2768 2124
rect 2452 2121 2519 2122
rect 2452 2089 2455 2121
rect 2487 2089 2519 2121
rect 2452 2088 2519 2089
rect 2701 2121 2768 2122
rect 2701 2089 2733 2121
rect 2765 2089 2768 2121
rect 2701 2088 2768 2089
rect 2452 2086 2490 2088
rect 2730 2086 2768 2088
rect 2800 2122 2838 2124
rect 3078 2122 3116 2124
rect 2800 2121 2867 2122
rect 2800 2089 2803 2121
rect 2835 2089 2867 2121
rect 2800 2088 2867 2089
rect 3049 2121 3116 2122
rect 3049 2089 3081 2121
rect 3113 2089 3116 2121
rect 3049 2088 3116 2089
rect 2800 2086 2838 2088
rect 3078 2086 3116 2088
rect 3148 2122 3186 2124
rect 3426 2122 3464 2124
rect 3148 2121 3215 2122
rect 3148 2089 3151 2121
rect 3183 2089 3215 2121
rect 3148 2088 3215 2089
rect 3397 2121 3464 2122
rect 3397 2089 3429 2121
rect 3461 2089 3464 2121
rect 3397 2088 3464 2089
rect 3148 2086 3186 2088
rect 3426 2086 3464 2088
rect 3496 2122 3534 2124
rect 3774 2122 3812 2124
rect 3496 2121 3563 2122
rect 3496 2089 3499 2121
rect 3531 2089 3563 2121
rect 3496 2088 3563 2089
rect 3745 2121 3812 2122
rect 3745 2089 3777 2121
rect 3809 2089 3812 2121
rect 3745 2088 3812 2089
rect 3496 2086 3534 2088
rect 3774 2086 3812 2088
rect 3844 2122 3882 2124
rect 4122 2122 4160 2124
rect 3844 2121 3911 2122
rect 3844 2089 3847 2121
rect 3879 2089 3911 2121
rect 3844 2088 3911 2089
rect 4093 2121 4160 2122
rect 4093 2089 4125 2121
rect 4157 2089 4160 2121
rect 4093 2088 4160 2089
rect 3844 2086 3882 2088
rect 4122 2086 4160 2088
rect 4192 2122 4230 2124
rect 4470 2122 4508 2124
rect 4192 2121 4259 2122
rect 4192 2089 4195 2121
rect 4227 2089 4259 2121
rect 4192 2088 4259 2089
rect 4441 2121 4508 2122
rect 4441 2089 4473 2121
rect 4505 2089 4508 2121
rect 4441 2088 4508 2089
rect 4192 2086 4230 2088
rect 4470 2086 4508 2088
rect 4540 2122 4578 2124
rect 4818 2122 4856 2124
rect 4540 2121 4607 2122
rect 4540 2089 4543 2121
rect 4575 2089 4607 2121
rect 4540 2088 4607 2089
rect 4789 2121 4856 2122
rect 4789 2089 4821 2121
rect 4853 2089 4856 2121
rect 4789 2088 4856 2089
rect 4540 2086 4578 2088
rect 4818 2086 4856 2088
rect 4888 2122 4926 2124
rect 5166 2122 5204 2124
rect 4888 2121 4955 2122
rect 4888 2089 4891 2121
rect 4923 2089 4955 2121
rect 4888 2088 4955 2089
rect 5137 2121 5204 2122
rect 5137 2089 5169 2121
rect 5201 2089 5204 2121
rect 5137 2088 5204 2089
rect 4888 2086 4926 2088
rect 5166 2086 5204 2088
rect 5236 2122 5274 2124
rect 5514 2122 5552 2124
rect 5236 2121 5303 2122
rect 5236 2089 5239 2121
rect 5271 2089 5303 2121
rect 5236 2088 5303 2089
rect 5485 2121 5552 2122
rect 5485 2089 5517 2121
rect 5549 2089 5552 2121
rect 5485 2088 5552 2089
rect 5236 2086 5274 2088
rect 5514 2086 5552 2088
rect 5584 2122 5622 2124
rect 5862 2122 5900 2124
rect 5584 2121 5651 2122
rect 5584 2089 5587 2121
rect 5619 2089 5651 2121
rect 5584 2088 5651 2089
rect 5833 2121 5900 2122
rect 5833 2089 5865 2121
rect 5897 2089 5900 2121
rect 5833 2088 5900 2089
rect 5584 2086 5622 2088
rect 5862 2086 5900 2088
rect 5932 2122 5970 2124
rect 6210 2122 6248 2124
rect 5932 2121 5999 2122
rect 5932 2089 5935 2121
rect 5967 2089 5999 2121
rect 5932 2088 5999 2089
rect 6181 2121 6248 2122
rect 6181 2089 6213 2121
rect 6245 2089 6248 2121
rect 6181 2088 6248 2089
rect 5932 2086 5970 2088
rect 6210 2086 6248 2088
rect 6280 2122 6318 2124
rect 6558 2122 6596 2124
rect 6280 2121 6347 2122
rect 6280 2089 6283 2121
rect 6315 2089 6347 2121
rect 6280 2088 6347 2089
rect 6529 2121 6596 2122
rect 6529 2089 6561 2121
rect 6593 2089 6596 2121
rect 6529 2088 6596 2089
rect 6280 2086 6318 2088
rect 6558 2086 6596 2088
rect 6628 2122 6666 2124
rect 6906 2122 6944 2124
rect 6628 2121 6695 2122
rect 6628 2089 6631 2121
rect 6663 2089 6695 2121
rect 6628 2088 6695 2089
rect 6877 2121 6944 2122
rect 6877 2089 6909 2121
rect 6941 2089 6944 2121
rect 6877 2088 6944 2089
rect 6628 2086 6666 2088
rect 6906 2086 6944 2088
rect 6976 2122 7014 2124
rect 7254 2122 7292 2124
rect 6976 2121 7043 2122
rect 6976 2089 6979 2121
rect 7011 2089 7043 2121
rect 6976 2088 7043 2089
rect 7225 2121 7292 2122
rect 7225 2089 7257 2121
rect 7289 2089 7292 2121
rect 7225 2088 7292 2089
rect 6976 2086 7014 2088
rect 7254 2086 7292 2088
rect 16 1998 54 2000
rect 294 1998 332 2000
rect 16 1997 83 1998
rect 16 1965 19 1997
rect 51 1965 83 1997
rect 16 1964 83 1965
rect 265 1997 332 1998
rect 265 1965 297 1997
rect 329 1965 332 1997
rect 265 1964 332 1965
rect 16 1962 54 1964
rect 294 1962 332 1964
rect 364 1998 402 2000
rect 642 1998 680 2000
rect 364 1997 431 1998
rect 364 1965 367 1997
rect 399 1965 431 1997
rect 364 1964 431 1965
rect 613 1997 680 1998
rect 613 1965 645 1997
rect 677 1965 680 1997
rect 613 1964 680 1965
rect 364 1962 402 1964
rect 642 1962 680 1964
rect 712 1998 750 2000
rect 990 1998 1028 2000
rect 712 1997 779 1998
rect 712 1965 715 1997
rect 747 1965 779 1997
rect 712 1964 779 1965
rect 961 1997 1028 1998
rect 961 1965 993 1997
rect 1025 1965 1028 1997
rect 961 1964 1028 1965
rect 712 1962 750 1964
rect 990 1962 1028 1964
rect 1060 1998 1098 2000
rect 1338 1998 1376 2000
rect 1060 1997 1127 1998
rect 1060 1965 1063 1997
rect 1095 1965 1127 1997
rect 1060 1964 1127 1965
rect 1309 1997 1376 1998
rect 1309 1965 1341 1997
rect 1373 1965 1376 1997
rect 1309 1964 1376 1965
rect 1060 1962 1098 1964
rect 1338 1962 1376 1964
rect 1408 1998 1446 2000
rect 1686 1998 1724 2000
rect 1408 1997 1475 1998
rect 1408 1965 1411 1997
rect 1443 1965 1475 1997
rect 1408 1964 1475 1965
rect 1657 1997 1724 1998
rect 1657 1965 1689 1997
rect 1721 1965 1724 1997
rect 1657 1964 1724 1965
rect 1408 1962 1446 1964
rect 1686 1962 1724 1964
rect 1756 1998 1794 2000
rect 2034 1998 2072 2000
rect 1756 1997 1823 1998
rect 1756 1965 1759 1997
rect 1791 1965 1823 1997
rect 1756 1964 1823 1965
rect 2005 1997 2072 1998
rect 2005 1965 2037 1997
rect 2069 1965 2072 1997
rect 2005 1964 2072 1965
rect 1756 1962 1794 1964
rect 2034 1962 2072 1964
rect 2104 1998 2142 2000
rect 2382 1998 2420 2000
rect 2104 1997 2171 1998
rect 2104 1965 2107 1997
rect 2139 1965 2171 1997
rect 2104 1964 2171 1965
rect 2353 1997 2420 1998
rect 2353 1965 2385 1997
rect 2417 1965 2420 1997
rect 2353 1964 2420 1965
rect 2104 1962 2142 1964
rect 2382 1962 2420 1964
rect 2452 1998 2490 2000
rect 2730 1998 2768 2000
rect 2452 1997 2519 1998
rect 2452 1965 2455 1997
rect 2487 1965 2519 1997
rect 2452 1964 2519 1965
rect 2701 1997 2768 1998
rect 2701 1965 2733 1997
rect 2765 1965 2768 1997
rect 2701 1964 2768 1965
rect 2452 1962 2490 1964
rect 2730 1962 2768 1964
rect 2800 1998 2838 2000
rect 3078 1998 3116 2000
rect 2800 1997 2867 1998
rect 2800 1965 2803 1997
rect 2835 1965 2867 1997
rect 2800 1964 2867 1965
rect 3049 1997 3116 1998
rect 3049 1965 3081 1997
rect 3113 1965 3116 1997
rect 3049 1964 3116 1965
rect 2800 1962 2838 1964
rect 3078 1962 3116 1964
rect 3148 1998 3186 2000
rect 3426 1998 3464 2000
rect 3148 1997 3215 1998
rect 3148 1965 3151 1997
rect 3183 1965 3215 1997
rect 3148 1964 3215 1965
rect 3397 1997 3464 1998
rect 3397 1965 3429 1997
rect 3461 1965 3464 1997
rect 3397 1964 3464 1965
rect 3148 1962 3186 1964
rect 3426 1962 3464 1964
rect 3496 1998 3534 2000
rect 3774 1998 3812 2000
rect 3496 1997 3563 1998
rect 3496 1965 3499 1997
rect 3531 1965 3563 1997
rect 3496 1964 3563 1965
rect 3745 1997 3812 1998
rect 3745 1965 3777 1997
rect 3809 1965 3812 1997
rect 3745 1964 3812 1965
rect 3496 1962 3534 1964
rect 3774 1962 3812 1964
rect 3844 1998 3882 2000
rect 4122 1998 4160 2000
rect 3844 1997 3911 1998
rect 3844 1965 3847 1997
rect 3879 1965 3911 1997
rect 3844 1964 3911 1965
rect 4093 1997 4160 1998
rect 4093 1965 4125 1997
rect 4157 1965 4160 1997
rect 4093 1964 4160 1965
rect 3844 1962 3882 1964
rect 4122 1962 4160 1964
rect 4192 1998 4230 2000
rect 4470 1998 4508 2000
rect 4192 1997 4259 1998
rect 4192 1965 4195 1997
rect 4227 1965 4259 1997
rect 4192 1964 4259 1965
rect 4441 1997 4508 1998
rect 4441 1965 4473 1997
rect 4505 1965 4508 1997
rect 4441 1964 4508 1965
rect 4192 1962 4230 1964
rect 4470 1962 4508 1964
rect 4540 1998 4578 2000
rect 4818 1998 4856 2000
rect 4540 1997 4607 1998
rect 4540 1965 4543 1997
rect 4575 1965 4607 1997
rect 4540 1964 4607 1965
rect 4789 1997 4856 1998
rect 4789 1965 4821 1997
rect 4853 1965 4856 1997
rect 4789 1964 4856 1965
rect 4540 1962 4578 1964
rect 4818 1962 4856 1964
rect 4888 1998 4926 2000
rect 5166 1998 5204 2000
rect 4888 1997 4955 1998
rect 4888 1965 4891 1997
rect 4923 1965 4955 1997
rect 4888 1964 4955 1965
rect 5137 1997 5204 1998
rect 5137 1965 5169 1997
rect 5201 1965 5204 1997
rect 5137 1964 5204 1965
rect 4888 1962 4926 1964
rect 5166 1962 5204 1964
rect 5236 1998 5274 2000
rect 5514 1998 5552 2000
rect 5236 1997 5303 1998
rect 5236 1965 5239 1997
rect 5271 1965 5303 1997
rect 5236 1964 5303 1965
rect 5485 1997 5552 1998
rect 5485 1965 5517 1997
rect 5549 1965 5552 1997
rect 5485 1964 5552 1965
rect 5236 1962 5274 1964
rect 5514 1962 5552 1964
rect 5584 1998 5622 2000
rect 5862 1998 5900 2000
rect 5584 1997 5651 1998
rect 5584 1965 5587 1997
rect 5619 1965 5651 1997
rect 5584 1964 5651 1965
rect 5833 1997 5900 1998
rect 5833 1965 5865 1997
rect 5897 1965 5900 1997
rect 5833 1964 5900 1965
rect 5584 1962 5622 1964
rect 5862 1962 5900 1964
rect 5932 1998 5970 2000
rect 6210 1998 6248 2000
rect 5932 1997 5999 1998
rect 5932 1965 5935 1997
rect 5967 1965 5999 1997
rect 5932 1964 5999 1965
rect 6181 1997 6248 1998
rect 6181 1965 6213 1997
rect 6245 1965 6248 1997
rect 6181 1964 6248 1965
rect 5932 1962 5970 1964
rect 6210 1962 6248 1964
rect 6280 1998 6318 2000
rect 6558 1998 6596 2000
rect 6280 1997 6347 1998
rect 6280 1965 6283 1997
rect 6315 1965 6347 1997
rect 6280 1964 6347 1965
rect 6529 1997 6596 1998
rect 6529 1965 6561 1997
rect 6593 1965 6596 1997
rect 6529 1964 6596 1965
rect 6280 1962 6318 1964
rect 6558 1962 6596 1964
rect 6628 1998 6666 2000
rect 6906 1998 6944 2000
rect 6628 1997 6695 1998
rect 6628 1965 6631 1997
rect 6663 1965 6695 1997
rect 6628 1964 6695 1965
rect 6877 1997 6944 1998
rect 6877 1965 6909 1997
rect 6941 1965 6944 1997
rect 6877 1964 6944 1965
rect 6628 1962 6666 1964
rect 6906 1962 6944 1964
rect 6976 1998 7014 2000
rect 7254 1998 7292 2000
rect 6976 1997 7043 1998
rect 6976 1965 6979 1997
rect 7011 1965 7043 1997
rect 6976 1964 7043 1965
rect 7225 1997 7292 1998
rect 7225 1965 7257 1997
rect 7289 1965 7292 1997
rect 7225 1964 7292 1965
rect 6976 1962 7014 1964
rect 7254 1962 7292 1964
rect 16 1874 54 1876
rect 294 1874 332 1876
rect 16 1873 83 1874
rect 16 1841 19 1873
rect 51 1841 83 1873
rect 16 1840 83 1841
rect 265 1873 332 1874
rect 265 1841 297 1873
rect 329 1841 332 1873
rect 265 1840 332 1841
rect 16 1838 54 1840
rect 294 1838 332 1840
rect 364 1874 402 1876
rect 642 1874 680 1876
rect 364 1873 431 1874
rect 364 1841 367 1873
rect 399 1841 431 1873
rect 364 1840 431 1841
rect 613 1873 680 1874
rect 613 1841 645 1873
rect 677 1841 680 1873
rect 613 1840 680 1841
rect 364 1838 402 1840
rect 642 1838 680 1840
rect 712 1874 750 1876
rect 990 1874 1028 1876
rect 712 1873 779 1874
rect 712 1841 715 1873
rect 747 1841 779 1873
rect 712 1840 779 1841
rect 961 1873 1028 1874
rect 961 1841 993 1873
rect 1025 1841 1028 1873
rect 961 1840 1028 1841
rect 712 1838 750 1840
rect 990 1838 1028 1840
rect 1060 1874 1098 1876
rect 1338 1874 1376 1876
rect 1060 1873 1127 1874
rect 1060 1841 1063 1873
rect 1095 1841 1127 1873
rect 1060 1840 1127 1841
rect 1309 1873 1376 1874
rect 1309 1841 1341 1873
rect 1373 1841 1376 1873
rect 1309 1840 1376 1841
rect 1060 1838 1098 1840
rect 1338 1838 1376 1840
rect 1408 1874 1446 1876
rect 1686 1874 1724 1876
rect 1408 1873 1475 1874
rect 1408 1841 1411 1873
rect 1443 1841 1475 1873
rect 1408 1840 1475 1841
rect 1657 1873 1724 1874
rect 1657 1841 1689 1873
rect 1721 1841 1724 1873
rect 1657 1840 1724 1841
rect 1408 1838 1446 1840
rect 1686 1838 1724 1840
rect 1756 1874 1794 1876
rect 2034 1874 2072 1876
rect 1756 1873 1823 1874
rect 1756 1841 1759 1873
rect 1791 1841 1823 1873
rect 1756 1840 1823 1841
rect 2005 1873 2072 1874
rect 2005 1841 2037 1873
rect 2069 1841 2072 1873
rect 2005 1840 2072 1841
rect 1756 1838 1794 1840
rect 2034 1838 2072 1840
rect 2104 1874 2142 1876
rect 2382 1874 2420 1876
rect 2104 1873 2171 1874
rect 2104 1841 2107 1873
rect 2139 1841 2171 1873
rect 2104 1840 2171 1841
rect 2353 1873 2420 1874
rect 2353 1841 2385 1873
rect 2417 1841 2420 1873
rect 2353 1840 2420 1841
rect 2104 1838 2142 1840
rect 2382 1838 2420 1840
rect 2452 1874 2490 1876
rect 2730 1874 2768 1876
rect 2452 1873 2519 1874
rect 2452 1841 2455 1873
rect 2487 1841 2519 1873
rect 2452 1840 2519 1841
rect 2701 1873 2768 1874
rect 2701 1841 2733 1873
rect 2765 1841 2768 1873
rect 2701 1840 2768 1841
rect 2452 1838 2490 1840
rect 2730 1838 2768 1840
rect 2800 1874 2838 1876
rect 3078 1874 3116 1876
rect 2800 1873 2867 1874
rect 2800 1841 2803 1873
rect 2835 1841 2867 1873
rect 2800 1840 2867 1841
rect 3049 1873 3116 1874
rect 3049 1841 3081 1873
rect 3113 1841 3116 1873
rect 3049 1840 3116 1841
rect 2800 1838 2838 1840
rect 3078 1838 3116 1840
rect 3148 1874 3186 1876
rect 3426 1874 3464 1876
rect 3148 1873 3215 1874
rect 3148 1841 3151 1873
rect 3183 1841 3215 1873
rect 3148 1840 3215 1841
rect 3397 1873 3464 1874
rect 3397 1841 3429 1873
rect 3461 1841 3464 1873
rect 3397 1840 3464 1841
rect 3148 1838 3186 1840
rect 3426 1838 3464 1840
rect 3496 1874 3534 1876
rect 3774 1874 3812 1876
rect 3496 1873 3563 1874
rect 3496 1841 3499 1873
rect 3531 1841 3563 1873
rect 3496 1840 3563 1841
rect 3745 1873 3812 1874
rect 3745 1841 3777 1873
rect 3809 1841 3812 1873
rect 3745 1840 3812 1841
rect 3496 1838 3534 1840
rect 3774 1838 3812 1840
rect 3844 1874 3882 1876
rect 4122 1874 4160 1876
rect 3844 1873 3911 1874
rect 3844 1841 3847 1873
rect 3879 1841 3911 1873
rect 3844 1840 3911 1841
rect 4093 1873 4160 1874
rect 4093 1841 4125 1873
rect 4157 1841 4160 1873
rect 4093 1840 4160 1841
rect 3844 1838 3882 1840
rect 4122 1838 4160 1840
rect 4192 1874 4230 1876
rect 4470 1874 4508 1876
rect 4192 1873 4259 1874
rect 4192 1841 4195 1873
rect 4227 1841 4259 1873
rect 4192 1840 4259 1841
rect 4441 1873 4508 1874
rect 4441 1841 4473 1873
rect 4505 1841 4508 1873
rect 4441 1840 4508 1841
rect 4192 1838 4230 1840
rect 4470 1838 4508 1840
rect 4540 1874 4578 1876
rect 4818 1874 4856 1876
rect 4540 1873 4607 1874
rect 4540 1841 4543 1873
rect 4575 1841 4607 1873
rect 4540 1840 4607 1841
rect 4789 1873 4856 1874
rect 4789 1841 4821 1873
rect 4853 1841 4856 1873
rect 4789 1840 4856 1841
rect 4540 1838 4578 1840
rect 4818 1838 4856 1840
rect 4888 1874 4926 1876
rect 5166 1874 5204 1876
rect 4888 1873 4955 1874
rect 4888 1841 4891 1873
rect 4923 1841 4955 1873
rect 4888 1840 4955 1841
rect 5137 1873 5204 1874
rect 5137 1841 5169 1873
rect 5201 1841 5204 1873
rect 5137 1840 5204 1841
rect 4888 1838 4926 1840
rect 5166 1838 5204 1840
rect 5236 1874 5274 1876
rect 5514 1874 5552 1876
rect 5236 1873 5303 1874
rect 5236 1841 5239 1873
rect 5271 1841 5303 1873
rect 5236 1840 5303 1841
rect 5485 1873 5552 1874
rect 5485 1841 5517 1873
rect 5549 1841 5552 1873
rect 5485 1840 5552 1841
rect 5236 1838 5274 1840
rect 5514 1838 5552 1840
rect 5584 1874 5622 1876
rect 5862 1874 5900 1876
rect 5584 1873 5651 1874
rect 5584 1841 5587 1873
rect 5619 1841 5651 1873
rect 5584 1840 5651 1841
rect 5833 1873 5900 1874
rect 5833 1841 5865 1873
rect 5897 1841 5900 1873
rect 5833 1840 5900 1841
rect 5584 1838 5622 1840
rect 5862 1838 5900 1840
rect 5932 1874 5970 1876
rect 6210 1874 6248 1876
rect 5932 1873 5999 1874
rect 5932 1841 5935 1873
rect 5967 1841 5999 1873
rect 5932 1840 5999 1841
rect 6181 1873 6248 1874
rect 6181 1841 6213 1873
rect 6245 1841 6248 1873
rect 6181 1840 6248 1841
rect 5932 1838 5970 1840
rect 6210 1838 6248 1840
rect 6280 1874 6318 1876
rect 6558 1874 6596 1876
rect 6280 1873 6347 1874
rect 6280 1841 6283 1873
rect 6315 1841 6347 1873
rect 6280 1840 6347 1841
rect 6529 1873 6596 1874
rect 6529 1841 6561 1873
rect 6593 1841 6596 1873
rect 6529 1840 6596 1841
rect 6280 1838 6318 1840
rect 6558 1838 6596 1840
rect 6628 1874 6666 1876
rect 6906 1874 6944 1876
rect 6628 1873 6695 1874
rect 6628 1841 6631 1873
rect 6663 1841 6695 1873
rect 6628 1840 6695 1841
rect 6877 1873 6944 1874
rect 6877 1841 6909 1873
rect 6941 1841 6944 1873
rect 6877 1840 6944 1841
rect 6628 1838 6666 1840
rect 6906 1838 6944 1840
rect 6976 1874 7014 1876
rect 7254 1874 7292 1876
rect 6976 1873 7043 1874
rect 6976 1841 6979 1873
rect 7011 1841 7043 1873
rect 6976 1840 7043 1841
rect 7225 1873 7292 1874
rect 7225 1841 7257 1873
rect 7289 1841 7292 1873
rect 7225 1840 7292 1841
rect 6976 1838 7014 1840
rect 7254 1838 7292 1840
rect 16 1750 54 1752
rect 294 1750 332 1752
rect 16 1749 83 1750
rect 16 1717 19 1749
rect 51 1717 83 1749
rect 16 1716 83 1717
rect 265 1749 332 1750
rect 265 1717 297 1749
rect 329 1717 332 1749
rect 265 1716 332 1717
rect 16 1714 54 1716
rect 294 1714 332 1716
rect 364 1750 402 1752
rect 642 1750 680 1752
rect 364 1749 431 1750
rect 364 1717 367 1749
rect 399 1717 431 1749
rect 364 1716 431 1717
rect 613 1749 680 1750
rect 613 1717 645 1749
rect 677 1717 680 1749
rect 613 1716 680 1717
rect 364 1714 402 1716
rect 642 1714 680 1716
rect 712 1750 750 1752
rect 990 1750 1028 1752
rect 712 1749 779 1750
rect 712 1717 715 1749
rect 747 1717 779 1749
rect 712 1716 779 1717
rect 961 1749 1028 1750
rect 961 1717 993 1749
rect 1025 1717 1028 1749
rect 961 1716 1028 1717
rect 712 1714 750 1716
rect 990 1714 1028 1716
rect 1060 1750 1098 1752
rect 1338 1750 1376 1752
rect 1060 1749 1127 1750
rect 1060 1717 1063 1749
rect 1095 1717 1127 1749
rect 1060 1716 1127 1717
rect 1309 1749 1376 1750
rect 1309 1717 1341 1749
rect 1373 1717 1376 1749
rect 1309 1716 1376 1717
rect 1060 1714 1098 1716
rect 1338 1714 1376 1716
rect 1408 1750 1446 1752
rect 1686 1750 1724 1752
rect 1408 1749 1475 1750
rect 1408 1717 1411 1749
rect 1443 1717 1475 1749
rect 1408 1716 1475 1717
rect 1657 1749 1724 1750
rect 1657 1717 1689 1749
rect 1721 1717 1724 1749
rect 1657 1716 1724 1717
rect 1408 1714 1446 1716
rect 1686 1714 1724 1716
rect 1756 1750 1794 1752
rect 2034 1750 2072 1752
rect 1756 1749 1823 1750
rect 1756 1717 1759 1749
rect 1791 1717 1823 1749
rect 1756 1716 1823 1717
rect 2005 1749 2072 1750
rect 2005 1717 2037 1749
rect 2069 1717 2072 1749
rect 2005 1716 2072 1717
rect 1756 1714 1794 1716
rect 2034 1714 2072 1716
rect 2104 1750 2142 1752
rect 2382 1750 2420 1752
rect 2104 1749 2171 1750
rect 2104 1717 2107 1749
rect 2139 1717 2171 1749
rect 2104 1716 2171 1717
rect 2353 1749 2420 1750
rect 2353 1717 2385 1749
rect 2417 1717 2420 1749
rect 2353 1716 2420 1717
rect 2104 1714 2142 1716
rect 2382 1714 2420 1716
rect 2452 1750 2490 1752
rect 2730 1750 2768 1752
rect 2452 1749 2519 1750
rect 2452 1717 2455 1749
rect 2487 1717 2519 1749
rect 2452 1716 2519 1717
rect 2701 1749 2768 1750
rect 2701 1717 2733 1749
rect 2765 1717 2768 1749
rect 2701 1716 2768 1717
rect 2452 1714 2490 1716
rect 2730 1714 2768 1716
rect 2800 1750 2838 1752
rect 3078 1750 3116 1752
rect 2800 1749 2867 1750
rect 2800 1717 2803 1749
rect 2835 1717 2867 1749
rect 2800 1716 2867 1717
rect 3049 1749 3116 1750
rect 3049 1717 3081 1749
rect 3113 1717 3116 1749
rect 3049 1716 3116 1717
rect 2800 1714 2838 1716
rect 3078 1714 3116 1716
rect 3148 1750 3186 1752
rect 3426 1750 3464 1752
rect 3148 1749 3215 1750
rect 3148 1717 3151 1749
rect 3183 1717 3215 1749
rect 3148 1716 3215 1717
rect 3397 1749 3464 1750
rect 3397 1717 3429 1749
rect 3461 1717 3464 1749
rect 3397 1716 3464 1717
rect 3148 1714 3186 1716
rect 3426 1714 3464 1716
rect 3496 1750 3534 1752
rect 3774 1750 3812 1752
rect 3496 1749 3563 1750
rect 3496 1717 3499 1749
rect 3531 1717 3563 1749
rect 3496 1716 3563 1717
rect 3745 1749 3812 1750
rect 3745 1717 3777 1749
rect 3809 1717 3812 1749
rect 3745 1716 3812 1717
rect 3496 1714 3534 1716
rect 3774 1714 3812 1716
rect 3844 1750 3882 1752
rect 4122 1750 4160 1752
rect 3844 1749 3911 1750
rect 3844 1717 3847 1749
rect 3879 1717 3911 1749
rect 3844 1716 3911 1717
rect 4093 1749 4160 1750
rect 4093 1717 4125 1749
rect 4157 1717 4160 1749
rect 4093 1716 4160 1717
rect 3844 1714 3882 1716
rect 4122 1714 4160 1716
rect 4192 1750 4230 1752
rect 4470 1750 4508 1752
rect 4192 1749 4259 1750
rect 4192 1717 4195 1749
rect 4227 1717 4259 1749
rect 4192 1716 4259 1717
rect 4441 1749 4508 1750
rect 4441 1717 4473 1749
rect 4505 1717 4508 1749
rect 4441 1716 4508 1717
rect 4192 1714 4230 1716
rect 4470 1714 4508 1716
rect 4540 1750 4578 1752
rect 4818 1750 4856 1752
rect 4540 1749 4607 1750
rect 4540 1717 4543 1749
rect 4575 1717 4607 1749
rect 4540 1716 4607 1717
rect 4789 1749 4856 1750
rect 4789 1717 4821 1749
rect 4853 1717 4856 1749
rect 4789 1716 4856 1717
rect 4540 1714 4578 1716
rect 4818 1714 4856 1716
rect 4888 1750 4926 1752
rect 5166 1750 5204 1752
rect 4888 1749 4955 1750
rect 4888 1717 4891 1749
rect 4923 1717 4955 1749
rect 4888 1716 4955 1717
rect 5137 1749 5204 1750
rect 5137 1717 5169 1749
rect 5201 1717 5204 1749
rect 5137 1716 5204 1717
rect 4888 1714 4926 1716
rect 5166 1714 5204 1716
rect 5236 1750 5274 1752
rect 5514 1750 5552 1752
rect 5236 1749 5303 1750
rect 5236 1717 5239 1749
rect 5271 1717 5303 1749
rect 5236 1716 5303 1717
rect 5485 1749 5552 1750
rect 5485 1717 5517 1749
rect 5549 1717 5552 1749
rect 5485 1716 5552 1717
rect 5236 1714 5274 1716
rect 5514 1714 5552 1716
rect 5584 1750 5622 1752
rect 5862 1750 5900 1752
rect 5584 1749 5651 1750
rect 5584 1717 5587 1749
rect 5619 1717 5651 1749
rect 5584 1716 5651 1717
rect 5833 1749 5900 1750
rect 5833 1717 5865 1749
rect 5897 1717 5900 1749
rect 5833 1716 5900 1717
rect 5584 1714 5622 1716
rect 5862 1714 5900 1716
rect 5932 1750 5970 1752
rect 6210 1750 6248 1752
rect 5932 1749 5999 1750
rect 5932 1717 5935 1749
rect 5967 1717 5999 1749
rect 5932 1716 5999 1717
rect 6181 1749 6248 1750
rect 6181 1717 6213 1749
rect 6245 1717 6248 1749
rect 6181 1716 6248 1717
rect 5932 1714 5970 1716
rect 6210 1714 6248 1716
rect 6280 1750 6318 1752
rect 6558 1750 6596 1752
rect 6280 1749 6347 1750
rect 6280 1717 6283 1749
rect 6315 1717 6347 1749
rect 6280 1716 6347 1717
rect 6529 1749 6596 1750
rect 6529 1717 6561 1749
rect 6593 1717 6596 1749
rect 6529 1716 6596 1717
rect 6280 1714 6318 1716
rect 6558 1714 6596 1716
rect 6628 1750 6666 1752
rect 6906 1750 6944 1752
rect 6628 1749 6695 1750
rect 6628 1717 6631 1749
rect 6663 1717 6695 1749
rect 6628 1716 6695 1717
rect 6877 1749 6944 1750
rect 6877 1717 6909 1749
rect 6941 1717 6944 1749
rect 6877 1716 6944 1717
rect 6628 1714 6666 1716
rect 6906 1714 6944 1716
rect 6976 1750 7014 1752
rect 7254 1750 7292 1752
rect 6976 1749 7043 1750
rect 6976 1717 6979 1749
rect 7011 1717 7043 1749
rect 6976 1716 7043 1717
rect 7225 1749 7292 1750
rect 7225 1717 7257 1749
rect 7289 1717 7292 1749
rect 7225 1716 7292 1717
rect 6976 1714 7014 1716
rect 7254 1714 7292 1716
rect 16 1680 54 1682
rect 294 1680 332 1682
rect 16 1679 83 1680
rect 16 1647 19 1679
rect 51 1647 83 1679
rect 16 1646 83 1647
rect 265 1679 332 1680
rect 265 1647 297 1679
rect 329 1647 332 1679
rect 265 1646 332 1647
rect 16 1644 54 1646
rect 294 1644 332 1646
rect 364 1680 402 1682
rect 642 1680 680 1682
rect 364 1679 431 1680
rect 364 1647 367 1679
rect 399 1647 431 1679
rect 364 1646 431 1647
rect 613 1679 680 1680
rect 613 1647 645 1679
rect 677 1647 680 1679
rect 613 1646 680 1647
rect 364 1644 402 1646
rect 642 1644 680 1646
rect 712 1680 750 1682
rect 990 1680 1028 1682
rect 712 1679 779 1680
rect 712 1647 715 1679
rect 747 1647 779 1679
rect 712 1646 779 1647
rect 961 1679 1028 1680
rect 961 1647 993 1679
rect 1025 1647 1028 1679
rect 961 1646 1028 1647
rect 712 1644 750 1646
rect 990 1644 1028 1646
rect 1060 1680 1098 1682
rect 1338 1680 1376 1682
rect 1060 1679 1127 1680
rect 1060 1647 1063 1679
rect 1095 1647 1127 1679
rect 1060 1646 1127 1647
rect 1309 1679 1376 1680
rect 1309 1647 1341 1679
rect 1373 1647 1376 1679
rect 1309 1646 1376 1647
rect 1060 1644 1098 1646
rect 1338 1644 1376 1646
rect 1408 1680 1446 1682
rect 1686 1680 1724 1682
rect 1408 1679 1475 1680
rect 1408 1647 1411 1679
rect 1443 1647 1475 1679
rect 1408 1646 1475 1647
rect 1657 1679 1724 1680
rect 1657 1647 1689 1679
rect 1721 1647 1724 1679
rect 1657 1646 1724 1647
rect 1408 1644 1446 1646
rect 1686 1644 1724 1646
rect 1756 1680 1794 1682
rect 2034 1680 2072 1682
rect 1756 1679 1823 1680
rect 1756 1647 1759 1679
rect 1791 1647 1823 1679
rect 1756 1646 1823 1647
rect 2005 1679 2072 1680
rect 2005 1647 2037 1679
rect 2069 1647 2072 1679
rect 2005 1646 2072 1647
rect 1756 1644 1794 1646
rect 2034 1644 2072 1646
rect 2104 1680 2142 1682
rect 2382 1680 2420 1682
rect 2104 1679 2171 1680
rect 2104 1647 2107 1679
rect 2139 1647 2171 1679
rect 2104 1646 2171 1647
rect 2353 1679 2420 1680
rect 2353 1647 2385 1679
rect 2417 1647 2420 1679
rect 2353 1646 2420 1647
rect 2104 1644 2142 1646
rect 2382 1644 2420 1646
rect 2452 1680 2490 1682
rect 2730 1680 2768 1682
rect 2452 1679 2519 1680
rect 2452 1647 2455 1679
rect 2487 1647 2519 1679
rect 2452 1646 2519 1647
rect 2701 1679 2768 1680
rect 2701 1647 2733 1679
rect 2765 1647 2768 1679
rect 2701 1646 2768 1647
rect 2452 1644 2490 1646
rect 2730 1644 2768 1646
rect 2800 1680 2838 1682
rect 3078 1680 3116 1682
rect 2800 1679 2867 1680
rect 2800 1647 2803 1679
rect 2835 1647 2867 1679
rect 2800 1646 2867 1647
rect 3049 1679 3116 1680
rect 3049 1647 3081 1679
rect 3113 1647 3116 1679
rect 3049 1646 3116 1647
rect 2800 1644 2838 1646
rect 3078 1644 3116 1646
rect 3148 1680 3186 1682
rect 3426 1680 3464 1682
rect 3148 1679 3215 1680
rect 3148 1647 3151 1679
rect 3183 1647 3215 1679
rect 3148 1646 3215 1647
rect 3397 1679 3464 1680
rect 3397 1647 3429 1679
rect 3461 1647 3464 1679
rect 3397 1646 3464 1647
rect 3148 1644 3186 1646
rect 3426 1644 3464 1646
rect 3496 1680 3534 1682
rect 3774 1680 3812 1682
rect 3496 1679 3563 1680
rect 3496 1647 3499 1679
rect 3531 1647 3563 1679
rect 3496 1646 3563 1647
rect 3745 1679 3812 1680
rect 3745 1647 3777 1679
rect 3809 1647 3812 1679
rect 3745 1646 3812 1647
rect 3496 1644 3534 1646
rect 3774 1644 3812 1646
rect 3844 1680 3882 1682
rect 4122 1680 4160 1682
rect 3844 1679 3911 1680
rect 3844 1647 3847 1679
rect 3879 1647 3911 1679
rect 3844 1646 3911 1647
rect 4093 1679 4160 1680
rect 4093 1647 4125 1679
rect 4157 1647 4160 1679
rect 4093 1646 4160 1647
rect 3844 1644 3882 1646
rect 4122 1644 4160 1646
rect 4192 1680 4230 1682
rect 4470 1680 4508 1682
rect 4192 1679 4259 1680
rect 4192 1647 4195 1679
rect 4227 1647 4259 1679
rect 4192 1646 4259 1647
rect 4441 1679 4508 1680
rect 4441 1647 4473 1679
rect 4505 1647 4508 1679
rect 4441 1646 4508 1647
rect 4192 1644 4230 1646
rect 4470 1644 4508 1646
rect 4540 1680 4578 1682
rect 4818 1680 4856 1682
rect 4540 1679 4607 1680
rect 4540 1647 4543 1679
rect 4575 1647 4607 1679
rect 4540 1646 4607 1647
rect 4789 1679 4856 1680
rect 4789 1647 4821 1679
rect 4853 1647 4856 1679
rect 4789 1646 4856 1647
rect 4540 1644 4578 1646
rect 4818 1644 4856 1646
rect 4888 1680 4926 1682
rect 5166 1680 5204 1682
rect 4888 1679 4955 1680
rect 4888 1647 4891 1679
rect 4923 1647 4955 1679
rect 4888 1646 4955 1647
rect 5137 1679 5204 1680
rect 5137 1647 5169 1679
rect 5201 1647 5204 1679
rect 5137 1646 5204 1647
rect 4888 1644 4926 1646
rect 5166 1644 5204 1646
rect 5236 1680 5274 1682
rect 5514 1680 5552 1682
rect 5236 1679 5303 1680
rect 5236 1647 5239 1679
rect 5271 1647 5303 1679
rect 5236 1646 5303 1647
rect 5485 1679 5552 1680
rect 5485 1647 5517 1679
rect 5549 1647 5552 1679
rect 5485 1646 5552 1647
rect 5236 1644 5274 1646
rect 5514 1644 5552 1646
rect 5584 1680 5622 1682
rect 5862 1680 5900 1682
rect 5584 1679 5651 1680
rect 5584 1647 5587 1679
rect 5619 1647 5651 1679
rect 5584 1646 5651 1647
rect 5833 1679 5900 1680
rect 5833 1647 5865 1679
rect 5897 1647 5900 1679
rect 5833 1646 5900 1647
rect 5584 1644 5622 1646
rect 5862 1644 5900 1646
rect 5932 1680 5970 1682
rect 6210 1680 6248 1682
rect 5932 1679 5999 1680
rect 5932 1647 5935 1679
rect 5967 1647 5999 1679
rect 5932 1646 5999 1647
rect 6181 1679 6248 1680
rect 6181 1647 6213 1679
rect 6245 1647 6248 1679
rect 6181 1646 6248 1647
rect 5932 1644 5970 1646
rect 6210 1644 6248 1646
rect 6280 1680 6318 1682
rect 6558 1680 6596 1682
rect 6280 1679 6347 1680
rect 6280 1647 6283 1679
rect 6315 1647 6347 1679
rect 6280 1646 6347 1647
rect 6529 1679 6596 1680
rect 6529 1647 6561 1679
rect 6593 1647 6596 1679
rect 6529 1646 6596 1647
rect 6280 1644 6318 1646
rect 6558 1644 6596 1646
rect 6628 1680 6666 1682
rect 6906 1680 6944 1682
rect 6628 1679 6695 1680
rect 6628 1647 6631 1679
rect 6663 1647 6695 1679
rect 6628 1646 6695 1647
rect 6877 1679 6944 1680
rect 6877 1647 6909 1679
rect 6941 1647 6944 1679
rect 6877 1646 6944 1647
rect 6628 1644 6666 1646
rect 6906 1644 6944 1646
rect 6976 1680 7014 1682
rect 7254 1680 7292 1682
rect 6976 1679 7043 1680
rect 6976 1647 6979 1679
rect 7011 1647 7043 1679
rect 6976 1646 7043 1647
rect 7225 1679 7292 1680
rect 7225 1647 7257 1679
rect 7289 1647 7292 1679
rect 7225 1646 7292 1647
rect 6976 1644 7014 1646
rect 7254 1644 7292 1646
rect 16 1556 54 1558
rect 294 1556 332 1558
rect 16 1555 83 1556
rect 16 1523 19 1555
rect 51 1523 83 1555
rect 16 1522 83 1523
rect 265 1555 332 1556
rect 265 1523 297 1555
rect 329 1523 332 1555
rect 265 1522 332 1523
rect 16 1520 54 1522
rect 294 1520 332 1522
rect 364 1556 402 1558
rect 642 1556 680 1558
rect 364 1555 431 1556
rect 364 1523 367 1555
rect 399 1523 431 1555
rect 364 1522 431 1523
rect 613 1555 680 1556
rect 613 1523 645 1555
rect 677 1523 680 1555
rect 613 1522 680 1523
rect 364 1520 402 1522
rect 642 1520 680 1522
rect 712 1556 750 1558
rect 990 1556 1028 1558
rect 712 1555 779 1556
rect 712 1523 715 1555
rect 747 1523 779 1555
rect 712 1522 779 1523
rect 961 1555 1028 1556
rect 961 1523 993 1555
rect 1025 1523 1028 1555
rect 961 1522 1028 1523
rect 712 1520 750 1522
rect 990 1520 1028 1522
rect 1060 1556 1098 1558
rect 1338 1556 1376 1558
rect 1060 1555 1127 1556
rect 1060 1523 1063 1555
rect 1095 1523 1127 1555
rect 1060 1522 1127 1523
rect 1309 1555 1376 1556
rect 1309 1523 1341 1555
rect 1373 1523 1376 1555
rect 1309 1522 1376 1523
rect 1060 1520 1098 1522
rect 1338 1520 1376 1522
rect 1408 1556 1446 1558
rect 1686 1556 1724 1558
rect 1408 1555 1475 1556
rect 1408 1523 1411 1555
rect 1443 1523 1475 1555
rect 1408 1522 1475 1523
rect 1657 1555 1724 1556
rect 1657 1523 1689 1555
rect 1721 1523 1724 1555
rect 1657 1522 1724 1523
rect 1408 1520 1446 1522
rect 1686 1520 1724 1522
rect 1756 1556 1794 1558
rect 2034 1556 2072 1558
rect 1756 1555 1823 1556
rect 1756 1523 1759 1555
rect 1791 1523 1823 1555
rect 1756 1522 1823 1523
rect 2005 1555 2072 1556
rect 2005 1523 2037 1555
rect 2069 1523 2072 1555
rect 2005 1522 2072 1523
rect 1756 1520 1794 1522
rect 2034 1520 2072 1522
rect 2104 1556 2142 1558
rect 2382 1556 2420 1558
rect 2104 1555 2171 1556
rect 2104 1523 2107 1555
rect 2139 1523 2171 1555
rect 2104 1522 2171 1523
rect 2353 1555 2420 1556
rect 2353 1523 2385 1555
rect 2417 1523 2420 1555
rect 2353 1522 2420 1523
rect 2104 1520 2142 1522
rect 2382 1520 2420 1522
rect 2452 1556 2490 1558
rect 2730 1556 2768 1558
rect 2452 1555 2519 1556
rect 2452 1523 2455 1555
rect 2487 1523 2519 1555
rect 2452 1522 2519 1523
rect 2701 1555 2768 1556
rect 2701 1523 2733 1555
rect 2765 1523 2768 1555
rect 2701 1522 2768 1523
rect 2452 1520 2490 1522
rect 2730 1520 2768 1522
rect 2800 1556 2838 1558
rect 3078 1556 3116 1558
rect 2800 1555 2867 1556
rect 2800 1523 2803 1555
rect 2835 1523 2867 1555
rect 2800 1522 2867 1523
rect 3049 1555 3116 1556
rect 3049 1523 3081 1555
rect 3113 1523 3116 1555
rect 3049 1522 3116 1523
rect 2800 1520 2838 1522
rect 3078 1520 3116 1522
rect 3148 1556 3186 1558
rect 3426 1556 3464 1558
rect 3148 1555 3215 1556
rect 3148 1523 3151 1555
rect 3183 1523 3215 1555
rect 3148 1522 3215 1523
rect 3397 1555 3464 1556
rect 3397 1523 3429 1555
rect 3461 1523 3464 1555
rect 3397 1522 3464 1523
rect 3148 1520 3186 1522
rect 3426 1520 3464 1522
rect 3496 1556 3534 1558
rect 3774 1556 3812 1558
rect 3496 1555 3563 1556
rect 3496 1523 3499 1555
rect 3531 1523 3563 1555
rect 3496 1522 3563 1523
rect 3745 1555 3812 1556
rect 3745 1523 3777 1555
rect 3809 1523 3812 1555
rect 3745 1522 3812 1523
rect 3496 1520 3534 1522
rect 3774 1520 3812 1522
rect 3844 1556 3882 1558
rect 4122 1556 4160 1558
rect 3844 1555 3911 1556
rect 3844 1523 3847 1555
rect 3879 1523 3911 1555
rect 3844 1522 3911 1523
rect 4093 1555 4160 1556
rect 4093 1523 4125 1555
rect 4157 1523 4160 1555
rect 4093 1522 4160 1523
rect 3844 1520 3882 1522
rect 4122 1520 4160 1522
rect 4192 1556 4230 1558
rect 4470 1556 4508 1558
rect 4192 1555 4259 1556
rect 4192 1523 4195 1555
rect 4227 1523 4259 1555
rect 4192 1522 4259 1523
rect 4441 1555 4508 1556
rect 4441 1523 4473 1555
rect 4505 1523 4508 1555
rect 4441 1522 4508 1523
rect 4192 1520 4230 1522
rect 4470 1520 4508 1522
rect 4540 1556 4578 1558
rect 4818 1556 4856 1558
rect 4540 1555 4607 1556
rect 4540 1523 4543 1555
rect 4575 1523 4607 1555
rect 4540 1522 4607 1523
rect 4789 1555 4856 1556
rect 4789 1523 4821 1555
rect 4853 1523 4856 1555
rect 4789 1522 4856 1523
rect 4540 1520 4578 1522
rect 4818 1520 4856 1522
rect 4888 1556 4926 1558
rect 5166 1556 5204 1558
rect 4888 1555 4955 1556
rect 4888 1523 4891 1555
rect 4923 1523 4955 1555
rect 4888 1522 4955 1523
rect 5137 1555 5204 1556
rect 5137 1523 5169 1555
rect 5201 1523 5204 1555
rect 5137 1522 5204 1523
rect 4888 1520 4926 1522
rect 5166 1520 5204 1522
rect 5236 1556 5274 1558
rect 5514 1556 5552 1558
rect 5236 1555 5303 1556
rect 5236 1523 5239 1555
rect 5271 1523 5303 1555
rect 5236 1522 5303 1523
rect 5485 1555 5552 1556
rect 5485 1523 5517 1555
rect 5549 1523 5552 1555
rect 5485 1522 5552 1523
rect 5236 1520 5274 1522
rect 5514 1520 5552 1522
rect 5584 1556 5622 1558
rect 5862 1556 5900 1558
rect 5584 1555 5651 1556
rect 5584 1523 5587 1555
rect 5619 1523 5651 1555
rect 5584 1522 5651 1523
rect 5833 1555 5900 1556
rect 5833 1523 5865 1555
rect 5897 1523 5900 1555
rect 5833 1522 5900 1523
rect 5584 1520 5622 1522
rect 5862 1520 5900 1522
rect 5932 1556 5970 1558
rect 6210 1556 6248 1558
rect 5932 1555 5999 1556
rect 5932 1523 5935 1555
rect 5967 1523 5999 1555
rect 5932 1522 5999 1523
rect 6181 1555 6248 1556
rect 6181 1523 6213 1555
rect 6245 1523 6248 1555
rect 6181 1522 6248 1523
rect 5932 1520 5970 1522
rect 6210 1520 6248 1522
rect 6280 1556 6318 1558
rect 6558 1556 6596 1558
rect 6280 1555 6347 1556
rect 6280 1523 6283 1555
rect 6315 1523 6347 1555
rect 6280 1522 6347 1523
rect 6529 1555 6596 1556
rect 6529 1523 6561 1555
rect 6593 1523 6596 1555
rect 6529 1522 6596 1523
rect 6280 1520 6318 1522
rect 6558 1520 6596 1522
rect 6628 1556 6666 1558
rect 6906 1556 6944 1558
rect 6628 1555 6695 1556
rect 6628 1523 6631 1555
rect 6663 1523 6695 1555
rect 6628 1522 6695 1523
rect 6877 1555 6944 1556
rect 6877 1523 6909 1555
rect 6941 1523 6944 1555
rect 6877 1522 6944 1523
rect 6628 1520 6666 1522
rect 6906 1520 6944 1522
rect 6976 1556 7014 1558
rect 7254 1556 7292 1558
rect 6976 1555 7043 1556
rect 6976 1523 6979 1555
rect 7011 1523 7043 1555
rect 6976 1522 7043 1523
rect 7225 1555 7292 1556
rect 7225 1523 7257 1555
rect 7289 1523 7292 1555
rect 7225 1522 7292 1523
rect 6976 1520 7014 1522
rect 7254 1520 7292 1522
rect 16 1432 54 1434
rect 294 1432 332 1434
rect 16 1431 83 1432
rect 16 1399 19 1431
rect 51 1399 83 1431
rect 16 1398 83 1399
rect 265 1431 332 1432
rect 265 1399 297 1431
rect 329 1399 332 1431
rect 265 1398 332 1399
rect 16 1396 54 1398
rect 294 1396 332 1398
rect 364 1432 402 1434
rect 642 1432 680 1434
rect 364 1431 431 1432
rect 364 1399 367 1431
rect 399 1399 431 1431
rect 364 1398 431 1399
rect 613 1431 680 1432
rect 613 1399 645 1431
rect 677 1399 680 1431
rect 613 1398 680 1399
rect 364 1396 402 1398
rect 642 1396 680 1398
rect 712 1432 750 1434
rect 990 1432 1028 1434
rect 712 1431 779 1432
rect 712 1399 715 1431
rect 747 1399 779 1431
rect 712 1398 779 1399
rect 961 1431 1028 1432
rect 961 1399 993 1431
rect 1025 1399 1028 1431
rect 961 1398 1028 1399
rect 712 1396 750 1398
rect 990 1396 1028 1398
rect 1060 1432 1098 1434
rect 1338 1432 1376 1434
rect 1060 1431 1127 1432
rect 1060 1399 1063 1431
rect 1095 1399 1127 1431
rect 1060 1398 1127 1399
rect 1309 1431 1376 1432
rect 1309 1399 1341 1431
rect 1373 1399 1376 1431
rect 1309 1398 1376 1399
rect 1060 1396 1098 1398
rect 1338 1396 1376 1398
rect 1408 1432 1446 1434
rect 1686 1432 1724 1434
rect 1408 1431 1475 1432
rect 1408 1399 1411 1431
rect 1443 1399 1475 1431
rect 1408 1398 1475 1399
rect 1657 1431 1724 1432
rect 1657 1399 1689 1431
rect 1721 1399 1724 1431
rect 1657 1398 1724 1399
rect 1408 1396 1446 1398
rect 1686 1396 1724 1398
rect 1756 1432 1794 1434
rect 2034 1432 2072 1434
rect 1756 1431 1823 1432
rect 1756 1399 1759 1431
rect 1791 1399 1823 1431
rect 1756 1398 1823 1399
rect 2005 1431 2072 1432
rect 2005 1399 2037 1431
rect 2069 1399 2072 1431
rect 2005 1398 2072 1399
rect 1756 1396 1794 1398
rect 2034 1396 2072 1398
rect 2104 1432 2142 1434
rect 2382 1432 2420 1434
rect 2104 1431 2171 1432
rect 2104 1399 2107 1431
rect 2139 1399 2171 1431
rect 2104 1398 2171 1399
rect 2353 1431 2420 1432
rect 2353 1399 2385 1431
rect 2417 1399 2420 1431
rect 2353 1398 2420 1399
rect 2104 1396 2142 1398
rect 2382 1396 2420 1398
rect 2452 1432 2490 1434
rect 2730 1432 2768 1434
rect 2452 1431 2519 1432
rect 2452 1399 2455 1431
rect 2487 1399 2519 1431
rect 2452 1398 2519 1399
rect 2701 1431 2768 1432
rect 2701 1399 2733 1431
rect 2765 1399 2768 1431
rect 2701 1398 2768 1399
rect 2452 1396 2490 1398
rect 2730 1396 2768 1398
rect 2800 1432 2838 1434
rect 3078 1432 3116 1434
rect 2800 1431 2867 1432
rect 2800 1399 2803 1431
rect 2835 1399 2867 1431
rect 2800 1398 2867 1399
rect 3049 1431 3116 1432
rect 3049 1399 3081 1431
rect 3113 1399 3116 1431
rect 3049 1398 3116 1399
rect 2800 1396 2838 1398
rect 3078 1396 3116 1398
rect 3148 1432 3186 1434
rect 3426 1432 3464 1434
rect 3148 1431 3215 1432
rect 3148 1399 3151 1431
rect 3183 1399 3215 1431
rect 3148 1398 3215 1399
rect 3397 1431 3464 1432
rect 3397 1399 3429 1431
rect 3461 1399 3464 1431
rect 3397 1398 3464 1399
rect 3148 1396 3186 1398
rect 3426 1396 3464 1398
rect 3496 1432 3534 1434
rect 3774 1432 3812 1434
rect 3496 1431 3563 1432
rect 3496 1399 3499 1431
rect 3531 1399 3563 1431
rect 3496 1398 3563 1399
rect 3745 1431 3812 1432
rect 3745 1399 3777 1431
rect 3809 1399 3812 1431
rect 3745 1398 3812 1399
rect 3496 1396 3534 1398
rect 3774 1396 3812 1398
rect 3844 1432 3882 1434
rect 4122 1432 4160 1434
rect 3844 1431 3911 1432
rect 3844 1399 3847 1431
rect 3879 1399 3911 1431
rect 3844 1398 3911 1399
rect 4093 1431 4160 1432
rect 4093 1399 4125 1431
rect 4157 1399 4160 1431
rect 4093 1398 4160 1399
rect 3844 1396 3882 1398
rect 4122 1396 4160 1398
rect 4192 1432 4230 1434
rect 4470 1432 4508 1434
rect 4192 1431 4259 1432
rect 4192 1399 4195 1431
rect 4227 1399 4259 1431
rect 4192 1398 4259 1399
rect 4441 1431 4508 1432
rect 4441 1399 4473 1431
rect 4505 1399 4508 1431
rect 4441 1398 4508 1399
rect 4192 1396 4230 1398
rect 4470 1396 4508 1398
rect 4540 1432 4578 1434
rect 4818 1432 4856 1434
rect 4540 1431 4607 1432
rect 4540 1399 4543 1431
rect 4575 1399 4607 1431
rect 4540 1398 4607 1399
rect 4789 1431 4856 1432
rect 4789 1399 4821 1431
rect 4853 1399 4856 1431
rect 4789 1398 4856 1399
rect 4540 1396 4578 1398
rect 4818 1396 4856 1398
rect 4888 1432 4926 1434
rect 5166 1432 5204 1434
rect 4888 1431 4955 1432
rect 4888 1399 4891 1431
rect 4923 1399 4955 1431
rect 4888 1398 4955 1399
rect 5137 1431 5204 1432
rect 5137 1399 5169 1431
rect 5201 1399 5204 1431
rect 5137 1398 5204 1399
rect 4888 1396 4926 1398
rect 5166 1396 5204 1398
rect 5236 1432 5274 1434
rect 5514 1432 5552 1434
rect 5236 1431 5303 1432
rect 5236 1399 5239 1431
rect 5271 1399 5303 1431
rect 5236 1398 5303 1399
rect 5485 1431 5552 1432
rect 5485 1399 5517 1431
rect 5549 1399 5552 1431
rect 5485 1398 5552 1399
rect 5236 1396 5274 1398
rect 5514 1396 5552 1398
rect 5584 1432 5622 1434
rect 5862 1432 5900 1434
rect 5584 1431 5651 1432
rect 5584 1399 5587 1431
rect 5619 1399 5651 1431
rect 5584 1398 5651 1399
rect 5833 1431 5900 1432
rect 5833 1399 5865 1431
rect 5897 1399 5900 1431
rect 5833 1398 5900 1399
rect 5584 1396 5622 1398
rect 5862 1396 5900 1398
rect 5932 1432 5970 1434
rect 6210 1432 6248 1434
rect 5932 1431 5999 1432
rect 5932 1399 5935 1431
rect 5967 1399 5999 1431
rect 5932 1398 5999 1399
rect 6181 1431 6248 1432
rect 6181 1399 6213 1431
rect 6245 1399 6248 1431
rect 6181 1398 6248 1399
rect 5932 1396 5970 1398
rect 6210 1396 6248 1398
rect 6280 1432 6318 1434
rect 6558 1432 6596 1434
rect 6280 1431 6347 1432
rect 6280 1399 6283 1431
rect 6315 1399 6347 1431
rect 6280 1398 6347 1399
rect 6529 1431 6596 1432
rect 6529 1399 6561 1431
rect 6593 1399 6596 1431
rect 6529 1398 6596 1399
rect 6280 1396 6318 1398
rect 6558 1396 6596 1398
rect 6628 1432 6666 1434
rect 6906 1432 6944 1434
rect 6628 1431 6695 1432
rect 6628 1399 6631 1431
rect 6663 1399 6695 1431
rect 6628 1398 6695 1399
rect 6877 1431 6944 1432
rect 6877 1399 6909 1431
rect 6941 1399 6944 1431
rect 6877 1398 6944 1399
rect 6628 1396 6666 1398
rect 6906 1396 6944 1398
rect 6976 1432 7014 1434
rect 7254 1432 7292 1434
rect 6976 1431 7043 1432
rect 6976 1399 6979 1431
rect 7011 1399 7043 1431
rect 6976 1398 7043 1399
rect 7225 1431 7292 1432
rect 7225 1399 7257 1431
rect 7289 1399 7292 1431
rect 7225 1398 7292 1399
rect 6976 1396 7014 1398
rect 7254 1396 7292 1398
rect 16 1308 54 1310
rect 294 1308 332 1310
rect 16 1307 83 1308
rect 16 1275 19 1307
rect 51 1275 83 1307
rect 16 1274 83 1275
rect 265 1307 332 1308
rect 265 1275 297 1307
rect 329 1275 332 1307
rect 265 1274 332 1275
rect 16 1272 54 1274
rect 294 1272 332 1274
rect 364 1308 402 1310
rect 642 1308 680 1310
rect 364 1307 431 1308
rect 364 1275 367 1307
rect 399 1275 431 1307
rect 364 1274 431 1275
rect 613 1307 680 1308
rect 613 1275 645 1307
rect 677 1275 680 1307
rect 613 1274 680 1275
rect 364 1272 402 1274
rect 642 1272 680 1274
rect 712 1308 750 1310
rect 990 1308 1028 1310
rect 712 1307 779 1308
rect 712 1275 715 1307
rect 747 1275 779 1307
rect 712 1274 779 1275
rect 961 1307 1028 1308
rect 961 1275 993 1307
rect 1025 1275 1028 1307
rect 961 1274 1028 1275
rect 712 1272 750 1274
rect 990 1272 1028 1274
rect 1060 1308 1098 1310
rect 1338 1308 1376 1310
rect 1060 1307 1127 1308
rect 1060 1275 1063 1307
rect 1095 1275 1127 1307
rect 1060 1274 1127 1275
rect 1309 1307 1376 1308
rect 1309 1275 1341 1307
rect 1373 1275 1376 1307
rect 1309 1274 1376 1275
rect 1060 1272 1098 1274
rect 1338 1272 1376 1274
rect 1408 1308 1446 1310
rect 1686 1308 1724 1310
rect 1408 1307 1475 1308
rect 1408 1275 1411 1307
rect 1443 1275 1475 1307
rect 1408 1274 1475 1275
rect 1657 1307 1724 1308
rect 1657 1275 1689 1307
rect 1721 1275 1724 1307
rect 1657 1274 1724 1275
rect 1408 1272 1446 1274
rect 1686 1272 1724 1274
rect 1756 1308 1794 1310
rect 2034 1308 2072 1310
rect 1756 1307 1823 1308
rect 1756 1275 1759 1307
rect 1791 1275 1823 1307
rect 1756 1274 1823 1275
rect 2005 1307 2072 1308
rect 2005 1275 2037 1307
rect 2069 1275 2072 1307
rect 2005 1274 2072 1275
rect 1756 1272 1794 1274
rect 2034 1272 2072 1274
rect 2104 1308 2142 1310
rect 2382 1308 2420 1310
rect 2104 1307 2171 1308
rect 2104 1275 2107 1307
rect 2139 1275 2171 1307
rect 2104 1274 2171 1275
rect 2353 1307 2420 1308
rect 2353 1275 2385 1307
rect 2417 1275 2420 1307
rect 2353 1274 2420 1275
rect 2104 1272 2142 1274
rect 2382 1272 2420 1274
rect 2452 1308 2490 1310
rect 2730 1308 2768 1310
rect 2452 1307 2519 1308
rect 2452 1275 2455 1307
rect 2487 1275 2519 1307
rect 2452 1274 2519 1275
rect 2701 1307 2768 1308
rect 2701 1275 2733 1307
rect 2765 1275 2768 1307
rect 2701 1274 2768 1275
rect 2452 1272 2490 1274
rect 2730 1272 2768 1274
rect 2800 1308 2838 1310
rect 3078 1308 3116 1310
rect 2800 1307 2867 1308
rect 2800 1275 2803 1307
rect 2835 1275 2867 1307
rect 2800 1274 2867 1275
rect 3049 1307 3116 1308
rect 3049 1275 3081 1307
rect 3113 1275 3116 1307
rect 3049 1274 3116 1275
rect 2800 1272 2838 1274
rect 3078 1272 3116 1274
rect 3148 1308 3186 1310
rect 3426 1308 3464 1310
rect 3148 1307 3215 1308
rect 3148 1275 3151 1307
rect 3183 1275 3215 1307
rect 3148 1274 3215 1275
rect 3397 1307 3464 1308
rect 3397 1275 3429 1307
rect 3461 1275 3464 1307
rect 3397 1274 3464 1275
rect 3148 1272 3186 1274
rect 3426 1272 3464 1274
rect 3496 1308 3534 1310
rect 3774 1308 3812 1310
rect 3496 1307 3563 1308
rect 3496 1275 3499 1307
rect 3531 1275 3563 1307
rect 3496 1274 3563 1275
rect 3745 1307 3812 1308
rect 3745 1275 3777 1307
rect 3809 1275 3812 1307
rect 3745 1274 3812 1275
rect 3496 1272 3534 1274
rect 3774 1272 3812 1274
rect 3844 1308 3882 1310
rect 4122 1308 4160 1310
rect 3844 1307 3911 1308
rect 3844 1275 3847 1307
rect 3879 1275 3911 1307
rect 3844 1274 3911 1275
rect 4093 1307 4160 1308
rect 4093 1275 4125 1307
rect 4157 1275 4160 1307
rect 4093 1274 4160 1275
rect 3844 1272 3882 1274
rect 4122 1272 4160 1274
rect 4192 1308 4230 1310
rect 4470 1308 4508 1310
rect 4192 1307 4259 1308
rect 4192 1275 4195 1307
rect 4227 1275 4259 1307
rect 4192 1274 4259 1275
rect 4441 1307 4508 1308
rect 4441 1275 4473 1307
rect 4505 1275 4508 1307
rect 4441 1274 4508 1275
rect 4192 1272 4230 1274
rect 4470 1272 4508 1274
rect 4540 1308 4578 1310
rect 4818 1308 4856 1310
rect 4540 1307 4607 1308
rect 4540 1275 4543 1307
rect 4575 1275 4607 1307
rect 4540 1274 4607 1275
rect 4789 1307 4856 1308
rect 4789 1275 4821 1307
rect 4853 1275 4856 1307
rect 4789 1274 4856 1275
rect 4540 1272 4578 1274
rect 4818 1272 4856 1274
rect 4888 1308 4926 1310
rect 5166 1308 5204 1310
rect 4888 1307 4955 1308
rect 4888 1275 4891 1307
rect 4923 1275 4955 1307
rect 4888 1274 4955 1275
rect 5137 1307 5204 1308
rect 5137 1275 5169 1307
rect 5201 1275 5204 1307
rect 5137 1274 5204 1275
rect 4888 1272 4926 1274
rect 5166 1272 5204 1274
rect 5236 1308 5274 1310
rect 5514 1308 5552 1310
rect 5236 1307 5303 1308
rect 5236 1275 5239 1307
rect 5271 1275 5303 1307
rect 5236 1274 5303 1275
rect 5485 1307 5552 1308
rect 5485 1275 5517 1307
rect 5549 1275 5552 1307
rect 5485 1274 5552 1275
rect 5236 1272 5274 1274
rect 5514 1272 5552 1274
rect 5584 1308 5622 1310
rect 5862 1308 5900 1310
rect 5584 1307 5651 1308
rect 5584 1275 5587 1307
rect 5619 1275 5651 1307
rect 5584 1274 5651 1275
rect 5833 1307 5900 1308
rect 5833 1275 5865 1307
rect 5897 1275 5900 1307
rect 5833 1274 5900 1275
rect 5584 1272 5622 1274
rect 5862 1272 5900 1274
rect 5932 1308 5970 1310
rect 6210 1308 6248 1310
rect 5932 1307 5999 1308
rect 5932 1275 5935 1307
rect 5967 1275 5999 1307
rect 5932 1274 5999 1275
rect 6181 1307 6248 1308
rect 6181 1275 6213 1307
rect 6245 1275 6248 1307
rect 6181 1274 6248 1275
rect 5932 1272 5970 1274
rect 6210 1272 6248 1274
rect 6280 1308 6318 1310
rect 6558 1308 6596 1310
rect 6280 1307 6347 1308
rect 6280 1275 6283 1307
rect 6315 1275 6347 1307
rect 6280 1274 6347 1275
rect 6529 1307 6596 1308
rect 6529 1275 6561 1307
rect 6593 1275 6596 1307
rect 6529 1274 6596 1275
rect 6280 1272 6318 1274
rect 6558 1272 6596 1274
rect 6628 1308 6666 1310
rect 6906 1308 6944 1310
rect 6628 1307 6695 1308
rect 6628 1275 6631 1307
rect 6663 1275 6695 1307
rect 6628 1274 6695 1275
rect 6877 1307 6944 1308
rect 6877 1275 6909 1307
rect 6941 1275 6944 1307
rect 6877 1274 6944 1275
rect 6628 1272 6666 1274
rect 6906 1272 6944 1274
rect 6976 1308 7014 1310
rect 7254 1308 7292 1310
rect 6976 1307 7043 1308
rect 6976 1275 6979 1307
rect 7011 1275 7043 1307
rect 6976 1274 7043 1275
rect 7225 1307 7292 1308
rect 7225 1275 7257 1307
rect 7289 1275 7292 1307
rect 7225 1274 7292 1275
rect 6976 1272 7014 1274
rect 7254 1272 7292 1274
rect 16 1184 54 1186
rect 294 1184 332 1186
rect 16 1183 83 1184
rect 16 1151 19 1183
rect 51 1151 83 1183
rect 16 1150 83 1151
rect 265 1183 332 1184
rect 265 1151 297 1183
rect 329 1151 332 1183
rect 265 1150 332 1151
rect 16 1148 54 1150
rect 294 1148 332 1150
rect 364 1184 402 1186
rect 642 1184 680 1186
rect 364 1183 431 1184
rect 364 1151 367 1183
rect 399 1151 431 1183
rect 364 1150 431 1151
rect 613 1183 680 1184
rect 613 1151 645 1183
rect 677 1151 680 1183
rect 613 1150 680 1151
rect 364 1148 402 1150
rect 642 1148 680 1150
rect 712 1184 750 1186
rect 990 1184 1028 1186
rect 712 1183 779 1184
rect 712 1151 715 1183
rect 747 1151 779 1183
rect 712 1150 779 1151
rect 961 1183 1028 1184
rect 961 1151 993 1183
rect 1025 1151 1028 1183
rect 961 1150 1028 1151
rect 712 1148 750 1150
rect 990 1148 1028 1150
rect 1060 1184 1098 1186
rect 1338 1184 1376 1186
rect 1060 1183 1127 1184
rect 1060 1151 1063 1183
rect 1095 1151 1127 1183
rect 1060 1150 1127 1151
rect 1309 1183 1376 1184
rect 1309 1151 1341 1183
rect 1373 1151 1376 1183
rect 1309 1150 1376 1151
rect 1060 1148 1098 1150
rect 1338 1148 1376 1150
rect 1408 1184 1446 1186
rect 1686 1184 1724 1186
rect 1408 1183 1475 1184
rect 1408 1151 1411 1183
rect 1443 1151 1475 1183
rect 1408 1150 1475 1151
rect 1657 1183 1724 1184
rect 1657 1151 1689 1183
rect 1721 1151 1724 1183
rect 1657 1150 1724 1151
rect 1408 1148 1446 1150
rect 1686 1148 1724 1150
rect 1756 1184 1794 1186
rect 2034 1184 2072 1186
rect 1756 1183 1823 1184
rect 1756 1151 1759 1183
rect 1791 1151 1823 1183
rect 1756 1150 1823 1151
rect 2005 1183 2072 1184
rect 2005 1151 2037 1183
rect 2069 1151 2072 1183
rect 2005 1150 2072 1151
rect 1756 1148 1794 1150
rect 2034 1148 2072 1150
rect 2104 1184 2142 1186
rect 2382 1184 2420 1186
rect 2104 1183 2171 1184
rect 2104 1151 2107 1183
rect 2139 1151 2171 1183
rect 2104 1150 2171 1151
rect 2353 1183 2420 1184
rect 2353 1151 2385 1183
rect 2417 1151 2420 1183
rect 2353 1150 2420 1151
rect 2104 1148 2142 1150
rect 2382 1148 2420 1150
rect 2452 1184 2490 1186
rect 2730 1184 2768 1186
rect 2452 1183 2519 1184
rect 2452 1151 2455 1183
rect 2487 1151 2519 1183
rect 2452 1150 2519 1151
rect 2701 1183 2768 1184
rect 2701 1151 2733 1183
rect 2765 1151 2768 1183
rect 2701 1150 2768 1151
rect 2452 1148 2490 1150
rect 2730 1148 2768 1150
rect 2800 1184 2838 1186
rect 3078 1184 3116 1186
rect 2800 1183 2867 1184
rect 2800 1151 2803 1183
rect 2835 1151 2867 1183
rect 2800 1150 2867 1151
rect 3049 1183 3116 1184
rect 3049 1151 3081 1183
rect 3113 1151 3116 1183
rect 3049 1150 3116 1151
rect 2800 1148 2838 1150
rect 3078 1148 3116 1150
rect 3148 1184 3186 1186
rect 3426 1184 3464 1186
rect 3148 1183 3215 1184
rect 3148 1151 3151 1183
rect 3183 1151 3215 1183
rect 3148 1150 3215 1151
rect 3397 1183 3464 1184
rect 3397 1151 3429 1183
rect 3461 1151 3464 1183
rect 3397 1150 3464 1151
rect 3148 1148 3186 1150
rect 3426 1148 3464 1150
rect 3496 1184 3534 1186
rect 3774 1184 3812 1186
rect 3496 1183 3563 1184
rect 3496 1151 3499 1183
rect 3531 1151 3563 1183
rect 3496 1150 3563 1151
rect 3745 1183 3812 1184
rect 3745 1151 3777 1183
rect 3809 1151 3812 1183
rect 3745 1150 3812 1151
rect 3496 1148 3534 1150
rect 3774 1148 3812 1150
rect 3844 1184 3882 1186
rect 4122 1184 4160 1186
rect 3844 1183 3911 1184
rect 3844 1151 3847 1183
rect 3879 1151 3911 1183
rect 3844 1150 3911 1151
rect 4093 1183 4160 1184
rect 4093 1151 4125 1183
rect 4157 1151 4160 1183
rect 4093 1150 4160 1151
rect 3844 1148 3882 1150
rect 4122 1148 4160 1150
rect 4192 1184 4230 1186
rect 4470 1184 4508 1186
rect 4192 1183 4259 1184
rect 4192 1151 4195 1183
rect 4227 1151 4259 1183
rect 4192 1150 4259 1151
rect 4441 1183 4508 1184
rect 4441 1151 4473 1183
rect 4505 1151 4508 1183
rect 4441 1150 4508 1151
rect 4192 1148 4230 1150
rect 4470 1148 4508 1150
rect 4540 1184 4578 1186
rect 4818 1184 4856 1186
rect 4540 1183 4607 1184
rect 4540 1151 4543 1183
rect 4575 1151 4607 1183
rect 4540 1150 4607 1151
rect 4789 1183 4856 1184
rect 4789 1151 4821 1183
rect 4853 1151 4856 1183
rect 4789 1150 4856 1151
rect 4540 1148 4578 1150
rect 4818 1148 4856 1150
rect 4888 1184 4926 1186
rect 5166 1184 5204 1186
rect 4888 1183 4955 1184
rect 4888 1151 4891 1183
rect 4923 1151 4955 1183
rect 4888 1150 4955 1151
rect 5137 1183 5204 1184
rect 5137 1151 5169 1183
rect 5201 1151 5204 1183
rect 5137 1150 5204 1151
rect 4888 1148 4926 1150
rect 5166 1148 5204 1150
rect 5236 1184 5274 1186
rect 5514 1184 5552 1186
rect 5236 1183 5303 1184
rect 5236 1151 5239 1183
rect 5271 1151 5303 1183
rect 5236 1150 5303 1151
rect 5485 1183 5552 1184
rect 5485 1151 5517 1183
rect 5549 1151 5552 1183
rect 5485 1150 5552 1151
rect 5236 1148 5274 1150
rect 5514 1148 5552 1150
rect 5584 1184 5622 1186
rect 5862 1184 5900 1186
rect 5584 1183 5651 1184
rect 5584 1151 5587 1183
rect 5619 1151 5651 1183
rect 5584 1150 5651 1151
rect 5833 1183 5900 1184
rect 5833 1151 5865 1183
rect 5897 1151 5900 1183
rect 5833 1150 5900 1151
rect 5584 1148 5622 1150
rect 5862 1148 5900 1150
rect 5932 1184 5970 1186
rect 6210 1184 6248 1186
rect 5932 1183 5999 1184
rect 5932 1151 5935 1183
rect 5967 1151 5999 1183
rect 5932 1150 5999 1151
rect 6181 1183 6248 1184
rect 6181 1151 6213 1183
rect 6245 1151 6248 1183
rect 6181 1150 6248 1151
rect 5932 1148 5970 1150
rect 6210 1148 6248 1150
rect 6280 1184 6318 1186
rect 6558 1184 6596 1186
rect 6280 1183 6347 1184
rect 6280 1151 6283 1183
rect 6315 1151 6347 1183
rect 6280 1150 6347 1151
rect 6529 1183 6596 1184
rect 6529 1151 6561 1183
rect 6593 1151 6596 1183
rect 6529 1150 6596 1151
rect 6280 1148 6318 1150
rect 6558 1148 6596 1150
rect 6628 1184 6666 1186
rect 6906 1184 6944 1186
rect 6628 1183 6695 1184
rect 6628 1151 6631 1183
rect 6663 1151 6695 1183
rect 6628 1150 6695 1151
rect 6877 1183 6944 1184
rect 6877 1151 6909 1183
rect 6941 1151 6944 1183
rect 6877 1150 6944 1151
rect 6628 1148 6666 1150
rect 6906 1148 6944 1150
rect 6976 1184 7014 1186
rect 7254 1184 7292 1186
rect 6976 1183 7043 1184
rect 6976 1151 6979 1183
rect 7011 1151 7043 1183
rect 6976 1150 7043 1151
rect 7225 1183 7292 1184
rect 7225 1151 7257 1183
rect 7289 1151 7292 1183
rect 7225 1150 7292 1151
rect 6976 1148 7014 1150
rect 7254 1148 7292 1150
rect 16 1114 54 1116
rect 294 1114 332 1116
rect 16 1113 83 1114
rect 16 1081 19 1113
rect 51 1081 83 1113
rect 16 1080 83 1081
rect 265 1113 332 1114
rect 265 1081 297 1113
rect 329 1081 332 1113
rect 265 1080 332 1081
rect 16 1078 54 1080
rect 294 1078 332 1080
rect 364 1114 402 1116
rect 642 1114 680 1116
rect 364 1113 431 1114
rect 364 1081 367 1113
rect 399 1081 431 1113
rect 364 1080 431 1081
rect 613 1113 680 1114
rect 613 1081 645 1113
rect 677 1081 680 1113
rect 613 1080 680 1081
rect 364 1078 402 1080
rect 642 1078 680 1080
rect 712 1114 750 1116
rect 990 1114 1028 1116
rect 712 1113 779 1114
rect 712 1081 715 1113
rect 747 1081 779 1113
rect 712 1080 779 1081
rect 961 1113 1028 1114
rect 961 1081 993 1113
rect 1025 1081 1028 1113
rect 961 1080 1028 1081
rect 712 1078 750 1080
rect 990 1078 1028 1080
rect 1060 1114 1098 1116
rect 1338 1114 1376 1116
rect 1060 1113 1127 1114
rect 1060 1081 1063 1113
rect 1095 1081 1127 1113
rect 1060 1080 1127 1081
rect 1309 1113 1376 1114
rect 1309 1081 1341 1113
rect 1373 1081 1376 1113
rect 1309 1080 1376 1081
rect 1060 1078 1098 1080
rect 1338 1078 1376 1080
rect 1408 1114 1446 1116
rect 1686 1114 1724 1116
rect 1408 1113 1475 1114
rect 1408 1081 1411 1113
rect 1443 1081 1475 1113
rect 1408 1080 1475 1081
rect 1657 1113 1724 1114
rect 1657 1081 1689 1113
rect 1721 1081 1724 1113
rect 1657 1080 1724 1081
rect 1408 1078 1446 1080
rect 1686 1078 1724 1080
rect 1756 1114 1794 1116
rect 2034 1114 2072 1116
rect 1756 1113 1823 1114
rect 1756 1081 1759 1113
rect 1791 1081 1823 1113
rect 1756 1080 1823 1081
rect 2005 1113 2072 1114
rect 2005 1081 2037 1113
rect 2069 1081 2072 1113
rect 2005 1080 2072 1081
rect 1756 1078 1794 1080
rect 2034 1078 2072 1080
rect 2104 1114 2142 1116
rect 2382 1114 2420 1116
rect 2104 1113 2171 1114
rect 2104 1081 2107 1113
rect 2139 1081 2171 1113
rect 2104 1080 2171 1081
rect 2353 1113 2420 1114
rect 2353 1081 2385 1113
rect 2417 1081 2420 1113
rect 2353 1080 2420 1081
rect 2104 1078 2142 1080
rect 2382 1078 2420 1080
rect 2452 1114 2490 1116
rect 2730 1114 2768 1116
rect 2452 1113 2519 1114
rect 2452 1081 2455 1113
rect 2487 1081 2519 1113
rect 2452 1080 2519 1081
rect 2701 1113 2768 1114
rect 2701 1081 2733 1113
rect 2765 1081 2768 1113
rect 2701 1080 2768 1081
rect 2452 1078 2490 1080
rect 2730 1078 2768 1080
rect 2800 1114 2838 1116
rect 3078 1114 3116 1116
rect 2800 1113 2867 1114
rect 2800 1081 2803 1113
rect 2835 1081 2867 1113
rect 2800 1080 2867 1081
rect 3049 1113 3116 1114
rect 3049 1081 3081 1113
rect 3113 1081 3116 1113
rect 3049 1080 3116 1081
rect 2800 1078 2838 1080
rect 3078 1078 3116 1080
rect 3148 1114 3186 1116
rect 3426 1114 3464 1116
rect 3148 1113 3215 1114
rect 3148 1081 3151 1113
rect 3183 1081 3215 1113
rect 3148 1080 3215 1081
rect 3397 1113 3464 1114
rect 3397 1081 3429 1113
rect 3461 1081 3464 1113
rect 3397 1080 3464 1081
rect 3148 1078 3186 1080
rect 3426 1078 3464 1080
rect 3496 1114 3534 1116
rect 3774 1114 3812 1116
rect 3496 1113 3563 1114
rect 3496 1081 3499 1113
rect 3531 1081 3563 1113
rect 3496 1080 3563 1081
rect 3745 1113 3812 1114
rect 3745 1081 3777 1113
rect 3809 1081 3812 1113
rect 3745 1080 3812 1081
rect 3496 1078 3534 1080
rect 3774 1078 3812 1080
rect 3844 1114 3882 1116
rect 4122 1114 4160 1116
rect 3844 1113 3911 1114
rect 3844 1081 3847 1113
rect 3879 1081 3911 1113
rect 3844 1080 3911 1081
rect 4093 1113 4160 1114
rect 4093 1081 4125 1113
rect 4157 1081 4160 1113
rect 4093 1080 4160 1081
rect 3844 1078 3882 1080
rect 4122 1078 4160 1080
rect 4192 1114 4230 1116
rect 4470 1114 4508 1116
rect 4192 1113 4259 1114
rect 4192 1081 4195 1113
rect 4227 1081 4259 1113
rect 4192 1080 4259 1081
rect 4441 1113 4508 1114
rect 4441 1081 4473 1113
rect 4505 1081 4508 1113
rect 4441 1080 4508 1081
rect 4192 1078 4230 1080
rect 4470 1078 4508 1080
rect 4540 1114 4578 1116
rect 4818 1114 4856 1116
rect 4540 1113 4607 1114
rect 4540 1081 4543 1113
rect 4575 1081 4607 1113
rect 4540 1080 4607 1081
rect 4789 1113 4856 1114
rect 4789 1081 4821 1113
rect 4853 1081 4856 1113
rect 4789 1080 4856 1081
rect 4540 1078 4578 1080
rect 4818 1078 4856 1080
rect 4888 1114 4926 1116
rect 5166 1114 5204 1116
rect 4888 1113 4955 1114
rect 4888 1081 4891 1113
rect 4923 1081 4955 1113
rect 4888 1080 4955 1081
rect 5137 1113 5204 1114
rect 5137 1081 5169 1113
rect 5201 1081 5204 1113
rect 5137 1080 5204 1081
rect 4888 1078 4926 1080
rect 5166 1078 5204 1080
rect 5236 1114 5274 1116
rect 5514 1114 5552 1116
rect 5236 1113 5303 1114
rect 5236 1081 5239 1113
rect 5271 1081 5303 1113
rect 5236 1080 5303 1081
rect 5485 1113 5552 1114
rect 5485 1081 5517 1113
rect 5549 1081 5552 1113
rect 5485 1080 5552 1081
rect 5236 1078 5274 1080
rect 5514 1078 5552 1080
rect 5584 1114 5622 1116
rect 5862 1114 5900 1116
rect 5584 1113 5651 1114
rect 5584 1081 5587 1113
rect 5619 1081 5651 1113
rect 5584 1080 5651 1081
rect 5833 1113 5900 1114
rect 5833 1081 5865 1113
rect 5897 1081 5900 1113
rect 5833 1080 5900 1081
rect 5584 1078 5622 1080
rect 5862 1078 5900 1080
rect 5932 1114 5970 1116
rect 6210 1114 6248 1116
rect 5932 1113 5999 1114
rect 5932 1081 5935 1113
rect 5967 1081 5999 1113
rect 5932 1080 5999 1081
rect 6181 1113 6248 1114
rect 6181 1081 6213 1113
rect 6245 1081 6248 1113
rect 6181 1080 6248 1081
rect 5932 1078 5970 1080
rect 6210 1078 6248 1080
rect 6280 1114 6318 1116
rect 6558 1114 6596 1116
rect 6280 1113 6347 1114
rect 6280 1081 6283 1113
rect 6315 1081 6347 1113
rect 6280 1080 6347 1081
rect 6529 1113 6596 1114
rect 6529 1081 6561 1113
rect 6593 1081 6596 1113
rect 6529 1080 6596 1081
rect 6280 1078 6318 1080
rect 6558 1078 6596 1080
rect 6628 1114 6666 1116
rect 6906 1114 6944 1116
rect 6628 1113 6695 1114
rect 6628 1081 6631 1113
rect 6663 1081 6695 1113
rect 6628 1080 6695 1081
rect 6877 1113 6944 1114
rect 6877 1081 6909 1113
rect 6941 1081 6944 1113
rect 6877 1080 6944 1081
rect 6628 1078 6666 1080
rect 6906 1078 6944 1080
rect 6976 1114 7014 1116
rect 7254 1114 7292 1116
rect 6976 1113 7043 1114
rect 6976 1081 6979 1113
rect 7011 1081 7043 1113
rect 6976 1080 7043 1081
rect 7225 1113 7292 1114
rect 7225 1081 7257 1113
rect 7289 1081 7292 1113
rect 7225 1080 7292 1081
rect 6976 1078 7014 1080
rect 7254 1078 7292 1080
rect 16 990 54 992
rect 294 990 332 992
rect 16 989 83 990
rect 16 957 19 989
rect 51 957 83 989
rect 16 956 83 957
rect 265 989 332 990
rect 265 957 297 989
rect 329 957 332 989
rect 265 956 332 957
rect 16 954 54 956
rect 294 954 332 956
rect 364 990 402 992
rect 642 990 680 992
rect 364 989 431 990
rect 364 957 367 989
rect 399 957 431 989
rect 364 956 431 957
rect 613 989 680 990
rect 613 957 645 989
rect 677 957 680 989
rect 613 956 680 957
rect 364 954 402 956
rect 642 954 680 956
rect 712 990 750 992
rect 990 990 1028 992
rect 712 989 779 990
rect 712 957 715 989
rect 747 957 779 989
rect 712 956 779 957
rect 961 989 1028 990
rect 961 957 993 989
rect 1025 957 1028 989
rect 961 956 1028 957
rect 712 954 750 956
rect 990 954 1028 956
rect 1060 990 1098 992
rect 1338 990 1376 992
rect 1060 989 1127 990
rect 1060 957 1063 989
rect 1095 957 1127 989
rect 1060 956 1127 957
rect 1309 989 1376 990
rect 1309 957 1341 989
rect 1373 957 1376 989
rect 1309 956 1376 957
rect 1060 954 1098 956
rect 1338 954 1376 956
rect 1408 990 1446 992
rect 1686 990 1724 992
rect 1408 989 1475 990
rect 1408 957 1411 989
rect 1443 957 1475 989
rect 1408 956 1475 957
rect 1657 989 1724 990
rect 1657 957 1689 989
rect 1721 957 1724 989
rect 1657 956 1724 957
rect 1408 954 1446 956
rect 1686 954 1724 956
rect 1756 990 1794 992
rect 2034 990 2072 992
rect 1756 989 1823 990
rect 1756 957 1759 989
rect 1791 957 1823 989
rect 1756 956 1823 957
rect 2005 989 2072 990
rect 2005 957 2037 989
rect 2069 957 2072 989
rect 2005 956 2072 957
rect 1756 954 1794 956
rect 2034 954 2072 956
rect 2104 990 2142 992
rect 2382 990 2420 992
rect 2104 989 2171 990
rect 2104 957 2107 989
rect 2139 957 2171 989
rect 2104 956 2171 957
rect 2353 989 2420 990
rect 2353 957 2385 989
rect 2417 957 2420 989
rect 2353 956 2420 957
rect 2104 954 2142 956
rect 2382 954 2420 956
rect 2452 990 2490 992
rect 2730 990 2768 992
rect 2452 989 2519 990
rect 2452 957 2455 989
rect 2487 957 2519 989
rect 2452 956 2519 957
rect 2701 989 2768 990
rect 2701 957 2733 989
rect 2765 957 2768 989
rect 2701 956 2768 957
rect 2452 954 2490 956
rect 2730 954 2768 956
rect 2800 990 2838 992
rect 3078 990 3116 992
rect 2800 989 2867 990
rect 2800 957 2803 989
rect 2835 957 2867 989
rect 2800 956 2867 957
rect 3049 989 3116 990
rect 3049 957 3081 989
rect 3113 957 3116 989
rect 3049 956 3116 957
rect 2800 954 2838 956
rect 3078 954 3116 956
rect 3148 990 3186 992
rect 3426 990 3464 992
rect 3148 989 3215 990
rect 3148 957 3151 989
rect 3183 957 3215 989
rect 3148 956 3215 957
rect 3397 989 3464 990
rect 3397 957 3429 989
rect 3461 957 3464 989
rect 3397 956 3464 957
rect 3148 954 3186 956
rect 3426 954 3464 956
rect 3496 990 3534 992
rect 3774 990 3812 992
rect 3496 989 3563 990
rect 3496 957 3499 989
rect 3531 957 3563 989
rect 3496 956 3563 957
rect 3745 989 3812 990
rect 3745 957 3777 989
rect 3809 957 3812 989
rect 3745 956 3812 957
rect 3496 954 3534 956
rect 3774 954 3812 956
rect 3844 990 3882 992
rect 4122 990 4160 992
rect 3844 989 3911 990
rect 3844 957 3847 989
rect 3879 957 3911 989
rect 3844 956 3911 957
rect 4093 989 4160 990
rect 4093 957 4125 989
rect 4157 957 4160 989
rect 4093 956 4160 957
rect 3844 954 3882 956
rect 4122 954 4160 956
rect 4192 990 4230 992
rect 4470 990 4508 992
rect 4192 989 4259 990
rect 4192 957 4195 989
rect 4227 957 4259 989
rect 4192 956 4259 957
rect 4441 989 4508 990
rect 4441 957 4473 989
rect 4505 957 4508 989
rect 4441 956 4508 957
rect 4192 954 4230 956
rect 4470 954 4508 956
rect 4540 990 4578 992
rect 4818 990 4856 992
rect 4540 989 4607 990
rect 4540 957 4543 989
rect 4575 957 4607 989
rect 4540 956 4607 957
rect 4789 989 4856 990
rect 4789 957 4821 989
rect 4853 957 4856 989
rect 4789 956 4856 957
rect 4540 954 4578 956
rect 4818 954 4856 956
rect 4888 990 4926 992
rect 5166 990 5204 992
rect 4888 989 4955 990
rect 4888 957 4891 989
rect 4923 957 4955 989
rect 4888 956 4955 957
rect 5137 989 5204 990
rect 5137 957 5169 989
rect 5201 957 5204 989
rect 5137 956 5204 957
rect 4888 954 4926 956
rect 5166 954 5204 956
rect 5236 990 5274 992
rect 5514 990 5552 992
rect 5236 989 5303 990
rect 5236 957 5239 989
rect 5271 957 5303 989
rect 5236 956 5303 957
rect 5485 989 5552 990
rect 5485 957 5517 989
rect 5549 957 5552 989
rect 5485 956 5552 957
rect 5236 954 5274 956
rect 5514 954 5552 956
rect 5584 990 5622 992
rect 5862 990 5900 992
rect 5584 989 5651 990
rect 5584 957 5587 989
rect 5619 957 5651 989
rect 5584 956 5651 957
rect 5833 989 5900 990
rect 5833 957 5865 989
rect 5897 957 5900 989
rect 5833 956 5900 957
rect 5584 954 5622 956
rect 5862 954 5900 956
rect 5932 990 5970 992
rect 6210 990 6248 992
rect 5932 989 5999 990
rect 5932 957 5935 989
rect 5967 957 5999 989
rect 5932 956 5999 957
rect 6181 989 6248 990
rect 6181 957 6213 989
rect 6245 957 6248 989
rect 6181 956 6248 957
rect 5932 954 5970 956
rect 6210 954 6248 956
rect 6280 990 6318 992
rect 6558 990 6596 992
rect 6280 989 6347 990
rect 6280 957 6283 989
rect 6315 957 6347 989
rect 6280 956 6347 957
rect 6529 989 6596 990
rect 6529 957 6561 989
rect 6593 957 6596 989
rect 6529 956 6596 957
rect 6280 954 6318 956
rect 6558 954 6596 956
rect 6628 990 6666 992
rect 6906 990 6944 992
rect 6628 989 6695 990
rect 6628 957 6631 989
rect 6663 957 6695 989
rect 6628 956 6695 957
rect 6877 989 6944 990
rect 6877 957 6909 989
rect 6941 957 6944 989
rect 6877 956 6944 957
rect 6628 954 6666 956
rect 6906 954 6944 956
rect 6976 990 7014 992
rect 7254 990 7292 992
rect 6976 989 7043 990
rect 6976 957 6979 989
rect 7011 957 7043 989
rect 6976 956 7043 957
rect 7225 989 7292 990
rect 7225 957 7257 989
rect 7289 957 7292 989
rect 7225 956 7292 957
rect 6976 954 7014 956
rect 7254 954 7292 956
rect 16 866 54 868
rect 294 866 332 868
rect 16 865 83 866
rect 16 833 19 865
rect 51 833 83 865
rect 16 832 83 833
rect 265 865 332 866
rect 265 833 297 865
rect 329 833 332 865
rect 265 832 332 833
rect 16 830 54 832
rect 294 830 332 832
rect 364 866 402 868
rect 642 866 680 868
rect 364 865 431 866
rect 364 833 367 865
rect 399 833 431 865
rect 364 832 431 833
rect 613 865 680 866
rect 613 833 645 865
rect 677 833 680 865
rect 613 832 680 833
rect 364 830 402 832
rect 642 830 680 832
rect 712 866 750 868
rect 990 866 1028 868
rect 712 865 779 866
rect 712 833 715 865
rect 747 833 779 865
rect 712 832 779 833
rect 961 865 1028 866
rect 961 833 993 865
rect 1025 833 1028 865
rect 961 832 1028 833
rect 712 830 750 832
rect 990 830 1028 832
rect 1060 866 1098 868
rect 1338 866 1376 868
rect 1060 865 1127 866
rect 1060 833 1063 865
rect 1095 833 1127 865
rect 1060 832 1127 833
rect 1309 865 1376 866
rect 1309 833 1341 865
rect 1373 833 1376 865
rect 1309 832 1376 833
rect 1060 830 1098 832
rect 1338 830 1376 832
rect 1408 866 1446 868
rect 1686 866 1724 868
rect 1408 865 1475 866
rect 1408 833 1411 865
rect 1443 833 1475 865
rect 1408 832 1475 833
rect 1657 865 1724 866
rect 1657 833 1689 865
rect 1721 833 1724 865
rect 1657 832 1724 833
rect 1408 830 1446 832
rect 1686 830 1724 832
rect 1756 866 1794 868
rect 2034 866 2072 868
rect 1756 865 1823 866
rect 1756 833 1759 865
rect 1791 833 1823 865
rect 1756 832 1823 833
rect 2005 865 2072 866
rect 2005 833 2037 865
rect 2069 833 2072 865
rect 2005 832 2072 833
rect 1756 830 1794 832
rect 2034 830 2072 832
rect 2104 866 2142 868
rect 2382 866 2420 868
rect 2104 865 2171 866
rect 2104 833 2107 865
rect 2139 833 2171 865
rect 2104 832 2171 833
rect 2353 865 2420 866
rect 2353 833 2385 865
rect 2417 833 2420 865
rect 2353 832 2420 833
rect 2104 830 2142 832
rect 2382 830 2420 832
rect 2452 866 2490 868
rect 2730 866 2768 868
rect 2452 865 2519 866
rect 2452 833 2455 865
rect 2487 833 2519 865
rect 2452 832 2519 833
rect 2701 865 2768 866
rect 2701 833 2733 865
rect 2765 833 2768 865
rect 2701 832 2768 833
rect 2452 830 2490 832
rect 2730 830 2768 832
rect 2800 866 2838 868
rect 3078 866 3116 868
rect 2800 865 2867 866
rect 2800 833 2803 865
rect 2835 833 2867 865
rect 2800 832 2867 833
rect 3049 865 3116 866
rect 3049 833 3081 865
rect 3113 833 3116 865
rect 3049 832 3116 833
rect 2800 830 2838 832
rect 3078 830 3116 832
rect 3148 866 3186 868
rect 3426 866 3464 868
rect 3148 865 3215 866
rect 3148 833 3151 865
rect 3183 833 3215 865
rect 3148 832 3215 833
rect 3397 865 3464 866
rect 3397 833 3429 865
rect 3461 833 3464 865
rect 3397 832 3464 833
rect 3148 830 3186 832
rect 3426 830 3464 832
rect 3496 866 3534 868
rect 3774 866 3812 868
rect 3496 865 3563 866
rect 3496 833 3499 865
rect 3531 833 3563 865
rect 3496 832 3563 833
rect 3745 865 3812 866
rect 3745 833 3777 865
rect 3809 833 3812 865
rect 3745 832 3812 833
rect 3496 830 3534 832
rect 3774 830 3812 832
rect 3844 866 3882 868
rect 4122 866 4160 868
rect 3844 865 3911 866
rect 3844 833 3847 865
rect 3879 833 3911 865
rect 3844 832 3911 833
rect 4093 865 4160 866
rect 4093 833 4125 865
rect 4157 833 4160 865
rect 4093 832 4160 833
rect 3844 830 3882 832
rect 4122 830 4160 832
rect 4192 866 4230 868
rect 4470 866 4508 868
rect 4192 865 4259 866
rect 4192 833 4195 865
rect 4227 833 4259 865
rect 4192 832 4259 833
rect 4441 865 4508 866
rect 4441 833 4473 865
rect 4505 833 4508 865
rect 4441 832 4508 833
rect 4192 830 4230 832
rect 4470 830 4508 832
rect 4540 866 4578 868
rect 4818 866 4856 868
rect 4540 865 4607 866
rect 4540 833 4543 865
rect 4575 833 4607 865
rect 4540 832 4607 833
rect 4789 865 4856 866
rect 4789 833 4821 865
rect 4853 833 4856 865
rect 4789 832 4856 833
rect 4540 830 4578 832
rect 4818 830 4856 832
rect 4888 866 4926 868
rect 5166 866 5204 868
rect 4888 865 4955 866
rect 4888 833 4891 865
rect 4923 833 4955 865
rect 4888 832 4955 833
rect 5137 865 5204 866
rect 5137 833 5169 865
rect 5201 833 5204 865
rect 5137 832 5204 833
rect 4888 830 4926 832
rect 5166 830 5204 832
rect 5236 866 5274 868
rect 5514 866 5552 868
rect 5236 865 5303 866
rect 5236 833 5239 865
rect 5271 833 5303 865
rect 5236 832 5303 833
rect 5485 865 5552 866
rect 5485 833 5517 865
rect 5549 833 5552 865
rect 5485 832 5552 833
rect 5236 830 5274 832
rect 5514 830 5552 832
rect 5584 866 5622 868
rect 5862 866 5900 868
rect 5584 865 5651 866
rect 5584 833 5587 865
rect 5619 833 5651 865
rect 5584 832 5651 833
rect 5833 865 5900 866
rect 5833 833 5865 865
rect 5897 833 5900 865
rect 5833 832 5900 833
rect 5584 830 5622 832
rect 5862 830 5900 832
rect 5932 866 5970 868
rect 6210 866 6248 868
rect 5932 865 5999 866
rect 5932 833 5935 865
rect 5967 833 5999 865
rect 5932 832 5999 833
rect 6181 865 6248 866
rect 6181 833 6213 865
rect 6245 833 6248 865
rect 6181 832 6248 833
rect 5932 830 5970 832
rect 6210 830 6248 832
rect 6280 866 6318 868
rect 6558 866 6596 868
rect 6280 865 6347 866
rect 6280 833 6283 865
rect 6315 833 6347 865
rect 6280 832 6347 833
rect 6529 865 6596 866
rect 6529 833 6561 865
rect 6593 833 6596 865
rect 6529 832 6596 833
rect 6280 830 6318 832
rect 6558 830 6596 832
rect 6628 866 6666 868
rect 6906 866 6944 868
rect 6628 865 6695 866
rect 6628 833 6631 865
rect 6663 833 6695 865
rect 6628 832 6695 833
rect 6877 865 6944 866
rect 6877 833 6909 865
rect 6941 833 6944 865
rect 6877 832 6944 833
rect 6628 830 6666 832
rect 6906 830 6944 832
rect 6976 866 7014 868
rect 7254 866 7292 868
rect 6976 865 7043 866
rect 6976 833 6979 865
rect 7011 833 7043 865
rect 6976 832 7043 833
rect 7225 865 7292 866
rect 7225 833 7257 865
rect 7289 833 7292 865
rect 7225 832 7292 833
rect 6976 830 7014 832
rect 7254 830 7292 832
rect 16 742 54 744
rect 294 742 332 744
rect 16 741 83 742
rect 16 709 19 741
rect 51 709 83 741
rect 16 708 83 709
rect 265 741 332 742
rect 265 709 297 741
rect 329 709 332 741
rect 265 708 332 709
rect 16 706 54 708
rect 294 706 332 708
rect 364 742 402 744
rect 642 742 680 744
rect 364 741 431 742
rect 364 709 367 741
rect 399 709 431 741
rect 364 708 431 709
rect 613 741 680 742
rect 613 709 645 741
rect 677 709 680 741
rect 613 708 680 709
rect 364 706 402 708
rect 642 706 680 708
rect 712 742 750 744
rect 990 742 1028 744
rect 712 741 779 742
rect 712 709 715 741
rect 747 709 779 741
rect 712 708 779 709
rect 961 741 1028 742
rect 961 709 993 741
rect 1025 709 1028 741
rect 961 708 1028 709
rect 712 706 750 708
rect 990 706 1028 708
rect 1060 742 1098 744
rect 1338 742 1376 744
rect 1060 741 1127 742
rect 1060 709 1063 741
rect 1095 709 1127 741
rect 1060 708 1127 709
rect 1309 741 1376 742
rect 1309 709 1341 741
rect 1373 709 1376 741
rect 1309 708 1376 709
rect 1060 706 1098 708
rect 1338 706 1376 708
rect 1408 742 1446 744
rect 1686 742 1724 744
rect 1408 741 1475 742
rect 1408 709 1411 741
rect 1443 709 1475 741
rect 1408 708 1475 709
rect 1657 741 1724 742
rect 1657 709 1689 741
rect 1721 709 1724 741
rect 1657 708 1724 709
rect 1408 706 1446 708
rect 1686 706 1724 708
rect 1756 742 1794 744
rect 2034 742 2072 744
rect 1756 741 1823 742
rect 1756 709 1759 741
rect 1791 709 1823 741
rect 1756 708 1823 709
rect 2005 741 2072 742
rect 2005 709 2037 741
rect 2069 709 2072 741
rect 2005 708 2072 709
rect 1756 706 1794 708
rect 2034 706 2072 708
rect 2104 742 2142 744
rect 2382 742 2420 744
rect 2104 741 2171 742
rect 2104 709 2107 741
rect 2139 709 2171 741
rect 2104 708 2171 709
rect 2353 741 2420 742
rect 2353 709 2385 741
rect 2417 709 2420 741
rect 2353 708 2420 709
rect 2104 706 2142 708
rect 2382 706 2420 708
rect 2452 742 2490 744
rect 2730 742 2768 744
rect 2452 741 2519 742
rect 2452 709 2455 741
rect 2487 709 2519 741
rect 2452 708 2519 709
rect 2701 741 2768 742
rect 2701 709 2733 741
rect 2765 709 2768 741
rect 2701 708 2768 709
rect 2452 706 2490 708
rect 2730 706 2768 708
rect 2800 742 2838 744
rect 3078 742 3116 744
rect 2800 741 2867 742
rect 2800 709 2803 741
rect 2835 709 2867 741
rect 2800 708 2867 709
rect 3049 741 3116 742
rect 3049 709 3081 741
rect 3113 709 3116 741
rect 3049 708 3116 709
rect 2800 706 2838 708
rect 3078 706 3116 708
rect 3148 742 3186 744
rect 3426 742 3464 744
rect 3148 741 3215 742
rect 3148 709 3151 741
rect 3183 709 3215 741
rect 3148 708 3215 709
rect 3397 741 3464 742
rect 3397 709 3429 741
rect 3461 709 3464 741
rect 3397 708 3464 709
rect 3148 706 3186 708
rect 3426 706 3464 708
rect 3496 742 3534 744
rect 3774 742 3812 744
rect 3496 741 3563 742
rect 3496 709 3499 741
rect 3531 709 3563 741
rect 3496 708 3563 709
rect 3745 741 3812 742
rect 3745 709 3777 741
rect 3809 709 3812 741
rect 3745 708 3812 709
rect 3496 706 3534 708
rect 3774 706 3812 708
rect 3844 742 3882 744
rect 4122 742 4160 744
rect 3844 741 3911 742
rect 3844 709 3847 741
rect 3879 709 3911 741
rect 3844 708 3911 709
rect 4093 741 4160 742
rect 4093 709 4125 741
rect 4157 709 4160 741
rect 4093 708 4160 709
rect 3844 706 3882 708
rect 4122 706 4160 708
rect 4192 742 4230 744
rect 4470 742 4508 744
rect 4192 741 4259 742
rect 4192 709 4195 741
rect 4227 709 4259 741
rect 4192 708 4259 709
rect 4441 741 4508 742
rect 4441 709 4473 741
rect 4505 709 4508 741
rect 4441 708 4508 709
rect 4192 706 4230 708
rect 4470 706 4508 708
rect 4540 742 4578 744
rect 4818 742 4856 744
rect 4540 741 4607 742
rect 4540 709 4543 741
rect 4575 709 4607 741
rect 4540 708 4607 709
rect 4789 741 4856 742
rect 4789 709 4821 741
rect 4853 709 4856 741
rect 4789 708 4856 709
rect 4540 706 4578 708
rect 4818 706 4856 708
rect 4888 742 4926 744
rect 5166 742 5204 744
rect 4888 741 4955 742
rect 4888 709 4891 741
rect 4923 709 4955 741
rect 4888 708 4955 709
rect 5137 741 5204 742
rect 5137 709 5169 741
rect 5201 709 5204 741
rect 5137 708 5204 709
rect 4888 706 4926 708
rect 5166 706 5204 708
rect 5236 742 5274 744
rect 5514 742 5552 744
rect 5236 741 5303 742
rect 5236 709 5239 741
rect 5271 709 5303 741
rect 5236 708 5303 709
rect 5485 741 5552 742
rect 5485 709 5517 741
rect 5549 709 5552 741
rect 5485 708 5552 709
rect 5236 706 5274 708
rect 5514 706 5552 708
rect 5584 742 5622 744
rect 5862 742 5900 744
rect 5584 741 5651 742
rect 5584 709 5587 741
rect 5619 709 5651 741
rect 5584 708 5651 709
rect 5833 741 5900 742
rect 5833 709 5865 741
rect 5897 709 5900 741
rect 5833 708 5900 709
rect 5584 706 5622 708
rect 5862 706 5900 708
rect 5932 742 5970 744
rect 6210 742 6248 744
rect 5932 741 5999 742
rect 5932 709 5935 741
rect 5967 709 5999 741
rect 5932 708 5999 709
rect 6181 741 6248 742
rect 6181 709 6213 741
rect 6245 709 6248 741
rect 6181 708 6248 709
rect 5932 706 5970 708
rect 6210 706 6248 708
rect 6280 742 6318 744
rect 6558 742 6596 744
rect 6280 741 6347 742
rect 6280 709 6283 741
rect 6315 709 6347 741
rect 6280 708 6347 709
rect 6529 741 6596 742
rect 6529 709 6561 741
rect 6593 709 6596 741
rect 6529 708 6596 709
rect 6280 706 6318 708
rect 6558 706 6596 708
rect 6628 742 6666 744
rect 6906 742 6944 744
rect 6628 741 6695 742
rect 6628 709 6631 741
rect 6663 709 6695 741
rect 6628 708 6695 709
rect 6877 741 6944 742
rect 6877 709 6909 741
rect 6941 709 6944 741
rect 6877 708 6944 709
rect 6628 706 6666 708
rect 6906 706 6944 708
rect 6976 742 7014 744
rect 7254 742 7292 744
rect 6976 741 7043 742
rect 6976 709 6979 741
rect 7011 709 7043 741
rect 6976 708 7043 709
rect 7225 741 7292 742
rect 7225 709 7257 741
rect 7289 709 7292 741
rect 7225 708 7292 709
rect 6976 706 7014 708
rect 7254 706 7292 708
rect 16 618 54 620
rect 294 618 332 620
rect 16 617 83 618
rect 16 585 19 617
rect 51 585 83 617
rect 16 584 83 585
rect 265 617 332 618
rect 265 585 297 617
rect 329 585 332 617
rect 265 584 332 585
rect 16 582 54 584
rect 294 582 332 584
rect 364 618 402 620
rect 642 618 680 620
rect 364 617 431 618
rect 364 585 367 617
rect 399 585 431 617
rect 364 584 431 585
rect 613 617 680 618
rect 613 585 645 617
rect 677 585 680 617
rect 613 584 680 585
rect 364 582 402 584
rect 642 582 680 584
rect 712 618 750 620
rect 990 618 1028 620
rect 712 617 779 618
rect 712 585 715 617
rect 747 585 779 617
rect 712 584 779 585
rect 961 617 1028 618
rect 961 585 993 617
rect 1025 585 1028 617
rect 961 584 1028 585
rect 712 582 750 584
rect 990 582 1028 584
rect 1060 618 1098 620
rect 1338 618 1376 620
rect 1060 617 1127 618
rect 1060 585 1063 617
rect 1095 585 1127 617
rect 1060 584 1127 585
rect 1309 617 1376 618
rect 1309 585 1341 617
rect 1373 585 1376 617
rect 1309 584 1376 585
rect 1060 582 1098 584
rect 1338 582 1376 584
rect 1408 618 1446 620
rect 1686 618 1724 620
rect 1408 617 1475 618
rect 1408 585 1411 617
rect 1443 585 1475 617
rect 1408 584 1475 585
rect 1657 617 1724 618
rect 1657 585 1689 617
rect 1721 585 1724 617
rect 1657 584 1724 585
rect 1408 582 1446 584
rect 1686 582 1724 584
rect 1756 618 1794 620
rect 2034 618 2072 620
rect 1756 617 1823 618
rect 1756 585 1759 617
rect 1791 585 1823 617
rect 1756 584 1823 585
rect 2005 617 2072 618
rect 2005 585 2037 617
rect 2069 585 2072 617
rect 2005 584 2072 585
rect 1756 582 1794 584
rect 2034 582 2072 584
rect 2104 618 2142 620
rect 2382 618 2420 620
rect 2104 617 2171 618
rect 2104 585 2107 617
rect 2139 585 2171 617
rect 2104 584 2171 585
rect 2353 617 2420 618
rect 2353 585 2385 617
rect 2417 585 2420 617
rect 2353 584 2420 585
rect 2104 582 2142 584
rect 2382 582 2420 584
rect 2452 618 2490 620
rect 2730 618 2768 620
rect 2452 617 2519 618
rect 2452 585 2455 617
rect 2487 585 2519 617
rect 2452 584 2519 585
rect 2701 617 2768 618
rect 2701 585 2733 617
rect 2765 585 2768 617
rect 2701 584 2768 585
rect 2452 582 2490 584
rect 2730 582 2768 584
rect 2800 618 2838 620
rect 3078 618 3116 620
rect 2800 617 2867 618
rect 2800 585 2803 617
rect 2835 585 2867 617
rect 2800 584 2867 585
rect 3049 617 3116 618
rect 3049 585 3081 617
rect 3113 585 3116 617
rect 3049 584 3116 585
rect 2800 582 2838 584
rect 3078 582 3116 584
rect 3148 618 3186 620
rect 3426 618 3464 620
rect 3148 617 3215 618
rect 3148 585 3151 617
rect 3183 585 3215 617
rect 3148 584 3215 585
rect 3397 617 3464 618
rect 3397 585 3429 617
rect 3461 585 3464 617
rect 3397 584 3464 585
rect 3148 582 3186 584
rect 3426 582 3464 584
rect 3496 618 3534 620
rect 3774 618 3812 620
rect 3496 617 3563 618
rect 3496 585 3499 617
rect 3531 585 3563 617
rect 3496 584 3563 585
rect 3745 617 3812 618
rect 3745 585 3777 617
rect 3809 585 3812 617
rect 3745 584 3812 585
rect 3496 582 3534 584
rect 3774 582 3812 584
rect 3844 618 3882 620
rect 4122 618 4160 620
rect 3844 617 3911 618
rect 3844 585 3847 617
rect 3879 585 3911 617
rect 3844 584 3911 585
rect 4093 617 4160 618
rect 4093 585 4125 617
rect 4157 585 4160 617
rect 4093 584 4160 585
rect 3844 582 3882 584
rect 4122 582 4160 584
rect 4192 618 4230 620
rect 4470 618 4508 620
rect 4192 617 4259 618
rect 4192 585 4195 617
rect 4227 585 4259 617
rect 4192 584 4259 585
rect 4441 617 4508 618
rect 4441 585 4473 617
rect 4505 585 4508 617
rect 4441 584 4508 585
rect 4192 582 4230 584
rect 4470 582 4508 584
rect 4540 618 4578 620
rect 4818 618 4856 620
rect 4540 617 4607 618
rect 4540 585 4543 617
rect 4575 585 4607 617
rect 4540 584 4607 585
rect 4789 617 4856 618
rect 4789 585 4821 617
rect 4853 585 4856 617
rect 4789 584 4856 585
rect 4540 582 4578 584
rect 4818 582 4856 584
rect 4888 618 4926 620
rect 5166 618 5204 620
rect 4888 617 4955 618
rect 4888 585 4891 617
rect 4923 585 4955 617
rect 4888 584 4955 585
rect 5137 617 5204 618
rect 5137 585 5169 617
rect 5201 585 5204 617
rect 5137 584 5204 585
rect 4888 582 4926 584
rect 5166 582 5204 584
rect 5236 618 5274 620
rect 5514 618 5552 620
rect 5236 617 5303 618
rect 5236 585 5239 617
rect 5271 585 5303 617
rect 5236 584 5303 585
rect 5485 617 5552 618
rect 5485 585 5517 617
rect 5549 585 5552 617
rect 5485 584 5552 585
rect 5236 582 5274 584
rect 5514 582 5552 584
rect 5584 618 5622 620
rect 5862 618 5900 620
rect 5584 617 5651 618
rect 5584 585 5587 617
rect 5619 585 5651 617
rect 5584 584 5651 585
rect 5833 617 5900 618
rect 5833 585 5865 617
rect 5897 585 5900 617
rect 5833 584 5900 585
rect 5584 582 5622 584
rect 5862 582 5900 584
rect 5932 618 5970 620
rect 6210 618 6248 620
rect 5932 617 5999 618
rect 5932 585 5935 617
rect 5967 585 5999 617
rect 5932 584 5999 585
rect 6181 617 6248 618
rect 6181 585 6213 617
rect 6245 585 6248 617
rect 6181 584 6248 585
rect 5932 582 5970 584
rect 6210 582 6248 584
rect 6280 618 6318 620
rect 6558 618 6596 620
rect 6280 617 6347 618
rect 6280 585 6283 617
rect 6315 585 6347 617
rect 6280 584 6347 585
rect 6529 617 6596 618
rect 6529 585 6561 617
rect 6593 585 6596 617
rect 6529 584 6596 585
rect 6280 582 6318 584
rect 6558 582 6596 584
rect 6628 618 6666 620
rect 6906 618 6944 620
rect 6628 617 6695 618
rect 6628 585 6631 617
rect 6663 585 6695 617
rect 6628 584 6695 585
rect 6877 617 6944 618
rect 6877 585 6909 617
rect 6941 585 6944 617
rect 6877 584 6944 585
rect 6628 582 6666 584
rect 6906 582 6944 584
rect 6976 618 7014 620
rect 7254 618 7292 620
rect 6976 617 7043 618
rect 6976 585 6979 617
rect 7011 585 7043 617
rect 6976 584 7043 585
rect 7225 617 7292 618
rect 7225 585 7257 617
rect 7289 585 7292 617
rect 7225 584 7292 585
rect 6976 582 7014 584
rect 7254 582 7292 584
rect 16 548 54 550
rect 294 548 332 550
rect 16 547 83 548
rect 16 515 19 547
rect 51 515 83 547
rect 16 514 83 515
rect 265 547 332 548
rect 265 515 297 547
rect 329 515 332 547
rect 265 514 332 515
rect 16 512 54 514
rect 294 512 332 514
rect 364 548 402 550
rect 642 548 680 550
rect 364 547 431 548
rect 364 515 367 547
rect 399 515 431 547
rect 364 514 431 515
rect 613 547 680 548
rect 613 515 645 547
rect 677 515 680 547
rect 613 514 680 515
rect 364 512 402 514
rect 642 512 680 514
rect 712 548 750 550
rect 990 548 1028 550
rect 712 547 779 548
rect 712 515 715 547
rect 747 515 779 547
rect 712 514 779 515
rect 961 547 1028 548
rect 961 515 993 547
rect 1025 515 1028 547
rect 961 514 1028 515
rect 712 512 750 514
rect 990 512 1028 514
rect 1060 548 1098 550
rect 1338 548 1376 550
rect 1060 547 1127 548
rect 1060 515 1063 547
rect 1095 515 1127 547
rect 1060 514 1127 515
rect 1309 547 1376 548
rect 1309 515 1341 547
rect 1373 515 1376 547
rect 1309 514 1376 515
rect 1060 512 1098 514
rect 1338 512 1376 514
rect 1408 548 1446 550
rect 1686 548 1724 550
rect 1408 547 1475 548
rect 1408 515 1411 547
rect 1443 515 1475 547
rect 1408 514 1475 515
rect 1657 547 1724 548
rect 1657 515 1689 547
rect 1721 515 1724 547
rect 1657 514 1724 515
rect 1408 512 1446 514
rect 1686 512 1724 514
rect 1756 548 1794 550
rect 2034 548 2072 550
rect 1756 547 1823 548
rect 1756 515 1759 547
rect 1791 515 1823 547
rect 1756 514 1823 515
rect 2005 547 2072 548
rect 2005 515 2037 547
rect 2069 515 2072 547
rect 2005 514 2072 515
rect 1756 512 1794 514
rect 2034 512 2072 514
rect 2104 548 2142 550
rect 2382 548 2420 550
rect 2104 547 2171 548
rect 2104 515 2107 547
rect 2139 515 2171 547
rect 2104 514 2171 515
rect 2353 547 2420 548
rect 2353 515 2385 547
rect 2417 515 2420 547
rect 2353 514 2420 515
rect 2104 512 2142 514
rect 2382 512 2420 514
rect 2452 548 2490 550
rect 2730 548 2768 550
rect 2452 547 2519 548
rect 2452 515 2455 547
rect 2487 515 2519 547
rect 2452 514 2519 515
rect 2701 547 2768 548
rect 2701 515 2733 547
rect 2765 515 2768 547
rect 2701 514 2768 515
rect 2452 512 2490 514
rect 2730 512 2768 514
rect 2800 548 2838 550
rect 3078 548 3116 550
rect 2800 547 2867 548
rect 2800 515 2803 547
rect 2835 515 2867 547
rect 2800 514 2867 515
rect 3049 547 3116 548
rect 3049 515 3081 547
rect 3113 515 3116 547
rect 3049 514 3116 515
rect 2800 512 2838 514
rect 3078 512 3116 514
rect 3148 548 3186 550
rect 3426 548 3464 550
rect 3148 547 3215 548
rect 3148 515 3151 547
rect 3183 515 3215 547
rect 3148 514 3215 515
rect 3397 547 3464 548
rect 3397 515 3429 547
rect 3461 515 3464 547
rect 3397 514 3464 515
rect 3148 512 3186 514
rect 3426 512 3464 514
rect 3496 548 3534 550
rect 3774 548 3812 550
rect 3496 547 3563 548
rect 3496 515 3499 547
rect 3531 515 3563 547
rect 3496 514 3563 515
rect 3745 547 3812 548
rect 3745 515 3777 547
rect 3809 515 3812 547
rect 3745 514 3812 515
rect 3496 512 3534 514
rect 3774 512 3812 514
rect 3844 548 3882 550
rect 4122 548 4160 550
rect 3844 547 3911 548
rect 3844 515 3847 547
rect 3879 515 3911 547
rect 3844 514 3911 515
rect 4093 547 4160 548
rect 4093 515 4125 547
rect 4157 515 4160 547
rect 4093 514 4160 515
rect 3844 512 3882 514
rect 4122 512 4160 514
rect 4192 548 4230 550
rect 4470 548 4508 550
rect 4192 547 4259 548
rect 4192 515 4195 547
rect 4227 515 4259 547
rect 4192 514 4259 515
rect 4441 547 4508 548
rect 4441 515 4473 547
rect 4505 515 4508 547
rect 4441 514 4508 515
rect 4192 512 4230 514
rect 4470 512 4508 514
rect 4540 548 4578 550
rect 4818 548 4856 550
rect 4540 547 4607 548
rect 4540 515 4543 547
rect 4575 515 4607 547
rect 4540 514 4607 515
rect 4789 547 4856 548
rect 4789 515 4821 547
rect 4853 515 4856 547
rect 4789 514 4856 515
rect 4540 512 4578 514
rect 4818 512 4856 514
rect 4888 548 4926 550
rect 5166 548 5204 550
rect 4888 547 4955 548
rect 4888 515 4891 547
rect 4923 515 4955 547
rect 4888 514 4955 515
rect 5137 547 5204 548
rect 5137 515 5169 547
rect 5201 515 5204 547
rect 5137 514 5204 515
rect 4888 512 4926 514
rect 5166 512 5204 514
rect 5236 548 5274 550
rect 5514 548 5552 550
rect 5236 547 5303 548
rect 5236 515 5239 547
rect 5271 515 5303 547
rect 5236 514 5303 515
rect 5485 547 5552 548
rect 5485 515 5517 547
rect 5549 515 5552 547
rect 5485 514 5552 515
rect 5236 512 5274 514
rect 5514 512 5552 514
rect 5584 548 5622 550
rect 5862 548 5900 550
rect 5584 547 5651 548
rect 5584 515 5587 547
rect 5619 515 5651 547
rect 5584 514 5651 515
rect 5833 547 5900 548
rect 5833 515 5865 547
rect 5897 515 5900 547
rect 5833 514 5900 515
rect 5584 512 5622 514
rect 5862 512 5900 514
rect 5932 548 5970 550
rect 6210 548 6248 550
rect 5932 547 5999 548
rect 5932 515 5935 547
rect 5967 515 5999 547
rect 5932 514 5999 515
rect 6181 547 6248 548
rect 6181 515 6213 547
rect 6245 515 6248 547
rect 6181 514 6248 515
rect 5932 512 5970 514
rect 6210 512 6248 514
rect 6280 548 6318 550
rect 6558 548 6596 550
rect 6280 547 6347 548
rect 6280 515 6283 547
rect 6315 515 6347 547
rect 6280 514 6347 515
rect 6529 547 6596 548
rect 6529 515 6561 547
rect 6593 515 6596 547
rect 6529 514 6596 515
rect 6280 512 6318 514
rect 6558 512 6596 514
rect 6628 548 6666 550
rect 6906 548 6944 550
rect 6628 547 6695 548
rect 6628 515 6631 547
rect 6663 515 6695 547
rect 6628 514 6695 515
rect 6877 547 6944 548
rect 6877 515 6909 547
rect 6941 515 6944 547
rect 6877 514 6944 515
rect 6628 512 6666 514
rect 6906 512 6944 514
rect 6976 548 7014 550
rect 7254 548 7292 550
rect 6976 547 7043 548
rect 6976 515 6979 547
rect 7011 515 7043 547
rect 6976 514 7043 515
rect 7225 547 7292 548
rect 7225 515 7257 547
rect 7289 515 7292 547
rect 7225 514 7292 515
rect 6976 512 7014 514
rect 7254 512 7292 514
rect 16 424 54 426
rect 294 424 332 426
rect 16 423 83 424
rect 16 391 19 423
rect 51 391 83 423
rect 16 390 83 391
rect 265 423 332 424
rect 265 391 297 423
rect 329 391 332 423
rect 265 390 332 391
rect 16 388 54 390
rect 294 388 332 390
rect 364 424 402 426
rect 642 424 680 426
rect 364 423 431 424
rect 364 391 367 423
rect 399 391 431 423
rect 364 390 431 391
rect 613 423 680 424
rect 613 391 645 423
rect 677 391 680 423
rect 613 390 680 391
rect 364 388 402 390
rect 642 388 680 390
rect 712 424 750 426
rect 990 424 1028 426
rect 712 423 779 424
rect 712 391 715 423
rect 747 391 779 423
rect 712 390 779 391
rect 961 423 1028 424
rect 961 391 993 423
rect 1025 391 1028 423
rect 961 390 1028 391
rect 712 388 750 390
rect 990 388 1028 390
rect 1060 424 1098 426
rect 1338 424 1376 426
rect 1060 423 1127 424
rect 1060 391 1063 423
rect 1095 391 1127 423
rect 1060 390 1127 391
rect 1309 423 1376 424
rect 1309 391 1341 423
rect 1373 391 1376 423
rect 1309 390 1376 391
rect 1060 388 1098 390
rect 1338 388 1376 390
rect 1408 424 1446 426
rect 1686 424 1724 426
rect 1408 423 1475 424
rect 1408 391 1411 423
rect 1443 391 1475 423
rect 1408 390 1475 391
rect 1657 423 1724 424
rect 1657 391 1689 423
rect 1721 391 1724 423
rect 1657 390 1724 391
rect 1408 388 1446 390
rect 1686 388 1724 390
rect 1756 424 1794 426
rect 2034 424 2072 426
rect 1756 423 1823 424
rect 1756 391 1759 423
rect 1791 391 1823 423
rect 1756 390 1823 391
rect 2005 423 2072 424
rect 2005 391 2037 423
rect 2069 391 2072 423
rect 2005 390 2072 391
rect 1756 388 1794 390
rect 2034 388 2072 390
rect 2104 424 2142 426
rect 2382 424 2420 426
rect 2104 423 2171 424
rect 2104 391 2107 423
rect 2139 391 2171 423
rect 2104 390 2171 391
rect 2353 423 2420 424
rect 2353 391 2385 423
rect 2417 391 2420 423
rect 2353 390 2420 391
rect 2104 388 2142 390
rect 2382 388 2420 390
rect 2452 424 2490 426
rect 2730 424 2768 426
rect 2452 423 2519 424
rect 2452 391 2455 423
rect 2487 391 2519 423
rect 2452 390 2519 391
rect 2701 423 2768 424
rect 2701 391 2733 423
rect 2765 391 2768 423
rect 2701 390 2768 391
rect 2452 388 2490 390
rect 2730 388 2768 390
rect 2800 424 2838 426
rect 3078 424 3116 426
rect 2800 423 2867 424
rect 2800 391 2803 423
rect 2835 391 2867 423
rect 2800 390 2867 391
rect 3049 423 3116 424
rect 3049 391 3081 423
rect 3113 391 3116 423
rect 3049 390 3116 391
rect 2800 388 2838 390
rect 3078 388 3116 390
rect 3148 424 3186 426
rect 3426 424 3464 426
rect 3148 423 3215 424
rect 3148 391 3151 423
rect 3183 391 3215 423
rect 3148 390 3215 391
rect 3397 423 3464 424
rect 3397 391 3429 423
rect 3461 391 3464 423
rect 3397 390 3464 391
rect 3148 388 3186 390
rect 3426 388 3464 390
rect 3496 424 3534 426
rect 3774 424 3812 426
rect 3496 423 3563 424
rect 3496 391 3499 423
rect 3531 391 3563 423
rect 3496 390 3563 391
rect 3745 423 3812 424
rect 3745 391 3777 423
rect 3809 391 3812 423
rect 3745 390 3812 391
rect 3496 388 3534 390
rect 3774 388 3812 390
rect 3844 424 3882 426
rect 4122 424 4160 426
rect 3844 423 3911 424
rect 3844 391 3847 423
rect 3879 391 3911 423
rect 3844 390 3911 391
rect 4093 423 4160 424
rect 4093 391 4125 423
rect 4157 391 4160 423
rect 4093 390 4160 391
rect 3844 388 3882 390
rect 4122 388 4160 390
rect 4192 424 4230 426
rect 4470 424 4508 426
rect 4192 423 4259 424
rect 4192 391 4195 423
rect 4227 391 4259 423
rect 4192 390 4259 391
rect 4441 423 4508 424
rect 4441 391 4473 423
rect 4505 391 4508 423
rect 4441 390 4508 391
rect 4192 388 4230 390
rect 4470 388 4508 390
rect 4540 424 4578 426
rect 4818 424 4856 426
rect 4540 423 4607 424
rect 4540 391 4543 423
rect 4575 391 4607 423
rect 4540 390 4607 391
rect 4789 423 4856 424
rect 4789 391 4821 423
rect 4853 391 4856 423
rect 4789 390 4856 391
rect 4540 388 4578 390
rect 4818 388 4856 390
rect 4888 424 4926 426
rect 5166 424 5204 426
rect 4888 423 4955 424
rect 4888 391 4891 423
rect 4923 391 4955 423
rect 4888 390 4955 391
rect 5137 423 5204 424
rect 5137 391 5169 423
rect 5201 391 5204 423
rect 5137 390 5204 391
rect 4888 388 4926 390
rect 5166 388 5204 390
rect 5236 424 5274 426
rect 5514 424 5552 426
rect 5236 423 5303 424
rect 5236 391 5239 423
rect 5271 391 5303 423
rect 5236 390 5303 391
rect 5485 423 5552 424
rect 5485 391 5517 423
rect 5549 391 5552 423
rect 5485 390 5552 391
rect 5236 388 5274 390
rect 5514 388 5552 390
rect 5584 424 5622 426
rect 5862 424 5900 426
rect 5584 423 5651 424
rect 5584 391 5587 423
rect 5619 391 5651 423
rect 5584 390 5651 391
rect 5833 423 5900 424
rect 5833 391 5865 423
rect 5897 391 5900 423
rect 5833 390 5900 391
rect 5584 388 5622 390
rect 5862 388 5900 390
rect 5932 424 5970 426
rect 6210 424 6248 426
rect 5932 423 5999 424
rect 5932 391 5935 423
rect 5967 391 5999 423
rect 5932 390 5999 391
rect 6181 423 6248 424
rect 6181 391 6213 423
rect 6245 391 6248 423
rect 6181 390 6248 391
rect 5932 388 5970 390
rect 6210 388 6248 390
rect 6280 424 6318 426
rect 6558 424 6596 426
rect 6280 423 6347 424
rect 6280 391 6283 423
rect 6315 391 6347 423
rect 6280 390 6347 391
rect 6529 423 6596 424
rect 6529 391 6561 423
rect 6593 391 6596 423
rect 6529 390 6596 391
rect 6280 388 6318 390
rect 6558 388 6596 390
rect 6628 424 6666 426
rect 6906 424 6944 426
rect 6628 423 6695 424
rect 6628 391 6631 423
rect 6663 391 6695 423
rect 6628 390 6695 391
rect 6877 423 6944 424
rect 6877 391 6909 423
rect 6941 391 6944 423
rect 6877 390 6944 391
rect 6628 388 6666 390
rect 6906 388 6944 390
rect 6976 424 7014 426
rect 7254 424 7292 426
rect 6976 423 7043 424
rect 6976 391 6979 423
rect 7011 391 7043 423
rect 6976 390 7043 391
rect 7225 423 7292 424
rect 7225 391 7257 423
rect 7289 391 7292 423
rect 7225 390 7292 391
rect 6976 388 7014 390
rect 7254 388 7292 390
rect 16 300 54 302
rect 294 300 332 302
rect 16 299 83 300
rect 16 267 19 299
rect 51 267 83 299
rect 16 266 83 267
rect 265 299 332 300
rect 265 267 297 299
rect 329 267 332 299
rect 265 266 332 267
rect 16 264 54 266
rect 294 264 332 266
rect 364 300 402 302
rect 642 300 680 302
rect 364 299 431 300
rect 364 267 367 299
rect 399 267 431 299
rect 364 266 431 267
rect 613 299 680 300
rect 613 267 645 299
rect 677 267 680 299
rect 613 266 680 267
rect 364 264 402 266
rect 642 264 680 266
rect 712 300 750 302
rect 990 300 1028 302
rect 712 299 779 300
rect 712 267 715 299
rect 747 267 779 299
rect 712 266 779 267
rect 961 299 1028 300
rect 961 267 993 299
rect 1025 267 1028 299
rect 961 266 1028 267
rect 712 264 750 266
rect 990 264 1028 266
rect 1060 300 1098 302
rect 1338 300 1376 302
rect 1060 299 1127 300
rect 1060 267 1063 299
rect 1095 267 1127 299
rect 1060 266 1127 267
rect 1309 299 1376 300
rect 1309 267 1341 299
rect 1373 267 1376 299
rect 1309 266 1376 267
rect 1060 264 1098 266
rect 1338 264 1376 266
rect 1408 300 1446 302
rect 1686 300 1724 302
rect 1408 299 1475 300
rect 1408 267 1411 299
rect 1443 267 1475 299
rect 1408 266 1475 267
rect 1657 299 1724 300
rect 1657 267 1689 299
rect 1721 267 1724 299
rect 1657 266 1724 267
rect 1408 264 1446 266
rect 1686 264 1724 266
rect 1756 300 1794 302
rect 2034 300 2072 302
rect 1756 299 1823 300
rect 1756 267 1759 299
rect 1791 267 1823 299
rect 1756 266 1823 267
rect 2005 299 2072 300
rect 2005 267 2037 299
rect 2069 267 2072 299
rect 2005 266 2072 267
rect 1756 264 1794 266
rect 2034 264 2072 266
rect 2104 300 2142 302
rect 2382 300 2420 302
rect 2104 299 2171 300
rect 2104 267 2107 299
rect 2139 267 2171 299
rect 2104 266 2171 267
rect 2353 299 2420 300
rect 2353 267 2385 299
rect 2417 267 2420 299
rect 2353 266 2420 267
rect 2104 264 2142 266
rect 2382 264 2420 266
rect 2452 300 2490 302
rect 2730 300 2768 302
rect 2452 299 2519 300
rect 2452 267 2455 299
rect 2487 267 2519 299
rect 2452 266 2519 267
rect 2701 299 2768 300
rect 2701 267 2733 299
rect 2765 267 2768 299
rect 2701 266 2768 267
rect 2452 264 2490 266
rect 2730 264 2768 266
rect 2800 300 2838 302
rect 3078 300 3116 302
rect 2800 299 2867 300
rect 2800 267 2803 299
rect 2835 267 2867 299
rect 2800 266 2867 267
rect 3049 299 3116 300
rect 3049 267 3081 299
rect 3113 267 3116 299
rect 3049 266 3116 267
rect 2800 264 2838 266
rect 3078 264 3116 266
rect 3148 300 3186 302
rect 3426 300 3464 302
rect 3148 299 3215 300
rect 3148 267 3151 299
rect 3183 267 3215 299
rect 3148 266 3215 267
rect 3397 299 3464 300
rect 3397 267 3429 299
rect 3461 267 3464 299
rect 3397 266 3464 267
rect 3148 264 3186 266
rect 3426 264 3464 266
rect 3496 300 3534 302
rect 3774 300 3812 302
rect 3496 299 3563 300
rect 3496 267 3499 299
rect 3531 267 3563 299
rect 3496 266 3563 267
rect 3745 299 3812 300
rect 3745 267 3777 299
rect 3809 267 3812 299
rect 3745 266 3812 267
rect 3496 264 3534 266
rect 3774 264 3812 266
rect 3844 300 3882 302
rect 4122 300 4160 302
rect 3844 299 3911 300
rect 3844 267 3847 299
rect 3879 267 3911 299
rect 3844 266 3911 267
rect 4093 299 4160 300
rect 4093 267 4125 299
rect 4157 267 4160 299
rect 4093 266 4160 267
rect 3844 264 3882 266
rect 4122 264 4160 266
rect 4192 300 4230 302
rect 4470 300 4508 302
rect 4192 299 4259 300
rect 4192 267 4195 299
rect 4227 267 4259 299
rect 4192 266 4259 267
rect 4441 299 4508 300
rect 4441 267 4473 299
rect 4505 267 4508 299
rect 4441 266 4508 267
rect 4192 264 4230 266
rect 4470 264 4508 266
rect 4540 300 4578 302
rect 4818 300 4856 302
rect 4540 299 4607 300
rect 4540 267 4543 299
rect 4575 267 4607 299
rect 4540 266 4607 267
rect 4789 299 4856 300
rect 4789 267 4821 299
rect 4853 267 4856 299
rect 4789 266 4856 267
rect 4540 264 4578 266
rect 4818 264 4856 266
rect 4888 300 4926 302
rect 5166 300 5204 302
rect 4888 299 4955 300
rect 4888 267 4891 299
rect 4923 267 4955 299
rect 4888 266 4955 267
rect 5137 299 5204 300
rect 5137 267 5169 299
rect 5201 267 5204 299
rect 5137 266 5204 267
rect 4888 264 4926 266
rect 5166 264 5204 266
rect 5236 300 5274 302
rect 5514 300 5552 302
rect 5236 299 5303 300
rect 5236 267 5239 299
rect 5271 267 5303 299
rect 5236 266 5303 267
rect 5485 299 5552 300
rect 5485 267 5517 299
rect 5549 267 5552 299
rect 5485 266 5552 267
rect 5236 264 5274 266
rect 5514 264 5552 266
rect 5584 300 5622 302
rect 5862 300 5900 302
rect 5584 299 5651 300
rect 5584 267 5587 299
rect 5619 267 5651 299
rect 5584 266 5651 267
rect 5833 299 5900 300
rect 5833 267 5865 299
rect 5897 267 5900 299
rect 5833 266 5900 267
rect 5584 264 5622 266
rect 5862 264 5900 266
rect 5932 300 5970 302
rect 6210 300 6248 302
rect 5932 299 5999 300
rect 5932 267 5935 299
rect 5967 267 5999 299
rect 5932 266 5999 267
rect 6181 299 6248 300
rect 6181 267 6213 299
rect 6245 267 6248 299
rect 6181 266 6248 267
rect 5932 264 5970 266
rect 6210 264 6248 266
rect 6280 300 6318 302
rect 6558 300 6596 302
rect 6280 299 6347 300
rect 6280 267 6283 299
rect 6315 267 6347 299
rect 6280 266 6347 267
rect 6529 299 6596 300
rect 6529 267 6561 299
rect 6593 267 6596 299
rect 6529 266 6596 267
rect 6280 264 6318 266
rect 6558 264 6596 266
rect 6628 300 6666 302
rect 6906 300 6944 302
rect 6628 299 6695 300
rect 6628 267 6631 299
rect 6663 267 6695 299
rect 6628 266 6695 267
rect 6877 299 6944 300
rect 6877 267 6909 299
rect 6941 267 6944 299
rect 6877 266 6944 267
rect 6628 264 6666 266
rect 6906 264 6944 266
rect 6976 300 7014 302
rect 7254 300 7292 302
rect 6976 299 7043 300
rect 6976 267 6979 299
rect 7011 267 7043 299
rect 6976 266 7043 267
rect 7225 299 7292 300
rect 7225 267 7257 299
rect 7289 267 7292 299
rect 7225 266 7292 267
rect 6976 264 7014 266
rect 7254 264 7292 266
rect 16 176 54 178
rect 294 176 332 178
rect 16 175 83 176
rect 16 143 19 175
rect 51 143 83 175
rect 16 142 83 143
rect 265 175 332 176
rect 265 143 297 175
rect 329 143 332 175
rect 265 142 332 143
rect 16 140 54 142
rect 294 140 332 142
rect 364 176 402 178
rect 642 176 680 178
rect 364 175 431 176
rect 364 143 367 175
rect 399 143 431 175
rect 364 142 431 143
rect 613 175 680 176
rect 613 143 645 175
rect 677 143 680 175
rect 613 142 680 143
rect 364 140 402 142
rect 642 140 680 142
rect 712 176 750 178
rect 990 176 1028 178
rect 712 175 779 176
rect 712 143 715 175
rect 747 143 779 175
rect 712 142 779 143
rect 961 175 1028 176
rect 961 143 993 175
rect 1025 143 1028 175
rect 961 142 1028 143
rect 712 140 750 142
rect 990 140 1028 142
rect 1060 176 1098 178
rect 1338 176 1376 178
rect 1060 175 1127 176
rect 1060 143 1063 175
rect 1095 143 1127 175
rect 1060 142 1127 143
rect 1309 175 1376 176
rect 1309 143 1341 175
rect 1373 143 1376 175
rect 1309 142 1376 143
rect 1060 140 1098 142
rect 1338 140 1376 142
rect 1408 176 1446 178
rect 1686 176 1724 178
rect 1408 175 1475 176
rect 1408 143 1411 175
rect 1443 143 1475 175
rect 1408 142 1475 143
rect 1657 175 1724 176
rect 1657 143 1689 175
rect 1721 143 1724 175
rect 1657 142 1724 143
rect 1408 140 1446 142
rect 1686 140 1724 142
rect 1756 176 1794 178
rect 2034 176 2072 178
rect 1756 175 1823 176
rect 1756 143 1759 175
rect 1791 143 1823 175
rect 1756 142 1823 143
rect 2005 175 2072 176
rect 2005 143 2037 175
rect 2069 143 2072 175
rect 2005 142 2072 143
rect 1756 140 1794 142
rect 2034 140 2072 142
rect 2104 176 2142 178
rect 2382 176 2420 178
rect 2104 175 2171 176
rect 2104 143 2107 175
rect 2139 143 2171 175
rect 2104 142 2171 143
rect 2353 175 2420 176
rect 2353 143 2385 175
rect 2417 143 2420 175
rect 2353 142 2420 143
rect 2104 140 2142 142
rect 2382 140 2420 142
rect 2452 176 2490 178
rect 2730 176 2768 178
rect 2452 175 2519 176
rect 2452 143 2455 175
rect 2487 143 2519 175
rect 2452 142 2519 143
rect 2701 175 2768 176
rect 2701 143 2733 175
rect 2765 143 2768 175
rect 2701 142 2768 143
rect 2452 140 2490 142
rect 2730 140 2768 142
rect 2800 176 2838 178
rect 3078 176 3116 178
rect 2800 175 2867 176
rect 2800 143 2803 175
rect 2835 143 2867 175
rect 2800 142 2867 143
rect 3049 175 3116 176
rect 3049 143 3081 175
rect 3113 143 3116 175
rect 3049 142 3116 143
rect 2800 140 2838 142
rect 3078 140 3116 142
rect 3148 176 3186 178
rect 3426 176 3464 178
rect 3148 175 3215 176
rect 3148 143 3151 175
rect 3183 143 3215 175
rect 3148 142 3215 143
rect 3397 175 3464 176
rect 3397 143 3429 175
rect 3461 143 3464 175
rect 3397 142 3464 143
rect 3148 140 3186 142
rect 3426 140 3464 142
rect 3496 176 3534 178
rect 3774 176 3812 178
rect 3496 175 3563 176
rect 3496 143 3499 175
rect 3531 143 3563 175
rect 3496 142 3563 143
rect 3745 175 3812 176
rect 3745 143 3777 175
rect 3809 143 3812 175
rect 3745 142 3812 143
rect 3496 140 3534 142
rect 3774 140 3812 142
rect 3844 176 3882 178
rect 4122 176 4160 178
rect 3844 175 3911 176
rect 3844 143 3847 175
rect 3879 143 3911 175
rect 3844 142 3911 143
rect 4093 175 4160 176
rect 4093 143 4125 175
rect 4157 143 4160 175
rect 4093 142 4160 143
rect 3844 140 3882 142
rect 4122 140 4160 142
rect 4192 176 4230 178
rect 4470 176 4508 178
rect 4192 175 4259 176
rect 4192 143 4195 175
rect 4227 143 4259 175
rect 4192 142 4259 143
rect 4441 175 4508 176
rect 4441 143 4473 175
rect 4505 143 4508 175
rect 4441 142 4508 143
rect 4192 140 4230 142
rect 4470 140 4508 142
rect 4540 176 4578 178
rect 4818 176 4856 178
rect 4540 175 4607 176
rect 4540 143 4543 175
rect 4575 143 4607 175
rect 4540 142 4607 143
rect 4789 175 4856 176
rect 4789 143 4821 175
rect 4853 143 4856 175
rect 4789 142 4856 143
rect 4540 140 4578 142
rect 4818 140 4856 142
rect 4888 176 4926 178
rect 5166 176 5204 178
rect 4888 175 4955 176
rect 4888 143 4891 175
rect 4923 143 4955 175
rect 4888 142 4955 143
rect 5137 175 5204 176
rect 5137 143 5169 175
rect 5201 143 5204 175
rect 5137 142 5204 143
rect 4888 140 4926 142
rect 5166 140 5204 142
rect 5236 176 5274 178
rect 5514 176 5552 178
rect 5236 175 5303 176
rect 5236 143 5239 175
rect 5271 143 5303 175
rect 5236 142 5303 143
rect 5485 175 5552 176
rect 5485 143 5517 175
rect 5549 143 5552 175
rect 5485 142 5552 143
rect 5236 140 5274 142
rect 5514 140 5552 142
rect 5584 176 5622 178
rect 5862 176 5900 178
rect 5584 175 5651 176
rect 5584 143 5587 175
rect 5619 143 5651 175
rect 5584 142 5651 143
rect 5833 175 5900 176
rect 5833 143 5865 175
rect 5897 143 5900 175
rect 5833 142 5900 143
rect 5584 140 5622 142
rect 5862 140 5900 142
rect 5932 176 5970 178
rect 6210 176 6248 178
rect 5932 175 5999 176
rect 5932 143 5935 175
rect 5967 143 5999 175
rect 5932 142 5999 143
rect 6181 175 6248 176
rect 6181 143 6213 175
rect 6245 143 6248 175
rect 6181 142 6248 143
rect 5932 140 5970 142
rect 6210 140 6248 142
rect 6280 176 6318 178
rect 6558 176 6596 178
rect 6280 175 6347 176
rect 6280 143 6283 175
rect 6315 143 6347 175
rect 6280 142 6347 143
rect 6529 175 6596 176
rect 6529 143 6561 175
rect 6593 143 6596 175
rect 6529 142 6596 143
rect 6280 140 6318 142
rect 6558 140 6596 142
rect 6628 176 6666 178
rect 6906 176 6944 178
rect 6628 175 6695 176
rect 6628 143 6631 175
rect 6663 143 6695 175
rect 6628 142 6695 143
rect 6877 175 6944 176
rect 6877 143 6909 175
rect 6941 143 6944 175
rect 6877 142 6944 143
rect 6628 140 6666 142
rect 6906 140 6944 142
rect 6976 176 7014 178
rect 7254 176 7292 178
rect 6976 175 7043 176
rect 6976 143 6979 175
rect 7011 143 7043 175
rect 6976 142 7043 143
rect 7225 175 7292 176
rect 7225 143 7257 175
rect 7289 143 7292 175
rect 7225 142 7292 143
rect 6976 140 7014 142
rect 7254 140 7292 142
rect 16 52 54 54
rect 294 52 332 54
rect 16 51 83 52
rect 16 19 19 51
rect 51 19 83 51
rect 16 18 83 19
rect 265 51 332 52
rect 265 19 297 51
rect 329 19 332 51
rect 265 18 332 19
rect 16 16 54 18
rect 294 16 332 18
rect 364 52 402 54
rect 642 52 680 54
rect 364 51 431 52
rect 364 19 367 51
rect 399 19 431 51
rect 364 18 431 19
rect 613 51 680 52
rect 613 19 645 51
rect 677 19 680 51
rect 613 18 680 19
rect 364 16 402 18
rect 642 16 680 18
rect 712 52 750 54
rect 990 52 1028 54
rect 712 51 779 52
rect 712 19 715 51
rect 747 19 779 51
rect 712 18 779 19
rect 961 51 1028 52
rect 961 19 993 51
rect 1025 19 1028 51
rect 961 18 1028 19
rect 712 16 750 18
rect 990 16 1028 18
rect 1060 52 1098 54
rect 1338 52 1376 54
rect 1060 51 1127 52
rect 1060 19 1063 51
rect 1095 19 1127 51
rect 1060 18 1127 19
rect 1309 51 1376 52
rect 1309 19 1341 51
rect 1373 19 1376 51
rect 1309 18 1376 19
rect 1060 16 1098 18
rect 1338 16 1376 18
rect 1408 52 1446 54
rect 1686 52 1724 54
rect 1408 51 1475 52
rect 1408 19 1411 51
rect 1443 19 1475 51
rect 1408 18 1475 19
rect 1657 51 1724 52
rect 1657 19 1689 51
rect 1721 19 1724 51
rect 1657 18 1724 19
rect 1408 16 1446 18
rect 1686 16 1724 18
rect 1756 52 1794 54
rect 2034 52 2072 54
rect 1756 51 1823 52
rect 1756 19 1759 51
rect 1791 19 1823 51
rect 1756 18 1823 19
rect 2005 51 2072 52
rect 2005 19 2037 51
rect 2069 19 2072 51
rect 2005 18 2072 19
rect 1756 16 1794 18
rect 2034 16 2072 18
rect 2104 52 2142 54
rect 2382 52 2420 54
rect 2104 51 2171 52
rect 2104 19 2107 51
rect 2139 19 2171 51
rect 2104 18 2171 19
rect 2353 51 2420 52
rect 2353 19 2385 51
rect 2417 19 2420 51
rect 2353 18 2420 19
rect 2104 16 2142 18
rect 2382 16 2420 18
rect 2452 52 2490 54
rect 2730 52 2768 54
rect 2452 51 2519 52
rect 2452 19 2455 51
rect 2487 19 2519 51
rect 2452 18 2519 19
rect 2701 51 2768 52
rect 2701 19 2733 51
rect 2765 19 2768 51
rect 2701 18 2768 19
rect 2452 16 2490 18
rect 2730 16 2768 18
rect 2800 52 2838 54
rect 3078 52 3116 54
rect 2800 51 2867 52
rect 2800 19 2803 51
rect 2835 19 2867 51
rect 2800 18 2867 19
rect 3049 51 3116 52
rect 3049 19 3081 51
rect 3113 19 3116 51
rect 3049 18 3116 19
rect 2800 16 2838 18
rect 3078 16 3116 18
rect 3148 52 3186 54
rect 3426 52 3464 54
rect 3148 51 3215 52
rect 3148 19 3151 51
rect 3183 19 3215 51
rect 3148 18 3215 19
rect 3397 51 3464 52
rect 3397 19 3429 51
rect 3461 19 3464 51
rect 3397 18 3464 19
rect 3148 16 3186 18
rect 3426 16 3464 18
rect 3496 52 3534 54
rect 3774 52 3812 54
rect 3496 51 3563 52
rect 3496 19 3499 51
rect 3531 19 3563 51
rect 3496 18 3563 19
rect 3745 51 3812 52
rect 3745 19 3777 51
rect 3809 19 3812 51
rect 3745 18 3812 19
rect 3496 16 3534 18
rect 3774 16 3812 18
rect 3844 52 3882 54
rect 4122 52 4160 54
rect 3844 51 3911 52
rect 3844 19 3847 51
rect 3879 19 3911 51
rect 3844 18 3911 19
rect 4093 51 4160 52
rect 4093 19 4125 51
rect 4157 19 4160 51
rect 4093 18 4160 19
rect 3844 16 3882 18
rect 4122 16 4160 18
rect 4192 52 4230 54
rect 4470 52 4508 54
rect 4192 51 4259 52
rect 4192 19 4195 51
rect 4227 19 4259 51
rect 4192 18 4259 19
rect 4441 51 4508 52
rect 4441 19 4473 51
rect 4505 19 4508 51
rect 4441 18 4508 19
rect 4192 16 4230 18
rect 4470 16 4508 18
rect 4540 52 4578 54
rect 4818 52 4856 54
rect 4540 51 4607 52
rect 4540 19 4543 51
rect 4575 19 4607 51
rect 4540 18 4607 19
rect 4789 51 4856 52
rect 4789 19 4821 51
rect 4853 19 4856 51
rect 4789 18 4856 19
rect 4540 16 4578 18
rect 4818 16 4856 18
rect 4888 52 4926 54
rect 5166 52 5204 54
rect 4888 51 4955 52
rect 4888 19 4891 51
rect 4923 19 4955 51
rect 4888 18 4955 19
rect 5137 51 5204 52
rect 5137 19 5169 51
rect 5201 19 5204 51
rect 5137 18 5204 19
rect 4888 16 4926 18
rect 5166 16 5204 18
rect 5236 52 5274 54
rect 5514 52 5552 54
rect 5236 51 5303 52
rect 5236 19 5239 51
rect 5271 19 5303 51
rect 5236 18 5303 19
rect 5485 51 5552 52
rect 5485 19 5517 51
rect 5549 19 5552 51
rect 5485 18 5552 19
rect 5236 16 5274 18
rect 5514 16 5552 18
rect 5584 52 5622 54
rect 5862 52 5900 54
rect 5584 51 5651 52
rect 5584 19 5587 51
rect 5619 19 5651 51
rect 5584 18 5651 19
rect 5833 51 5900 52
rect 5833 19 5865 51
rect 5897 19 5900 51
rect 5833 18 5900 19
rect 5584 16 5622 18
rect 5862 16 5900 18
rect 5932 52 5970 54
rect 6210 52 6248 54
rect 5932 51 5999 52
rect 5932 19 5935 51
rect 5967 19 5999 51
rect 5932 18 5999 19
rect 6181 51 6248 52
rect 6181 19 6213 51
rect 6245 19 6248 51
rect 6181 18 6248 19
rect 5932 16 5970 18
rect 6210 16 6248 18
rect 6280 52 6318 54
rect 6558 52 6596 54
rect 6280 51 6347 52
rect 6280 19 6283 51
rect 6315 19 6347 51
rect 6280 18 6347 19
rect 6529 51 6596 52
rect 6529 19 6561 51
rect 6593 19 6596 51
rect 6529 18 6596 19
rect 6280 16 6318 18
rect 6558 16 6596 18
rect 6628 52 6666 54
rect 6906 52 6944 54
rect 6628 51 6695 52
rect 6628 19 6631 51
rect 6663 19 6695 51
rect 6628 18 6695 19
rect 6877 51 6944 52
rect 6877 19 6909 51
rect 6941 19 6944 51
rect 6877 18 6944 19
rect 6628 16 6666 18
rect 6906 16 6944 18
rect 6976 52 7014 54
rect 7254 52 7292 54
rect 6976 51 7043 52
rect 6976 19 6979 51
rect 7011 19 7043 51
rect 6976 18 7043 19
rect 7225 51 7292 52
rect 7225 19 7257 51
rect 7289 19 7292 51
rect 7225 18 7292 19
rect 6976 16 7014 18
rect 7254 16 7292 18
<< via3 >>
rect 19 2213 51 2245
rect 297 2213 329 2245
rect 367 2213 399 2245
rect 645 2213 677 2245
rect 715 2213 747 2245
rect 993 2213 1025 2245
rect 1063 2213 1095 2245
rect 1341 2213 1373 2245
rect 1411 2213 1443 2245
rect 1689 2213 1721 2245
rect 1759 2213 1791 2245
rect 2037 2213 2069 2245
rect 2107 2213 2139 2245
rect 2385 2213 2417 2245
rect 2455 2213 2487 2245
rect 2733 2213 2765 2245
rect 2803 2213 2835 2245
rect 3081 2213 3113 2245
rect 3151 2213 3183 2245
rect 3429 2213 3461 2245
rect 3499 2213 3531 2245
rect 3777 2213 3809 2245
rect 3847 2213 3879 2245
rect 4125 2213 4157 2245
rect 4195 2213 4227 2245
rect 4473 2213 4505 2245
rect 4543 2213 4575 2245
rect 4821 2213 4853 2245
rect 4891 2213 4923 2245
rect 5169 2213 5201 2245
rect 5239 2213 5271 2245
rect 5517 2213 5549 2245
rect 5587 2213 5619 2245
rect 5865 2213 5897 2245
rect 5935 2213 5967 2245
rect 6213 2213 6245 2245
rect 6283 2213 6315 2245
rect 6561 2213 6593 2245
rect 6631 2213 6663 2245
rect 6909 2213 6941 2245
rect 6979 2213 7011 2245
rect 7257 2213 7289 2245
rect 19 2089 51 2121
rect 297 2089 329 2121
rect 367 2089 399 2121
rect 645 2089 677 2121
rect 715 2089 747 2121
rect 993 2089 1025 2121
rect 1063 2089 1095 2121
rect 1341 2089 1373 2121
rect 1411 2089 1443 2121
rect 1689 2089 1721 2121
rect 1759 2089 1791 2121
rect 2037 2089 2069 2121
rect 2107 2089 2139 2121
rect 2385 2089 2417 2121
rect 2455 2089 2487 2121
rect 2733 2089 2765 2121
rect 2803 2089 2835 2121
rect 3081 2089 3113 2121
rect 3151 2089 3183 2121
rect 3429 2089 3461 2121
rect 3499 2089 3531 2121
rect 3777 2089 3809 2121
rect 3847 2089 3879 2121
rect 4125 2089 4157 2121
rect 4195 2089 4227 2121
rect 4473 2089 4505 2121
rect 4543 2089 4575 2121
rect 4821 2089 4853 2121
rect 4891 2089 4923 2121
rect 5169 2089 5201 2121
rect 5239 2089 5271 2121
rect 5517 2089 5549 2121
rect 5587 2089 5619 2121
rect 5865 2089 5897 2121
rect 5935 2089 5967 2121
rect 6213 2089 6245 2121
rect 6283 2089 6315 2121
rect 6561 2089 6593 2121
rect 6631 2089 6663 2121
rect 6909 2089 6941 2121
rect 6979 2089 7011 2121
rect 7257 2089 7289 2121
rect 19 1965 51 1997
rect 297 1965 329 1997
rect 367 1965 399 1997
rect 645 1965 677 1997
rect 715 1965 747 1997
rect 993 1965 1025 1997
rect 1063 1965 1095 1997
rect 1341 1965 1373 1997
rect 1411 1965 1443 1997
rect 1689 1965 1721 1997
rect 1759 1965 1791 1997
rect 2037 1965 2069 1997
rect 2107 1965 2139 1997
rect 2385 1965 2417 1997
rect 2455 1965 2487 1997
rect 2733 1965 2765 1997
rect 2803 1965 2835 1997
rect 3081 1965 3113 1997
rect 3151 1965 3183 1997
rect 3429 1965 3461 1997
rect 3499 1965 3531 1997
rect 3777 1965 3809 1997
rect 3847 1965 3879 1997
rect 4125 1965 4157 1997
rect 4195 1965 4227 1997
rect 4473 1965 4505 1997
rect 4543 1965 4575 1997
rect 4821 1965 4853 1997
rect 4891 1965 4923 1997
rect 5169 1965 5201 1997
rect 5239 1965 5271 1997
rect 5517 1965 5549 1997
rect 5587 1965 5619 1997
rect 5865 1965 5897 1997
rect 5935 1965 5967 1997
rect 6213 1965 6245 1997
rect 6283 1965 6315 1997
rect 6561 1965 6593 1997
rect 6631 1965 6663 1997
rect 6909 1965 6941 1997
rect 6979 1965 7011 1997
rect 7257 1965 7289 1997
rect 19 1841 51 1873
rect 297 1841 329 1873
rect 367 1841 399 1873
rect 645 1841 677 1873
rect 715 1841 747 1873
rect 993 1841 1025 1873
rect 1063 1841 1095 1873
rect 1341 1841 1373 1873
rect 1411 1841 1443 1873
rect 1689 1841 1721 1873
rect 1759 1841 1791 1873
rect 2037 1841 2069 1873
rect 2107 1841 2139 1873
rect 2385 1841 2417 1873
rect 2455 1841 2487 1873
rect 2733 1841 2765 1873
rect 2803 1841 2835 1873
rect 3081 1841 3113 1873
rect 3151 1841 3183 1873
rect 3429 1841 3461 1873
rect 3499 1841 3531 1873
rect 3777 1841 3809 1873
rect 3847 1841 3879 1873
rect 4125 1841 4157 1873
rect 4195 1841 4227 1873
rect 4473 1841 4505 1873
rect 4543 1841 4575 1873
rect 4821 1841 4853 1873
rect 4891 1841 4923 1873
rect 5169 1841 5201 1873
rect 5239 1841 5271 1873
rect 5517 1841 5549 1873
rect 5587 1841 5619 1873
rect 5865 1841 5897 1873
rect 5935 1841 5967 1873
rect 6213 1841 6245 1873
rect 6283 1841 6315 1873
rect 6561 1841 6593 1873
rect 6631 1841 6663 1873
rect 6909 1841 6941 1873
rect 6979 1841 7011 1873
rect 7257 1841 7289 1873
rect 19 1717 51 1749
rect 297 1717 329 1749
rect 367 1717 399 1749
rect 645 1717 677 1749
rect 715 1717 747 1749
rect 993 1717 1025 1749
rect 1063 1717 1095 1749
rect 1341 1717 1373 1749
rect 1411 1717 1443 1749
rect 1689 1717 1721 1749
rect 1759 1717 1791 1749
rect 2037 1717 2069 1749
rect 2107 1717 2139 1749
rect 2385 1717 2417 1749
rect 2455 1717 2487 1749
rect 2733 1717 2765 1749
rect 2803 1717 2835 1749
rect 3081 1717 3113 1749
rect 3151 1717 3183 1749
rect 3429 1717 3461 1749
rect 3499 1717 3531 1749
rect 3777 1717 3809 1749
rect 3847 1717 3879 1749
rect 4125 1717 4157 1749
rect 4195 1717 4227 1749
rect 4473 1717 4505 1749
rect 4543 1717 4575 1749
rect 4821 1717 4853 1749
rect 4891 1717 4923 1749
rect 5169 1717 5201 1749
rect 5239 1717 5271 1749
rect 5517 1717 5549 1749
rect 5587 1717 5619 1749
rect 5865 1717 5897 1749
rect 5935 1717 5967 1749
rect 6213 1717 6245 1749
rect 6283 1717 6315 1749
rect 6561 1717 6593 1749
rect 6631 1717 6663 1749
rect 6909 1717 6941 1749
rect 6979 1717 7011 1749
rect 7257 1717 7289 1749
rect 19 1647 51 1679
rect 297 1647 329 1679
rect 367 1647 399 1679
rect 645 1647 677 1679
rect 715 1647 747 1679
rect 993 1647 1025 1679
rect 1063 1647 1095 1679
rect 1341 1647 1373 1679
rect 1411 1647 1443 1679
rect 1689 1647 1721 1679
rect 1759 1647 1791 1679
rect 2037 1647 2069 1679
rect 2107 1647 2139 1679
rect 2385 1647 2417 1679
rect 2455 1647 2487 1679
rect 2733 1647 2765 1679
rect 2803 1647 2835 1679
rect 3081 1647 3113 1679
rect 3151 1647 3183 1679
rect 3429 1647 3461 1679
rect 3499 1647 3531 1679
rect 3777 1647 3809 1679
rect 3847 1647 3879 1679
rect 4125 1647 4157 1679
rect 4195 1647 4227 1679
rect 4473 1647 4505 1679
rect 4543 1647 4575 1679
rect 4821 1647 4853 1679
rect 4891 1647 4923 1679
rect 5169 1647 5201 1679
rect 5239 1647 5271 1679
rect 5517 1647 5549 1679
rect 5587 1647 5619 1679
rect 5865 1647 5897 1679
rect 5935 1647 5967 1679
rect 6213 1647 6245 1679
rect 6283 1647 6315 1679
rect 6561 1647 6593 1679
rect 6631 1647 6663 1679
rect 6909 1647 6941 1679
rect 6979 1647 7011 1679
rect 7257 1647 7289 1679
rect 19 1523 51 1555
rect 297 1523 329 1555
rect 367 1523 399 1555
rect 645 1523 677 1555
rect 715 1523 747 1555
rect 993 1523 1025 1555
rect 1063 1523 1095 1555
rect 1341 1523 1373 1555
rect 1411 1523 1443 1555
rect 1689 1523 1721 1555
rect 1759 1523 1791 1555
rect 2037 1523 2069 1555
rect 2107 1523 2139 1555
rect 2385 1523 2417 1555
rect 2455 1523 2487 1555
rect 2733 1523 2765 1555
rect 2803 1523 2835 1555
rect 3081 1523 3113 1555
rect 3151 1523 3183 1555
rect 3429 1523 3461 1555
rect 3499 1523 3531 1555
rect 3777 1523 3809 1555
rect 3847 1523 3879 1555
rect 4125 1523 4157 1555
rect 4195 1523 4227 1555
rect 4473 1523 4505 1555
rect 4543 1523 4575 1555
rect 4821 1523 4853 1555
rect 4891 1523 4923 1555
rect 5169 1523 5201 1555
rect 5239 1523 5271 1555
rect 5517 1523 5549 1555
rect 5587 1523 5619 1555
rect 5865 1523 5897 1555
rect 5935 1523 5967 1555
rect 6213 1523 6245 1555
rect 6283 1523 6315 1555
rect 6561 1523 6593 1555
rect 6631 1523 6663 1555
rect 6909 1523 6941 1555
rect 6979 1523 7011 1555
rect 7257 1523 7289 1555
rect 19 1399 51 1431
rect 297 1399 329 1431
rect 367 1399 399 1431
rect 645 1399 677 1431
rect 715 1399 747 1431
rect 993 1399 1025 1431
rect 1063 1399 1095 1431
rect 1341 1399 1373 1431
rect 1411 1399 1443 1431
rect 1689 1399 1721 1431
rect 1759 1399 1791 1431
rect 2037 1399 2069 1431
rect 2107 1399 2139 1431
rect 2385 1399 2417 1431
rect 2455 1399 2487 1431
rect 2733 1399 2765 1431
rect 2803 1399 2835 1431
rect 3081 1399 3113 1431
rect 3151 1399 3183 1431
rect 3429 1399 3461 1431
rect 3499 1399 3531 1431
rect 3777 1399 3809 1431
rect 3847 1399 3879 1431
rect 4125 1399 4157 1431
rect 4195 1399 4227 1431
rect 4473 1399 4505 1431
rect 4543 1399 4575 1431
rect 4821 1399 4853 1431
rect 4891 1399 4923 1431
rect 5169 1399 5201 1431
rect 5239 1399 5271 1431
rect 5517 1399 5549 1431
rect 5587 1399 5619 1431
rect 5865 1399 5897 1431
rect 5935 1399 5967 1431
rect 6213 1399 6245 1431
rect 6283 1399 6315 1431
rect 6561 1399 6593 1431
rect 6631 1399 6663 1431
rect 6909 1399 6941 1431
rect 6979 1399 7011 1431
rect 7257 1399 7289 1431
rect 19 1275 51 1307
rect 297 1275 329 1307
rect 367 1275 399 1307
rect 645 1275 677 1307
rect 715 1275 747 1307
rect 993 1275 1025 1307
rect 1063 1275 1095 1307
rect 1341 1275 1373 1307
rect 1411 1275 1443 1307
rect 1689 1275 1721 1307
rect 1759 1275 1791 1307
rect 2037 1275 2069 1307
rect 2107 1275 2139 1307
rect 2385 1275 2417 1307
rect 2455 1275 2487 1307
rect 2733 1275 2765 1307
rect 2803 1275 2835 1307
rect 3081 1275 3113 1307
rect 3151 1275 3183 1307
rect 3429 1275 3461 1307
rect 3499 1275 3531 1307
rect 3777 1275 3809 1307
rect 3847 1275 3879 1307
rect 4125 1275 4157 1307
rect 4195 1275 4227 1307
rect 4473 1275 4505 1307
rect 4543 1275 4575 1307
rect 4821 1275 4853 1307
rect 4891 1275 4923 1307
rect 5169 1275 5201 1307
rect 5239 1275 5271 1307
rect 5517 1275 5549 1307
rect 5587 1275 5619 1307
rect 5865 1275 5897 1307
rect 5935 1275 5967 1307
rect 6213 1275 6245 1307
rect 6283 1275 6315 1307
rect 6561 1275 6593 1307
rect 6631 1275 6663 1307
rect 6909 1275 6941 1307
rect 6979 1275 7011 1307
rect 7257 1275 7289 1307
rect 19 1151 51 1183
rect 297 1151 329 1183
rect 367 1151 399 1183
rect 645 1151 677 1183
rect 715 1151 747 1183
rect 993 1151 1025 1183
rect 1063 1151 1095 1183
rect 1341 1151 1373 1183
rect 1411 1151 1443 1183
rect 1689 1151 1721 1183
rect 1759 1151 1791 1183
rect 2037 1151 2069 1183
rect 2107 1151 2139 1183
rect 2385 1151 2417 1183
rect 2455 1151 2487 1183
rect 2733 1151 2765 1183
rect 2803 1151 2835 1183
rect 3081 1151 3113 1183
rect 3151 1151 3183 1183
rect 3429 1151 3461 1183
rect 3499 1151 3531 1183
rect 3777 1151 3809 1183
rect 3847 1151 3879 1183
rect 4125 1151 4157 1183
rect 4195 1151 4227 1183
rect 4473 1151 4505 1183
rect 4543 1151 4575 1183
rect 4821 1151 4853 1183
rect 4891 1151 4923 1183
rect 5169 1151 5201 1183
rect 5239 1151 5271 1183
rect 5517 1151 5549 1183
rect 5587 1151 5619 1183
rect 5865 1151 5897 1183
rect 5935 1151 5967 1183
rect 6213 1151 6245 1183
rect 6283 1151 6315 1183
rect 6561 1151 6593 1183
rect 6631 1151 6663 1183
rect 6909 1151 6941 1183
rect 6979 1151 7011 1183
rect 7257 1151 7289 1183
rect 19 1081 51 1113
rect 297 1081 329 1113
rect 367 1081 399 1113
rect 645 1081 677 1113
rect 715 1081 747 1113
rect 993 1081 1025 1113
rect 1063 1081 1095 1113
rect 1341 1081 1373 1113
rect 1411 1081 1443 1113
rect 1689 1081 1721 1113
rect 1759 1081 1791 1113
rect 2037 1081 2069 1113
rect 2107 1081 2139 1113
rect 2385 1081 2417 1113
rect 2455 1081 2487 1113
rect 2733 1081 2765 1113
rect 2803 1081 2835 1113
rect 3081 1081 3113 1113
rect 3151 1081 3183 1113
rect 3429 1081 3461 1113
rect 3499 1081 3531 1113
rect 3777 1081 3809 1113
rect 3847 1081 3879 1113
rect 4125 1081 4157 1113
rect 4195 1081 4227 1113
rect 4473 1081 4505 1113
rect 4543 1081 4575 1113
rect 4821 1081 4853 1113
rect 4891 1081 4923 1113
rect 5169 1081 5201 1113
rect 5239 1081 5271 1113
rect 5517 1081 5549 1113
rect 5587 1081 5619 1113
rect 5865 1081 5897 1113
rect 5935 1081 5967 1113
rect 6213 1081 6245 1113
rect 6283 1081 6315 1113
rect 6561 1081 6593 1113
rect 6631 1081 6663 1113
rect 6909 1081 6941 1113
rect 6979 1081 7011 1113
rect 7257 1081 7289 1113
rect 19 957 51 989
rect 297 957 329 989
rect 367 957 399 989
rect 645 957 677 989
rect 715 957 747 989
rect 993 957 1025 989
rect 1063 957 1095 989
rect 1341 957 1373 989
rect 1411 957 1443 989
rect 1689 957 1721 989
rect 1759 957 1791 989
rect 2037 957 2069 989
rect 2107 957 2139 989
rect 2385 957 2417 989
rect 2455 957 2487 989
rect 2733 957 2765 989
rect 2803 957 2835 989
rect 3081 957 3113 989
rect 3151 957 3183 989
rect 3429 957 3461 989
rect 3499 957 3531 989
rect 3777 957 3809 989
rect 3847 957 3879 989
rect 4125 957 4157 989
rect 4195 957 4227 989
rect 4473 957 4505 989
rect 4543 957 4575 989
rect 4821 957 4853 989
rect 4891 957 4923 989
rect 5169 957 5201 989
rect 5239 957 5271 989
rect 5517 957 5549 989
rect 5587 957 5619 989
rect 5865 957 5897 989
rect 5935 957 5967 989
rect 6213 957 6245 989
rect 6283 957 6315 989
rect 6561 957 6593 989
rect 6631 957 6663 989
rect 6909 957 6941 989
rect 6979 957 7011 989
rect 7257 957 7289 989
rect 19 833 51 865
rect 297 833 329 865
rect 367 833 399 865
rect 645 833 677 865
rect 715 833 747 865
rect 993 833 1025 865
rect 1063 833 1095 865
rect 1341 833 1373 865
rect 1411 833 1443 865
rect 1689 833 1721 865
rect 1759 833 1791 865
rect 2037 833 2069 865
rect 2107 833 2139 865
rect 2385 833 2417 865
rect 2455 833 2487 865
rect 2733 833 2765 865
rect 2803 833 2835 865
rect 3081 833 3113 865
rect 3151 833 3183 865
rect 3429 833 3461 865
rect 3499 833 3531 865
rect 3777 833 3809 865
rect 3847 833 3879 865
rect 4125 833 4157 865
rect 4195 833 4227 865
rect 4473 833 4505 865
rect 4543 833 4575 865
rect 4821 833 4853 865
rect 4891 833 4923 865
rect 5169 833 5201 865
rect 5239 833 5271 865
rect 5517 833 5549 865
rect 5587 833 5619 865
rect 5865 833 5897 865
rect 5935 833 5967 865
rect 6213 833 6245 865
rect 6283 833 6315 865
rect 6561 833 6593 865
rect 6631 833 6663 865
rect 6909 833 6941 865
rect 6979 833 7011 865
rect 7257 833 7289 865
rect 19 709 51 741
rect 297 709 329 741
rect 367 709 399 741
rect 645 709 677 741
rect 715 709 747 741
rect 993 709 1025 741
rect 1063 709 1095 741
rect 1341 709 1373 741
rect 1411 709 1443 741
rect 1689 709 1721 741
rect 1759 709 1791 741
rect 2037 709 2069 741
rect 2107 709 2139 741
rect 2385 709 2417 741
rect 2455 709 2487 741
rect 2733 709 2765 741
rect 2803 709 2835 741
rect 3081 709 3113 741
rect 3151 709 3183 741
rect 3429 709 3461 741
rect 3499 709 3531 741
rect 3777 709 3809 741
rect 3847 709 3879 741
rect 4125 709 4157 741
rect 4195 709 4227 741
rect 4473 709 4505 741
rect 4543 709 4575 741
rect 4821 709 4853 741
rect 4891 709 4923 741
rect 5169 709 5201 741
rect 5239 709 5271 741
rect 5517 709 5549 741
rect 5587 709 5619 741
rect 5865 709 5897 741
rect 5935 709 5967 741
rect 6213 709 6245 741
rect 6283 709 6315 741
rect 6561 709 6593 741
rect 6631 709 6663 741
rect 6909 709 6941 741
rect 6979 709 7011 741
rect 7257 709 7289 741
rect 19 585 51 617
rect 297 585 329 617
rect 367 585 399 617
rect 645 585 677 617
rect 715 585 747 617
rect 993 585 1025 617
rect 1063 585 1095 617
rect 1341 585 1373 617
rect 1411 585 1443 617
rect 1689 585 1721 617
rect 1759 585 1791 617
rect 2037 585 2069 617
rect 2107 585 2139 617
rect 2385 585 2417 617
rect 2455 585 2487 617
rect 2733 585 2765 617
rect 2803 585 2835 617
rect 3081 585 3113 617
rect 3151 585 3183 617
rect 3429 585 3461 617
rect 3499 585 3531 617
rect 3777 585 3809 617
rect 3847 585 3879 617
rect 4125 585 4157 617
rect 4195 585 4227 617
rect 4473 585 4505 617
rect 4543 585 4575 617
rect 4821 585 4853 617
rect 4891 585 4923 617
rect 5169 585 5201 617
rect 5239 585 5271 617
rect 5517 585 5549 617
rect 5587 585 5619 617
rect 5865 585 5897 617
rect 5935 585 5967 617
rect 6213 585 6245 617
rect 6283 585 6315 617
rect 6561 585 6593 617
rect 6631 585 6663 617
rect 6909 585 6941 617
rect 6979 585 7011 617
rect 7257 585 7289 617
rect 19 515 51 547
rect 297 515 329 547
rect 367 515 399 547
rect 645 515 677 547
rect 715 515 747 547
rect 993 515 1025 547
rect 1063 515 1095 547
rect 1341 515 1373 547
rect 1411 515 1443 547
rect 1689 515 1721 547
rect 1759 515 1791 547
rect 2037 515 2069 547
rect 2107 515 2139 547
rect 2385 515 2417 547
rect 2455 515 2487 547
rect 2733 515 2765 547
rect 2803 515 2835 547
rect 3081 515 3113 547
rect 3151 515 3183 547
rect 3429 515 3461 547
rect 3499 515 3531 547
rect 3777 515 3809 547
rect 3847 515 3879 547
rect 4125 515 4157 547
rect 4195 515 4227 547
rect 4473 515 4505 547
rect 4543 515 4575 547
rect 4821 515 4853 547
rect 4891 515 4923 547
rect 5169 515 5201 547
rect 5239 515 5271 547
rect 5517 515 5549 547
rect 5587 515 5619 547
rect 5865 515 5897 547
rect 5935 515 5967 547
rect 6213 515 6245 547
rect 6283 515 6315 547
rect 6561 515 6593 547
rect 6631 515 6663 547
rect 6909 515 6941 547
rect 6979 515 7011 547
rect 7257 515 7289 547
rect 19 391 51 423
rect 297 391 329 423
rect 367 391 399 423
rect 645 391 677 423
rect 715 391 747 423
rect 993 391 1025 423
rect 1063 391 1095 423
rect 1341 391 1373 423
rect 1411 391 1443 423
rect 1689 391 1721 423
rect 1759 391 1791 423
rect 2037 391 2069 423
rect 2107 391 2139 423
rect 2385 391 2417 423
rect 2455 391 2487 423
rect 2733 391 2765 423
rect 2803 391 2835 423
rect 3081 391 3113 423
rect 3151 391 3183 423
rect 3429 391 3461 423
rect 3499 391 3531 423
rect 3777 391 3809 423
rect 3847 391 3879 423
rect 4125 391 4157 423
rect 4195 391 4227 423
rect 4473 391 4505 423
rect 4543 391 4575 423
rect 4821 391 4853 423
rect 4891 391 4923 423
rect 5169 391 5201 423
rect 5239 391 5271 423
rect 5517 391 5549 423
rect 5587 391 5619 423
rect 5865 391 5897 423
rect 5935 391 5967 423
rect 6213 391 6245 423
rect 6283 391 6315 423
rect 6561 391 6593 423
rect 6631 391 6663 423
rect 6909 391 6941 423
rect 6979 391 7011 423
rect 7257 391 7289 423
rect 19 267 51 299
rect 297 267 329 299
rect 367 267 399 299
rect 645 267 677 299
rect 715 267 747 299
rect 993 267 1025 299
rect 1063 267 1095 299
rect 1341 267 1373 299
rect 1411 267 1443 299
rect 1689 267 1721 299
rect 1759 267 1791 299
rect 2037 267 2069 299
rect 2107 267 2139 299
rect 2385 267 2417 299
rect 2455 267 2487 299
rect 2733 267 2765 299
rect 2803 267 2835 299
rect 3081 267 3113 299
rect 3151 267 3183 299
rect 3429 267 3461 299
rect 3499 267 3531 299
rect 3777 267 3809 299
rect 3847 267 3879 299
rect 4125 267 4157 299
rect 4195 267 4227 299
rect 4473 267 4505 299
rect 4543 267 4575 299
rect 4821 267 4853 299
rect 4891 267 4923 299
rect 5169 267 5201 299
rect 5239 267 5271 299
rect 5517 267 5549 299
rect 5587 267 5619 299
rect 5865 267 5897 299
rect 5935 267 5967 299
rect 6213 267 6245 299
rect 6283 267 6315 299
rect 6561 267 6593 299
rect 6631 267 6663 299
rect 6909 267 6941 299
rect 6979 267 7011 299
rect 7257 267 7289 299
rect 19 143 51 175
rect 297 143 329 175
rect 367 143 399 175
rect 645 143 677 175
rect 715 143 747 175
rect 993 143 1025 175
rect 1063 143 1095 175
rect 1341 143 1373 175
rect 1411 143 1443 175
rect 1689 143 1721 175
rect 1759 143 1791 175
rect 2037 143 2069 175
rect 2107 143 2139 175
rect 2385 143 2417 175
rect 2455 143 2487 175
rect 2733 143 2765 175
rect 2803 143 2835 175
rect 3081 143 3113 175
rect 3151 143 3183 175
rect 3429 143 3461 175
rect 3499 143 3531 175
rect 3777 143 3809 175
rect 3847 143 3879 175
rect 4125 143 4157 175
rect 4195 143 4227 175
rect 4473 143 4505 175
rect 4543 143 4575 175
rect 4821 143 4853 175
rect 4891 143 4923 175
rect 5169 143 5201 175
rect 5239 143 5271 175
rect 5517 143 5549 175
rect 5587 143 5619 175
rect 5865 143 5897 175
rect 5935 143 5967 175
rect 6213 143 6245 175
rect 6283 143 6315 175
rect 6561 143 6593 175
rect 6631 143 6663 175
rect 6909 143 6941 175
rect 6979 143 7011 175
rect 7257 143 7289 175
rect 19 19 51 51
rect 297 19 329 51
rect 367 19 399 51
rect 645 19 677 51
rect 715 19 747 51
rect 993 19 1025 51
rect 1063 19 1095 51
rect 1341 19 1373 51
rect 1411 19 1443 51
rect 1689 19 1721 51
rect 1759 19 1791 51
rect 2037 19 2069 51
rect 2107 19 2139 51
rect 2385 19 2417 51
rect 2455 19 2487 51
rect 2733 19 2765 51
rect 2803 19 2835 51
rect 3081 19 3113 51
rect 3151 19 3183 51
rect 3429 19 3461 51
rect 3499 19 3531 51
rect 3777 19 3809 51
rect 3847 19 3879 51
rect 4125 19 4157 51
rect 4195 19 4227 51
rect 4473 19 4505 51
rect 4543 19 4575 51
rect 4821 19 4853 51
rect 4891 19 4923 51
rect 5169 19 5201 51
rect 5239 19 5271 51
rect 5517 19 5549 51
rect 5587 19 5619 51
rect 5865 19 5897 51
rect 5935 19 5967 51
rect 6213 19 6245 51
rect 6283 19 6315 51
rect 6561 19 6593 51
rect 6631 19 6663 51
rect 6909 19 6941 51
rect 6979 19 7011 51
rect 7257 19 7289 51
<< metal4 >>
rect 18 2245 52 2246
rect 18 2244 19 2245
rect 16 2214 19 2244
rect 18 2213 19 2214
rect 51 2244 52 2245
rect 51 2214 130 2244
rect 51 2213 52 2214
rect 18 2212 52 2213
rect 160 2182 190 2264
rect 296 2245 330 2246
rect 296 2244 297 2245
rect 220 2214 297 2244
rect 296 2213 297 2214
rect 329 2244 330 2245
rect 366 2245 400 2246
rect 366 2244 367 2245
rect 329 2214 332 2244
rect 364 2214 367 2244
rect 329 2213 330 2214
rect 296 2212 330 2213
rect 366 2213 367 2214
rect 399 2244 400 2245
rect 399 2214 478 2244
rect 399 2213 400 2214
rect 366 2212 400 2213
rect 508 2182 538 2264
rect 644 2245 678 2246
rect 644 2244 645 2245
rect 568 2214 645 2244
rect 644 2213 645 2214
rect 677 2244 678 2245
rect 714 2245 748 2246
rect 714 2244 715 2245
rect 677 2214 680 2244
rect 712 2214 715 2244
rect 677 2213 678 2214
rect 644 2212 678 2213
rect 714 2213 715 2214
rect 747 2244 748 2245
rect 747 2214 826 2244
rect 747 2213 748 2214
rect 714 2212 748 2213
rect 856 2182 886 2264
rect 992 2245 1026 2246
rect 992 2244 993 2245
rect 916 2214 993 2244
rect 992 2213 993 2214
rect 1025 2244 1026 2245
rect 1062 2245 1096 2246
rect 1062 2244 1063 2245
rect 1025 2214 1028 2244
rect 1060 2214 1063 2244
rect 1025 2213 1026 2214
rect 992 2212 1026 2213
rect 1062 2213 1063 2214
rect 1095 2244 1096 2245
rect 1095 2214 1174 2244
rect 1095 2213 1096 2214
rect 1062 2212 1096 2213
rect 1204 2182 1234 2264
rect 1340 2245 1374 2246
rect 1340 2244 1341 2245
rect 1264 2214 1341 2244
rect 1340 2213 1341 2214
rect 1373 2244 1374 2245
rect 1410 2245 1444 2246
rect 1410 2244 1411 2245
rect 1373 2214 1376 2244
rect 1408 2214 1411 2244
rect 1373 2213 1374 2214
rect 1340 2212 1374 2213
rect 1410 2213 1411 2214
rect 1443 2244 1444 2245
rect 1443 2214 1522 2244
rect 1443 2213 1444 2214
rect 1410 2212 1444 2213
rect 1552 2182 1582 2264
rect 1688 2245 1722 2246
rect 1688 2244 1689 2245
rect 1612 2214 1689 2244
rect 1688 2213 1689 2214
rect 1721 2244 1722 2245
rect 1758 2245 1792 2246
rect 1758 2244 1759 2245
rect 1721 2214 1724 2244
rect 1756 2214 1759 2244
rect 1721 2213 1722 2214
rect 1688 2212 1722 2213
rect 1758 2213 1759 2214
rect 1791 2244 1792 2245
rect 1791 2214 1870 2244
rect 1791 2213 1792 2214
rect 1758 2212 1792 2213
rect 1900 2182 1930 2264
rect 2036 2245 2070 2246
rect 2036 2244 2037 2245
rect 1960 2214 2037 2244
rect 2036 2213 2037 2214
rect 2069 2244 2070 2245
rect 2106 2245 2140 2246
rect 2106 2244 2107 2245
rect 2069 2214 2072 2244
rect 2104 2214 2107 2244
rect 2069 2213 2070 2214
rect 2036 2212 2070 2213
rect 2106 2213 2107 2214
rect 2139 2244 2140 2245
rect 2139 2214 2218 2244
rect 2139 2213 2140 2214
rect 2106 2212 2140 2213
rect 2248 2182 2278 2264
rect 2384 2245 2418 2246
rect 2384 2244 2385 2245
rect 2308 2214 2385 2244
rect 2384 2213 2385 2214
rect 2417 2244 2418 2245
rect 2454 2245 2488 2246
rect 2454 2244 2455 2245
rect 2417 2214 2420 2244
rect 2452 2214 2455 2244
rect 2417 2213 2418 2214
rect 2384 2212 2418 2213
rect 2454 2213 2455 2214
rect 2487 2244 2488 2245
rect 2487 2214 2566 2244
rect 2487 2213 2488 2214
rect 2454 2212 2488 2213
rect 2596 2182 2626 2264
rect 2732 2245 2766 2246
rect 2732 2244 2733 2245
rect 2656 2214 2733 2244
rect 2732 2213 2733 2214
rect 2765 2244 2766 2245
rect 2802 2245 2836 2246
rect 2802 2244 2803 2245
rect 2765 2214 2768 2244
rect 2800 2214 2803 2244
rect 2765 2213 2766 2214
rect 2732 2212 2766 2213
rect 2802 2213 2803 2214
rect 2835 2244 2836 2245
rect 2835 2214 2914 2244
rect 2835 2213 2836 2214
rect 2802 2212 2836 2213
rect 2944 2182 2974 2264
rect 3080 2245 3114 2246
rect 3080 2244 3081 2245
rect 3004 2214 3081 2244
rect 3080 2213 3081 2214
rect 3113 2244 3114 2245
rect 3150 2245 3184 2246
rect 3150 2244 3151 2245
rect 3113 2214 3116 2244
rect 3148 2214 3151 2244
rect 3113 2213 3114 2214
rect 3080 2212 3114 2213
rect 3150 2213 3151 2214
rect 3183 2244 3184 2245
rect 3183 2214 3262 2244
rect 3183 2213 3184 2214
rect 3150 2212 3184 2213
rect 3292 2182 3322 2264
rect 3428 2245 3462 2246
rect 3428 2244 3429 2245
rect 3352 2214 3429 2244
rect 3428 2213 3429 2214
rect 3461 2244 3462 2245
rect 3498 2245 3532 2246
rect 3498 2244 3499 2245
rect 3461 2214 3464 2244
rect 3496 2214 3499 2244
rect 3461 2213 3462 2214
rect 3428 2212 3462 2213
rect 3498 2213 3499 2214
rect 3531 2244 3532 2245
rect 3531 2214 3610 2244
rect 3531 2213 3532 2214
rect 3498 2212 3532 2213
rect 3640 2182 3670 2264
rect 3776 2245 3810 2246
rect 3776 2244 3777 2245
rect 3700 2214 3777 2244
rect 3776 2213 3777 2214
rect 3809 2244 3810 2245
rect 3846 2245 3880 2246
rect 3846 2244 3847 2245
rect 3809 2214 3812 2244
rect 3844 2214 3847 2244
rect 3809 2213 3810 2214
rect 3776 2212 3810 2213
rect 3846 2213 3847 2214
rect 3879 2244 3880 2245
rect 3879 2214 3958 2244
rect 3879 2213 3880 2214
rect 3846 2212 3880 2213
rect 3988 2182 4018 2264
rect 4124 2245 4158 2246
rect 4124 2244 4125 2245
rect 4048 2214 4125 2244
rect 4124 2213 4125 2214
rect 4157 2244 4158 2245
rect 4194 2245 4228 2246
rect 4194 2244 4195 2245
rect 4157 2214 4160 2244
rect 4192 2214 4195 2244
rect 4157 2213 4158 2214
rect 4124 2212 4158 2213
rect 4194 2213 4195 2214
rect 4227 2244 4228 2245
rect 4227 2214 4306 2244
rect 4227 2213 4228 2214
rect 4194 2212 4228 2213
rect 4336 2182 4366 2264
rect 4472 2245 4506 2246
rect 4472 2244 4473 2245
rect 4396 2214 4473 2244
rect 4472 2213 4473 2214
rect 4505 2244 4506 2245
rect 4542 2245 4576 2246
rect 4542 2244 4543 2245
rect 4505 2214 4508 2244
rect 4540 2214 4543 2244
rect 4505 2213 4506 2214
rect 4472 2212 4506 2213
rect 4542 2213 4543 2214
rect 4575 2244 4576 2245
rect 4575 2214 4654 2244
rect 4575 2213 4576 2214
rect 4542 2212 4576 2213
rect 4684 2182 4714 2264
rect 4820 2245 4854 2246
rect 4820 2244 4821 2245
rect 4744 2214 4821 2244
rect 4820 2213 4821 2214
rect 4853 2244 4854 2245
rect 4890 2245 4924 2246
rect 4890 2244 4891 2245
rect 4853 2214 4856 2244
rect 4888 2214 4891 2244
rect 4853 2213 4854 2214
rect 4820 2212 4854 2213
rect 4890 2213 4891 2214
rect 4923 2244 4924 2245
rect 4923 2214 5002 2244
rect 4923 2213 4924 2214
rect 4890 2212 4924 2213
rect 5032 2182 5062 2264
rect 5168 2245 5202 2246
rect 5168 2244 5169 2245
rect 5092 2214 5169 2244
rect 5168 2213 5169 2214
rect 5201 2244 5202 2245
rect 5238 2245 5272 2246
rect 5238 2244 5239 2245
rect 5201 2214 5204 2244
rect 5236 2214 5239 2244
rect 5201 2213 5202 2214
rect 5168 2212 5202 2213
rect 5238 2213 5239 2214
rect 5271 2244 5272 2245
rect 5271 2214 5350 2244
rect 5271 2213 5272 2214
rect 5238 2212 5272 2213
rect 5380 2182 5410 2264
rect 5516 2245 5550 2246
rect 5516 2244 5517 2245
rect 5440 2214 5517 2244
rect 5516 2213 5517 2214
rect 5549 2244 5550 2245
rect 5586 2245 5620 2246
rect 5586 2244 5587 2245
rect 5549 2214 5552 2244
rect 5584 2214 5587 2244
rect 5549 2213 5550 2214
rect 5516 2212 5550 2213
rect 5586 2213 5587 2214
rect 5619 2244 5620 2245
rect 5619 2214 5698 2244
rect 5619 2213 5620 2214
rect 5586 2212 5620 2213
rect 5728 2182 5758 2264
rect 5864 2245 5898 2246
rect 5864 2244 5865 2245
rect 5788 2214 5865 2244
rect 5864 2213 5865 2214
rect 5897 2244 5898 2245
rect 5934 2245 5968 2246
rect 5934 2244 5935 2245
rect 5897 2214 5900 2244
rect 5932 2214 5935 2244
rect 5897 2213 5898 2214
rect 5864 2212 5898 2213
rect 5934 2213 5935 2214
rect 5967 2244 5968 2245
rect 5967 2214 6046 2244
rect 5967 2213 5968 2214
rect 5934 2212 5968 2213
rect 6076 2182 6106 2264
rect 6212 2245 6246 2246
rect 6212 2244 6213 2245
rect 6136 2214 6213 2244
rect 6212 2213 6213 2214
rect 6245 2244 6246 2245
rect 6282 2245 6316 2246
rect 6282 2244 6283 2245
rect 6245 2214 6248 2244
rect 6280 2214 6283 2244
rect 6245 2213 6246 2214
rect 6212 2212 6246 2213
rect 6282 2213 6283 2214
rect 6315 2244 6316 2245
rect 6315 2214 6394 2244
rect 6315 2213 6316 2214
rect 6282 2212 6316 2213
rect 6424 2182 6454 2264
rect 6560 2245 6594 2246
rect 6560 2244 6561 2245
rect 6484 2214 6561 2244
rect 6560 2213 6561 2214
rect 6593 2244 6594 2245
rect 6630 2245 6664 2246
rect 6630 2244 6631 2245
rect 6593 2214 6596 2244
rect 6628 2214 6631 2244
rect 6593 2213 6594 2214
rect 6560 2212 6594 2213
rect 6630 2213 6631 2214
rect 6663 2244 6664 2245
rect 6663 2214 6742 2244
rect 6663 2213 6664 2214
rect 6630 2212 6664 2213
rect 6772 2182 6802 2264
rect 6908 2245 6942 2246
rect 6908 2244 6909 2245
rect 6832 2214 6909 2244
rect 6908 2213 6909 2214
rect 6941 2244 6942 2245
rect 6978 2245 7012 2246
rect 6978 2244 6979 2245
rect 6941 2214 6944 2244
rect 6976 2214 6979 2244
rect 6941 2213 6942 2214
rect 6908 2212 6942 2213
rect 6978 2213 6979 2214
rect 7011 2244 7012 2245
rect 7011 2214 7090 2244
rect 7011 2213 7012 2214
rect 6978 2212 7012 2213
rect 7120 2182 7150 2264
rect 7256 2245 7290 2246
rect 7256 2244 7257 2245
rect 7180 2214 7257 2244
rect 7256 2213 7257 2214
rect 7289 2244 7290 2245
rect 7289 2214 7292 2244
rect 7289 2213 7290 2214
rect 7256 2212 7290 2213
rect 0 2152 7307 2182
rect 18 2121 52 2122
rect 18 2120 19 2121
rect 16 2090 19 2120
rect 18 2089 19 2090
rect 51 2120 52 2121
rect 51 2090 130 2120
rect 51 2089 52 2090
rect 18 2088 52 2089
rect 160 2058 190 2152
rect 296 2121 330 2122
rect 296 2120 297 2121
rect 220 2090 297 2120
rect 296 2089 297 2090
rect 329 2120 330 2121
rect 366 2121 400 2122
rect 366 2120 367 2121
rect 329 2090 332 2120
rect 364 2090 367 2120
rect 329 2089 330 2090
rect 296 2088 330 2089
rect 366 2089 367 2090
rect 399 2120 400 2121
rect 399 2090 478 2120
rect 399 2089 400 2090
rect 366 2088 400 2089
rect 508 2058 538 2152
rect 644 2121 678 2122
rect 644 2120 645 2121
rect 568 2090 645 2120
rect 644 2089 645 2090
rect 677 2120 678 2121
rect 714 2121 748 2122
rect 714 2120 715 2121
rect 677 2090 680 2120
rect 712 2090 715 2120
rect 677 2089 678 2090
rect 644 2088 678 2089
rect 714 2089 715 2090
rect 747 2120 748 2121
rect 747 2090 826 2120
rect 747 2089 748 2090
rect 714 2088 748 2089
rect 856 2058 886 2152
rect 992 2121 1026 2122
rect 992 2120 993 2121
rect 916 2090 993 2120
rect 992 2089 993 2090
rect 1025 2120 1026 2121
rect 1062 2121 1096 2122
rect 1062 2120 1063 2121
rect 1025 2090 1028 2120
rect 1060 2090 1063 2120
rect 1025 2089 1026 2090
rect 992 2088 1026 2089
rect 1062 2089 1063 2090
rect 1095 2120 1096 2121
rect 1095 2090 1174 2120
rect 1095 2089 1096 2090
rect 1062 2088 1096 2089
rect 1204 2058 1234 2152
rect 1340 2121 1374 2122
rect 1340 2120 1341 2121
rect 1264 2090 1341 2120
rect 1340 2089 1341 2090
rect 1373 2120 1374 2121
rect 1410 2121 1444 2122
rect 1410 2120 1411 2121
rect 1373 2090 1376 2120
rect 1408 2090 1411 2120
rect 1373 2089 1374 2090
rect 1340 2088 1374 2089
rect 1410 2089 1411 2090
rect 1443 2120 1444 2121
rect 1443 2090 1522 2120
rect 1443 2089 1444 2090
rect 1410 2088 1444 2089
rect 1552 2058 1582 2152
rect 1688 2121 1722 2122
rect 1688 2120 1689 2121
rect 1612 2090 1689 2120
rect 1688 2089 1689 2090
rect 1721 2120 1722 2121
rect 1758 2121 1792 2122
rect 1758 2120 1759 2121
rect 1721 2090 1724 2120
rect 1756 2090 1759 2120
rect 1721 2089 1722 2090
rect 1688 2088 1722 2089
rect 1758 2089 1759 2090
rect 1791 2120 1792 2121
rect 1791 2090 1870 2120
rect 1791 2089 1792 2090
rect 1758 2088 1792 2089
rect 1900 2058 1930 2152
rect 2036 2121 2070 2122
rect 2036 2120 2037 2121
rect 1960 2090 2037 2120
rect 2036 2089 2037 2090
rect 2069 2120 2070 2121
rect 2106 2121 2140 2122
rect 2106 2120 2107 2121
rect 2069 2090 2072 2120
rect 2104 2090 2107 2120
rect 2069 2089 2070 2090
rect 2036 2088 2070 2089
rect 2106 2089 2107 2090
rect 2139 2120 2140 2121
rect 2139 2090 2218 2120
rect 2139 2089 2140 2090
rect 2106 2088 2140 2089
rect 2248 2058 2278 2152
rect 2384 2121 2418 2122
rect 2384 2120 2385 2121
rect 2308 2090 2385 2120
rect 2384 2089 2385 2090
rect 2417 2120 2418 2121
rect 2454 2121 2488 2122
rect 2454 2120 2455 2121
rect 2417 2090 2420 2120
rect 2452 2090 2455 2120
rect 2417 2089 2418 2090
rect 2384 2088 2418 2089
rect 2454 2089 2455 2090
rect 2487 2120 2488 2121
rect 2487 2090 2566 2120
rect 2487 2089 2488 2090
rect 2454 2088 2488 2089
rect 2596 2058 2626 2152
rect 2732 2121 2766 2122
rect 2732 2120 2733 2121
rect 2656 2090 2733 2120
rect 2732 2089 2733 2090
rect 2765 2120 2766 2121
rect 2802 2121 2836 2122
rect 2802 2120 2803 2121
rect 2765 2090 2768 2120
rect 2800 2090 2803 2120
rect 2765 2089 2766 2090
rect 2732 2088 2766 2089
rect 2802 2089 2803 2090
rect 2835 2120 2836 2121
rect 2835 2090 2914 2120
rect 2835 2089 2836 2090
rect 2802 2088 2836 2089
rect 2944 2058 2974 2152
rect 3080 2121 3114 2122
rect 3080 2120 3081 2121
rect 3004 2090 3081 2120
rect 3080 2089 3081 2090
rect 3113 2120 3114 2121
rect 3150 2121 3184 2122
rect 3150 2120 3151 2121
rect 3113 2090 3116 2120
rect 3148 2090 3151 2120
rect 3113 2089 3114 2090
rect 3080 2088 3114 2089
rect 3150 2089 3151 2090
rect 3183 2120 3184 2121
rect 3183 2090 3262 2120
rect 3183 2089 3184 2090
rect 3150 2088 3184 2089
rect 3292 2058 3322 2152
rect 3428 2121 3462 2122
rect 3428 2120 3429 2121
rect 3352 2090 3429 2120
rect 3428 2089 3429 2090
rect 3461 2120 3462 2121
rect 3498 2121 3532 2122
rect 3498 2120 3499 2121
rect 3461 2090 3464 2120
rect 3496 2090 3499 2120
rect 3461 2089 3462 2090
rect 3428 2088 3462 2089
rect 3498 2089 3499 2090
rect 3531 2120 3532 2121
rect 3531 2090 3610 2120
rect 3531 2089 3532 2090
rect 3498 2088 3532 2089
rect 3640 2058 3670 2152
rect 3776 2121 3810 2122
rect 3776 2120 3777 2121
rect 3700 2090 3777 2120
rect 3776 2089 3777 2090
rect 3809 2120 3810 2121
rect 3846 2121 3880 2122
rect 3846 2120 3847 2121
rect 3809 2090 3812 2120
rect 3844 2090 3847 2120
rect 3809 2089 3810 2090
rect 3776 2088 3810 2089
rect 3846 2089 3847 2090
rect 3879 2120 3880 2121
rect 3879 2090 3958 2120
rect 3879 2089 3880 2090
rect 3846 2088 3880 2089
rect 3988 2058 4018 2152
rect 4124 2121 4158 2122
rect 4124 2120 4125 2121
rect 4048 2090 4125 2120
rect 4124 2089 4125 2090
rect 4157 2120 4158 2121
rect 4194 2121 4228 2122
rect 4194 2120 4195 2121
rect 4157 2090 4160 2120
rect 4192 2090 4195 2120
rect 4157 2089 4158 2090
rect 4124 2088 4158 2089
rect 4194 2089 4195 2090
rect 4227 2120 4228 2121
rect 4227 2090 4306 2120
rect 4227 2089 4228 2090
rect 4194 2088 4228 2089
rect 4336 2058 4366 2152
rect 4472 2121 4506 2122
rect 4472 2120 4473 2121
rect 4396 2090 4473 2120
rect 4472 2089 4473 2090
rect 4505 2120 4506 2121
rect 4542 2121 4576 2122
rect 4542 2120 4543 2121
rect 4505 2090 4508 2120
rect 4540 2090 4543 2120
rect 4505 2089 4506 2090
rect 4472 2088 4506 2089
rect 4542 2089 4543 2090
rect 4575 2120 4576 2121
rect 4575 2090 4654 2120
rect 4575 2089 4576 2090
rect 4542 2088 4576 2089
rect 4684 2058 4714 2152
rect 4820 2121 4854 2122
rect 4820 2120 4821 2121
rect 4744 2090 4821 2120
rect 4820 2089 4821 2090
rect 4853 2120 4854 2121
rect 4890 2121 4924 2122
rect 4890 2120 4891 2121
rect 4853 2090 4856 2120
rect 4888 2090 4891 2120
rect 4853 2089 4854 2090
rect 4820 2088 4854 2089
rect 4890 2089 4891 2090
rect 4923 2120 4924 2121
rect 4923 2090 5002 2120
rect 4923 2089 4924 2090
rect 4890 2088 4924 2089
rect 5032 2058 5062 2152
rect 5168 2121 5202 2122
rect 5168 2120 5169 2121
rect 5092 2090 5169 2120
rect 5168 2089 5169 2090
rect 5201 2120 5202 2121
rect 5238 2121 5272 2122
rect 5238 2120 5239 2121
rect 5201 2090 5204 2120
rect 5236 2090 5239 2120
rect 5201 2089 5202 2090
rect 5168 2088 5202 2089
rect 5238 2089 5239 2090
rect 5271 2120 5272 2121
rect 5271 2090 5350 2120
rect 5271 2089 5272 2090
rect 5238 2088 5272 2089
rect 5380 2058 5410 2152
rect 5516 2121 5550 2122
rect 5516 2120 5517 2121
rect 5440 2090 5517 2120
rect 5516 2089 5517 2090
rect 5549 2120 5550 2121
rect 5586 2121 5620 2122
rect 5586 2120 5587 2121
rect 5549 2090 5552 2120
rect 5584 2090 5587 2120
rect 5549 2089 5550 2090
rect 5516 2088 5550 2089
rect 5586 2089 5587 2090
rect 5619 2120 5620 2121
rect 5619 2090 5698 2120
rect 5619 2089 5620 2090
rect 5586 2088 5620 2089
rect 5728 2058 5758 2152
rect 5864 2121 5898 2122
rect 5864 2120 5865 2121
rect 5788 2090 5865 2120
rect 5864 2089 5865 2090
rect 5897 2120 5898 2121
rect 5934 2121 5968 2122
rect 5934 2120 5935 2121
rect 5897 2090 5900 2120
rect 5932 2090 5935 2120
rect 5897 2089 5898 2090
rect 5864 2088 5898 2089
rect 5934 2089 5935 2090
rect 5967 2120 5968 2121
rect 5967 2090 6046 2120
rect 5967 2089 5968 2090
rect 5934 2088 5968 2089
rect 6076 2058 6106 2152
rect 6212 2121 6246 2122
rect 6212 2120 6213 2121
rect 6136 2090 6213 2120
rect 6212 2089 6213 2090
rect 6245 2120 6246 2121
rect 6282 2121 6316 2122
rect 6282 2120 6283 2121
rect 6245 2090 6248 2120
rect 6280 2090 6283 2120
rect 6245 2089 6246 2090
rect 6212 2088 6246 2089
rect 6282 2089 6283 2090
rect 6315 2120 6316 2121
rect 6315 2090 6394 2120
rect 6315 2089 6316 2090
rect 6282 2088 6316 2089
rect 6424 2058 6454 2152
rect 6560 2121 6594 2122
rect 6560 2120 6561 2121
rect 6484 2090 6561 2120
rect 6560 2089 6561 2090
rect 6593 2120 6594 2121
rect 6630 2121 6664 2122
rect 6630 2120 6631 2121
rect 6593 2090 6596 2120
rect 6628 2090 6631 2120
rect 6593 2089 6594 2090
rect 6560 2088 6594 2089
rect 6630 2089 6631 2090
rect 6663 2120 6664 2121
rect 6663 2090 6742 2120
rect 6663 2089 6664 2090
rect 6630 2088 6664 2089
rect 6772 2058 6802 2152
rect 6908 2121 6942 2122
rect 6908 2120 6909 2121
rect 6832 2090 6909 2120
rect 6908 2089 6909 2090
rect 6941 2120 6942 2121
rect 6978 2121 7012 2122
rect 6978 2120 6979 2121
rect 6941 2090 6944 2120
rect 6976 2090 6979 2120
rect 6941 2089 6942 2090
rect 6908 2088 6942 2089
rect 6978 2089 6979 2090
rect 7011 2120 7012 2121
rect 7011 2090 7090 2120
rect 7011 2089 7012 2090
rect 6978 2088 7012 2089
rect 7120 2058 7150 2152
rect 7256 2121 7290 2122
rect 7256 2120 7257 2121
rect 7180 2090 7257 2120
rect 7256 2089 7257 2090
rect 7289 2120 7290 2121
rect 7289 2090 7292 2120
rect 7289 2089 7290 2090
rect 7256 2088 7290 2089
rect 0 2028 7307 2058
rect 18 1997 52 1998
rect 18 1996 19 1997
rect 16 1966 19 1996
rect 18 1965 19 1966
rect 51 1996 52 1997
rect 51 1966 130 1996
rect 51 1965 52 1966
rect 18 1964 52 1965
rect 160 1934 190 2028
rect 296 1997 330 1998
rect 296 1996 297 1997
rect 220 1966 297 1996
rect 296 1965 297 1966
rect 329 1996 330 1997
rect 366 1997 400 1998
rect 366 1996 367 1997
rect 329 1966 332 1996
rect 364 1966 367 1996
rect 329 1965 330 1966
rect 296 1964 330 1965
rect 366 1965 367 1966
rect 399 1996 400 1997
rect 399 1966 478 1996
rect 399 1965 400 1966
rect 366 1964 400 1965
rect 508 1934 538 2028
rect 644 1997 678 1998
rect 644 1996 645 1997
rect 568 1966 645 1996
rect 644 1965 645 1966
rect 677 1996 678 1997
rect 714 1997 748 1998
rect 714 1996 715 1997
rect 677 1966 680 1996
rect 712 1966 715 1996
rect 677 1965 678 1966
rect 644 1964 678 1965
rect 714 1965 715 1966
rect 747 1996 748 1997
rect 747 1966 826 1996
rect 747 1965 748 1966
rect 714 1964 748 1965
rect 856 1934 886 2028
rect 992 1997 1026 1998
rect 992 1996 993 1997
rect 916 1966 993 1996
rect 992 1965 993 1966
rect 1025 1996 1026 1997
rect 1062 1997 1096 1998
rect 1062 1996 1063 1997
rect 1025 1966 1028 1996
rect 1060 1966 1063 1996
rect 1025 1965 1026 1966
rect 992 1964 1026 1965
rect 1062 1965 1063 1966
rect 1095 1996 1096 1997
rect 1095 1966 1174 1996
rect 1095 1965 1096 1966
rect 1062 1964 1096 1965
rect 1204 1934 1234 2028
rect 1340 1997 1374 1998
rect 1340 1996 1341 1997
rect 1264 1966 1341 1996
rect 1340 1965 1341 1966
rect 1373 1996 1374 1997
rect 1410 1997 1444 1998
rect 1410 1996 1411 1997
rect 1373 1966 1376 1996
rect 1408 1966 1411 1996
rect 1373 1965 1374 1966
rect 1340 1964 1374 1965
rect 1410 1965 1411 1966
rect 1443 1996 1444 1997
rect 1443 1966 1522 1996
rect 1443 1965 1444 1966
rect 1410 1964 1444 1965
rect 1552 1934 1582 2028
rect 1688 1997 1722 1998
rect 1688 1996 1689 1997
rect 1612 1966 1689 1996
rect 1688 1965 1689 1966
rect 1721 1996 1722 1997
rect 1758 1997 1792 1998
rect 1758 1996 1759 1997
rect 1721 1966 1724 1996
rect 1756 1966 1759 1996
rect 1721 1965 1722 1966
rect 1688 1964 1722 1965
rect 1758 1965 1759 1966
rect 1791 1996 1792 1997
rect 1791 1966 1870 1996
rect 1791 1965 1792 1966
rect 1758 1964 1792 1965
rect 1900 1934 1930 2028
rect 2036 1997 2070 1998
rect 2036 1996 2037 1997
rect 1960 1966 2037 1996
rect 2036 1965 2037 1966
rect 2069 1996 2070 1997
rect 2106 1997 2140 1998
rect 2106 1996 2107 1997
rect 2069 1966 2072 1996
rect 2104 1966 2107 1996
rect 2069 1965 2070 1966
rect 2036 1964 2070 1965
rect 2106 1965 2107 1966
rect 2139 1996 2140 1997
rect 2139 1966 2218 1996
rect 2139 1965 2140 1966
rect 2106 1964 2140 1965
rect 2248 1934 2278 2028
rect 2384 1997 2418 1998
rect 2384 1996 2385 1997
rect 2308 1966 2385 1996
rect 2384 1965 2385 1966
rect 2417 1996 2418 1997
rect 2454 1997 2488 1998
rect 2454 1996 2455 1997
rect 2417 1966 2420 1996
rect 2452 1966 2455 1996
rect 2417 1965 2418 1966
rect 2384 1964 2418 1965
rect 2454 1965 2455 1966
rect 2487 1996 2488 1997
rect 2487 1966 2566 1996
rect 2487 1965 2488 1966
rect 2454 1964 2488 1965
rect 2596 1934 2626 2028
rect 2732 1997 2766 1998
rect 2732 1996 2733 1997
rect 2656 1966 2733 1996
rect 2732 1965 2733 1966
rect 2765 1996 2766 1997
rect 2802 1997 2836 1998
rect 2802 1996 2803 1997
rect 2765 1966 2768 1996
rect 2800 1966 2803 1996
rect 2765 1965 2766 1966
rect 2732 1964 2766 1965
rect 2802 1965 2803 1966
rect 2835 1996 2836 1997
rect 2835 1966 2914 1996
rect 2835 1965 2836 1966
rect 2802 1964 2836 1965
rect 2944 1934 2974 2028
rect 3080 1997 3114 1998
rect 3080 1996 3081 1997
rect 3004 1966 3081 1996
rect 3080 1965 3081 1966
rect 3113 1996 3114 1997
rect 3150 1997 3184 1998
rect 3150 1996 3151 1997
rect 3113 1966 3116 1996
rect 3148 1966 3151 1996
rect 3113 1965 3114 1966
rect 3080 1964 3114 1965
rect 3150 1965 3151 1966
rect 3183 1996 3184 1997
rect 3183 1966 3262 1996
rect 3183 1965 3184 1966
rect 3150 1964 3184 1965
rect 3292 1934 3322 2028
rect 3428 1997 3462 1998
rect 3428 1996 3429 1997
rect 3352 1966 3429 1996
rect 3428 1965 3429 1966
rect 3461 1996 3462 1997
rect 3498 1997 3532 1998
rect 3498 1996 3499 1997
rect 3461 1966 3464 1996
rect 3496 1966 3499 1996
rect 3461 1965 3462 1966
rect 3428 1964 3462 1965
rect 3498 1965 3499 1966
rect 3531 1996 3532 1997
rect 3531 1966 3610 1996
rect 3531 1965 3532 1966
rect 3498 1964 3532 1965
rect 3640 1934 3670 2028
rect 3776 1997 3810 1998
rect 3776 1996 3777 1997
rect 3700 1966 3777 1996
rect 3776 1965 3777 1966
rect 3809 1996 3810 1997
rect 3846 1997 3880 1998
rect 3846 1996 3847 1997
rect 3809 1966 3812 1996
rect 3844 1966 3847 1996
rect 3809 1965 3810 1966
rect 3776 1964 3810 1965
rect 3846 1965 3847 1966
rect 3879 1996 3880 1997
rect 3879 1966 3958 1996
rect 3879 1965 3880 1966
rect 3846 1964 3880 1965
rect 3988 1934 4018 2028
rect 4124 1997 4158 1998
rect 4124 1996 4125 1997
rect 4048 1966 4125 1996
rect 4124 1965 4125 1966
rect 4157 1996 4158 1997
rect 4194 1997 4228 1998
rect 4194 1996 4195 1997
rect 4157 1966 4160 1996
rect 4192 1966 4195 1996
rect 4157 1965 4158 1966
rect 4124 1964 4158 1965
rect 4194 1965 4195 1966
rect 4227 1996 4228 1997
rect 4227 1966 4306 1996
rect 4227 1965 4228 1966
rect 4194 1964 4228 1965
rect 4336 1934 4366 2028
rect 4472 1997 4506 1998
rect 4472 1996 4473 1997
rect 4396 1966 4473 1996
rect 4472 1965 4473 1966
rect 4505 1996 4506 1997
rect 4542 1997 4576 1998
rect 4542 1996 4543 1997
rect 4505 1966 4508 1996
rect 4540 1966 4543 1996
rect 4505 1965 4506 1966
rect 4472 1964 4506 1965
rect 4542 1965 4543 1966
rect 4575 1996 4576 1997
rect 4575 1966 4654 1996
rect 4575 1965 4576 1966
rect 4542 1964 4576 1965
rect 4684 1934 4714 2028
rect 4820 1997 4854 1998
rect 4820 1996 4821 1997
rect 4744 1966 4821 1996
rect 4820 1965 4821 1966
rect 4853 1996 4854 1997
rect 4890 1997 4924 1998
rect 4890 1996 4891 1997
rect 4853 1966 4856 1996
rect 4888 1966 4891 1996
rect 4853 1965 4854 1966
rect 4820 1964 4854 1965
rect 4890 1965 4891 1966
rect 4923 1996 4924 1997
rect 4923 1966 5002 1996
rect 4923 1965 4924 1966
rect 4890 1964 4924 1965
rect 5032 1934 5062 2028
rect 5168 1997 5202 1998
rect 5168 1996 5169 1997
rect 5092 1966 5169 1996
rect 5168 1965 5169 1966
rect 5201 1996 5202 1997
rect 5238 1997 5272 1998
rect 5238 1996 5239 1997
rect 5201 1966 5204 1996
rect 5236 1966 5239 1996
rect 5201 1965 5202 1966
rect 5168 1964 5202 1965
rect 5238 1965 5239 1966
rect 5271 1996 5272 1997
rect 5271 1966 5350 1996
rect 5271 1965 5272 1966
rect 5238 1964 5272 1965
rect 5380 1934 5410 2028
rect 5516 1997 5550 1998
rect 5516 1996 5517 1997
rect 5440 1966 5517 1996
rect 5516 1965 5517 1966
rect 5549 1996 5550 1997
rect 5586 1997 5620 1998
rect 5586 1996 5587 1997
rect 5549 1966 5552 1996
rect 5584 1966 5587 1996
rect 5549 1965 5550 1966
rect 5516 1964 5550 1965
rect 5586 1965 5587 1966
rect 5619 1996 5620 1997
rect 5619 1966 5698 1996
rect 5619 1965 5620 1966
rect 5586 1964 5620 1965
rect 5728 1934 5758 2028
rect 5864 1997 5898 1998
rect 5864 1996 5865 1997
rect 5788 1966 5865 1996
rect 5864 1965 5865 1966
rect 5897 1996 5898 1997
rect 5934 1997 5968 1998
rect 5934 1996 5935 1997
rect 5897 1966 5900 1996
rect 5932 1966 5935 1996
rect 5897 1965 5898 1966
rect 5864 1964 5898 1965
rect 5934 1965 5935 1966
rect 5967 1996 5968 1997
rect 5967 1966 6046 1996
rect 5967 1965 5968 1966
rect 5934 1964 5968 1965
rect 6076 1934 6106 2028
rect 6212 1997 6246 1998
rect 6212 1996 6213 1997
rect 6136 1966 6213 1996
rect 6212 1965 6213 1966
rect 6245 1996 6246 1997
rect 6282 1997 6316 1998
rect 6282 1996 6283 1997
rect 6245 1966 6248 1996
rect 6280 1966 6283 1996
rect 6245 1965 6246 1966
rect 6212 1964 6246 1965
rect 6282 1965 6283 1966
rect 6315 1996 6316 1997
rect 6315 1966 6394 1996
rect 6315 1965 6316 1966
rect 6282 1964 6316 1965
rect 6424 1934 6454 2028
rect 6560 1997 6594 1998
rect 6560 1996 6561 1997
rect 6484 1966 6561 1996
rect 6560 1965 6561 1966
rect 6593 1996 6594 1997
rect 6630 1997 6664 1998
rect 6630 1996 6631 1997
rect 6593 1966 6596 1996
rect 6628 1966 6631 1996
rect 6593 1965 6594 1966
rect 6560 1964 6594 1965
rect 6630 1965 6631 1966
rect 6663 1996 6664 1997
rect 6663 1966 6742 1996
rect 6663 1965 6664 1966
rect 6630 1964 6664 1965
rect 6772 1934 6802 2028
rect 6908 1997 6942 1998
rect 6908 1996 6909 1997
rect 6832 1966 6909 1996
rect 6908 1965 6909 1966
rect 6941 1996 6942 1997
rect 6978 1997 7012 1998
rect 6978 1996 6979 1997
rect 6941 1966 6944 1996
rect 6976 1966 6979 1996
rect 6941 1965 6942 1966
rect 6908 1964 6942 1965
rect 6978 1965 6979 1966
rect 7011 1996 7012 1997
rect 7011 1966 7090 1996
rect 7011 1965 7012 1966
rect 6978 1964 7012 1965
rect 7120 1934 7150 2028
rect 7256 1997 7290 1998
rect 7256 1996 7257 1997
rect 7180 1966 7257 1996
rect 7256 1965 7257 1966
rect 7289 1996 7290 1997
rect 7289 1966 7292 1996
rect 7289 1965 7290 1966
rect 7256 1964 7290 1965
rect 0 1904 7307 1934
rect 18 1873 52 1874
rect 18 1872 19 1873
rect 16 1842 19 1872
rect 18 1841 19 1842
rect 51 1872 52 1873
rect 51 1842 130 1872
rect 51 1841 52 1842
rect 18 1840 52 1841
rect 160 1810 190 1904
rect 296 1873 330 1874
rect 296 1872 297 1873
rect 220 1842 297 1872
rect 296 1841 297 1842
rect 329 1872 330 1873
rect 366 1873 400 1874
rect 366 1872 367 1873
rect 329 1842 332 1872
rect 364 1842 367 1872
rect 329 1841 330 1842
rect 296 1840 330 1841
rect 366 1841 367 1842
rect 399 1872 400 1873
rect 399 1842 478 1872
rect 399 1841 400 1842
rect 366 1840 400 1841
rect 508 1810 538 1904
rect 644 1873 678 1874
rect 644 1872 645 1873
rect 568 1842 645 1872
rect 644 1841 645 1842
rect 677 1872 678 1873
rect 714 1873 748 1874
rect 714 1872 715 1873
rect 677 1842 680 1872
rect 712 1842 715 1872
rect 677 1841 678 1842
rect 644 1840 678 1841
rect 714 1841 715 1842
rect 747 1872 748 1873
rect 747 1842 826 1872
rect 747 1841 748 1842
rect 714 1840 748 1841
rect 856 1810 886 1904
rect 992 1873 1026 1874
rect 992 1872 993 1873
rect 916 1842 993 1872
rect 992 1841 993 1842
rect 1025 1872 1026 1873
rect 1062 1873 1096 1874
rect 1062 1872 1063 1873
rect 1025 1842 1028 1872
rect 1060 1842 1063 1872
rect 1025 1841 1026 1842
rect 992 1840 1026 1841
rect 1062 1841 1063 1842
rect 1095 1872 1096 1873
rect 1095 1842 1174 1872
rect 1095 1841 1096 1842
rect 1062 1840 1096 1841
rect 1204 1810 1234 1904
rect 1340 1873 1374 1874
rect 1340 1872 1341 1873
rect 1264 1842 1341 1872
rect 1340 1841 1341 1842
rect 1373 1872 1374 1873
rect 1410 1873 1444 1874
rect 1410 1872 1411 1873
rect 1373 1842 1376 1872
rect 1408 1842 1411 1872
rect 1373 1841 1374 1842
rect 1340 1840 1374 1841
rect 1410 1841 1411 1842
rect 1443 1872 1444 1873
rect 1443 1842 1522 1872
rect 1443 1841 1444 1842
rect 1410 1840 1444 1841
rect 1552 1810 1582 1904
rect 1688 1873 1722 1874
rect 1688 1872 1689 1873
rect 1612 1842 1689 1872
rect 1688 1841 1689 1842
rect 1721 1872 1722 1873
rect 1758 1873 1792 1874
rect 1758 1872 1759 1873
rect 1721 1842 1724 1872
rect 1756 1842 1759 1872
rect 1721 1841 1722 1842
rect 1688 1840 1722 1841
rect 1758 1841 1759 1842
rect 1791 1872 1792 1873
rect 1791 1842 1870 1872
rect 1791 1841 1792 1842
rect 1758 1840 1792 1841
rect 1900 1810 1930 1904
rect 2036 1873 2070 1874
rect 2036 1872 2037 1873
rect 1960 1842 2037 1872
rect 2036 1841 2037 1842
rect 2069 1872 2070 1873
rect 2106 1873 2140 1874
rect 2106 1872 2107 1873
rect 2069 1842 2072 1872
rect 2104 1842 2107 1872
rect 2069 1841 2070 1842
rect 2036 1840 2070 1841
rect 2106 1841 2107 1842
rect 2139 1872 2140 1873
rect 2139 1842 2218 1872
rect 2139 1841 2140 1842
rect 2106 1840 2140 1841
rect 2248 1810 2278 1904
rect 2384 1873 2418 1874
rect 2384 1872 2385 1873
rect 2308 1842 2385 1872
rect 2384 1841 2385 1842
rect 2417 1872 2418 1873
rect 2454 1873 2488 1874
rect 2454 1872 2455 1873
rect 2417 1842 2420 1872
rect 2452 1842 2455 1872
rect 2417 1841 2418 1842
rect 2384 1840 2418 1841
rect 2454 1841 2455 1842
rect 2487 1872 2488 1873
rect 2487 1842 2566 1872
rect 2487 1841 2488 1842
rect 2454 1840 2488 1841
rect 2596 1810 2626 1904
rect 2732 1873 2766 1874
rect 2732 1872 2733 1873
rect 2656 1842 2733 1872
rect 2732 1841 2733 1842
rect 2765 1872 2766 1873
rect 2802 1873 2836 1874
rect 2802 1872 2803 1873
rect 2765 1842 2768 1872
rect 2800 1842 2803 1872
rect 2765 1841 2766 1842
rect 2732 1840 2766 1841
rect 2802 1841 2803 1842
rect 2835 1872 2836 1873
rect 2835 1842 2914 1872
rect 2835 1841 2836 1842
rect 2802 1840 2836 1841
rect 2944 1810 2974 1904
rect 3080 1873 3114 1874
rect 3080 1872 3081 1873
rect 3004 1842 3081 1872
rect 3080 1841 3081 1842
rect 3113 1872 3114 1873
rect 3150 1873 3184 1874
rect 3150 1872 3151 1873
rect 3113 1842 3116 1872
rect 3148 1842 3151 1872
rect 3113 1841 3114 1842
rect 3080 1840 3114 1841
rect 3150 1841 3151 1842
rect 3183 1872 3184 1873
rect 3183 1842 3262 1872
rect 3183 1841 3184 1842
rect 3150 1840 3184 1841
rect 3292 1810 3322 1904
rect 3428 1873 3462 1874
rect 3428 1872 3429 1873
rect 3352 1842 3429 1872
rect 3428 1841 3429 1842
rect 3461 1872 3462 1873
rect 3498 1873 3532 1874
rect 3498 1872 3499 1873
rect 3461 1842 3464 1872
rect 3496 1842 3499 1872
rect 3461 1841 3462 1842
rect 3428 1840 3462 1841
rect 3498 1841 3499 1842
rect 3531 1872 3532 1873
rect 3531 1842 3610 1872
rect 3531 1841 3532 1842
rect 3498 1840 3532 1841
rect 3640 1810 3670 1904
rect 3776 1873 3810 1874
rect 3776 1872 3777 1873
rect 3700 1842 3777 1872
rect 3776 1841 3777 1842
rect 3809 1872 3810 1873
rect 3846 1873 3880 1874
rect 3846 1872 3847 1873
rect 3809 1842 3812 1872
rect 3844 1842 3847 1872
rect 3809 1841 3810 1842
rect 3776 1840 3810 1841
rect 3846 1841 3847 1842
rect 3879 1872 3880 1873
rect 3879 1842 3958 1872
rect 3879 1841 3880 1842
rect 3846 1840 3880 1841
rect 3988 1810 4018 1904
rect 4124 1873 4158 1874
rect 4124 1872 4125 1873
rect 4048 1842 4125 1872
rect 4124 1841 4125 1842
rect 4157 1872 4158 1873
rect 4194 1873 4228 1874
rect 4194 1872 4195 1873
rect 4157 1842 4160 1872
rect 4192 1842 4195 1872
rect 4157 1841 4158 1842
rect 4124 1840 4158 1841
rect 4194 1841 4195 1842
rect 4227 1872 4228 1873
rect 4227 1842 4306 1872
rect 4227 1841 4228 1842
rect 4194 1840 4228 1841
rect 4336 1810 4366 1904
rect 4472 1873 4506 1874
rect 4472 1872 4473 1873
rect 4396 1842 4473 1872
rect 4472 1841 4473 1842
rect 4505 1872 4506 1873
rect 4542 1873 4576 1874
rect 4542 1872 4543 1873
rect 4505 1842 4508 1872
rect 4540 1842 4543 1872
rect 4505 1841 4506 1842
rect 4472 1840 4506 1841
rect 4542 1841 4543 1842
rect 4575 1872 4576 1873
rect 4575 1842 4654 1872
rect 4575 1841 4576 1842
rect 4542 1840 4576 1841
rect 4684 1810 4714 1904
rect 4820 1873 4854 1874
rect 4820 1872 4821 1873
rect 4744 1842 4821 1872
rect 4820 1841 4821 1842
rect 4853 1872 4854 1873
rect 4890 1873 4924 1874
rect 4890 1872 4891 1873
rect 4853 1842 4856 1872
rect 4888 1842 4891 1872
rect 4853 1841 4854 1842
rect 4820 1840 4854 1841
rect 4890 1841 4891 1842
rect 4923 1872 4924 1873
rect 4923 1842 5002 1872
rect 4923 1841 4924 1842
rect 4890 1840 4924 1841
rect 5032 1810 5062 1904
rect 5168 1873 5202 1874
rect 5168 1872 5169 1873
rect 5092 1842 5169 1872
rect 5168 1841 5169 1842
rect 5201 1872 5202 1873
rect 5238 1873 5272 1874
rect 5238 1872 5239 1873
rect 5201 1842 5204 1872
rect 5236 1842 5239 1872
rect 5201 1841 5202 1842
rect 5168 1840 5202 1841
rect 5238 1841 5239 1842
rect 5271 1872 5272 1873
rect 5271 1842 5350 1872
rect 5271 1841 5272 1842
rect 5238 1840 5272 1841
rect 5380 1810 5410 1904
rect 5516 1873 5550 1874
rect 5516 1872 5517 1873
rect 5440 1842 5517 1872
rect 5516 1841 5517 1842
rect 5549 1872 5550 1873
rect 5586 1873 5620 1874
rect 5586 1872 5587 1873
rect 5549 1842 5552 1872
rect 5584 1842 5587 1872
rect 5549 1841 5550 1842
rect 5516 1840 5550 1841
rect 5586 1841 5587 1842
rect 5619 1872 5620 1873
rect 5619 1842 5698 1872
rect 5619 1841 5620 1842
rect 5586 1840 5620 1841
rect 5728 1810 5758 1904
rect 5864 1873 5898 1874
rect 5864 1872 5865 1873
rect 5788 1842 5865 1872
rect 5864 1841 5865 1842
rect 5897 1872 5898 1873
rect 5934 1873 5968 1874
rect 5934 1872 5935 1873
rect 5897 1842 5900 1872
rect 5932 1842 5935 1872
rect 5897 1841 5898 1842
rect 5864 1840 5898 1841
rect 5934 1841 5935 1842
rect 5967 1872 5968 1873
rect 5967 1842 6046 1872
rect 5967 1841 5968 1842
rect 5934 1840 5968 1841
rect 6076 1810 6106 1904
rect 6212 1873 6246 1874
rect 6212 1872 6213 1873
rect 6136 1842 6213 1872
rect 6212 1841 6213 1842
rect 6245 1872 6246 1873
rect 6282 1873 6316 1874
rect 6282 1872 6283 1873
rect 6245 1842 6248 1872
rect 6280 1842 6283 1872
rect 6245 1841 6246 1842
rect 6212 1840 6246 1841
rect 6282 1841 6283 1842
rect 6315 1872 6316 1873
rect 6315 1842 6394 1872
rect 6315 1841 6316 1842
rect 6282 1840 6316 1841
rect 6424 1810 6454 1904
rect 6560 1873 6594 1874
rect 6560 1872 6561 1873
rect 6484 1842 6561 1872
rect 6560 1841 6561 1842
rect 6593 1872 6594 1873
rect 6630 1873 6664 1874
rect 6630 1872 6631 1873
rect 6593 1842 6596 1872
rect 6628 1842 6631 1872
rect 6593 1841 6594 1842
rect 6560 1840 6594 1841
rect 6630 1841 6631 1842
rect 6663 1872 6664 1873
rect 6663 1842 6742 1872
rect 6663 1841 6664 1842
rect 6630 1840 6664 1841
rect 6772 1810 6802 1904
rect 6908 1873 6942 1874
rect 6908 1872 6909 1873
rect 6832 1842 6909 1872
rect 6908 1841 6909 1842
rect 6941 1872 6942 1873
rect 6978 1873 7012 1874
rect 6978 1872 6979 1873
rect 6941 1842 6944 1872
rect 6976 1842 6979 1872
rect 6941 1841 6942 1842
rect 6908 1840 6942 1841
rect 6978 1841 6979 1842
rect 7011 1872 7012 1873
rect 7011 1842 7090 1872
rect 7011 1841 7012 1842
rect 6978 1840 7012 1841
rect 7120 1810 7150 1904
rect 7256 1873 7290 1874
rect 7256 1872 7257 1873
rect 7180 1842 7257 1872
rect 7256 1841 7257 1842
rect 7289 1872 7290 1873
rect 7289 1842 7292 1872
rect 7289 1841 7290 1842
rect 7256 1840 7290 1841
rect 0 1780 7307 1810
rect 18 1749 52 1750
rect 18 1748 19 1749
rect 16 1718 19 1748
rect 18 1717 19 1718
rect 51 1748 52 1749
rect 51 1718 130 1748
rect 51 1717 52 1718
rect 18 1716 52 1717
rect 18 1679 52 1680
rect 18 1678 19 1679
rect 16 1648 19 1678
rect 18 1647 19 1648
rect 51 1678 52 1679
rect 51 1648 130 1678
rect 51 1647 52 1648
rect 18 1646 52 1647
rect 160 1616 190 1780
rect 296 1749 330 1750
rect 296 1748 297 1749
rect 220 1718 297 1748
rect 296 1717 297 1718
rect 329 1748 330 1749
rect 366 1749 400 1750
rect 366 1748 367 1749
rect 329 1718 332 1748
rect 364 1718 367 1748
rect 329 1717 330 1718
rect 296 1716 330 1717
rect 366 1717 367 1718
rect 399 1748 400 1749
rect 399 1718 478 1748
rect 508 1728 538 1780
rect 644 1749 678 1750
rect 644 1748 645 1749
rect 568 1718 645 1748
rect 399 1717 400 1718
rect 366 1716 400 1717
rect 644 1717 645 1718
rect 677 1748 678 1749
rect 714 1749 748 1750
rect 714 1748 715 1749
rect 677 1718 680 1748
rect 712 1718 715 1748
rect 677 1717 678 1718
rect 644 1716 678 1717
rect 714 1717 715 1718
rect 747 1748 748 1749
rect 747 1718 826 1748
rect 856 1728 886 1780
rect 992 1749 1026 1750
rect 992 1748 993 1749
rect 916 1718 993 1748
rect 747 1717 748 1718
rect 714 1716 748 1717
rect 992 1717 993 1718
rect 1025 1748 1026 1749
rect 1062 1749 1096 1750
rect 1062 1748 1063 1749
rect 1025 1718 1028 1748
rect 1060 1718 1063 1748
rect 1025 1717 1026 1718
rect 992 1716 1026 1717
rect 1062 1717 1063 1718
rect 1095 1748 1096 1749
rect 1095 1718 1174 1748
rect 1204 1728 1234 1780
rect 1340 1749 1374 1750
rect 1340 1748 1341 1749
rect 1264 1718 1341 1748
rect 1095 1717 1096 1718
rect 1062 1716 1096 1717
rect 1340 1717 1341 1718
rect 1373 1748 1374 1749
rect 1410 1749 1444 1750
rect 1410 1748 1411 1749
rect 1373 1718 1376 1748
rect 1408 1718 1411 1748
rect 1373 1717 1374 1718
rect 1340 1716 1374 1717
rect 1410 1717 1411 1718
rect 1443 1748 1444 1749
rect 1443 1718 1522 1748
rect 1443 1717 1444 1718
rect 1410 1716 1444 1717
rect 296 1679 330 1680
rect 296 1678 297 1679
rect 220 1648 297 1678
rect 296 1647 297 1648
rect 329 1678 330 1679
rect 366 1679 400 1680
rect 366 1678 367 1679
rect 329 1648 332 1678
rect 364 1648 367 1678
rect 329 1647 330 1648
rect 296 1646 330 1647
rect 366 1647 367 1648
rect 399 1678 400 1679
rect 399 1648 478 1678
rect 399 1647 400 1648
rect 366 1646 400 1647
rect 508 1616 538 1698
rect 644 1679 678 1680
rect 644 1678 645 1679
rect 568 1648 645 1678
rect 644 1647 645 1648
rect 677 1678 678 1679
rect 714 1679 748 1680
rect 714 1678 715 1679
rect 677 1648 680 1678
rect 712 1648 715 1678
rect 677 1647 678 1648
rect 644 1646 678 1647
rect 714 1647 715 1648
rect 747 1678 748 1679
rect 747 1648 826 1678
rect 747 1647 748 1648
rect 714 1646 748 1647
rect 856 1616 886 1698
rect 992 1679 1026 1680
rect 992 1678 993 1679
rect 916 1648 993 1678
rect 992 1647 993 1648
rect 1025 1678 1026 1679
rect 1062 1679 1096 1680
rect 1062 1678 1063 1679
rect 1025 1648 1028 1678
rect 1060 1648 1063 1678
rect 1025 1647 1026 1648
rect 992 1646 1026 1647
rect 1062 1647 1063 1648
rect 1095 1678 1096 1679
rect 1095 1648 1174 1678
rect 1095 1647 1096 1648
rect 1062 1646 1096 1647
rect 1204 1616 1234 1698
rect 1340 1679 1374 1680
rect 1340 1678 1341 1679
rect 1264 1648 1341 1678
rect 1340 1647 1341 1648
rect 1373 1678 1374 1679
rect 1410 1679 1444 1680
rect 1410 1678 1411 1679
rect 1373 1648 1376 1678
rect 1408 1648 1411 1678
rect 1373 1647 1374 1648
rect 1340 1646 1374 1647
rect 1410 1647 1411 1648
rect 1443 1678 1444 1679
rect 1443 1648 1522 1678
rect 1443 1647 1444 1648
rect 1410 1646 1444 1647
rect 1552 1616 1582 1780
rect 1688 1749 1722 1750
rect 1688 1748 1689 1749
rect 1612 1718 1689 1748
rect 1688 1717 1689 1718
rect 1721 1748 1722 1749
rect 1758 1749 1792 1750
rect 1758 1748 1759 1749
rect 1721 1718 1724 1748
rect 1756 1718 1759 1748
rect 1721 1717 1722 1718
rect 1688 1716 1722 1717
rect 1758 1717 1759 1718
rect 1791 1748 1792 1749
rect 1791 1718 1870 1748
rect 1791 1717 1792 1718
rect 1758 1716 1792 1717
rect 1688 1679 1722 1680
rect 1688 1678 1689 1679
rect 1612 1648 1689 1678
rect 1688 1647 1689 1648
rect 1721 1678 1722 1679
rect 1758 1679 1792 1680
rect 1758 1678 1759 1679
rect 1721 1648 1724 1678
rect 1756 1648 1759 1678
rect 1721 1647 1722 1648
rect 1688 1646 1722 1647
rect 1758 1647 1759 1648
rect 1791 1678 1792 1679
rect 1791 1648 1870 1678
rect 1791 1647 1792 1648
rect 1758 1646 1792 1647
rect 1900 1616 1930 1780
rect 2036 1749 2070 1750
rect 2036 1748 2037 1749
rect 1960 1718 2037 1748
rect 2036 1717 2037 1718
rect 2069 1748 2070 1749
rect 2106 1749 2140 1750
rect 2106 1748 2107 1749
rect 2069 1718 2072 1748
rect 2104 1718 2107 1748
rect 2069 1717 2070 1718
rect 2036 1716 2070 1717
rect 2106 1717 2107 1718
rect 2139 1748 2140 1749
rect 2139 1718 2218 1748
rect 2248 1728 2278 1780
rect 2384 1749 2418 1750
rect 2384 1748 2385 1749
rect 2308 1718 2385 1748
rect 2139 1717 2140 1718
rect 2106 1716 2140 1717
rect 2384 1717 2385 1718
rect 2417 1748 2418 1749
rect 2454 1749 2488 1750
rect 2454 1748 2455 1749
rect 2417 1718 2420 1748
rect 2452 1718 2455 1748
rect 2417 1717 2418 1718
rect 2384 1716 2418 1717
rect 2454 1717 2455 1718
rect 2487 1748 2488 1749
rect 2487 1718 2566 1748
rect 2596 1728 2626 1780
rect 2732 1749 2766 1750
rect 2732 1748 2733 1749
rect 2656 1718 2733 1748
rect 2487 1717 2488 1718
rect 2454 1716 2488 1717
rect 2732 1717 2733 1718
rect 2765 1748 2766 1749
rect 2802 1749 2836 1750
rect 2802 1748 2803 1749
rect 2765 1718 2768 1748
rect 2800 1718 2803 1748
rect 2765 1717 2766 1718
rect 2732 1716 2766 1717
rect 2802 1717 2803 1718
rect 2835 1748 2836 1749
rect 2835 1718 2914 1748
rect 2944 1728 2974 1780
rect 3080 1749 3114 1750
rect 3080 1748 3081 1749
rect 3004 1718 3081 1748
rect 2835 1717 2836 1718
rect 2802 1716 2836 1717
rect 3080 1717 3081 1718
rect 3113 1748 3114 1749
rect 3150 1749 3184 1750
rect 3150 1748 3151 1749
rect 3113 1718 3116 1748
rect 3148 1718 3151 1748
rect 3113 1717 3114 1718
rect 3080 1716 3114 1717
rect 3150 1717 3151 1718
rect 3183 1748 3184 1749
rect 3183 1718 3262 1748
rect 3183 1717 3184 1718
rect 3150 1716 3184 1717
rect 2036 1679 2070 1680
rect 2036 1678 2037 1679
rect 1960 1648 2037 1678
rect 2036 1647 2037 1648
rect 2069 1678 2070 1679
rect 2106 1679 2140 1680
rect 2106 1678 2107 1679
rect 2069 1648 2072 1678
rect 2104 1648 2107 1678
rect 2069 1647 2070 1648
rect 2036 1646 2070 1647
rect 2106 1647 2107 1648
rect 2139 1678 2140 1679
rect 2139 1648 2218 1678
rect 2139 1647 2140 1648
rect 2106 1646 2140 1647
rect 2248 1616 2278 1698
rect 2384 1679 2418 1680
rect 2384 1678 2385 1679
rect 2308 1648 2385 1678
rect 2384 1647 2385 1648
rect 2417 1678 2418 1679
rect 2454 1679 2488 1680
rect 2454 1678 2455 1679
rect 2417 1648 2420 1678
rect 2452 1648 2455 1678
rect 2417 1647 2418 1648
rect 2384 1646 2418 1647
rect 2454 1647 2455 1648
rect 2487 1678 2488 1679
rect 2487 1648 2566 1678
rect 2487 1647 2488 1648
rect 2454 1646 2488 1647
rect 2596 1616 2626 1698
rect 2732 1679 2766 1680
rect 2732 1678 2733 1679
rect 2656 1648 2733 1678
rect 2732 1647 2733 1648
rect 2765 1678 2766 1679
rect 2802 1679 2836 1680
rect 2802 1678 2803 1679
rect 2765 1648 2768 1678
rect 2800 1648 2803 1678
rect 2765 1647 2766 1648
rect 2732 1646 2766 1647
rect 2802 1647 2803 1648
rect 2835 1678 2836 1679
rect 2835 1648 2914 1678
rect 2835 1647 2836 1648
rect 2802 1646 2836 1647
rect 2944 1616 2974 1698
rect 3080 1679 3114 1680
rect 3080 1678 3081 1679
rect 3004 1648 3081 1678
rect 3080 1647 3081 1648
rect 3113 1678 3114 1679
rect 3150 1679 3184 1680
rect 3150 1678 3151 1679
rect 3113 1648 3116 1678
rect 3148 1648 3151 1678
rect 3113 1647 3114 1648
rect 3080 1646 3114 1647
rect 3150 1647 3151 1648
rect 3183 1678 3184 1679
rect 3183 1648 3262 1678
rect 3183 1647 3184 1648
rect 3150 1646 3184 1647
rect 3292 1616 3322 1780
rect 3428 1749 3462 1750
rect 3428 1748 3429 1749
rect 3352 1718 3429 1748
rect 3428 1717 3429 1718
rect 3461 1748 3462 1749
rect 3498 1749 3532 1750
rect 3498 1748 3499 1749
rect 3461 1718 3464 1748
rect 3496 1718 3499 1748
rect 3461 1717 3462 1718
rect 3428 1716 3462 1717
rect 3498 1717 3499 1718
rect 3531 1748 3532 1749
rect 3531 1718 3610 1748
rect 3531 1717 3532 1718
rect 3498 1716 3532 1717
rect 3428 1679 3462 1680
rect 3428 1678 3429 1679
rect 3352 1648 3429 1678
rect 3428 1647 3429 1648
rect 3461 1678 3462 1679
rect 3498 1679 3532 1680
rect 3498 1678 3499 1679
rect 3461 1648 3464 1678
rect 3496 1648 3499 1678
rect 3461 1647 3462 1648
rect 3428 1646 3462 1647
rect 3498 1647 3499 1648
rect 3531 1678 3532 1679
rect 3531 1648 3610 1678
rect 3531 1647 3532 1648
rect 3498 1646 3532 1647
rect 3640 1616 3670 1780
rect 3776 1749 3810 1750
rect 3776 1748 3777 1749
rect 3700 1718 3777 1748
rect 3776 1717 3777 1718
rect 3809 1748 3810 1749
rect 3846 1749 3880 1750
rect 3846 1748 3847 1749
rect 3809 1718 3812 1748
rect 3844 1718 3847 1748
rect 3809 1717 3810 1718
rect 3776 1716 3810 1717
rect 3846 1717 3847 1718
rect 3879 1748 3880 1749
rect 3879 1718 3958 1748
rect 3988 1728 4018 1780
rect 4124 1749 4158 1750
rect 4124 1748 4125 1749
rect 4048 1718 4125 1748
rect 3879 1717 3880 1718
rect 3846 1716 3880 1717
rect 4124 1717 4125 1718
rect 4157 1748 4158 1749
rect 4194 1749 4228 1750
rect 4194 1748 4195 1749
rect 4157 1718 4160 1748
rect 4192 1718 4195 1748
rect 4157 1717 4158 1718
rect 4124 1716 4158 1717
rect 4194 1717 4195 1718
rect 4227 1748 4228 1749
rect 4227 1718 4306 1748
rect 4336 1728 4366 1780
rect 4472 1749 4506 1750
rect 4472 1748 4473 1749
rect 4396 1718 4473 1748
rect 4227 1717 4228 1718
rect 4194 1716 4228 1717
rect 4472 1717 4473 1718
rect 4505 1748 4506 1749
rect 4542 1749 4576 1750
rect 4542 1748 4543 1749
rect 4505 1718 4508 1748
rect 4540 1718 4543 1748
rect 4505 1717 4506 1718
rect 4472 1716 4506 1717
rect 4542 1717 4543 1718
rect 4575 1748 4576 1749
rect 4575 1718 4654 1748
rect 4684 1728 4714 1780
rect 4820 1749 4854 1750
rect 4820 1748 4821 1749
rect 4744 1718 4821 1748
rect 4575 1717 4576 1718
rect 4542 1716 4576 1717
rect 4820 1717 4821 1718
rect 4853 1748 4854 1749
rect 4890 1749 4924 1750
rect 4890 1748 4891 1749
rect 4853 1718 4856 1748
rect 4888 1718 4891 1748
rect 4853 1717 4854 1718
rect 4820 1716 4854 1717
rect 4890 1717 4891 1718
rect 4923 1748 4924 1749
rect 4923 1718 5002 1748
rect 4923 1717 4924 1718
rect 4890 1716 4924 1717
rect 3776 1679 3810 1680
rect 3776 1678 3777 1679
rect 3700 1648 3777 1678
rect 3776 1647 3777 1648
rect 3809 1678 3810 1679
rect 3846 1679 3880 1680
rect 3846 1678 3847 1679
rect 3809 1648 3812 1678
rect 3844 1648 3847 1678
rect 3809 1647 3810 1648
rect 3776 1646 3810 1647
rect 3846 1647 3847 1648
rect 3879 1678 3880 1679
rect 3879 1648 3958 1678
rect 3879 1647 3880 1648
rect 3846 1646 3880 1647
rect 3988 1616 4018 1698
rect 4124 1679 4158 1680
rect 4124 1678 4125 1679
rect 4048 1648 4125 1678
rect 4124 1647 4125 1648
rect 4157 1678 4158 1679
rect 4194 1679 4228 1680
rect 4194 1678 4195 1679
rect 4157 1648 4160 1678
rect 4192 1648 4195 1678
rect 4157 1647 4158 1648
rect 4124 1646 4158 1647
rect 4194 1647 4195 1648
rect 4227 1678 4228 1679
rect 4227 1648 4306 1678
rect 4227 1647 4228 1648
rect 4194 1646 4228 1647
rect 4336 1616 4366 1698
rect 4472 1679 4506 1680
rect 4472 1678 4473 1679
rect 4396 1648 4473 1678
rect 4472 1647 4473 1648
rect 4505 1678 4506 1679
rect 4542 1679 4576 1680
rect 4542 1678 4543 1679
rect 4505 1648 4508 1678
rect 4540 1648 4543 1678
rect 4505 1647 4506 1648
rect 4472 1646 4506 1647
rect 4542 1647 4543 1648
rect 4575 1678 4576 1679
rect 4575 1648 4654 1678
rect 4575 1647 4576 1648
rect 4542 1646 4576 1647
rect 4684 1616 4714 1698
rect 4820 1679 4854 1680
rect 4820 1678 4821 1679
rect 4744 1648 4821 1678
rect 4820 1647 4821 1648
rect 4853 1678 4854 1679
rect 4890 1679 4924 1680
rect 4890 1678 4891 1679
rect 4853 1648 4856 1678
rect 4888 1648 4891 1678
rect 4853 1647 4854 1648
rect 4820 1646 4854 1647
rect 4890 1647 4891 1648
rect 4923 1678 4924 1679
rect 4923 1648 5002 1678
rect 4923 1647 4924 1648
rect 4890 1646 4924 1647
rect 5032 1616 5062 1780
rect 5168 1749 5202 1750
rect 5168 1748 5169 1749
rect 5092 1718 5169 1748
rect 5168 1717 5169 1718
rect 5201 1748 5202 1749
rect 5238 1749 5272 1750
rect 5238 1748 5239 1749
rect 5201 1718 5204 1748
rect 5236 1718 5239 1748
rect 5201 1717 5202 1718
rect 5168 1716 5202 1717
rect 5238 1717 5239 1718
rect 5271 1748 5272 1749
rect 5271 1718 5350 1748
rect 5271 1717 5272 1718
rect 5238 1716 5272 1717
rect 5168 1679 5202 1680
rect 5168 1678 5169 1679
rect 5092 1648 5169 1678
rect 5168 1647 5169 1648
rect 5201 1678 5202 1679
rect 5238 1679 5272 1680
rect 5238 1678 5239 1679
rect 5201 1648 5204 1678
rect 5236 1648 5239 1678
rect 5201 1647 5202 1648
rect 5168 1646 5202 1647
rect 5238 1647 5239 1648
rect 5271 1678 5272 1679
rect 5271 1648 5350 1678
rect 5271 1647 5272 1648
rect 5238 1646 5272 1647
rect 5380 1616 5410 1780
rect 5516 1749 5550 1750
rect 5516 1748 5517 1749
rect 5440 1718 5517 1748
rect 5516 1717 5517 1718
rect 5549 1748 5550 1749
rect 5586 1749 5620 1750
rect 5586 1748 5587 1749
rect 5549 1718 5552 1748
rect 5584 1718 5587 1748
rect 5549 1717 5550 1718
rect 5516 1716 5550 1717
rect 5586 1717 5587 1718
rect 5619 1748 5620 1749
rect 5619 1718 5698 1748
rect 5728 1728 5758 1780
rect 5864 1749 5898 1750
rect 5864 1748 5865 1749
rect 5788 1718 5865 1748
rect 5619 1717 5620 1718
rect 5586 1716 5620 1717
rect 5864 1717 5865 1718
rect 5897 1748 5898 1749
rect 5934 1749 5968 1750
rect 5934 1748 5935 1749
rect 5897 1718 5900 1748
rect 5932 1718 5935 1748
rect 5897 1717 5898 1718
rect 5864 1716 5898 1717
rect 5934 1717 5935 1718
rect 5967 1748 5968 1749
rect 5967 1718 6046 1748
rect 6076 1728 6106 1780
rect 6212 1749 6246 1750
rect 6212 1748 6213 1749
rect 6136 1718 6213 1748
rect 5967 1717 5968 1718
rect 5934 1716 5968 1717
rect 6212 1717 6213 1718
rect 6245 1748 6246 1749
rect 6282 1749 6316 1750
rect 6282 1748 6283 1749
rect 6245 1718 6248 1748
rect 6280 1718 6283 1748
rect 6245 1717 6246 1718
rect 6212 1716 6246 1717
rect 6282 1717 6283 1718
rect 6315 1748 6316 1749
rect 6315 1718 6394 1748
rect 6424 1728 6454 1780
rect 6560 1749 6594 1750
rect 6560 1748 6561 1749
rect 6484 1718 6561 1748
rect 6315 1717 6316 1718
rect 6282 1716 6316 1717
rect 6560 1717 6561 1718
rect 6593 1748 6594 1749
rect 6630 1749 6664 1750
rect 6630 1748 6631 1749
rect 6593 1718 6596 1748
rect 6628 1718 6631 1748
rect 6593 1717 6594 1718
rect 6560 1716 6594 1717
rect 6630 1717 6631 1718
rect 6663 1748 6664 1749
rect 6663 1718 6742 1748
rect 6663 1717 6664 1718
rect 6630 1716 6664 1717
rect 5516 1679 5550 1680
rect 5516 1678 5517 1679
rect 5440 1648 5517 1678
rect 5516 1647 5517 1648
rect 5549 1678 5550 1679
rect 5586 1679 5620 1680
rect 5586 1678 5587 1679
rect 5549 1648 5552 1678
rect 5584 1648 5587 1678
rect 5549 1647 5550 1648
rect 5516 1646 5550 1647
rect 5586 1647 5587 1648
rect 5619 1678 5620 1679
rect 5619 1648 5698 1678
rect 5619 1647 5620 1648
rect 5586 1646 5620 1647
rect 5728 1616 5758 1698
rect 5864 1679 5898 1680
rect 5864 1678 5865 1679
rect 5788 1648 5865 1678
rect 5864 1647 5865 1648
rect 5897 1678 5898 1679
rect 5934 1679 5968 1680
rect 5934 1678 5935 1679
rect 5897 1648 5900 1678
rect 5932 1648 5935 1678
rect 5897 1647 5898 1648
rect 5864 1646 5898 1647
rect 5934 1647 5935 1648
rect 5967 1678 5968 1679
rect 5967 1648 6046 1678
rect 5967 1647 5968 1648
rect 5934 1646 5968 1647
rect 6076 1616 6106 1698
rect 6212 1679 6246 1680
rect 6212 1678 6213 1679
rect 6136 1648 6213 1678
rect 6212 1647 6213 1648
rect 6245 1678 6246 1679
rect 6282 1679 6316 1680
rect 6282 1678 6283 1679
rect 6245 1648 6248 1678
rect 6280 1648 6283 1678
rect 6245 1647 6246 1648
rect 6212 1646 6246 1647
rect 6282 1647 6283 1648
rect 6315 1678 6316 1679
rect 6315 1648 6394 1678
rect 6315 1647 6316 1648
rect 6282 1646 6316 1647
rect 6424 1616 6454 1698
rect 6560 1679 6594 1680
rect 6560 1678 6561 1679
rect 6484 1648 6561 1678
rect 6560 1647 6561 1648
rect 6593 1678 6594 1679
rect 6630 1679 6664 1680
rect 6630 1678 6631 1679
rect 6593 1648 6596 1678
rect 6628 1648 6631 1678
rect 6593 1647 6594 1648
rect 6560 1646 6594 1647
rect 6630 1647 6631 1648
rect 6663 1678 6664 1679
rect 6663 1648 6742 1678
rect 6663 1647 6664 1648
rect 6630 1646 6664 1647
rect 6772 1616 6802 1780
rect 6908 1749 6942 1750
rect 6908 1748 6909 1749
rect 6832 1718 6909 1748
rect 6908 1717 6909 1718
rect 6941 1748 6942 1749
rect 6978 1749 7012 1750
rect 6978 1748 6979 1749
rect 6941 1718 6944 1748
rect 6976 1718 6979 1748
rect 6941 1717 6942 1718
rect 6908 1716 6942 1717
rect 6978 1717 6979 1718
rect 7011 1748 7012 1749
rect 7011 1718 7090 1748
rect 7011 1717 7012 1718
rect 6978 1716 7012 1717
rect 6908 1679 6942 1680
rect 6908 1678 6909 1679
rect 6832 1648 6909 1678
rect 6908 1647 6909 1648
rect 6941 1678 6942 1679
rect 6978 1679 7012 1680
rect 6978 1678 6979 1679
rect 6941 1648 6944 1678
rect 6976 1648 6979 1678
rect 6941 1647 6942 1648
rect 6908 1646 6942 1647
rect 6978 1647 6979 1648
rect 7011 1678 7012 1679
rect 7011 1648 7090 1678
rect 7011 1647 7012 1648
rect 6978 1646 7012 1647
rect 7120 1616 7150 1780
rect 7256 1749 7290 1750
rect 7256 1748 7257 1749
rect 7180 1718 7257 1748
rect 7256 1717 7257 1718
rect 7289 1748 7290 1749
rect 7289 1718 7292 1748
rect 7289 1717 7290 1718
rect 7256 1716 7290 1717
rect 7256 1679 7290 1680
rect 7256 1678 7257 1679
rect 7180 1648 7257 1678
rect 7256 1647 7257 1648
rect 7289 1678 7290 1679
rect 7289 1648 7292 1678
rect 7289 1647 7290 1648
rect 7256 1646 7290 1647
rect 0 1586 318 1616
rect 348 1586 1392 1616
rect 1422 1586 2058 1616
rect 2088 1586 3132 1616
rect 3162 1586 3798 1616
rect 3828 1586 4872 1616
rect 4902 1586 5538 1616
rect 5568 1586 6612 1616
rect 6642 1586 7278 1616
rect 18 1555 52 1556
rect 18 1554 19 1555
rect 16 1524 19 1554
rect 18 1523 19 1524
rect 51 1554 52 1555
rect 51 1524 130 1554
rect 51 1523 52 1524
rect 18 1522 52 1523
rect 160 1492 190 1586
rect 296 1555 330 1556
rect 296 1554 297 1555
rect 220 1524 297 1554
rect 296 1523 297 1524
rect 329 1554 330 1555
rect 366 1555 400 1556
rect 366 1554 367 1555
rect 329 1524 332 1554
rect 364 1524 367 1554
rect 329 1523 330 1524
rect 296 1522 330 1523
rect 366 1523 367 1524
rect 399 1554 400 1555
rect 399 1524 478 1554
rect 399 1523 400 1524
rect 366 1522 400 1523
rect 508 1492 538 1586
rect 644 1555 678 1556
rect 644 1554 645 1555
rect 568 1524 645 1554
rect 644 1523 645 1524
rect 677 1554 678 1555
rect 714 1555 748 1556
rect 714 1554 715 1555
rect 677 1524 680 1554
rect 712 1524 715 1554
rect 677 1523 678 1524
rect 644 1522 678 1523
rect 714 1523 715 1524
rect 747 1554 748 1555
rect 747 1524 826 1554
rect 747 1523 748 1524
rect 714 1522 748 1523
rect 856 1492 886 1586
rect 992 1555 1026 1556
rect 992 1554 993 1555
rect 916 1524 993 1554
rect 992 1523 993 1524
rect 1025 1554 1026 1555
rect 1062 1555 1096 1556
rect 1062 1554 1063 1555
rect 1025 1524 1028 1554
rect 1060 1524 1063 1554
rect 1025 1523 1026 1524
rect 992 1522 1026 1523
rect 1062 1523 1063 1524
rect 1095 1554 1096 1555
rect 1095 1524 1174 1554
rect 1095 1523 1096 1524
rect 1062 1522 1096 1523
rect 1204 1492 1234 1586
rect 1340 1555 1374 1556
rect 1340 1554 1341 1555
rect 1264 1524 1341 1554
rect 1340 1523 1341 1524
rect 1373 1554 1374 1555
rect 1410 1555 1444 1556
rect 1410 1554 1411 1555
rect 1373 1524 1376 1554
rect 1408 1524 1411 1554
rect 1373 1523 1374 1524
rect 1340 1522 1374 1523
rect 1410 1523 1411 1524
rect 1443 1554 1444 1555
rect 1443 1524 1522 1554
rect 1443 1523 1444 1524
rect 1410 1522 1444 1523
rect 1552 1492 1582 1586
rect 1688 1555 1722 1556
rect 1688 1554 1689 1555
rect 1612 1524 1689 1554
rect 1688 1523 1689 1524
rect 1721 1554 1722 1555
rect 1758 1555 1792 1556
rect 1758 1554 1759 1555
rect 1721 1524 1724 1554
rect 1756 1524 1759 1554
rect 1721 1523 1722 1524
rect 1688 1522 1722 1523
rect 1758 1523 1759 1524
rect 1791 1554 1792 1555
rect 1791 1524 1870 1554
rect 1791 1523 1792 1524
rect 1758 1522 1792 1523
rect 1900 1492 1930 1586
rect 2036 1555 2070 1556
rect 2036 1554 2037 1555
rect 1960 1524 2037 1554
rect 2036 1523 2037 1524
rect 2069 1554 2070 1555
rect 2106 1555 2140 1556
rect 2106 1554 2107 1555
rect 2069 1524 2072 1554
rect 2104 1524 2107 1554
rect 2069 1523 2070 1524
rect 2036 1522 2070 1523
rect 2106 1523 2107 1524
rect 2139 1554 2140 1555
rect 2139 1524 2218 1554
rect 2139 1523 2140 1524
rect 2106 1522 2140 1523
rect 2248 1492 2278 1586
rect 2384 1555 2418 1556
rect 2384 1554 2385 1555
rect 2308 1524 2385 1554
rect 2384 1523 2385 1524
rect 2417 1554 2418 1555
rect 2454 1555 2488 1556
rect 2454 1554 2455 1555
rect 2417 1524 2420 1554
rect 2452 1524 2455 1554
rect 2417 1523 2418 1524
rect 2384 1522 2418 1523
rect 2454 1523 2455 1524
rect 2487 1554 2488 1555
rect 2487 1524 2566 1554
rect 2487 1523 2488 1524
rect 2454 1522 2488 1523
rect 2596 1492 2626 1586
rect 2732 1555 2766 1556
rect 2732 1554 2733 1555
rect 2656 1524 2733 1554
rect 2732 1523 2733 1524
rect 2765 1554 2766 1555
rect 2802 1555 2836 1556
rect 2802 1554 2803 1555
rect 2765 1524 2768 1554
rect 2800 1524 2803 1554
rect 2765 1523 2766 1524
rect 2732 1522 2766 1523
rect 2802 1523 2803 1524
rect 2835 1554 2836 1555
rect 2835 1524 2914 1554
rect 2835 1523 2836 1524
rect 2802 1522 2836 1523
rect 2944 1492 2974 1586
rect 3080 1555 3114 1556
rect 3080 1554 3081 1555
rect 3004 1524 3081 1554
rect 3080 1523 3081 1524
rect 3113 1554 3114 1555
rect 3150 1555 3184 1556
rect 3150 1554 3151 1555
rect 3113 1524 3116 1554
rect 3148 1524 3151 1554
rect 3113 1523 3114 1524
rect 3080 1522 3114 1523
rect 3150 1523 3151 1524
rect 3183 1554 3184 1555
rect 3183 1524 3262 1554
rect 3183 1523 3184 1524
rect 3150 1522 3184 1523
rect 3292 1492 3322 1586
rect 3428 1555 3462 1556
rect 3428 1554 3429 1555
rect 3352 1524 3429 1554
rect 3428 1523 3429 1524
rect 3461 1554 3462 1555
rect 3498 1555 3532 1556
rect 3498 1554 3499 1555
rect 3461 1524 3464 1554
rect 3496 1524 3499 1554
rect 3461 1523 3462 1524
rect 3428 1522 3462 1523
rect 3498 1523 3499 1524
rect 3531 1554 3532 1555
rect 3531 1524 3610 1554
rect 3531 1523 3532 1524
rect 3498 1522 3532 1523
rect 3640 1492 3670 1586
rect 3776 1555 3810 1556
rect 3776 1554 3777 1555
rect 3700 1524 3777 1554
rect 3776 1523 3777 1524
rect 3809 1554 3810 1555
rect 3846 1555 3880 1556
rect 3846 1554 3847 1555
rect 3809 1524 3812 1554
rect 3844 1524 3847 1554
rect 3809 1523 3810 1524
rect 3776 1522 3810 1523
rect 3846 1523 3847 1524
rect 3879 1554 3880 1555
rect 3879 1524 3958 1554
rect 3879 1523 3880 1524
rect 3846 1522 3880 1523
rect 3988 1492 4018 1586
rect 4124 1555 4158 1556
rect 4124 1554 4125 1555
rect 4048 1524 4125 1554
rect 4124 1523 4125 1524
rect 4157 1554 4158 1555
rect 4194 1555 4228 1556
rect 4194 1554 4195 1555
rect 4157 1524 4160 1554
rect 4192 1524 4195 1554
rect 4157 1523 4158 1524
rect 4124 1522 4158 1523
rect 4194 1523 4195 1524
rect 4227 1554 4228 1555
rect 4227 1524 4306 1554
rect 4227 1523 4228 1524
rect 4194 1522 4228 1523
rect 4336 1492 4366 1586
rect 4472 1555 4506 1556
rect 4472 1554 4473 1555
rect 4396 1524 4473 1554
rect 4472 1523 4473 1524
rect 4505 1554 4506 1555
rect 4542 1555 4576 1556
rect 4542 1554 4543 1555
rect 4505 1524 4508 1554
rect 4540 1524 4543 1554
rect 4505 1523 4506 1524
rect 4472 1522 4506 1523
rect 4542 1523 4543 1524
rect 4575 1554 4576 1555
rect 4575 1524 4654 1554
rect 4575 1523 4576 1524
rect 4542 1522 4576 1523
rect 4684 1492 4714 1586
rect 4820 1555 4854 1556
rect 4820 1554 4821 1555
rect 4744 1524 4821 1554
rect 4820 1523 4821 1524
rect 4853 1554 4854 1555
rect 4890 1555 4924 1556
rect 4890 1554 4891 1555
rect 4853 1524 4856 1554
rect 4888 1524 4891 1554
rect 4853 1523 4854 1524
rect 4820 1522 4854 1523
rect 4890 1523 4891 1524
rect 4923 1554 4924 1555
rect 4923 1524 5002 1554
rect 4923 1523 4924 1524
rect 4890 1522 4924 1523
rect 5032 1492 5062 1586
rect 5168 1555 5202 1556
rect 5168 1554 5169 1555
rect 5092 1524 5169 1554
rect 5168 1523 5169 1524
rect 5201 1554 5202 1555
rect 5238 1555 5272 1556
rect 5238 1554 5239 1555
rect 5201 1524 5204 1554
rect 5236 1524 5239 1554
rect 5201 1523 5202 1524
rect 5168 1522 5202 1523
rect 5238 1523 5239 1524
rect 5271 1554 5272 1555
rect 5271 1524 5350 1554
rect 5271 1523 5272 1524
rect 5238 1522 5272 1523
rect 5380 1492 5410 1586
rect 5516 1555 5550 1556
rect 5516 1554 5517 1555
rect 5440 1524 5517 1554
rect 5516 1523 5517 1524
rect 5549 1554 5550 1555
rect 5586 1555 5620 1556
rect 5586 1554 5587 1555
rect 5549 1524 5552 1554
rect 5584 1524 5587 1554
rect 5549 1523 5550 1524
rect 5516 1522 5550 1523
rect 5586 1523 5587 1524
rect 5619 1554 5620 1555
rect 5619 1524 5698 1554
rect 5619 1523 5620 1524
rect 5586 1522 5620 1523
rect 5728 1492 5758 1586
rect 5864 1555 5898 1556
rect 5864 1554 5865 1555
rect 5788 1524 5865 1554
rect 5864 1523 5865 1524
rect 5897 1554 5898 1555
rect 5934 1555 5968 1556
rect 5934 1554 5935 1555
rect 5897 1524 5900 1554
rect 5932 1524 5935 1554
rect 5897 1523 5898 1524
rect 5864 1522 5898 1523
rect 5934 1523 5935 1524
rect 5967 1554 5968 1555
rect 5967 1524 6046 1554
rect 5967 1523 5968 1524
rect 5934 1522 5968 1523
rect 6076 1492 6106 1586
rect 6212 1555 6246 1556
rect 6212 1554 6213 1555
rect 6136 1524 6213 1554
rect 6212 1523 6213 1524
rect 6245 1554 6246 1555
rect 6282 1555 6316 1556
rect 6282 1554 6283 1555
rect 6245 1524 6248 1554
rect 6280 1524 6283 1554
rect 6245 1523 6246 1524
rect 6212 1522 6246 1523
rect 6282 1523 6283 1524
rect 6315 1554 6316 1555
rect 6315 1524 6394 1554
rect 6315 1523 6316 1524
rect 6282 1522 6316 1523
rect 6424 1492 6454 1586
rect 6560 1555 6594 1556
rect 6560 1554 6561 1555
rect 6484 1524 6561 1554
rect 6560 1523 6561 1524
rect 6593 1554 6594 1555
rect 6630 1555 6664 1556
rect 6630 1554 6631 1555
rect 6593 1524 6596 1554
rect 6628 1524 6631 1554
rect 6593 1523 6594 1524
rect 6560 1522 6594 1523
rect 6630 1523 6631 1524
rect 6663 1554 6664 1555
rect 6663 1524 6742 1554
rect 6663 1523 6664 1524
rect 6630 1522 6664 1523
rect 6772 1492 6802 1586
rect 6908 1555 6942 1556
rect 6908 1554 6909 1555
rect 6832 1524 6909 1554
rect 6908 1523 6909 1524
rect 6941 1554 6942 1555
rect 6978 1555 7012 1556
rect 6978 1554 6979 1555
rect 6941 1524 6944 1554
rect 6976 1524 6979 1554
rect 6941 1523 6942 1524
rect 6908 1522 6942 1523
rect 6978 1523 6979 1524
rect 7011 1554 7012 1555
rect 7011 1524 7090 1554
rect 7011 1523 7012 1524
rect 6978 1522 7012 1523
rect 7120 1492 7150 1586
rect 7256 1555 7290 1556
rect 7256 1554 7257 1555
rect 7180 1524 7257 1554
rect 7256 1523 7257 1524
rect 7289 1554 7290 1555
rect 7289 1524 7292 1554
rect 7289 1523 7290 1524
rect 7256 1522 7290 1523
rect 0 1462 318 1492
rect 348 1462 1392 1492
rect 1422 1462 2058 1492
rect 2088 1462 3132 1492
rect 3162 1462 3798 1492
rect 3828 1462 4872 1492
rect 4902 1462 5538 1492
rect 5568 1462 6612 1492
rect 6642 1462 7278 1492
rect 18 1431 52 1432
rect 18 1430 19 1431
rect 16 1400 19 1430
rect 18 1399 19 1400
rect 51 1430 52 1431
rect 51 1400 130 1430
rect 51 1399 52 1400
rect 18 1398 52 1399
rect 160 1368 190 1462
rect 296 1431 330 1432
rect 296 1430 297 1431
rect 220 1400 297 1430
rect 296 1399 297 1400
rect 329 1430 330 1431
rect 366 1431 400 1432
rect 366 1430 367 1431
rect 329 1400 332 1430
rect 364 1400 367 1430
rect 329 1399 330 1400
rect 296 1398 330 1399
rect 366 1399 367 1400
rect 399 1430 400 1431
rect 399 1400 478 1430
rect 399 1399 400 1400
rect 366 1398 400 1399
rect 508 1368 538 1462
rect 644 1431 678 1432
rect 644 1430 645 1431
rect 568 1400 645 1430
rect 644 1399 645 1400
rect 677 1430 678 1431
rect 714 1431 748 1432
rect 714 1430 715 1431
rect 677 1400 680 1430
rect 712 1400 715 1430
rect 677 1399 678 1400
rect 644 1398 678 1399
rect 714 1399 715 1400
rect 747 1430 748 1431
rect 747 1400 826 1430
rect 747 1399 748 1400
rect 714 1398 748 1399
rect 856 1368 886 1462
rect 992 1431 1026 1432
rect 992 1430 993 1431
rect 916 1400 993 1430
rect 992 1399 993 1400
rect 1025 1430 1026 1431
rect 1062 1431 1096 1432
rect 1062 1430 1063 1431
rect 1025 1400 1028 1430
rect 1060 1400 1063 1430
rect 1025 1399 1026 1400
rect 992 1398 1026 1399
rect 1062 1399 1063 1400
rect 1095 1430 1096 1431
rect 1095 1400 1174 1430
rect 1095 1399 1096 1400
rect 1062 1398 1096 1399
rect 1204 1368 1234 1462
rect 1340 1431 1374 1432
rect 1340 1430 1341 1431
rect 1264 1400 1341 1430
rect 1340 1399 1341 1400
rect 1373 1430 1374 1431
rect 1410 1431 1444 1432
rect 1410 1430 1411 1431
rect 1373 1400 1376 1430
rect 1408 1400 1411 1430
rect 1373 1399 1374 1400
rect 1340 1398 1374 1399
rect 1410 1399 1411 1400
rect 1443 1430 1444 1431
rect 1443 1400 1522 1430
rect 1443 1399 1444 1400
rect 1410 1398 1444 1399
rect 1552 1368 1582 1462
rect 1688 1431 1722 1432
rect 1688 1430 1689 1431
rect 1612 1400 1689 1430
rect 1688 1399 1689 1400
rect 1721 1430 1722 1431
rect 1758 1431 1792 1432
rect 1758 1430 1759 1431
rect 1721 1400 1724 1430
rect 1756 1400 1759 1430
rect 1721 1399 1722 1400
rect 1688 1398 1722 1399
rect 1758 1399 1759 1400
rect 1791 1430 1792 1431
rect 1791 1400 1870 1430
rect 1791 1399 1792 1400
rect 1758 1398 1792 1399
rect 1900 1368 1930 1462
rect 2036 1431 2070 1432
rect 2036 1430 2037 1431
rect 1960 1400 2037 1430
rect 2036 1399 2037 1400
rect 2069 1430 2070 1431
rect 2106 1431 2140 1432
rect 2106 1430 2107 1431
rect 2069 1400 2072 1430
rect 2104 1400 2107 1430
rect 2069 1399 2070 1400
rect 2036 1398 2070 1399
rect 2106 1399 2107 1400
rect 2139 1430 2140 1431
rect 2139 1400 2218 1430
rect 2139 1399 2140 1400
rect 2106 1398 2140 1399
rect 2248 1368 2278 1462
rect 2384 1431 2418 1432
rect 2384 1430 2385 1431
rect 2308 1400 2385 1430
rect 2384 1399 2385 1400
rect 2417 1430 2418 1431
rect 2454 1431 2488 1432
rect 2454 1430 2455 1431
rect 2417 1400 2420 1430
rect 2452 1400 2455 1430
rect 2417 1399 2418 1400
rect 2384 1398 2418 1399
rect 2454 1399 2455 1400
rect 2487 1430 2488 1431
rect 2487 1400 2566 1430
rect 2487 1399 2488 1400
rect 2454 1398 2488 1399
rect 2596 1368 2626 1462
rect 2732 1431 2766 1432
rect 2732 1430 2733 1431
rect 2656 1400 2733 1430
rect 2732 1399 2733 1400
rect 2765 1430 2766 1431
rect 2802 1431 2836 1432
rect 2802 1430 2803 1431
rect 2765 1400 2768 1430
rect 2800 1400 2803 1430
rect 2765 1399 2766 1400
rect 2732 1398 2766 1399
rect 2802 1399 2803 1400
rect 2835 1430 2836 1431
rect 2835 1400 2914 1430
rect 2835 1399 2836 1400
rect 2802 1398 2836 1399
rect 2944 1368 2974 1462
rect 3080 1431 3114 1432
rect 3080 1430 3081 1431
rect 3004 1400 3081 1430
rect 3080 1399 3081 1400
rect 3113 1430 3114 1431
rect 3150 1431 3184 1432
rect 3150 1430 3151 1431
rect 3113 1400 3116 1430
rect 3148 1400 3151 1430
rect 3113 1399 3114 1400
rect 3080 1398 3114 1399
rect 3150 1399 3151 1400
rect 3183 1430 3184 1431
rect 3183 1400 3262 1430
rect 3183 1399 3184 1400
rect 3150 1398 3184 1399
rect 3292 1368 3322 1462
rect 3428 1431 3462 1432
rect 3428 1430 3429 1431
rect 3352 1400 3429 1430
rect 3428 1399 3429 1400
rect 3461 1430 3462 1431
rect 3498 1431 3532 1432
rect 3498 1430 3499 1431
rect 3461 1400 3464 1430
rect 3496 1400 3499 1430
rect 3461 1399 3462 1400
rect 3428 1398 3462 1399
rect 3498 1399 3499 1400
rect 3531 1430 3532 1431
rect 3531 1400 3610 1430
rect 3531 1399 3532 1400
rect 3498 1398 3532 1399
rect 3640 1368 3670 1462
rect 3776 1431 3810 1432
rect 3776 1430 3777 1431
rect 3700 1400 3777 1430
rect 3776 1399 3777 1400
rect 3809 1430 3810 1431
rect 3846 1431 3880 1432
rect 3846 1430 3847 1431
rect 3809 1400 3812 1430
rect 3844 1400 3847 1430
rect 3809 1399 3810 1400
rect 3776 1398 3810 1399
rect 3846 1399 3847 1400
rect 3879 1430 3880 1431
rect 3879 1400 3958 1430
rect 3879 1399 3880 1400
rect 3846 1398 3880 1399
rect 3988 1368 4018 1462
rect 4124 1431 4158 1432
rect 4124 1430 4125 1431
rect 4048 1400 4125 1430
rect 4124 1399 4125 1400
rect 4157 1430 4158 1431
rect 4194 1431 4228 1432
rect 4194 1430 4195 1431
rect 4157 1400 4160 1430
rect 4192 1400 4195 1430
rect 4157 1399 4158 1400
rect 4124 1398 4158 1399
rect 4194 1399 4195 1400
rect 4227 1430 4228 1431
rect 4227 1400 4306 1430
rect 4227 1399 4228 1400
rect 4194 1398 4228 1399
rect 4336 1368 4366 1462
rect 4472 1431 4506 1432
rect 4472 1430 4473 1431
rect 4396 1400 4473 1430
rect 4472 1399 4473 1400
rect 4505 1430 4506 1431
rect 4542 1431 4576 1432
rect 4542 1430 4543 1431
rect 4505 1400 4508 1430
rect 4540 1400 4543 1430
rect 4505 1399 4506 1400
rect 4472 1398 4506 1399
rect 4542 1399 4543 1400
rect 4575 1430 4576 1431
rect 4575 1400 4654 1430
rect 4575 1399 4576 1400
rect 4542 1398 4576 1399
rect 4684 1368 4714 1462
rect 4820 1431 4854 1432
rect 4820 1430 4821 1431
rect 4744 1400 4821 1430
rect 4820 1399 4821 1400
rect 4853 1430 4854 1431
rect 4890 1431 4924 1432
rect 4890 1430 4891 1431
rect 4853 1400 4856 1430
rect 4888 1400 4891 1430
rect 4853 1399 4854 1400
rect 4820 1398 4854 1399
rect 4890 1399 4891 1400
rect 4923 1430 4924 1431
rect 4923 1400 5002 1430
rect 4923 1399 4924 1400
rect 4890 1398 4924 1399
rect 5032 1368 5062 1462
rect 5168 1431 5202 1432
rect 5168 1430 5169 1431
rect 5092 1400 5169 1430
rect 5168 1399 5169 1400
rect 5201 1430 5202 1431
rect 5238 1431 5272 1432
rect 5238 1430 5239 1431
rect 5201 1400 5204 1430
rect 5236 1400 5239 1430
rect 5201 1399 5202 1400
rect 5168 1398 5202 1399
rect 5238 1399 5239 1400
rect 5271 1430 5272 1431
rect 5271 1400 5350 1430
rect 5271 1399 5272 1400
rect 5238 1398 5272 1399
rect 5380 1368 5410 1462
rect 5516 1431 5550 1432
rect 5516 1430 5517 1431
rect 5440 1400 5517 1430
rect 5516 1399 5517 1400
rect 5549 1430 5550 1431
rect 5586 1431 5620 1432
rect 5586 1430 5587 1431
rect 5549 1400 5552 1430
rect 5584 1400 5587 1430
rect 5549 1399 5550 1400
rect 5516 1398 5550 1399
rect 5586 1399 5587 1400
rect 5619 1430 5620 1431
rect 5619 1400 5698 1430
rect 5619 1399 5620 1400
rect 5586 1398 5620 1399
rect 5728 1368 5758 1462
rect 5864 1431 5898 1432
rect 5864 1430 5865 1431
rect 5788 1400 5865 1430
rect 5864 1399 5865 1400
rect 5897 1430 5898 1431
rect 5934 1431 5968 1432
rect 5934 1430 5935 1431
rect 5897 1400 5900 1430
rect 5932 1400 5935 1430
rect 5897 1399 5898 1400
rect 5864 1398 5898 1399
rect 5934 1399 5935 1400
rect 5967 1430 5968 1431
rect 5967 1400 6046 1430
rect 5967 1399 5968 1400
rect 5934 1398 5968 1399
rect 6076 1368 6106 1462
rect 6212 1431 6246 1432
rect 6212 1430 6213 1431
rect 6136 1400 6213 1430
rect 6212 1399 6213 1400
rect 6245 1430 6246 1431
rect 6282 1431 6316 1432
rect 6282 1430 6283 1431
rect 6245 1400 6248 1430
rect 6280 1400 6283 1430
rect 6245 1399 6246 1400
rect 6212 1398 6246 1399
rect 6282 1399 6283 1400
rect 6315 1430 6316 1431
rect 6315 1400 6394 1430
rect 6315 1399 6316 1400
rect 6282 1398 6316 1399
rect 6424 1368 6454 1462
rect 6560 1431 6594 1432
rect 6560 1430 6561 1431
rect 6484 1400 6561 1430
rect 6560 1399 6561 1400
rect 6593 1430 6594 1431
rect 6630 1431 6664 1432
rect 6630 1430 6631 1431
rect 6593 1400 6596 1430
rect 6628 1400 6631 1430
rect 6593 1399 6594 1400
rect 6560 1398 6594 1399
rect 6630 1399 6631 1400
rect 6663 1430 6664 1431
rect 6663 1400 6742 1430
rect 6663 1399 6664 1400
rect 6630 1398 6664 1399
rect 6772 1368 6802 1462
rect 6908 1431 6942 1432
rect 6908 1430 6909 1431
rect 6832 1400 6909 1430
rect 6908 1399 6909 1400
rect 6941 1430 6942 1431
rect 6978 1431 7012 1432
rect 6978 1430 6979 1431
rect 6941 1400 6944 1430
rect 6976 1400 6979 1430
rect 6941 1399 6942 1400
rect 6908 1398 6942 1399
rect 6978 1399 6979 1400
rect 7011 1430 7012 1431
rect 7011 1400 7090 1430
rect 7011 1399 7012 1400
rect 6978 1398 7012 1399
rect 7120 1368 7150 1462
rect 7256 1431 7290 1432
rect 7256 1430 7257 1431
rect 7180 1400 7257 1430
rect 7256 1399 7257 1400
rect 7289 1430 7290 1431
rect 7289 1400 7292 1430
rect 7289 1399 7290 1400
rect 7256 1398 7290 1399
rect 0 1338 318 1368
rect 348 1338 1392 1368
rect 1422 1338 2058 1368
rect 2088 1338 3132 1368
rect 3162 1338 3798 1368
rect 3828 1338 4872 1368
rect 4902 1338 5538 1368
rect 5568 1338 6612 1368
rect 6642 1338 7278 1368
rect 18 1307 52 1308
rect 18 1306 19 1307
rect 16 1276 19 1306
rect 18 1275 19 1276
rect 51 1306 52 1307
rect 51 1276 130 1306
rect 51 1275 52 1276
rect 18 1274 52 1275
rect 160 1244 190 1338
rect 296 1307 330 1308
rect 296 1306 297 1307
rect 220 1276 297 1306
rect 296 1275 297 1276
rect 329 1306 330 1307
rect 366 1307 400 1308
rect 366 1306 367 1307
rect 329 1276 332 1306
rect 364 1276 367 1306
rect 329 1275 330 1276
rect 296 1274 330 1275
rect 366 1275 367 1276
rect 399 1306 400 1307
rect 399 1276 478 1306
rect 399 1275 400 1276
rect 366 1274 400 1275
rect 508 1244 538 1338
rect 644 1307 678 1308
rect 644 1306 645 1307
rect 568 1276 645 1306
rect 644 1275 645 1276
rect 677 1306 678 1307
rect 714 1307 748 1308
rect 714 1306 715 1307
rect 677 1276 680 1306
rect 712 1276 715 1306
rect 677 1275 678 1276
rect 644 1274 678 1275
rect 714 1275 715 1276
rect 747 1306 748 1307
rect 747 1276 826 1306
rect 747 1275 748 1276
rect 714 1274 748 1275
rect 856 1244 886 1338
rect 992 1307 1026 1308
rect 992 1306 993 1307
rect 916 1276 993 1306
rect 992 1275 993 1276
rect 1025 1306 1026 1307
rect 1062 1307 1096 1308
rect 1062 1306 1063 1307
rect 1025 1276 1028 1306
rect 1060 1276 1063 1306
rect 1025 1275 1026 1276
rect 992 1274 1026 1275
rect 1062 1275 1063 1276
rect 1095 1306 1096 1307
rect 1095 1276 1174 1306
rect 1095 1275 1096 1276
rect 1062 1274 1096 1275
rect 1204 1244 1234 1338
rect 1340 1307 1374 1308
rect 1340 1306 1341 1307
rect 1264 1276 1341 1306
rect 1340 1275 1341 1276
rect 1373 1306 1374 1307
rect 1410 1307 1444 1308
rect 1410 1306 1411 1307
rect 1373 1276 1376 1306
rect 1408 1276 1411 1306
rect 1373 1275 1374 1276
rect 1340 1274 1374 1275
rect 1410 1275 1411 1276
rect 1443 1306 1444 1307
rect 1443 1276 1522 1306
rect 1443 1275 1444 1276
rect 1410 1274 1444 1275
rect 1552 1244 1582 1338
rect 1688 1307 1722 1308
rect 1688 1306 1689 1307
rect 1612 1276 1689 1306
rect 1688 1275 1689 1276
rect 1721 1306 1722 1307
rect 1758 1307 1792 1308
rect 1758 1306 1759 1307
rect 1721 1276 1724 1306
rect 1756 1276 1759 1306
rect 1721 1275 1722 1276
rect 1688 1274 1722 1275
rect 1758 1275 1759 1276
rect 1791 1306 1792 1307
rect 1791 1276 1870 1306
rect 1791 1275 1792 1276
rect 1758 1274 1792 1275
rect 1900 1244 1930 1338
rect 2036 1307 2070 1308
rect 2036 1306 2037 1307
rect 1960 1276 2037 1306
rect 2036 1275 2037 1276
rect 2069 1306 2070 1307
rect 2106 1307 2140 1308
rect 2106 1306 2107 1307
rect 2069 1276 2072 1306
rect 2104 1276 2107 1306
rect 2069 1275 2070 1276
rect 2036 1274 2070 1275
rect 2106 1275 2107 1276
rect 2139 1306 2140 1307
rect 2139 1276 2218 1306
rect 2139 1275 2140 1276
rect 2106 1274 2140 1275
rect 2248 1244 2278 1338
rect 2384 1307 2418 1308
rect 2384 1306 2385 1307
rect 2308 1276 2385 1306
rect 2384 1275 2385 1276
rect 2417 1306 2418 1307
rect 2454 1307 2488 1308
rect 2454 1306 2455 1307
rect 2417 1276 2420 1306
rect 2452 1276 2455 1306
rect 2417 1275 2418 1276
rect 2384 1274 2418 1275
rect 2454 1275 2455 1276
rect 2487 1306 2488 1307
rect 2487 1276 2566 1306
rect 2487 1275 2488 1276
rect 2454 1274 2488 1275
rect 2596 1244 2626 1338
rect 2732 1307 2766 1308
rect 2732 1306 2733 1307
rect 2656 1276 2733 1306
rect 2732 1275 2733 1276
rect 2765 1306 2766 1307
rect 2802 1307 2836 1308
rect 2802 1306 2803 1307
rect 2765 1276 2768 1306
rect 2800 1276 2803 1306
rect 2765 1275 2766 1276
rect 2732 1274 2766 1275
rect 2802 1275 2803 1276
rect 2835 1306 2836 1307
rect 2835 1276 2914 1306
rect 2835 1275 2836 1276
rect 2802 1274 2836 1275
rect 2944 1244 2974 1338
rect 3080 1307 3114 1308
rect 3080 1306 3081 1307
rect 3004 1276 3081 1306
rect 3080 1275 3081 1276
rect 3113 1306 3114 1307
rect 3150 1307 3184 1308
rect 3150 1306 3151 1307
rect 3113 1276 3116 1306
rect 3148 1276 3151 1306
rect 3113 1275 3114 1276
rect 3080 1274 3114 1275
rect 3150 1275 3151 1276
rect 3183 1306 3184 1307
rect 3183 1276 3262 1306
rect 3183 1275 3184 1276
rect 3150 1274 3184 1275
rect 3292 1244 3322 1338
rect 3428 1307 3462 1308
rect 3428 1306 3429 1307
rect 3352 1276 3429 1306
rect 3428 1275 3429 1276
rect 3461 1306 3462 1307
rect 3498 1307 3532 1308
rect 3498 1306 3499 1307
rect 3461 1276 3464 1306
rect 3496 1276 3499 1306
rect 3461 1275 3462 1276
rect 3428 1274 3462 1275
rect 3498 1275 3499 1276
rect 3531 1306 3532 1307
rect 3531 1276 3610 1306
rect 3531 1275 3532 1276
rect 3498 1274 3532 1275
rect 3640 1244 3670 1338
rect 3776 1307 3810 1308
rect 3776 1306 3777 1307
rect 3700 1276 3777 1306
rect 3776 1275 3777 1276
rect 3809 1306 3810 1307
rect 3846 1307 3880 1308
rect 3846 1306 3847 1307
rect 3809 1276 3812 1306
rect 3844 1276 3847 1306
rect 3809 1275 3810 1276
rect 3776 1274 3810 1275
rect 3846 1275 3847 1276
rect 3879 1306 3880 1307
rect 3879 1276 3958 1306
rect 3879 1275 3880 1276
rect 3846 1274 3880 1275
rect 3988 1244 4018 1338
rect 4124 1307 4158 1308
rect 4124 1306 4125 1307
rect 4048 1276 4125 1306
rect 4124 1275 4125 1276
rect 4157 1306 4158 1307
rect 4194 1307 4228 1308
rect 4194 1306 4195 1307
rect 4157 1276 4160 1306
rect 4192 1276 4195 1306
rect 4157 1275 4158 1276
rect 4124 1274 4158 1275
rect 4194 1275 4195 1276
rect 4227 1306 4228 1307
rect 4227 1276 4306 1306
rect 4227 1275 4228 1276
rect 4194 1274 4228 1275
rect 4336 1244 4366 1338
rect 4472 1307 4506 1308
rect 4472 1306 4473 1307
rect 4396 1276 4473 1306
rect 4472 1275 4473 1276
rect 4505 1306 4506 1307
rect 4542 1307 4576 1308
rect 4542 1306 4543 1307
rect 4505 1276 4508 1306
rect 4540 1276 4543 1306
rect 4505 1275 4506 1276
rect 4472 1274 4506 1275
rect 4542 1275 4543 1276
rect 4575 1306 4576 1307
rect 4575 1276 4654 1306
rect 4575 1275 4576 1276
rect 4542 1274 4576 1275
rect 4684 1244 4714 1338
rect 4820 1307 4854 1308
rect 4820 1306 4821 1307
rect 4744 1276 4821 1306
rect 4820 1275 4821 1276
rect 4853 1306 4854 1307
rect 4890 1307 4924 1308
rect 4890 1306 4891 1307
rect 4853 1276 4856 1306
rect 4888 1276 4891 1306
rect 4853 1275 4854 1276
rect 4820 1274 4854 1275
rect 4890 1275 4891 1276
rect 4923 1306 4924 1307
rect 4923 1276 5002 1306
rect 4923 1275 4924 1276
rect 4890 1274 4924 1275
rect 5032 1244 5062 1338
rect 5168 1307 5202 1308
rect 5168 1306 5169 1307
rect 5092 1276 5169 1306
rect 5168 1275 5169 1276
rect 5201 1306 5202 1307
rect 5238 1307 5272 1308
rect 5238 1306 5239 1307
rect 5201 1276 5204 1306
rect 5236 1276 5239 1306
rect 5201 1275 5202 1276
rect 5168 1274 5202 1275
rect 5238 1275 5239 1276
rect 5271 1306 5272 1307
rect 5271 1276 5350 1306
rect 5271 1275 5272 1276
rect 5238 1274 5272 1275
rect 5380 1244 5410 1338
rect 5516 1307 5550 1308
rect 5516 1306 5517 1307
rect 5440 1276 5517 1306
rect 5516 1275 5517 1276
rect 5549 1306 5550 1307
rect 5586 1307 5620 1308
rect 5586 1306 5587 1307
rect 5549 1276 5552 1306
rect 5584 1276 5587 1306
rect 5549 1275 5550 1276
rect 5516 1274 5550 1275
rect 5586 1275 5587 1276
rect 5619 1306 5620 1307
rect 5619 1276 5698 1306
rect 5619 1275 5620 1276
rect 5586 1274 5620 1275
rect 5728 1244 5758 1338
rect 5864 1307 5898 1308
rect 5864 1306 5865 1307
rect 5788 1276 5865 1306
rect 5864 1275 5865 1276
rect 5897 1306 5898 1307
rect 5934 1307 5968 1308
rect 5934 1306 5935 1307
rect 5897 1276 5900 1306
rect 5932 1276 5935 1306
rect 5897 1275 5898 1276
rect 5864 1274 5898 1275
rect 5934 1275 5935 1276
rect 5967 1306 5968 1307
rect 5967 1276 6046 1306
rect 5967 1275 5968 1276
rect 5934 1274 5968 1275
rect 6076 1244 6106 1338
rect 6212 1307 6246 1308
rect 6212 1306 6213 1307
rect 6136 1276 6213 1306
rect 6212 1275 6213 1276
rect 6245 1306 6246 1307
rect 6282 1307 6316 1308
rect 6282 1306 6283 1307
rect 6245 1276 6248 1306
rect 6280 1276 6283 1306
rect 6245 1275 6246 1276
rect 6212 1274 6246 1275
rect 6282 1275 6283 1276
rect 6315 1306 6316 1307
rect 6315 1276 6394 1306
rect 6315 1275 6316 1276
rect 6282 1274 6316 1275
rect 6424 1244 6454 1338
rect 6560 1307 6594 1308
rect 6560 1306 6561 1307
rect 6484 1276 6561 1306
rect 6560 1275 6561 1276
rect 6593 1306 6594 1307
rect 6630 1307 6664 1308
rect 6630 1306 6631 1307
rect 6593 1276 6596 1306
rect 6628 1276 6631 1306
rect 6593 1275 6594 1276
rect 6560 1274 6594 1275
rect 6630 1275 6631 1276
rect 6663 1306 6664 1307
rect 6663 1276 6742 1306
rect 6663 1275 6664 1276
rect 6630 1274 6664 1275
rect 6772 1244 6802 1338
rect 6908 1307 6942 1308
rect 6908 1306 6909 1307
rect 6832 1276 6909 1306
rect 6908 1275 6909 1276
rect 6941 1306 6942 1307
rect 6978 1307 7012 1308
rect 6978 1306 6979 1307
rect 6941 1276 6944 1306
rect 6976 1276 6979 1306
rect 6941 1275 6942 1276
rect 6908 1274 6942 1275
rect 6978 1275 6979 1276
rect 7011 1306 7012 1307
rect 7011 1276 7090 1306
rect 7011 1275 7012 1276
rect 6978 1274 7012 1275
rect 7120 1244 7150 1338
rect 7256 1307 7290 1308
rect 7256 1306 7257 1307
rect 7180 1276 7257 1306
rect 7256 1275 7257 1276
rect 7289 1306 7290 1307
rect 7289 1276 7292 1306
rect 7289 1275 7290 1276
rect 7256 1274 7290 1275
rect 0 1214 318 1244
rect 348 1214 1392 1244
rect 1422 1214 2058 1244
rect 2088 1214 3132 1244
rect 3162 1214 3798 1244
rect 3828 1214 4872 1244
rect 4902 1214 5538 1244
rect 5568 1214 6612 1244
rect 6642 1214 7278 1244
rect 18 1183 52 1184
rect 18 1182 19 1183
rect 16 1152 19 1182
rect 18 1151 19 1152
rect 51 1182 52 1183
rect 51 1152 130 1182
rect 51 1151 52 1152
rect 18 1150 52 1151
rect 18 1113 52 1114
rect 18 1112 19 1113
rect 16 1082 19 1112
rect 18 1081 19 1082
rect 51 1112 52 1113
rect 51 1082 130 1112
rect 51 1081 52 1082
rect 18 1080 52 1081
rect 160 1050 190 1214
rect 296 1183 330 1184
rect 296 1182 297 1183
rect 220 1152 297 1182
rect 296 1151 297 1152
rect 329 1182 330 1183
rect 366 1183 400 1184
rect 366 1182 367 1183
rect 329 1152 332 1182
rect 364 1152 367 1182
rect 329 1151 330 1152
rect 296 1150 330 1151
rect 366 1151 367 1152
rect 399 1182 400 1183
rect 399 1152 478 1182
rect 399 1151 400 1152
rect 366 1150 400 1151
rect 296 1113 330 1114
rect 296 1112 297 1113
rect 220 1082 297 1112
rect 296 1081 297 1082
rect 329 1112 330 1113
rect 366 1113 400 1114
rect 366 1112 367 1113
rect 329 1082 332 1112
rect 364 1082 367 1112
rect 329 1081 330 1082
rect 296 1080 330 1081
rect 366 1081 367 1082
rect 399 1112 400 1113
rect 399 1082 478 1112
rect 399 1081 400 1082
rect 366 1080 400 1081
rect 508 1050 538 1214
rect 644 1183 678 1184
rect 644 1182 645 1183
rect 568 1152 645 1182
rect 644 1151 645 1152
rect 677 1182 678 1183
rect 714 1183 748 1184
rect 714 1182 715 1183
rect 677 1152 680 1182
rect 712 1152 715 1182
rect 677 1151 678 1152
rect 644 1150 678 1151
rect 714 1151 715 1152
rect 747 1182 748 1183
rect 747 1152 826 1182
rect 747 1151 748 1152
rect 714 1150 748 1151
rect 644 1113 678 1114
rect 644 1112 645 1113
rect 568 1082 645 1112
rect 644 1081 645 1082
rect 677 1112 678 1113
rect 714 1113 748 1114
rect 714 1112 715 1113
rect 677 1082 680 1112
rect 712 1082 715 1112
rect 677 1081 678 1082
rect 644 1080 678 1081
rect 714 1081 715 1082
rect 747 1112 748 1113
rect 747 1082 826 1112
rect 747 1081 748 1082
rect 714 1080 748 1081
rect 856 1050 886 1214
rect 992 1183 1026 1184
rect 992 1182 993 1183
rect 916 1152 993 1182
rect 992 1151 993 1152
rect 1025 1182 1026 1183
rect 1062 1183 1096 1184
rect 1062 1182 1063 1183
rect 1025 1152 1028 1182
rect 1060 1152 1063 1182
rect 1025 1151 1026 1152
rect 992 1150 1026 1151
rect 1062 1151 1063 1152
rect 1095 1182 1096 1183
rect 1095 1152 1174 1182
rect 1095 1151 1096 1152
rect 1062 1150 1096 1151
rect 992 1113 1026 1114
rect 992 1112 993 1113
rect 916 1082 993 1112
rect 992 1081 993 1082
rect 1025 1112 1026 1113
rect 1062 1113 1096 1114
rect 1062 1112 1063 1113
rect 1025 1082 1028 1112
rect 1060 1082 1063 1112
rect 1025 1081 1026 1082
rect 992 1080 1026 1081
rect 1062 1081 1063 1082
rect 1095 1112 1096 1113
rect 1095 1082 1174 1112
rect 1095 1081 1096 1082
rect 1062 1080 1096 1081
rect 1204 1050 1234 1214
rect 1340 1183 1374 1184
rect 1340 1182 1341 1183
rect 1264 1152 1341 1182
rect 1340 1151 1341 1152
rect 1373 1182 1374 1183
rect 1410 1183 1444 1184
rect 1410 1182 1411 1183
rect 1373 1152 1376 1182
rect 1408 1152 1411 1182
rect 1373 1151 1374 1152
rect 1340 1150 1374 1151
rect 1410 1151 1411 1152
rect 1443 1182 1444 1183
rect 1443 1152 1522 1182
rect 1443 1151 1444 1152
rect 1410 1150 1444 1151
rect 1340 1113 1374 1114
rect 1340 1112 1341 1113
rect 1264 1082 1341 1112
rect 1340 1081 1341 1082
rect 1373 1112 1374 1113
rect 1410 1113 1444 1114
rect 1410 1112 1411 1113
rect 1373 1082 1376 1112
rect 1408 1082 1411 1112
rect 1373 1081 1374 1082
rect 1340 1080 1374 1081
rect 1410 1081 1411 1082
rect 1443 1112 1444 1113
rect 1443 1082 1522 1112
rect 1443 1081 1444 1082
rect 1410 1080 1444 1081
rect 1552 1050 1582 1214
rect 1688 1183 1722 1184
rect 1688 1182 1689 1183
rect 1612 1152 1689 1182
rect 1688 1151 1689 1152
rect 1721 1182 1722 1183
rect 1758 1183 1792 1184
rect 1758 1182 1759 1183
rect 1721 1152 1724 1182
rect 1756 1152 1759 1182
rect 1721 1151 1722 1152
rect 1688 1150 1722 1151
rect 1758 1151 1759 1152
rect 1791 1182 1792 1183
rect 1791 1152 1870 1182
rect 1791 1151 1792 1152
rect 1758 1150 1792 1151
rect 1688 1113 1722 1114
rect 1688 1112 1689 1113
rect 1612 1082 1689 1112
rect 1688 1081 1689 1082
rect 1721 1112 1722 1113
rect 1758 1113 1792 1114
rect 1758 1112 1759 1113
rect 1721 1082 1724 1112
rect 1756 1082 1759 1112
rect 1721 1081 1722 1082
rect 1688 1080 1722 1081
rect 1758 1081 1759 1082
rect 1791 1112 1792 1113
rect 1791 1082 1870 1112
rect 1791 1081 1792 1082
rect 1758 1080 1792 1081
rect 1900 1050 1930 1214
rect 2036 1183 2070 1184
rect 2036 1182 2037 1183
rect 1960 1152 2037 1182
rect 2036 1151 2037 1152
rect 2069 1182 2070 1183
rect 2106 1183 2140 1184
rect 2106 1182 2107 1183
rect 2069 1152 2072 1182
rect 2104 1152 2107 1182
rect 2069 1151 2070 1152
rect 2036 1150 2070 1151
rect 2106 1151 2107 1152
rect 2139 1182 2140 1183
rect 2139 1152 2218 1182
rect 2139 1151 2140 1152
rect 2106 1150 2140 1151
rect 2036 1113 2070 1114
rect 2036 1112 2037 1113
rect 1960 1082 2037 1112
rect 2036 1081 2037 1082
rect 2069 1112 2070 1113
rect 2106 1113 2140 1114
rect 2106 1112 2107 1113
rect 2069 1082 2072 1112
rect 2104 1082 2107 1112
rect 2069 1081 2070 1082
rect 2036 1080 2070 1081
rect 2106 1081 2107 1082
rect 2139 1112 2140 1113
rect 2139 1082 2218 1112
rect 2139 1081 2140 1082
rect 2106 1080 2140 1081
rect 2248 1050 2278 1214
rect 2384 1183 2418 1184
rect 2384 1182 2385 1183
rect 2308 1152 2385 1182
rect 2384 1151 2385 1152
rect 2417 1182 2418 1183
rect 2454 1183 2488 1184
rect 2454 1182 2455 1183
rect 2417 1152 2420 1182
rect 2452 1152 2455 1182
rect 2417 1151 2418 1152
rect 2384 1150 2418 1151
rect 2454 1151 2455 1152
rect 2487 1182 2488 1183
rect 2487 1152 2566 1182
rect 2487 1151 2488 1152
rect 2454 1150 2488 1151
rect 2384 1113 2418 1114
rect 2384 1112 2385 1113
rect 2308 1082 2385 1112
rect 2384 1081 2385 1082
rect 2417 1112 2418 1113
rect 2454 1113 2488 1114
rect 2454 1112 2455 1113
rect 2417 1082 2420 1112
rect 2452 1082 2455 1112
rect 2417 1081 2418 1082
rect 2384 1080 2418 1081
rect 2454 1081 2455 1082
rect 2487 1112 2488 1113
rect 2487 1082 2566 1112
rect 2487 1081 2488 1082
rect 2454 1080 2488 1081
rect 2596 1050 2626 1214
rect 2732 1183 2766 1184
rect 2732 1182 2733 1183
rect 2656 1152 2733 1182
rect 2732 1151 2733 1152
rect 2765 1182 2766 1183
rect 2802 1183 2836 1184
rect 2802 1182 2803 1183
rect 2765 1152 2768 1182
rect 2800 1152 2803 1182
rect 2765 1151 2766 1152
rect 2732 1150 2766 1151
rect 2802 1151 2803 1152
rect 2835 1182 2836 1183
rect 2835 1152 2914 1182
rect 2835 1151 2836 1152
rect 2802 1150 2836 1151
rect 2732 1113 2766 1114
rect 2732 1112 2733 1113
rect 2656 1082 2733 1112
rect 2732 1081 2733 1082
rect 2765 1112 2766 1113
rect 2802 1113 2836 1114
rect 2802 1112 2803 1113
rect 2765 1082 2768 1112
rect 2800 1082 2803 1112
rect 2765 1081 2766 1082
rect 2732 1080 2766 1081
rect 2802 1081 2803 1082
rect 2835 1112 2836 1113
rect 2835 1082 2914 1112
rect 2835 1081 2836 1082
rect 2802 1080 2836 1081
rect 2944 1050 2974 1214
rect 3080 1183 3114 1184
rect 3080 1182 3081 1183
rect 3004 1152 3081 1182
rect 3080 1151 3081 1152
rect 3113 1182 3114 1183
rect 3150 1183 3184 1184
rect 3150 1182 3151 1183
rect 3113 1152 3116 1182
rect 3148 1152 3151 1182
rect 3113 1151 3114 1152
rect 3080 1150 3114 1151
rect 3150 1151 3151 1152
rect 3183 1182 3184 1183
rect 3183 1152 3262 1182
rect 3183 1151 3184 1152
rect 3150 1150 3184 1151
rect 3080 1113 3114 1114
rect 3080 1112 3081 1113
rect 3004 1082 3081 1112
rect 3080 1081 3081 1082
rect 3113 1112 3114 1113
rect 3150 1113 3184 1114
rect 3150 1112 3151 1113
rect 3113 1082 3116 1112
rect 3148 1082 3151 1112
rect 3113 1081 3114 1082
rect 3080 1080 3114 1081
rect 3150 1081 3151 1082
rect 3183 1112 3184 1113
rect 3183 1082 3262 1112
rect 3183 1081 3184 1082
rect 3150 1080 3184 1081
rect 3292 1050 3322 1214
rect 3428 1183 3462 1184
rect 3428 1182 3429 1183
rect 3352 1152 3429 1182
rect 3428 1151 3429 1152
rect 3461 1182 3462 1183
rect 3498 1183 3532 1184
rect 3498 1182 3499 1183
rect 3461 1152 3464 1182
rect 3496 1152 3499 1182
rect 3461 1151 3462 1152
rect 3428 1150 3462 1151
rect 3498 1151 3499 1152
rect 3531 1182 3532 1183
rect 3531 1152 3610 1182
rect 3531 1151 3532 1152
rect 3498 1150 3532 1151
rect 3428 1113 3462 1114
rect 3428 1112 3429 1113
rect 3352 1082 3429 1112
rect 3428 1081 3429 1082
rect 3461 1112 3462 1113
rect 3498 1113 3532 1114
rect 3498 1112 3499 1113
rect 3461 1082 3464 1112
rect 3496 1082 3499 1112
rect 3461 1081 3462 1082
rect 3428 1080 3462 1081
rect 3498 1081 3499 1082
rect 3531 1112 3532 1113
rect 3531 1082 3610 1112
rect 3531 1081 3532 1082
rect 3498 1080 3532 1081
rect 3640 1050 3670 1214
rect 3776 1183 3810 1184
rect 3776 1182 3777 1183
rect 3700 1152 3777 1182
rect 3776 1151 3777 1152
rect 3809 1182 3810 1183
rect 3846 1183 3880 1184
rect 3846 1182 3847 1183
rect 3809 1152 3812 1182
rect 3844 1152 3847 1182
rect 3809 1151 3810 1152
rect 3776 1150 3810 1151
rect 3846 1151 3847 1152
rect 3879 1182 3880 1183
rect 3879 1152 3958 1182
rect 3879 1151 3880 1152
rect 3846 1150 3880 1151
rect 3776 1113 3810 1114
rect 3776 1112 3777 1113
rect 3700 1082 3777 1112
rect 3776 1081 3777 1082
rect 3809 1112 3810 1113
rect 3846 1113 3880 1114
rect 3846 1112 3847 1113
rect 3809 1082 3812 1112
rect 3844 1082 3847 1112
rect 3809 1081 3810 1082
rect 3776 1080 3810 1081
rect 3846 1081 3847 1082
rect 3879 1112 3880 1113
rect 3879 1082 3958 1112
rect 3879 1081 3880 1082
rect 3846 1080 3880 1081
rect 3988 1050 4018 1214
rect 4124 1183 4158 1184
rect 4124 1182 4125 1183
rect 4048 1152 4125 1182
rect 4124 1151 4125 1152
rect 4157 1182 4158 1183
rect 4194 1183 4228 1184
rect 4194 1182 4195 1183
rect 4157 1152 4160 1182
rect 4192 1152 4195 1182
rect 4157 1151 4158 1152
rect 4124 1150 4158 1151
rect 4194 1151 4195 1152
rect 4227 1182 4228 1183
rect 4227 1152 4306 1182
rect 4227 1151 4228 1152
rect 4194 1150 4228 1151
rect 4124 1113 4158 1114
rect 4124 1112 4125 1113
rect 4048 1082 4125 1112
rect 4124 1081 4125 1082
rect 4157 1112 4158 1113
rect 4194 1113 4228 1114
rect 4194 1112 4195 1113
rect 4157 1082 4160 1112
rect 4192 1082 4195 1112
rect 4157 1081 4158 1082
rect 4124 1080 4158 1081
rect 4194 1081 4195 1082
rect 4227 1112 4228 1113
rect 4227 1082 4306 1112
rect 4227 1081 4228 1082
rect 4194 1080 4228 1081
rect 4336 1050 4366 1214
rect 4472 1183 4506 1184
rect 4472 1182 4473 1183
rect 4396 1152 4473 1182
rect 4472 1151 4473 1152
rect 4505 1182 4506 1183
rect 4542 1183 4576 1184
rect 4542 1182 4543 1183
rect 4505 1152 4508 1182
rect 4540 1152 4543 1182
rect 4505 1151 4506 1152
rect 4472 1150 4506 1151
rect 4542 1151 4543 1152
rect 4575 1182 4576 1183
rect 4575 1152 4654 1182
rect 4575 1151 4576 1152
rect 4542 1150 4576 1151
rect 4472 1113 4506 1114
rect 4472 1112 4473 1113
rect 4396 1082 4473 1112
rect 4472 1081 4473 1082
rect 4505 1112 4506 1113
rect 4542 1113 4576 1114
rect 4542 1112 4543 1113
rect 4505 1082 4508 1112
rect 4540 1082 4543 1112
rect 4505 1081 4506 1082
rect 4472 1080 4506 1081
rect 4542 1081 4543 1082
rect 4575 1112 4576 1113
rect 4575 1082 4654 1112
rect 4575 1081 4576 1082
rect 4542 1080 4576 1081
rect 4684 1050 4714 1214
rect 4820 1183 4854 1184
rect 4820 1182 4821 1183
rect 4744 1152 4821 1182
rect 4820 1151 4821 1152
rect 4853 1182 4854 1183
rect 4890 1183 4924 1184
rect 4890 1182 4891 1183
rect 4853 1152 4856 1182
rect 4888 1152 4891 1182
rect 4853 1151 4854 1152
rect 4820 1150 4854 1151
rect 4890 1151 4891 1152
rect 4923 1182 4924 1183
rect 4923 1152 5002 1182
rect 4923 1151 4924 1152
rect 4890 1150 4924 1151
rect 4820 1113 4854 1114
rect 4820 1112 4821 1113
rect 4744 1082 4821 1112
rect 4820 1081 4821 1082
rect 4853 1112 4854 1113
rect 4890 1113 4924 1114
rect 4890 1112 4891 1113
rect 4853 1082 4856 1112
rect 4888 1082 4891 1112
rect 4853 1081 4854 1082
rect 4820 1080 4854 1081
rect 4890 1081 4891 1082
rect 4923 1112 4924 1113
rect 4923 1082 5002 1112
rect 4923 1081 4924 1082
rect 4890 1080 4924 1081
rect 5032 1050 5062 1214
rect 5168 1183 5202 1184
rect 5168 1182 5169 1183
rect 5092 1152 5169 1182
rect 5168 1151 5169 1152
rect 5201 1182 5202 1183
rect 5238 1183 5272 1184
rect 5238 1182 5239 1183
rect 5201 1152 5204 1182
rect 5236 1152 5239 1182
rect 5201 1151 5202 1152
rect 5168 1150 5202 1151
rect 5238 1151 5239 1152
rect 5271 1182 5272 1183
rect 5271 1152 5350 1182
rect 5271 1151 5272 1152
rect 5238 1150 5272 1151
rect 5168 1113 5202 1114
rect 5168 1112 5169 1113
rect 5092 1082 5169 1112
rect 5168 1081 5169 1082
rect 5201 1112 5202 1113
rect 5238 1113 5272 1114
rect 5238 1112 5239 1113
rect 5201 1082 5204 1112
rect 5236 1082 5239 1112
rect 5201 1081 5202 1082
rect 5168 1080 5202 1081
rect 5238 1081 5239 1082
rect 5271 1112 5272 1113
rect 5271 1082 5350 1112
rect 5271 1081 5272 1082
rect 5238 1080 5272 1081
rect 5380 1050 5410 1214
rect 5516 1183 5550 1184
rect 5516 1182 5517 1183
rect 5440 1152 5517 1182
rect 5516 1151 5517 1152
rect 5549 1182 5550 1183
rect 5586 1183 5620 1184
rect 5586 1182 5587 1183
rect 5549 1152 5552 1182
rect 5584 1152 5587 1182
rect 5549 1151 5550 1152
rect 5516 1150 5550 1151
rect 5586 1151 5587 1152
rect 5619 1182 5620 1183
rect 5619 1152 5698 1182
rect 5619 1151 5620 1152
rect 5586 1150 5620 1151
rect 5516 1113 5550 1114
rect 5516 1112 5517 1113
rect 5440 1082 5517 1112
rect 5516 1081 5517 1082
rect 5549 1112 5550 1113
rect 5586 1113 5620 1114
rect 5586 1112 5587 1113
rect 5549 1082 5552 1112
rect 5584 1082 5587 1112
rect 5549 1081 5550 1082
rect 5516 1080 5550 1081
rect 5586 1081 5587 1082
rect 5619 1112 5620 1113
rect 5619 1082 5698 1112
rect 5619 1081 5620 1082
rect 5586 1080 5620 1081
rect 5728 1050 5758 1214
rect 5864 1183 5898 1184
rect 5864 1182 5865 1183
rect 5788 1152 5865 1182
rect 5864 1151 5865 1152
rect 5897 1182 5898 1183
rect 5934 1183 5968 1184
rect 5934 1182 5935 1183
rect 5897 1152 5900 1182
rect 5932 1152 5935 1182
rect 5897 1151 5898 1152
rect 5864 1150 5898 1151
rect 5934 1151 5935 1152
rect 5967 1182 5968 1183
rect 5967 1152 6046 1182
rect 5967 1151 5968 1152
rect 5934 1150 5968 1151
rect 5864 1113 5898 1114
rect 5864 1112 5865 1113
rect 5788 1082 5865 1112
rect 5864 1081 5865 1082
rect 5897 1112 5898 1113
rect 5934 1113 5968 1114
rect 5934 1112 5935 1113
rect 5897 1082 5900 1112
rect 5932 1082 5935 1112
rect 5897 1081 5898 1082
rect 5864 1080 5898 1081
rect 5934 1081 5935 1082
rect 5967 1112 5968 1113
rect 5967 1082 6046 1112
rect 5967 1081 5968 1082
rect 5934 1080 5968 1081
rect 6076 1050 6106 1214
rect 6212 1183 6246 1184
rect 6212 1182 6213 1183
rect 6136 1152 6213 1182
rect 6212 1151 6213 1152
rect 6245 1182 6246 1183
rect 6282 1183 6316 1184
rect 6282 1182 6283 1183
rect 6245 1152 6248 1182
rect 6280 1152 6283 1182
rect 6245 1151 6246 1152
rect 6212 1150 6246 1151
rect 6282 1151 6283 1152
rect 6315 1182 6316 1183
rect 6315 1152 6394 1182
rect 6315 1151 6316 1152
rect 6282 1150 6316 1151
rect 6212 1113 6246 1114
rect 6212 1112 6213 1113
rect 6136 1082 6213 1112
rect 6212 1081 6213 1082
rect 6245 1112 6246 1113
rect 6282 1113 6316 1114
rect 6282 1112 6283 1113
rect 6245 1082 6248 1112
rect 6280 1082 6283 1112
rect 6245 1081 6246 1082
rect 6212 1080 6246 1081
rect 6282 1081 6283 1082
rect 6315 1112 6316 1113
rect 6315 1082 6394 1112
rect 6315 1081 6316 1082
rect 6282 1080 6316 1081
rect 6424 1050 6454 1214
rect 6560 1183 6594 1184
rect 6560 1182 6561 1183
rect 6484 1152 6561 1182
rect 6560 1151 6561 1152
rect 6593 1182 6594 1183
rect 6630 1183 6664 1184
rect 6630 1182 6631 1183
rect 6593 1152 6596 1182
rect 6628 1152 6631 1182
rect 6593 1151 6594 1152
rect 6560 1150 6594 1151
rect 6630 1151 6631 1152
rect 6663 1182 6664 1183
rect 6663 1152 6742 1182
rect 6663 1151 6664 1152
rect 6630 1150 6664 1151
rect 6560 1113 6594 1114
rect 6560 1112 6561 1113
rect 6484 1082 6561 1112
rect 6560 1081 6561 1082
rect 6593 1112 6594 1113
rect 6630 1113 6664 1114
rect 6630 1112 6631 1113
rect 6593 1082 6596 1112
rect 6628 1082 6631 1112
rect 6593 1081 6594 1082
rect 6560 1080 6594 1081
rect 6630 1081 6631 1082
rect 6663 1112 6664 1113
rect 6663 1082 6742 1112
rect 6663 1081 6664 1082
rect 6630 1080 6664 1081
rect 6772 1051 6802 1214
rect 6908 1183 6942 1184
rect 6908 1182 6909 1183
rect 6832 1152 6909 1182
rect 6908 1151 6909 1152
rect 6941 1182 6942 1183
rect 6978 1183 7012 1184
rect 6978 1182 6979 1183
rect 6941 1152 6944 1182
rect 6976 1152 6979 1182
rect 6941 1151 6942 1152
rect 6908 1150 6942 1151
rect 6978 1151 6979 1152
rect 7011 1182 7012 1183
rect 7011 1152 7090 1182
rect 7011 1151 7012 1152
rect 6978 1150 7012 1151
rect 6908 1113 6942 1114
rect 6908 1112 6909 1113
rect 6832 1082 6909 1112
rect 6908 1081 6909 1082
rect 6941 1112 6942 1113
rect 6978 1113 7012 1114
rect 6978 1112 6979 1113
rect 6941 1082 6944 1112
rect 6976 1082 6979 1112
rect 6941 1081 6942 1082
rect 6908 1080 6942 1081
rect 6978 1081 6979 1082
rect 7011 1112 7012 1113
rect 7011 1082 7090 1112
rect 7011 1081 7012 1082
rect 6978 1080 7012 1081
rect 6756 1050 6865 1051
rect 7120 1050 7150 1214
rect 7256 1183 7290 1184
rect 7256 1182 7257 1183
rect 7180 1152 7257 1182
rect 7256 1151 7257 1152
rect 7289 1182 7290 1183
rect 7289 1152 7292 1182
rect 7289 1151 7290 1152
rect 7256 1150 7290 1151
rect 7256 1113 7290 1114
rect 7256 1112 7257 1113
rect 7180 1082 7257 1112
rect 7256 1081 7257 1082
rect 7289 1112 7290 1113
rect 7289 1082 7292 1112
rect 7289 1081 7290 1082
rect 7256 1080 7290 1081
rect 0 1020 318 1050
rect 348 1020 1392 1050
rect 1422 1020 2058 1050
rect 2088 1020 3131 1050
rect 3161 1020 3480 1050
rect 3510 1020 3798 1050
rect 3828 1020 4872 1050
rect 4902 1020 5220 1050
rect 5250 1020 5538 1050
rect 5568 1020 6612 1050
rect 6642 1020 6960 1050
rect 6990 1020 7278 1050
rect 18 989 52 990
rect 18 988 19 989
rect 16 958 19 988
rect 18 957 19 958
rect 51 988 52 989
rect 51 958 130 988
rect 51 957 52 958
rect 18 956 52 957
rect 160 926 190 1020
rect 296 989 330 990
rect 296 988 297 989
rect 220 958 297 988
rect 296 957 297 958
rect 329 988 330 989
rect 366 989 400 990
rect 366 988 367 989
rect 329 958 332 988
rect 364 958 367 988
rect 329 957 330 958
rect 296 956 330 957
rect 366 957 367 958
rect 399 988 400 989
rect 399 958 478 988
rect 399 957 400 958
rect 366 956 400 957
rect 508 926 538 1020
rect 644 989 678 990
rect 644 988 645 989
rect 568 958 645 988
rect 644 957 645 958
rect 677 988 678 989
rect 714 989 748 990
rect 714 988 715 989
rect 677 958 680 988
rect 712 958 715 988
rect 677 957 678 958
rect 644 956 678 957
rect 714 957 715 958
rect 747 988 748 989
rect 747 958 826 988
rect 747 957 748 958
rect 714 956 748 957
rect 856 926 886 1020
rect 992 989 1026 990
rect 992 988 993 989
rect 916 958 993 988
rect 992 957 993 958
rect 1025 988 1026 989
rect 1062 989 1096 990
rect 1062 988 1063 989
rect 1025 958 1028 988
rect 1060 958 1063 988
rect 1025 957 1026 958
rect 992 956 1026 957
rect 1062 957 1063 958
rect 1095 988 1096 989
rect 1095 958 1174 988
rect 1095 957 1096 958
rect 1062 956 1096 957
rect 1204 926 1234 1020
rect 1340 989 1374 990
rect 1340 988 1341 989
rect 1264 958 1341 988
rect 1340 957 1341 958
rect 1373 988 1374 989
rect 1410 989 1444 990
rect 1410 988 1411 989
rect 1373 958 1376 988
rect 1408 958 1411 988
rect 1373 957 1374 958
rect 1340 956 1374 957
rect 1410 957 1411 958
rect 1443 988 1444 989
rect 1443 958 1522 988
rect 1443 957 1444 958
rect 1410 956 1444 957
rect 1552 926 1582 1020
rect 1688 989 1722 990
rect 1688 988 1689 989
rect 1612 958 1689 988
rect 1688 957 1689 958
rect 1721 988 1722 989
rect 1758 989 1792 990
rect 1758 988 1759 989
rect 1721 958 1724 988
rect 1756 958 1759 988
rect 1721 957 1722 958
rect 1688 956 1722 957
rect 1758 957 1759 958
rect 1791 988 1792 989
rect 1791 958 1870 988
rect 1791 957 1792 958
rect 1758 956 1792 957
rect 1900 926 1930 1020
rect 2036 989 2070 990
rect 2036 988 2037 989
rect 1960 958 2037 988
rect 2036 957 2037 958
rect 2069 988 2070 989
rect 2106 989 2140 990
rect 2106 988 2107 989
rect 2069 958 2072 988
rect 2104 958 2107 988
rect 2069 957 2070 958
rect 2036 956 2070 957
rect 2106 957 2107 958
rect 2139 988 2140 989
rect 2139 958 2218 988
rect 2139 957 2140 958
rect 2106 956 2140 957
rect 2248 926 2278 1020
rect 2384 989 2418 990
rect 2384 988 2385 989
rect 2308 958 2385 988
rect 2384 957 2385 958
rect 2417 988 2418 989
rect 2454 989 2488 990
rect 2454 988 2455 989
rect 2417 958 2420 988
rect 2452 958 2455 988
rect 2417 957 2418 958
rect 2384 956 2418 957
rect 2454 957 2455 958
rect 2487 988 2488 989
rect 2487 958 2566 988
rect 2487 957 2488 958
rect 2454 956 2488 957
rect 2596 926 2626 1020
rect 2732 989 2766 990
rect 2732 988 2733 989
rect 2656 958 2733 988
rect 2732 957 2733 958
rect 2765 988 2766 989
rect 2802 989 2836 990
rect 2802 988 2803 989
rect 2765 958 2768 988
rect 2800 958 2803 988
rect 2765 957 2766 958
rect 2732 956 2766 957
rect 2802 957 2803 958
rect 2835 988 2836 989
rect 2835 958 2914 988
rect 2835 957 2836 958
rect 2802 956 2836 957
rect 2944 926 2974 1020
rect 3080 989 3114 990
rect 3080 988 3081 989
rect 3004 958 3081 988
rect 3080 957 3081 958
rect 3113 988 3114 989
rect 3150 989 3184 990
rect 3150 988 3151 989
rect 3113 958 3116 988
rect 3148 958 3151 988
rect 3113 957 3114 958
rect 3080 956 3114 957
rect 3150 957 3151 958
rect 3183 988 3184 989
rect 3183 958 3262 988
rect 3183 957 3184 958
rect 3150 956 3184 957
rect 3292 926 3322 1020
rect 3428 989 3462 990
rect 3428 988 3429 989
rect 3352 958 3429 988
rect 3428 957 3429 958
rect 3461 988 3462 989
rect 3498 989 3532 990
rect 3498 988 3499 989
rect 3461 958 3464 988
rect 3496 958 3499 988
rect 3461 957 3462 958
rect 3428 956 3462 957
rect 3498 957 3499 958
rect 3531 988 3532 989
rect 3531 958 3610 988
rect 3531 957 3532 958
rect 3498 956 3532 957
rect 3640 926 3670 1020
rect 3776 989 3810 990
rect 3776 988 3777 989
rect 3700 958 3777 988
rect 3776 957 3777 958
rect 3809 988 3810 989
rect 3846 989 3880 990
rect 3846 988 3847 989
rect 3809 958 3812 988
rect 3844 958 3847 988
rect 3809 957 3810 958
rect 3776 956 3810 957
rect 3846 957 3847 958
rect 3879 988 3880 989
rect 3879 958 3958 988
rect 3879 957 3880 958
rect 3846 956 3880 957
rect 3988 926 4018 1020
rect 4124 989 4158 990
rect 4124 988 4125 989
rect 4048 958 4125 988
rect 4124 957 4125 958
rect 4157 988 4158 989
rect 4194 989 4228 990
rect 4194 988 4195 989
rect 4157 958 4160 988
rect 4192 958 4195 988
rect 4157 957 4158 958
rect 4124 956 4158 957
rect 4194 957 4195 958
rect 4227 988 4228 989
rect 4227 958 4306 988
rect 4227 957 4228 958
rect 4194 956 4228 957
rect 4336 926 4366 1020
rect 4472 989 4506 990
rect 4472 988 4473 989
rect 4396 958 4473 988
rect 4472 957 4473 958
rect 4505 988 4506 989
rect 4542 989 4576 990
rect 4542 988 4543 989
rect 4505 958 4508 988
rect 4540 958 4543 988
rect 4505 957 4506 958
rect 4472 956 4506 957
rect 4542 957 4543 958
rect 4575 988 4576 989
rect 4575 958 4654 988
rect 4575 957 4576 958
rect 4542 956 4576 957
rect 4684 926 4714 1020
rect 4820 989 4854 990
rect 4820 988 4821 989
rect 4744 958 4821 988
rect 4820 957 4821 958
rect 4853 988 4854 989
rect 4890 989 4924 990
rect 4890 988 4891 989
rect 4853 958 4856 988
rect 4888 958 4891 988
rect 4853 957 4854 958
rect 4820 956 4854 957
rect 4890 957 4891 958
rect 4923 988 4924 989
rect 4923 958 5002 988
rect 4923 957 4924 958
rect 4890 956 4924 957
rect 5032 926 5062 1020
rect 5168 989 5202 990
rect 5168 988 5169 989
rect 5092 958 5169 988
rect 5168 957 5169 958
rect 5201 988 5202 989
rect 5238 989 5272 990
rect 5238 988 5239 989
rect 5201 958 5204 988
rect 5236 958 5239 988
rect 5201 957 5202 958
rect 5168 956 5202 957
rect 5238 957 5239 958
rect 5271 988 5272 989
rect 5271 958 5350 988
rect 5271 957 5272 958
rect 5238 956 5272 957
rect 5380 926 5410 1020
rect 5516 989 5550 990
rect 5516 988 5517 989
rect 5440 958 5517 988
rect 5516 957 5517 958
rect 5549 988 5550 989
rect 5586 989 5620 990
rect 5586 988 5587 989
rect 5549 958 5552 988
rect 5584 958 5587 988
rect 5549 957 5550 958
rect 5516 956 5550 957
rect 5586 957 5587 958
rect 5619 988 5620 989
rect 5619 958 5698 988
rect 5619 957 5620 958
rect 5586 956 5620 957
rect 5728 926 5758 1020
rect 5864 989 5898 990
rect 5864 988 5865 989
rect 5788 958 5865 988
rect 5864 957 5865 958
rect 5897 988 5898 989
rect 5934 989 5968 990
rect 5934 988 5935 989
rect 5897 958 5900 988
rect 5932 958 5935 988
rect 5897 957 5898 958
rect 5864 956 5898 957
rect 5934 957 5935 958
rect 5967 988 5968 989
rect 5967 958 6046 988
rect 5967 957 5968 958
rect 5934 956 5968 957
rect 6076 926 6106 1020
rect 6212 989 6246 990
rect 6212 988 6213 989
rect 6136 958 6213 988
rect 6212 957 6213 958
rect 6245 988 6246 989
rect 6282 989 6316 990
rect 6282 988 6283 989
rect 6245 958 6248 988
rect 6280 958 6283 988
rect 6245 957 6246 958
rect 6212 956 6246 957
rect 6282 957 6283 958
rect 6315 988 6316 989
rect 6315 958 6394 988
rect 6315 957 6316 958
rect 6282 956 6316 957
rect 6424 926 6454 1020
rect 6560 989 6594 990
rect 6560 988 6561 989
rect 6484 958 6561 988
rect 6560 957 6561 958
rect 6593 988 6594 989
rect 6630 989 6664 990
rect 6630 988 6631 989
rect 6593 958 6596 988
rect 6628 958 6631 988
rect 6593 957 6594 958
rect 6560 956 6594 957
rect 6630 957 6631 958
rect 6663 988 6664 989
rect 6663 958 6742 988
rect 6663 957 6664 958
rect 6630 956 6664 957
rect 6772 926 6802 1020
rect 6908 989 6942 990
rect 6908 988 6909 989
rect 6832 958 6909 988
rect 6908 957 6909 958
rect 6941 988 6942 989
rect 6978 989 7012 990
rect 6978 988 6979 989
rect 6941 958 6944 988
rect 6976 958 6979 988
rect 6941 957 6942 958
rect 6908 956 6942 957
rect 6978 957 6979 958
rect 7011 988 7012 989
rect 7011 958 7090 988
rect 7011 957 7012 958
rect 6978 956 7012 957
rect 7120 926 7150 1020
rect 7256 989 7290 990
rect 7256 988 7257 989
rect 7180 958 7257 988
rect 7256 957 7257 958
rect 7289 988 7290 989
rect 7289 958 7292 988
rect 7289 957 7290 958
rect 7256 956 7290 957
rect 0 896 318 926
rect 348 896 1392 926
rect 1422 896 2058 926
rect 2088 896 3130 926
rect 3160 896 3480 926
rect 3510 896 3798 926
rect 3828 896 4872 926
rect 4902 896 5220 926
rect 5250 896 5538 926
rect 5568 896 6612 926
rect 6642 896 6960 926
rect 6990 896 7278 926
rect 18 865 52 866
rect 18 864 19 865
rect 16 834 19 864
rect 18 833 19 834
rect 51 864 52 865
rect 51 834 130 864
rect 51 833 52 834
rect 18 832 52 833
rect 160 802 190 896
rect 296 865 330 866
rect 296 864 297 865
rect 220 834 297 864
rect 296 833 297 834
rect 329 864 330 865
rect 366 865 400 866
rect 366 864 367 865
rect 329 834 332 864
rect 364 834 367 864
rect 329 833 330 834
rect 296 832 330 833
rect 366 833 367 834
rect 399 864 400 865
rect 399 834 478 864
rect 399 833 400 834
rect 366 832 400 833
rect 508 802 538 896
rect 644 865 678 866
rect 644 864 645 865
rect 568 834 645 864
rect 644 833 645 834
rect 677 864 678 865
rect 714 865 748 866
rect 714 864 715 865
rect 677 834 680 864
rect 712 834 715 864
rect 677 833 678 834
rect 644 832 678 833
rect 714 833 715 834
rect 747 864 748 865
rect 747 834 826 864
rect 747 833 748 834
rect 714 832 748 833
rect 856 802 886 896
rect 992 865 1026 866
rect 992 864 993 865
rect 916 834 993 864
rect 992 833 993 834
rect 1025 864 1026 865
rect 1062 865 1096 866
rect 1062 864 1063 865
rect 1025 834 1028 864
rect 1060 834 1063 864
rect 1025 833 1026 834
rect 992 832 1026 833
rect 1062 833 1063 834
rect 1095 864 1096 865
rect 1095 834 1174 864
rect 1095 833 1096 834
rect 1062 832 1096 833
rect 1204 802 1234 896
rect 1340 865 1374 866
rect 1340 864 1341 865
rect 1264 834 1341 864
rect 1340 833 1341 834
rect 1373 864 1374 865
rect 1410 865 1444 866
rect 1410 864 1411 865
rect 1373 834 1376 864
rect 1408 834 1411 864
rect 1373 833 1374 834
rect 1340 832 1374 833
rect 1410 833 1411 834
rect 1443 864 1444 865
rect 1443 834 1522 864
rect 1443 833 1444 834
rect 1410 832 1444 833
rect 1552 802 1582 896
rect 1688 865 1722 866
rect 1688 864 1689 865
rect 1612 834 1689 864
rect 1688 833 1689 834
rect 1721 864 1722 865
rect 1758 865 1792 866
rect 1758 864 1759 865
rect 1721 834 1724 864
rect 1756 834 1759 864
rect 1721 833 1722 834
rect 1688 832 1722 833
rect 1758 833 1759 834
rect 1791 864 1792 865
rect 1791 834 1870 864
rect 1791 833 1792 834
rect 1758 832 1792 833
rect 1900 802 1930 896
rect 2036 865 2070 866
rect 2036 864 2037 865
rect 1960 834 2037 864
rect 2036 833 2037 834
rect 2069 864 2070 865
rect 2106 865 2140 866
rect 2106 864 2107 865
rect 2069 834 2072 864
rect 2104 834 2107 864
rect 2069 833 2070 834
rect 2036 832 2070 833
rect 2106 833 2107 834
rect 2139 864 2140 865
rect 2139 834 2218 864
rect 2139 833 2140 834
rect 2106 832 2140 833
rect 2248 802 2278 896
rect 2384 865 2418 866
rect 2384 864 2385 865
rect 2308 834 2385 864
rect 2384 833 2385 834
rect 2417 864 2418 865
rect 2454 865 2488 866
rect 2454 864 2455 865
rect 2417 834 2420 864
rect 2452 834 2455 864
rect 2417 833 2418 834
rect 2384 832 2418 833
rect 2454 833 2455 834
rect 2487 864 2488 865
rect 2487 834 2566 864
rect 2487 833 2488 834
rect 2454 832 2488 833
rect 2596 802 2626 896
rect 2732 865 2766 866
rect 2732 864 2733 865
rect 2656 834 2733 864
rect 2732 833 2733 834
rect 2765 864 2766 865
rect 2802 865 2836 866
rect 2802 864 2803 865
rect 2765 834 2768 864
rect 2800 834 2803 864
rect 2765 833 2766 834
rect 2732 832 2766 833
rect 2802 833 2803 834
rect 2835 864 2836 865
rect 2835 834 2914 864
rect 2835 833 2836 834
rect 2802 832 2836 833
rect 2944 802 2974 896
rect 3080 865 3114 866
rect 3080 864 3081 865
rect 3004 834 3081 864
rect 3080 833 3081 834
rect 3113 864 3114 865
rect 3150 865 3184 866
rect 3150 864 3151 865
rect 3113 834 3116 864
rect 3148 834 3151 864
rect 3113 833 3114 834
rect 3080 832 3114 833
rect 3150 833 3151 834
rect 3183 864 3184 865
rect 3183 834 3262 864
rect 3183 833 3184 834
rect 3150 832 3184 833
rect 3292 802 3322 896
rect 3428 865 3462 866
rect 3428 864 3429 865
rect 3352 834 3429 864
rect 3428 833 3429 834
rect 3461 864 3462 865
rect 3498 865 3532 866
rect 3498 864 3499 865
rect 3461 834 3464 864
rect 3496 834 3499 864
rect 3461 833 3462 834
rect 3428 832 3462 833
rect 3498 833 3499 834
rect 3531 864 3532 865
rect 3531 834 3610 864
rect 3531 833 3532 834
rect 3498 832 3532 833
rect 3640 802 3670 896
rect 3776 865 3810 866
rect 3776 864 3777 865
rect 3700 834 3777 864
rect 3776 833 3777 834
rect 3809 864 3810 865
rect 3846 865 3880 866
rect 3846 864 3847 865
rect 3809 834 3812 864
rect 3844 834 3847 864
rect 3809 833 3810 834
rect 3776 832 3810 833
rect 3846 833 3847 834
rect 3879 864 3880 865
rect 3879 834 3958 864
rect 3879 833 3880 834
rect 3846 832 3880 833
rect 3988 802 4018 896
rect 4124 865 4158 866
rect 4124 864 4125 865
rect 4048 834 4125 864
rect 4124 833 4125 834
rect 4157 864 4158 865
rect 4194 865 4228 866
rect 4194 864 4195 865
rect 4157 834 4160 864
rect 4192 834 4195 864
rect 4157 833 4158 834
rect 4124 832 4158 833
rect 4194 833 4195 834
rect 4227 864 4228 865
rect 4227 834 4306 864
rect 4227 833 4228 834
rect 4194 832 4228 833
rect 4336 802 4366 896
rect 4472 865 4506 866
rect 4472 864 4473 865
rect 4396 834 4473 864
rect 4472 833 4473 834
rect 4505 864 4506 865
rect 4542 865 4576 866
rect 4542 864 4543 865
rect 4505 834 4508 864
rect 4540 834 4543 864
rect 4505 833 4506 834
rect 4472 832 4506 833
rect 4542 833 4543 834
rect 4575 864 4576 865
rect 4575 834 4654 864
rect 4575 833 4576 834
rect 4542 832 4576 833
rect 4684 802 4714 896
rect 4820 865 4854 866
rect 4820 864 4821 865
rect 4744 834 4821 864
rect 4820 833 4821 834
rect 4853 864 4854 865
rect 4890 865 4924 866
rect 4890 864 4891 865
rect 4853 834 4856 864
rect 4888 834 4891 864
rect 4853 833 4854 834
rect 4820 832 4854 833
rect 4890 833 4891 834
rect 4923 864 4924 865
rect 4923 834 5002 864
rect 4923 833 4924 834
rect 4890 832 4924 833
rect 5032 802 5062 896
rect 5168 865 5202 866
rect 5168 864 5169 865
rect 5092 834 5169 864
rect 5168 833 5169 834
rect 5201 864 5202 865
rect 5238 865 5272 866
rect 5238 864 5239 865
rect 5201 834 5204 864
rect 5236 834 5239 864
rect 5201 833 5202 834
rect 5168 832 5202 833
rect 5238 833 5239 834
rect 5271 864 5272 865
rect 5271 834 5350 864
rect 5271 833 5272 834
rect 5238 832 5272 833
rect 5380 802 5410 896
rect 5516 865 5550 866
rect 5516 864 5517 865
rect 5440 834 5517 864
rect 5516 833 5517 834
rect 5549 864 5550 865
rect 5586 865 5620 866
rect 5586 864 5587 865
rect 5549 834 5552 864
rect 5584 834 5587 864
rect 5549 833 5550 834
rect 5516 832 5550 833
rect 5586 833 5587 834
rect 5619 864 5620 865
rect 5619 834 5698 864
rect 5619 833 5620 834
rect 5586 832 5620 833
rect 5728 802 5758 896
rect 5864 865 5898 866
rect 5864 864 5865 865
rect 5788 834 5865 864
rect 5864 833 5865 834
rect 5897 864 5898 865
rect 5934 865 5968 866
rect 5934 864 5935 865
rect 5897 834 5900 864
rect 5932 834 5935 864
rect 5897 833 5898 834
rect 5864 832 5898 833
rect 5934 833 5935 834
rect 5967 864 5968 865
rect 5967 834 6046 864
rect 5967 833 5968 834
rect 5934 832 5968 833
rect 6076 802 6106 896
rect 6212 865 6246 866
rect 6212 864 6213 865
rect 6136 834 6213 864
rect 6212 833 6213 834
rect 6245 864 6246 865
rect 6282 865 6316 866
rect 6282 864 6283 865
rect 6245 834 6248 864
rect 6280 834 6283 864
rect 6245 833 6246 834
rect 6212 832 6246 833
rect 6282 833 6283 834
rect 6315 864 6316 865
rect 6315 834 6394 864
rect 6315 833 6316 834
rect 6282 832 6316 833
rect 6424 802 6454 896
rect 6560 865 6594 866
rect 6560 864 6561 865
rect 6484 834 6561 864
rect 6560 833 6561 834
rect 6593 864 6594 865
rect 6630 865 6664 866
rect 6630 864 6631 865
rect 6593 834 6596 864
rect 6628 834 6631 864
rect 6593 833 6594 834
rect 6560 832 6594 833
rect 6630 833 6631 834
rect 6663 864 6664 865
rect 6663 834 6742 864
rect 6663 833 6664 834
rect 6630 832 6664 833
rect 6772 802 6802 896
rect 6908 865 6942 866
rect 6908 864 6909 865
rect 6832 834 6909 864
rect 6908 833 6909 834
rect 6941 864 6942 865
rect 6978 865 7012 866
rect 6978 864 6979 865
rect 6941 834 6944 864
rect 6976 834 6979 864
rect 6941 833 6942 834
rect 6908 832 6942 833
rect 6978 833 6979 834
rect 7011 864 7012 865
rect 7011 834 7090 864
rect 7011 833 7012 834
rect 6978 832 7012 833
rect 7120 802 7150 896
rect 7256 865 7290 866
rect 7256 864 7257 865
rect 7180 834 7257 864
rect 7256 833 7257 834
rect 7289 864 7290 865
rect 7289 834 7292 864
rect 7289 833 7290 834
rect 7256 832 7290 833
rect 0 772 318 802
rect 348 772 1392 802
rect 1422 772 2058 802
rect 2088 772 3131 802
rect 3162 772 3480 802
rect 3510 772 3798 802
rect 3828 772 4872 802
rect 4902 772 5220 802
rect 5250 772 5538 802
rect 5568 772 6612 802
rect 6642 772 6960 802
rect 6990 772 7278 802
rect 18 741 52 742
rect 18 740 19 741
rect 16 710 19 740
rect 18 709 19 710
rect 51 740 52 741
rect 51 710 130 740
rect 51 709 52 710
rect 18 708 52 709
rect 160 678 190 772
rect 296 741 330 742
rect 296 740 297 741
rect 220 710 297 740
rect 296 709 297 710
rect 329 740 330 741
rect 366 741 400 742
rect 366 740 367 741
rect 329 710 332 740
rect 364 710 367 740
rect 329 709 330 710
rect 296 708 330 709
rect 366 709 367 710
rect 399 740 400 741
rect 399 710 478 740
rect 399 709 400 710
rect 366 708 400 709
rect 508 678 538 772
rect 644 741 678 742
rect 644 740 645 741
rect 568 710 645 740
rect 644 709 645 710
rect 677 740 678 741
rect 714 741 748 742
rect 714 740 715 741
rect 677 710 680 740
rect 712 710 715 740
rect 677 709 678 710
rect 644 708 678 709
rect 714 709 715 710
rect 747 740 748 741
rect 747 710 826 740
rect 747 709 748 710
rect 714 708 748 709
rect 856 678 886 772
rect 992 741 1026 742
rect 992 740 993 741
rect 916 710 993 740
rect 992 709 993 710
rect 1025 740 1026 741
rect 1062 741 1096 742
rect 1062 740 1063 741
rect 1025 710 1028 740
rect 1060 710 1063 740
rect 1025 709 1026 710
rect 992 708 1026 709
rect 1062 709 1063 710
rect 1095 740 1096 741
rect 1095 710 1174 740
rect 1095 709 1096 710
rect 1062 708 1096 709
rect 1204 678 1234 772
rect 1340 741 1374 742
rect 1340 740 1341 741
rect 1264 710 1341 740
rect 1340 709 1341 710
rect 1373 740 1374 741
rect 1410 741 1444 742
rect 1410 740 1411 741
rect 1373 710 1376 740
rect 1408 710 1411 740
rect 1373 709 1374 710
rect 1340 708 1374 709
rect 1410 709 1411 710
rect 1443 740 1444 741
rect 1443 710 1522 740
rect 1443 709 1444 710
rect 1410 708 1444 709
rect 1552 678 1582 772
rect 1688 741 1722 742
rect 1688 740 1689 741
rect 1612 710 1689 740
rect 1688 709 1689 710
rect 1721 740 1722 741
rect 1758 741 1792 742
rect 1758 740 1759 741
rect 1721 710 1724 740
rect 1756 710 1759 740
rect 1721 709 1722 710
rect 1688 708 1722 709
rect 1758 709 1759 710
rect 1791 740 1792 741
rect 1791 710 1870 740
rect 1791 709 1792 710
rect 1758 708 1792 709
rect 1900 678 1930 772
rect 2036 741 2070 742
rect 2036 740 2037 741
rect 1960 710 2037 740
rect 2036 709 2037 710
rect 2069 740 2070 741
rect 2106 741 2140 742
rect 2106 740 2107 741
rect 2069 710 2072 740
rect 2104 710 2107 740
rect 2069 709 2070 710
rect 2036 708 2070 709
rect 2106 709 2107 710
rect 2139 740 2140 741
rect 2139 710 2218 740
rect 2139 709 2140 710
rect 2106 708 2140 709
rect 2248 678 2278 772
rect 2384 741 2418 742
rect 2384 740 2385 741
rect 2308 710 2385 740
rect 2384 709 2385 710
rect 2417 740 2418 741
rect 2454 741 2488 742
rect 2454 740 2455 741
rect 2417 710 2420 740
rect 2452 710 2455 740
rect 2417 709 2418 710
rect 2384 708 2418 709
rect 2454 709 2455 710
rect 2487 740 2488 741
rect 2487 710 2566 740
rect 2487 709 2488 710
rect 2454 708 2488 709
rect 2596 678 2626 772
rect 2732 741 2766 742
rect 2732 740 2733 741
rect 2656 710 2733 740
rect 2732 709 2733 710
rect 2765 740 2766 741
rect 2802 741 2836 742
rect 2802 740 2803 741
rect 2765 710 2768 740
rect 2800 710 2803 740
rect 2765 709 2766 710
rect 2732 708 2766 709
rect 2802 709 2803 710
rect 2835 740 2836 741
rect 2835 710 2914 740
rect 2835 709 2836 710
rect 2802 708 2836 709
rect 2944 678 2974 772
rect 3080 741 3114 742
rect 3080 740 3081 741
rect 3004 710 3081 740
rect 3080 709 3081 710
rect 3113 740 3114 741
rect 3150 741 3184 742
rect 3150 740 3151 741
rect 3113 710 3116 740
rect 3148 710 3151 740
rect 3113 709 3114 710
rect 3080 708 3114 709
rect 3150 709 3151 710
rect 3183 740 3184 741
rect 3183 710 3262 740
rect 3183 709 3184 710
rect 3150 708 3184 709
rect 3292 678 3322 772
rect 3428 741 3462 742
rect 3428 740 3429 741
rect 3352 710 3429 740
rect 3428 709 3429 710
rect 3461 740 3462 741
rect 3498 741 3532 742
rect 3498 740 3499 741
rect 3461 710 3464 740
rect 3496 710 3499 740
rect 3461 709 3462 710
rect 3428 708 3462 709
rect 3498 709 3499 710
rect 3531 740 3532 741
rect 3531 710 3610 740
rect 3531 709 3532 710
rect 3498 708 3532 709
rect 3640 678 3670 772
rect 3776 741 3810 742
rect 3776 740 3777 741
rect 3700 710 3777 740
rect 3776 709 3777 710
rect 3809 740 3810 741
rect 3846 741 3880 742
rect 3846 740 3847 741
rect 3809 710 3812 740
rect 3844 710 3847 740
rect 3809 709 3810 710
rect 3776 708 3810 709
rect 3846 709 3847 710
rect 3879 740 3880 741
rect 3879 710 3958 740
rect 3879 709 3880 710
rect 3846 708 3880 709
rect 3988 678 4018 772
rect 4124 741 4158 742
rect 4124 740 4125 741
rect 4048 710 4125 740
rect 4124 709 4125 710
rect 4157 740 4158 741
rect 4194 741 4228 742
rect 4194 740 4195 741
rect 4157 710 4160 740
rect 4192 710 4195 740
rect 4157 709 4158 710
rect 4124 708 4158 709
rect 4194 709 4195 710
rect 4227 740 4228 741
rect 4227 710 4306 740
rect 4227 709 4228 710
rect 4194 708 4228 709
rect 4336 678 4366 772
rect 4472 741 4506 742
rect 4472 740 4473 741
rect 4396 710 4473 740
rect 4472 709 4473 710
rect 4505 740 4506 741
rect 4542 741 4576 742
rect 4542 740 4543 741
rect 4505 710 4508 740
rect 4540 710 4543 740
rect 4505 709 4506 710
rect 4472 708 4506 709
rect 4542 709 4543 710
rect 4575 740 4576 741
rect 4575 710 4654 740
rect 4575 709 4576 710
rect 4542 708 4576 709
rect 4684 678 4714 772
rect 4820 741 4854 742
rect 4820 740 4821 741
rect 4744 710 4821 740
rect 4820 709 4821 710
rect 4853 740 4854 741
rect 4890 741 4924 742
rect 4890 740 4891 741
rect 4853 710 4856 740
rect 4888 710 4891 740
rect 4853 709 4854 710
rect 4820 708 4854 709
rect 4890 709 4891 710
rect 4923 740 4924 741
rect 4923 710 5002 740
rect 4923 709 4924 710
rect 4890 708 4924 709
rect 5032 678 5062 772
rect 5168 741 5202 742
rect 5168 740 5169 741
rect 5092 710 5169 740
rect 5168 709 5169 710
rect 5201 740 5202 741
rect 5238 741 5272 742
rect 5238 740 5239 741
rect 5201 710 5204 740
rect 5236 710 5239 740
rect 5201 709 5202 710
rect 5168 708 5202 709
rect 5238 709 5239 710
rect 5271 740 5272 741
rect 5271 710 5350 740
rect 5271 709 5272 710
rect 5238 708 5272 709
rect 5380 678 5410 772
rect 5516 741 5550 742
rect 5516 740 5517 741
rect 5440 710 5517 740
rect 5516 709 5517 710
rect 5549 740 5550 741
rect 5586 741 5620 742
rect 5586 740 5587 741
rect 5549 710 5552 740
rect 5584 710 5587 740
rect 5549 709 5550 710
rect 5516 708 5550 709
rect 5586 709 5587 710
rect 5619 740 5620 741
rect 5619 710 5698 740
rect 5619 709 5620 710
rect 5586 708 5620 709
rect 5728 678 5758 772
rect 5864 741 5898 742
rect 5864 740 5865 741
rect 5788 710 5865 740
rect 5864 709 5865 710
rect 5897 740 5898 741
rect 5934 741 5968 742
rect 5934 740 5935 741
rect 5897 710 5900 740
rect 5932 710 5935 740
rect 5897 709 5898 710
rect 5864 708 5898 709
rect 5934 709 5935 710
rect 5967 740 5968 741
rect 5967 710 6046 740
rect 5967 709 5968 710
rect 5934 708 5968 709
rect 6076 678 6106 772
rect 6212 741 6246 742
rect 6212 740 6213 741
rect 6136 710 6213 740
rect 6212 709 6213 710
rect 6245 740 6246 741
rect 6282 741 6316 742
rect 6282 740 6283 741
rect 6245 710 6248 740
rect 6280 710 6283 740
rect 6245 709 6246 710
rect 6212 708 6246 709
rect 6282 709 6283 710
rect 6315 740 6316 741
rect 6315 710 6394 740
rect 6315 709 6316 710
rect 6282 708 6316 709
rect 6424 678 6454 772
rect 6560 741 6594 742
rect 6560 740 6561 741
rect 6484 710 6561 740
rect 6560 709 6561 710
rect 6593 740 6594 741
rect 6630 741 6664 742
rect 6630 740 6631 741
rect 6593 710 6596 740
rect 6628 710 6631 740
rect 6593 709 6594 710
rect 6560 708 6594 709
rect 6630 709 6631 710
rect 6663 740 6664 741
rect 6663 710 6742 740
rect 6663 709 6664 710
rect 6630 708 6664 709
rect 6772 678 6802 772
rect 6908 741 6942 742
rect 6908 740 6909 741
rect 6832 710 6909 740
rect 6908 709 6909 710
rect 6941 740 6942 741
rect 6978 741 7012 742
rect 6978 740 6979 741
rect 6941 710 6944 740
rect 6976 710 6979 740
rect 6941 709 6942 710
rect 6908 708 6942 709
rect 6978 709 6979 710
rect 7011 740 7012 741
rect 7011 710 7090 740
rect 7011 709 7012 710
rect 6978 708 7012 709
rect 7120 678 7150 772
rect 7256 741 7290 742
rect 7256 740 7257 741
rect 7180 710 7257 740
rect 7256 709 7257 710
rect 7289 740 7290 741
rect 7289 710 7292 740
rect 7289 709 7290 710
rect 7256 708 7290 709
rect 0 648 318 678
rect 348 648 1392 678
rect 1422 648 2058 678
rect 2088 648 3132 678
rect 3162 648 3480 678
rect 3510 648 3798 678
rect 3828 648 4872 678
rect 4902 648 5220 678
rect 5250 648 5538 678
rect 5568 648 6612 678
rect 6642 648 6960 678
rect 6990 648 7278 678
rect 18 617 52 618
rect 18 616 19 617
rect 16 586 19 616
rect 18 585 19 586
rect 51 616 52 617
rect 51 586 130 616
rect 51 585 52 586
rect 18 584 52 585
rect 18 547 52 548
rect 18 546 19 547
rect 16 516 19 546
rect 18 515 19 516
rect 51 546 52 547
rect 51 516 130 546
rect 51 515 52 516
rect 18 514 52 515
rect 160 484 190 648
rect 296 617 330 618
rect 296 616 297 617
rect 220 586 297 616
rect 296 585 297 586
rect 329 616 330 617
rect 366 617 400 618
rect 366 616 367 617
rect 329 586 332 616
rect 364 586 367 616
rect 329 585 330 586
rect 296 584 330 585
rect 366 585 367 586
rect 399 616 400 617
rect 399 586 478 616
rect 399 585 400 586
rect 366 584 400 585
rect 508 566 538 648
rect 644 617 678 618
rect 644 616 645 617
rect 568 586 645 616
rect 644 585 645 586
rect 677 616 678 617
rect 714 617 748 618
rect 714 616 715 617
rect 677 586 680 616
rect 712 586 715 616
rect 677 585 678 586
rect 644 584 678 585
rect 714 585 715 586
rect 747 616 748 617
rect 747 586 826 616
rect 747 585 748 586
rect 714 584 748 585
rect 856 566 886 648
rect 992 617 1026 618
rect 992 616 993 617
rect 916 586 993 616
rect 992 585 993 586
rect 1025 616 1026 617
rect 1062 617 1096 618
rect 1062 616 1063 617
rect 1025 586 1028 616
rect 1060 586 1063 616
rect 1025 585 1026 586
rect 992 584 1026 585
rect 1062 585 1063 586
rect 1095 616 1096 617
rect 1095 586 1174 616
rect 1095 585 1096 586
rect 1062 584 1096 585
rect 1204 566 1234 648
rect 1340 617 1374 618
rect 1340 616 1341 617
rect 1264 586 1341 616
rect 1340 585 1341 586
rect 1373 616 1374 617
rect 1410 617 1444 618
rect 1410 616 1411 617
rect 1373 586 1376 616
rect 1408 586 1411 616
rect 1373 585 1374 586
rect 1340 584 1374 585
rect 1410 585 1411 586
rect 1443 616 1444 617
rect 1443 586 1522 616
rect 1443 585 1444 586
rect 1410 584 1444 585
rect 296 547 330 548
rect 296 546 297 547
rect 220 516 297 546
rect 296 515 297 516
rect 329 546 330 547
rect 366 547 400 548
rect 366 546 367 547
rect 329 516 332 546
rect 364 516 367 546
rect 329 515 330 516
rect 296 514 330 515
rect 366 515 367 516
rect 399 546 400 547
rect 644 547 678 548
rect 644 546 645 547
rect 399 516 478 546
rect 399 515 400 516
rect 366 514 400 515
rect 508 484 538 536
rect 568 516 645 546
rect 644 515 645 516
rect 677 546 678 547
rect 714 547 748 548
rect 714 546 715 547
rect 677 516 680 546
rect 712 516 715 546
rect 677 515 678 516
rect 644 514 678 515
rect 714 515 715 516
rect 747 546 748 547
rect 992 547 1026 548
rect 992 546 993 547
rect 747 516 826 546
rect 747 515 748 516
rect 714 514 748 515
rect 856 484 886 536
rect 916 516 993 546
rect 992 515 993 516
rect 1025 546 1026 547
rect 1062 547 1096 548
rect 1062 546 1063 547
rect 1025 516 1028 546
rect 1060 516 1063 546
rect 1025 515 1026 516
rect 992 514 1026 515
rect 1062 515 1063 516
rect 1095 546 1096 547
rect 1340 547 1374 548
rect 1340 546 1341 547
rect 1095 516 1174 546
rect 1095 515 1096 516
rect 1062 514 1096 515
rect 1204 484 1234 536
rect 1264 516 1341 546
rect 1340 515 1341 516
rect 1373 546 1374 547
rect 1410 547 1444 548
rect 1410 546 1411 547
rect 1373 516 1376 546
rect 1408 516 1411 546
rect 1373 515 1374 516
rect 1340 514 1374 515
rect 1410 515 1411 516
rect 1443 546 1444 547
rect 1443 516 1522 546
rect 1443 515 1444 516
rect 1410 514 1444 515
rect 1552 484 1582 648
rect 1688 617 1722 618
rect 1688 616 1689 617
rect 1612 586 1689 616
rect 1688 585 1689 586
rect 1721 616 1722 617
rect 1758 617 1792 618
rect 1758 616 1759 617
rect 1721 586 1724 616
rect 1756 586 1759 616
rect 1721 585 1722 586
rect 1688 584 1722 585
rect 1758 585 1759 586
rect 1791 616 1792 617
rect 1791 586 1870 616
rect 1791 585 1792 586
rect 1758 584 1792 585
rect 1688 547 1722 548
rect 1688 546 1689 547
rect 1612 516 1689 546
rect 1688 515 1689 516
rect 1721 546 1722 547
rect 1758 547 1792 548
rect 1758 546 1759 547
rect 1721 516 1724 546
rect 1756 516 1759 546
rect 1721 515 1722 516
rect 1688 514 1722 515
rect 1758 515 1759 516
rect 1791 546 1792 547
rect 1791 516 1870 546
rect 1791 515 1792 516
rect 1758 514 1792 515
rect 1900 484 1930 648
rect 2036 617 2070 618
rect 2036 616 2037 617
rect 1960 586 2037 616
rect 2036 585 2037 586
rect 2069 616 2070 617
rect 2106 617 2140 618
rect 2106 616 2107 617
rect 2069 586 2072 616
rect 2104 586 2107 616
rect 2069 585 2070 586
rect 2036 584 2070 585
rect 2106 585 2107 586
rect 2139 616 2140 617
rect 2139 586 2218 616
rect 2139 585 2140 586
rect 2106 584 2140 585
rect 2248 566 2278 648
rect 2384 617 2418 618
rect 2384 616 2385 617
rect 2308 586 2385 616
rect 2384 585 2385 586
rect 2417 616 2418 617
rect 2454 617 2488 618
rect 2454 616 2455 617
rect 2417 586 2420 616
rect 2452 586 2455 616
rect 2417 585 2418 586
rect 2384 584 2418 585
rect 2454 585 2455 586
rect 2487 616 2488 617
rect 2487 586 2566 616
rect 2487 585 2488 586
rect 2454 584 2488 585
rect 2036 547 2070 548
rect 2036 546 2037 547
rect 1960 516 2037 546
rect 2036 515 2037 516
rect 2069 546 2070 547
rect 2106 547 2140 548
rect 2106 546 2107 547
rect 2069 516 2072 546
rect 2104 516 2107 546
rect 2069 515 2070 516
rect 2036 514 2070 515
rect 2106 515 2107 516
rect 2139 546 2140 547
rect 2384 547 2418 548
rect 2384 546 2385 547
rect 2139 516 2218 546
rect 2139 515 2140 516
rect 2106 514 2140 515
rect 2248 484 2278 536
rect 2308 516 2385 546
rect 2384 515 2385 516
rect 2417 546 2418 547
rect 2454 547 2488 548
rect 2454 546 2455 547
rect 2417 516 2420 546
rect 2452 516 2455 546
rect 2417 515 2418 516
rect 2384 514 2418 515
rect 2454 515 2455 516
rect 2487 546 2488 547
rect 2487 516 2566 546
rect 2487 515 2488 516
rect 2454 514 2488 515
rect 2596 484 2626 648
rect 2732 617 2766 618
rect 2732 616 2733 617
rect 2656 586 2733 616
rect 2732 585 2733 586
rect 2765 616 2766 617
rect 2802 617 2836 618
rect 2802 616 2803 617
rect 2765 586 2768 616
rect 2800 586 2803 616
rect 2765 585 2766 586
rect 2732 584 2766 585
rect 2802 585 2803 586
rect 2835 616 2836 617
rect 2835 586 2914 616
rect 2835 585 2836 586
rect 2802 584 2836 585
rect 2944 566 2974 648
rect 3080 617 3114 618
rect 3080 616 3081 617
rect 3004 586 3081 616
rect 3080 585 3081 586
rect 3113 616 3114 617
rect 3150 617 3184 618
rect 3150 616 3151 617
rect 3113 586 3116 616
rect 3148 586 3151 616
rect 3113 585 3114 586
rect 3080 584 3114 585
rect 3150 585 3151 586
rect 3183 616 3184 617
rect 3183 586 3262 616
rect 3183 585 3184 586
rect 3150 584 3184 585
rect 2732 547 2766 548
rect 2732 546 2733 547
rect 2656 516 2733 546
rect 2732 515 2733 516
rect 2765 546 2766 547
rect 2802 547 2836 548
rect 2802 546 2803 547
rect 2765 516 2768 546
rect 2800 516 2803 546
rect 2765 515 2766 516
rect 2732 514 2766 515
rect 2802 515 2803 516
rect 2835 546 2836 547
rect 3080 547 3114 548
rect 3080 546 3081 547
rect 2835 516 2914 546
rect 2835 515 2836 516
rect 2802 514 2836 515
rect 2944 484 2974 536
rect 3004 516 3081 546
rect 3080 515 3081 516
rect 3113 546 3114 547
rect 3150 547 3184 548
rect 3150 546 3151 547
rect 3113 516 3116 546
rect 3148 516 3151 546
rect 3113 515 3114 516
rect 3080 514 3114 515
rect 3150 515 3151 516
rect 3183 546 3184 547
rect 3183 516 3262 546
rect 3183 515 3184 516
rect 3150 514 3184 515
rect 3292 484 3322 648
rect 3428 617 3462 618
rect 3428 616 3429 617
rect 3352 586 3429 616
rect 3428 585 3429 586
rect 3461 616 3462 617
rect 3498 617 3532 618
rect 3498 616 3499 617
rect 3461 586 3464 616
rect 3496 586 3499 616
rect 3461 585 3462 586
rect 3428 584 3462 585
rect 3498 585 3499 586
rect 3531 616 3532 617
rect 3531 586 3610 616
rect 3531 585 3532 586
rect 3498 584 3532 585
rect 3428 547 3462 548
rect 3428 546 3429 547
rect 3352 516 3429 546
rect 3428 515 3429 516
rect 3461 546 3462 547
rect 3498 547 3532 548
rect 3498 546 3499 547
rect 3461 516 3464 546
rect 3496 516 3499 546
rect 3461 515 3462 516
rect 3428 514 3462 515
rect 3498 515 3499 516
rect 3531 546 3532 547
rect 3531 516 3610 546
rect 3531 515 3532 516
rect 3498 514 3532 515
rect 3640 484 3670 648
rect 3776 617 3810 618
rect 3776 616 3777 617
rect 3700 586 3777 616
rect 3776 585 3777 586
rect 3809 616 3810 617
rect 3846 617 3880 618
rect 3846 616 3847 617
rect 3809 586 3812 616
rect 3844 586 3847 616
rect 3809 585 3810 586
rect 3776 584 3810 585
rect 3846 585 3847 586
rect 3879 616 3880 617
rect 3879 586 3958 616
rect 3879 585 3880 586
rect 3846 584 3880 585
rect 3988 566 4018 648
rect 4124 617 4158 618
rect 4124 616 4125 617
rect 4048 586 4125 616
rect 4124 585 4125 586
rect 4157 616 4158 617
rect 4194 617 4228 618
rect 4194 616 4195 617
rect 4157 586 4160 616
rect 4192 586 4195 616
rect 4157 585 4158 586
rect 4124 584 4158 585
rect 4194 585 4195 586
rect 4227 616 4228 617
rect 4227 586 4306 616
rect 4227 585 4228 586
rect 4194 584 4228 585
rect 3776 547 3810 548
rect 3776 546 3777 547
rect 3700 516 3777 546
rect 3776 515 3777 516
rect 3809 546 3810 547
rect 3846 547 3880 548
rect 3846 546 3847 547
rect 3809 516 3812 546
rect 3844 516 3847 546
rect 3809 515 3810 516
rect 3776 514 3810 515
rect 3846 515 3847 516
rect 3879 546 3880 547
rect 4124 547 4158 548
rect 4124 546 4125 547
rect 3879 516 3958 546
rect 3879 515 3880 516
rect 3846 514 3880 515
rect 3988 484 4018 536
rect 4048 516 4125 546
rect 4124 515 4125 516
rect 4157 546 4158 547
rect 4194 547 4228 548
rect 4194 546 4195 547
rect 4157 516 4160 546
rect 4192 516 4195 546
rect 4157 515 4158 516
rect 4124 514 4158 515
rect 4194 515 4195 516
rect 4227 546 4228 547
rect 4227 516 4306 546
rect 4227 515 4228 516
rect 4194 514 4228 515
rect 4336 484 4366 648
rect 4472 617 4506 618
rect 4472 616 4473 617
rect 4396 586 4473 616
rect 4472 585 4473 586
rect 4505 616 4506 617
rect 4542 617 4576 618
rect 4542 616 4543 617
rect 4505 586 4508 616
rect 4540 586 4543 616
rect 4505 585 4506 586
rect 4472 584 4506 585
rect 4542 585 4543 586
rect 4575 616 4576 617
rect 4575 586 4654 616
rect 4575 585 4576 586
rect 4542 584 4576 585
rect 4684 566 4714 648
rect 4820 617 4854 618
rect 4820 616 4821 617
rect 4744 586 4821 616
rect 4820 585 4821 586
rect 4853 616 4854 617
rect 4890 617 4924 618
rect 4890 616 4891 617
rect 4853 586 4856 616
rect 4888 586 4891 616
rect 4853 585 4854 586
rect 4820 584 4854 585
rect 4890 585 4891 586
rect 4923 616 4924 617
rect 4923 586 5002 616
rect 4923 585 4924 586
rect 4890 584 4924 585
rect 4472 547 4506 548
rect 4472 546 4473 547
rect 4396 516 4473 546
rect 4472 515 4473 516
rect 4505 546 4506 547
rect 4542 547 4576 548
rect 4542 546 4543 547
rect 4505 516 4508 546
rect 4540 516 4543 546
rect 4505 515 4506 516
rect 4472 514 4506 515
rect 4542 515 4543 516
rect 4575 546 4576 547
rect 4820 547 4854 548
rect 4820 546 4821 547
rect 4575 516 4654 546
rect 4575 515 4576 516
rect 4542 514 4576 515
rect 4684 484 4714 536
rect 4744 516 4821 546
rect 4820 515 4821 516
rect 4853 546 4854 547
rect 4890 547 4924 548
rect 4890 546 4891 547
rect 4853 516 4856 546
rect 4888 516 4891 546
rect 4853 515 4854 516
rect 4820 514 4854 515
rect 4890 515 4891 516
rect 4923 546 4924 547
rect 4923 516 5002 546
rect 4923 515 4924 516
rect 4890 514 4924 515
rect 5032 484 5062 648
rect 5168 617 5202 618
rect 5168 616 5169 617
rect 5092 586 5169 616
rect 5168 585 5169 586
rect 5201 616 5202 617
rect 5238 617 5272 618
rect 5238 616 5239 617
rect 5201 586 5204 616
rect 5236 586 5239 616
rect 5201 585 5202 586
rect 5168 584 5202 585
rect 5238 585 5239 586
rect 5271 616 5272 617
rect 5271 586 5350 616
rect 5271 585 5272 586
rect 5238 584 5272 585
rect 5168 547 5202 548
rect 5168 546 5169 547
rect 5092 516 5169 546
rect 5168 515 5169 516
rect 5201 546 5202 547
rect 5238 547 5272 548
rect 5238 546 5239 547
rect 5201 516 5204 546
rect 5236 516 5239 546
rect 5201 515 5202 516
rect 5168 514 5202 515
rect 5238 515 5239 516
rect 5271 546 5272 547
rect 5271 516 5350 546
rect 5271 515 5272 516
rect 5238 514 5272 515
rect 5380 484 5410 648
rect 5516 617 5550 618
rect 5516 616 5517 617
rect 5440 586 5517 616
rect 5516 585 5517 586
rect 5549 616 5550 617
rect 5586 617 5620 618
rect 5586 616 5587 617
rect 5549 586 5552 616
rect 5584 586 5587 616
rect 5549 585 5550 586
rect 5516 584 5550 585
rect 5586 585 5587 586
rect 5619 616 5620 617
rect 5619 586 5698 616
rect 5619 585 5620 586
rect 5586 584 5620 585
rect 5728 566 5758 648
rect 5864 617 5898 618
rect 5864 616 5865 617
rect 5788 586 5865 616
rect 5864 585 5865 586
rect 5897 616 5898 617
rect 5934 617 5968 618
rect 5934 616 5935 617
rect 5897 586 5900 616
rect 5932 586 5935 616
rect 5897 585 5898 586
rect 5864 584 5898 585
rect 5934 585 5935 586
rect 5967 616 5968 617
rect 5967 586 6046 616
rect 5967 585 5968 586
rect 5934 584 5968 585
rect 5516 547 5550 548
rect 5516 546 5517 547
rect 5440 516 5517 546
rect 5516 515 5517 516
rect 5549 546 5550 547
rect 5586 547 5620 548
rect 5586 546 5587 547
rect 5549 516 5552 546
rect 5584 516 5587 546
rect 5549 515 5550 516
rect 5516 514 5550 515
rect 5586 515 5587 516
rect 5619 546 5620 547
rect 5864 547 5898 548
rect 5864 546 5865 547
rect 5619 516 5698 546
rect 5619 515 5620 516
rect 5586 514 5620 515
rect 5728 484 5758 536
rect 5788 516 5865 546
rect 5864 515 5865 516
rect 5897 546 5898 547
rect 5934 547 5968 548
rect 5934 546 5935 547
rect 5897 516 5900 546
rect 5932 516 5935 546
rect 5897 515 5898 516
rect 5864 514 5898 515
rect 5934 515 5935 516
rect 5967 546 5968 547
rect 5967 516 6046 546
rect 5967 515 5968 516
rect 5934 514 5968 515
rect 6076 484 6106 648
rect 6212 617 6246 618
rect 6212 616 6213 617
rect 6136 586 6213 616
rect 6212 585 6213 586
rect 6245 616 6246 617
rect 6282 617 6316 618
rect 6282 616 6283 617
rect 6245 586 6248 616
rect 6280 586 6283 616
rect 6245 585 6246 586
rect 6212 584 6246 585
rect 6282 585 6283 586
rect 6315 616 6316 617
rect 6315 586 6394 616
rect 6315 585 6316 586
rect 6282 584 6316 585
rect 6424 566 6454 648
rect 6560 617 6594 618
rect 6560 616 6561 617
rect 6484 586 6561 616
rect 6560 585 6561 586
rect 6593 616 6594 617
rect 6630 617 6664 618
rect 6630 616 6631 617
rect 6593 586 6596 616
rect 6628 586 6631 616
rect 6593 585 6594 586
rect 6560 584 6594 585
rect 6630 585 6631 586
rect 6663 616 6664 617
rect 6663 586 6742 616
rect 6663 585 6664 586
rect 6630 584 6664 585
rect 6212 547 6246 548
rect 6212 546 6213 547
rect 6136 516 6213 546
rect 6212 515 6213 516
rect 6245 546 6246 547
rect 6282 547 6316 548
rect 6282 546 6283 547
rect 6245 516 6248 546
rect 6280 516 6283 546
rect 6245 515 6246 516
rect 6212 514 6246 515
rect 6282 515 6283 516
rect 6315 546 6316 547
rect 6560 547 6594 548
rect 6560 546 6561 547
rect 6315 516 6394 546
rect 6315 515 6316 516
rect 6282 514 6316 515
rect 6424 484 6454 536
rect 6484 516 6561 546
rect 6560 515 6561 516
rect 6593 546 6594 547
rect 6630 547 6664 548
rect 6630 546 6631 547
rect 6593 516 6596 546
rect 6628 516 6631 546
rect 6593 515 6594 516
rect 6560 514 6594 515
rect 6630 515 6631 516
rect 6663 546 6664 547
rect 6663 516 6742 546
rect 6663 515 6664 516
rect 6630 514 6664 515
rect 6772 484 6802 648
rect 6908 617 6942 618
rect 6908 616 6909 617
rect 6832 586 6909 616
rect 6908 585 6909 586
rect 6941 616 6942 617
rect 6978 617 7012 618
rect 6978 616 6979 617
rect 6941 586 6944 616
rect 6976 586 6979 616
rect 6941 585 6942 586
rect 6908 584 6942 585
rect 6978 585 6979 586
rect 7011 616 7012 617
rect 7011 586 7090 616
rect 7011 585 7012 586
rect 6978 584 7012 585
rect 6908 547 6942 548
rect 6908 546 6909 547
rect 6832 516 6909 546
rect 6908 515 6909 516
rect 6941 546 6942 547
rect 6978 547 7012 548
rect 6978 546 6979 547
rect 6941 516 6944 546
rect 6976 516 6979 546
rect 6941 515 6942 516
rect 6908 514 6942 515
rect 6978 515 6979 516
rect 7011 546 7012 547
rect 7011 516 7090 546
rect 7011 515 7012 516
rect 6978 514 7012 515
rect 7120 484 7150 648
rect 7256 617 7290 618
rect 7256 616 7257 617
rect 7180 586 7257 616
rect 7256 585 7257 586
rect 7289 616 7290 617
rect 7289 586 7292 616
rect 7289 585 7290 586
rect 7256 584 7290 585
rect 7256 547 7290 548
rect 7256 546 7257 547
rect 7180 516 7257 546
rect 7256 515 7257 516
rect 7289 546 7290 547
rect 7289 516 7292 546
rect 7289 515 7290 516
rect 7256 514 7290 515
rect 0 454 2406 484
rect 2436 454 2784 484
rect 2814 454 4146 484
rect 4176 454 4524 484
rect 4554 454 5886 484
rect 5916 454 6106 484
rect 6165 454 6264 484
rect 6294 454 7307 484
rect 18 423 52 424
rect 18 422 19 423
rect 16 392 19 422
rect 18 391 19 392
rect 51 422 52 423
rect 51 392 130 422
rect 51 391 52 392
rect 18 390 52 391
rect 160 360 190 454
rect 296 423 330 424
rect 296 422 297 423
rect 220 392 297 422
rect 296 391 297 392
rect 329 422 330 423
rect 366 423 400 424
rect 366 422 367 423
rect 329 392 332 422
rect 364 392 367 422
rect 329 391 330 392
rect 296 390 330 391
rect 366 391 367 392
rect 399 422 400 423
rect 399 392 478 422
rect 399 391 400 392
rect 366 390 400 391
rect 508 360 538 454
rect 644 423 678 424
rect 644 422 645 423
rect 568 392 645 422
rect 644 391 645 392
rect 677 422 678 423
rect 714 423 748 424
rect 714 422 715 423
rect 677 392 680 422
rect 712 392 715 422
rect 677 391 678 392
rect 644 390 678 391
rect 714 391 715 392
rect 747 422 748 423
rect 747 392 826 422
rect 747 391 748 392
rect 714 390 748 391
rect 856 360 886 454
rect 992 423 1026 424
rect 992 422 993 423
rect 916 392 993 422
rect 992 391 993 392
rect 1025 422 1026 423
rect 1062 423 1096 424
rect 1062 422 1063 423
rect 1025 392 1028 422
rect 1060 392 1063 422
rect 1025 391 1026 392
rect 992 390 1026 391
rect 1062 391 1063 392
rect 1095 422 1096 423
rect 1095 392 1174 422
rect 1095 391 1096 392
rect 1062 390 1096 391
rect 1204 360 1234 454
rect 1340 423 1374 424
rect 1340 422 1341 423
rect 1264 392 1341 422
rect 1340 391 1341 392
rect 1373 422 1374 423
rect 1410 423 1444 424
rect 1410 422 1411 423
rect 1373 392 1376 422
rect 1408 392 1411 422
rect 1373 391 1374 392
rect 1340 390 1374 391
rect 1410 391 1411 392
rect 1443 422 1444 423
rect 1443 392 1522 422
rect 1443 391 1444 392
rect 1410 390 1444 391
rect 1552 360 1582 454
rect 1688 423 1722 424
rect 1688 422 1689 423
rect 1612 392 1689 422
rect 1688 391 1689 392
rect 1721 422 1722 423
rect 1758 423 1792 424
rect 1758 422 1759 423
rect 1721 392 1724 422
rect 1756 392 1759 422
rect 1721 391 1722 392
rect 1688 390 1722 391
rect 1758 391 1759 392
rect 1791 422 1792 423
rect 1791 392 1870 422
rect 1791 391 1792 392
rect 1758 390 1792 391
rect 1900 360 1930 454
rect 2036 423 2070 424
rect 2036 422 2037 423
rect 1960 392 2037 422
rect 2036 391 2037 392
rect 2069 422 2070 423
rect 2106 423 2140 424
rect 2106 422 2107 423
rect 2069 392 2072 422
rect 2104 392 2107 422
rect 2069 391 2070 392
rect 2036 390 2070 391
rect 2106 391 2107 392
rect 2139 422 2140 423
rect 2139 392 2218 422
rect 2139 391 2140 392
rect 2106 390 2140 391
rect 2248 360 2278 454
rect 2384 423 2418 424
rect 2384 422 2385 423
rect 2308 392 2385 422
rect 2384 391 2385 392
rect 2417 422 2418 423
rect 2454 423 2488 424
rect 2454 422 2455 423
rect 2417 392 2420 422
rect 2452 392 2455 422
rect 2417 391 2418 392
rect 2384 390 2418 391
rect 2454 391 2455 392
rect 2487 422 2488 423
rect 2487 392 2566 422
rect 2487 391 2488 392
rect 2454 390 2488 391
rect 2596 360 2626 454
rect 2732 423 2766 424
rect 2732 422 2733 423
rect 2656 392 2733 422
rect 2732 391 2733 392
rect 2765 422 2766 423
rect 2802 423 2836 424
rect 2802 422 2803 423
rect 2765 392 2768 422
rect 2800 392 2803 422
rect 2765 391 2766 392
rect 2732 390 2766 391
rect 2802 391 2803 392
rect 2835 422 2836 423
rect 2835 392 2914 422
rect 2835 391 2836 392
rect 2802 390 2836 391
rect 2944 360 2974 454
rect 3080 423 3114 424
rect 3080 422 3081 423
rect 3004 392 3081 422
rect 3080 391 3081 392
rect 3113 422 3114 423
rect 3150 423 3184 424
rect 3150 422 3151 423
rect 3113 392 3116 422
rect 3148 392 3151 422
rect 3113 391 3114 392
rect 3080 390 3114 391
rect 3150 391 3151 392
rect 3183 422 3184 423
rect 3183 392 3262 422
rect 3183 391 3184 392
rect 3150 390 3184 391
rect 3292 360 3322 454
rect 3428 423 3462 424
rect 3428 422 3429 423
rect 3352 392 3429 422
rect 3428 391 3429 392
rect 3461 422 3462 423
rect 3498 423 3532 424
rect 3498 422 3499 423
rect 3461 392 3464 422
rect 3496 392 3499 422
rect 3461 391 3462 392
rect 3428 390 3462 391
rect 3498 391 3499 392
rect 3531 422 3532 423
rect 3531 392 3610 422
rect 3531 391 3532 392
rect 3498 390 3532 391
rect 3640 360 3670 454
rect 3776 423 3810 424
rect 3776 422 3777 423
rect 3700 392 3777 422
rect 3776 391 3777 392
rect 3809 422 3810 423
rect 3846 423 3880 424
rect 3846 422 3847 423
rect 3809 392 3812 422
rect 3844 392 3847 422
rect 3809 391 3810 392
rect 3776 390 3810 391
rect 3846 391 3847 392
rect 3879 422 3880 423
rect 3879 392 3958 422
rect 3879 391 3880 392
rect 3846 390 3880 391
rect 3988 360 4018 454
rect 4124 423 4158 424
rect 4124 422 4125 423
rect 4048 392 4125 422
rect 4124 391 4125 392
rect 4157 422 4158 423
rect 4194 423 4228 424
rect 4194 422 4195 423
rect 4157 392 4160 422
rect 4192 392 4195 422
rect 4157 391 4158 392
rect 4124 390 4158 391
rect 4194 391 4195 392
rect 4227 422 4228 423
rect 4227 392 4306 422
rect 4336 407 4366 454
rect 4472 423 4506 424
rect 4472 422 4473 423
rect 4396 392 4473 422
rect 4227 391 4228 392
rect 4194 390 4228 391
rect 4472 391 4473 392
rect 4505 422 4506 423
rect 4542 423 4576 424
rect 4542 422 4543 423
rect 4505 392 4508 422
rect 4540 392 4543 422
rect 4505 391 4506 392
rect 4472 390 4506 391
rect 4542 391 4543 392
rect 4575 422 4576 423
rect 4575 392 4654 422
rect 4575 391 4576 392
rect 4542 390 4576 391
rect 4684 360 4714 454
rect 4820 423 4854 424
rect 4820 422 4821 423
rect 4744 392 4821 422
rect 4820 391 4821 392
rect 4853 422 4854 423
rect 4890 423 4924 424
rect 4890 422 4891 423
rect 4853 392 4856 422
rect 4888 392 4891 422
rect 4853 391 4854 392
rect 4820 390 4854 391
rect 4890 391 4891 392
rect 4923 422 4924 423
rect 4923 392 5002 422
rect 4923 391 4924 392
rect 4890 390 4924 391
rect 5032 360 5062 454
rect 5168 423 5202 424
rect 5168 422 5169 423
rect 5092 392 5169 422
rect 5168 391 5169 392
rect 5201 422 5202 423
rect 5238 423 5272 424
rect 5238 422 5239 423
rect 5201 392 5204 422
rect 5236 392 5239 422
rect 5201 391 5202 392
rect 5168 390 5202 391
rect 5238 391 5239 392
rect 5271 422 5272 423
rect 5271 392 5350 422
rect 5271 391 5272 392
rect 5238 390 5272 391
rect 5380 360 5410 454
rect 5516 423 5550 424
rect 5516 422 5517 423
rect 5440 392 5517 422
rect 5516 391 5517 392
rect 5549 422 5550 423
rect 5586 423 5620 424
rect 5586 422 5587 423
rect 5549 392 5552 422
rect 5584 392 5587 422
rect 5549 391 5550 392
rect 5516 390 5550 391
rect 5586 391 5587 392
rect 5619 422 5620 423
rect 5619 392 5698 422
rect 5619 391 5620 392
rect 5586 390 5620 391
rect 5728 360 5758 454
rect 5864 423 5898 424
rect 5864 422 5865 423
rect 5788 392 5865 422
rect 5864 391 5865 392
rect 5897 422 5898 423
rect 5934 423 5968 424
rect 5934 422 5935 423
rect 5897 392 5900 422
rect 5932 392 5935 422
rect 5897 391 5898 392
rect 5864 390 5898 391
rect 5934 391 5935 392
rect 5967 422 5968 423
rect 6212 423 6246 424
rect 6212 422 6213 423
rect 5967 392 6046 422
rect 5967 391 5968 392
rect 5934 390 5968 391
rect 6076 360 6106 407
rect 6136 392 6213 422
rect 6212 391 6213 392
rect 6245 422 6246 423
rect 6282 423 6316 424
rect 6282 422 6283 423
rect 6245 392 6248 422
rect 6280 392 6283 422
rect 6245 391 6246 392
rect 6212 390 6246 391
rect 6282 391 6283 392
rect 6315 422 6316 423
rect 6315 392 6394 422
rect 6315 391 6316 392
rect 6282 390 6316 391
rect 6424 360 6454 454
rect 6560 423 6594 424
rect 6560 422 6561 423
rect 6484 392 6561 422
rect 6560 391 6561 392
rect 6593 422 6594 423
rect 6630 423 6664 424
rect 6630 422 6631 423
rect 6593 392 6596 422
rect 6628 392 6631 422
rect 6593 391 6594 392
rect 6560 390 6594 391
rect 6630 391 6631 392
rect 6663 422 6664 423
rect 6663 392 6742 422
rect 6663 391 6664 392
rect 6630 390 6664 391
rect 6772 360 6802 454
rect 6908 423 6942 424
rect 6908 422 6909 423
rect 6832 392 6909 422
rect 6908 391 6909 392
rect 6941 422 6942 423
rect 6978 423 7012 424
rect 6978 422 6979 423
rect 6941 392 6944 422
rect 6976 392 6979 422
rect 6941 391 6942 392
rect 6908 390 6942 391
rect 6978 391 6979 392
rect 7011 422 7012 423
rect 7011 392 7090 422
rect 7011 391 7012 392
rect 6978 390 7012 391
rect 7120 360 7150 454
rect 7256 423 7290 424
rect 7256 422 7257 423
rect 7180 392 7257 422
rect 7256 391 7257 392
rect 7289 422 7290 423
rect 7289 392 7292 422
rect 7289 391 7290 392
rect 7256 390 7290 391
rect 0 330 2406 360
rect 2436 330 2784 360
rect 2814 330 4146 360
rect 4176 330 4524 360
rect 4554 330 5886 360
rect 5916 330 6264 360
rect 6294 330 7307 360
rect 18 299 52 300
rect 18 298 19 299
rect 16 268 19 298
rect 18 267 19 268
rect 51 298 52 299
rect 51 268 130 298
rect 51 267 52 268
rect 18 266 52 267
rect 160 236 190 330
rect 296 299 330 300
rect 296 298 297 299
rect 220 268 297 298
rect 296 267 297 268
rect 329 298 330 299
rect 366 299 400 300
rect 366 298 367 299
rect 329 268 332 298
rect 364 268 367 298
rect 329 267 330 268
rect 296 266 330 267
rect 366 267 367 268
rect 399 298 400 299
rect 399 268 478 298
rect 399 267 400 268
rect 366 266 400 267
rect 508 236 538 330
rect 644 299 678 300
rect 644 298 645 299
rect 568 268 645 298
rect 644 267 645 268
rect 677 298 678 299
rect 714 299 748 300
rect 714 298 715 299
rect 677 268 680 298
rect 712 268 715 298
rect 677 267 678 268
rect 644 266 678 267
rect 714 267 715 268
rect 747 298 748 299
rect 747 268 826 298
rect 747 267 748 268
rect 714 266 748 267
rect 856 236 886 330
rect 992 299 1026 300
rect 992 298 993 299
rect 916 268 993 298
rect 992 267 993 268
rect 1025 298 1026 299
rect 1062 299 1096 300
rect 1062 298 1063 299
rect 1025 268 1028 298
rect 1060 268 1063 298
rect 1025 267 1026 268
rect 992 266 1026 267
rect 1062 267 1063 268
rect 1095 298 1096 299
rect 1095 268 1174 298
rect 1095 267 1096 268
rect 1062 266 1096 267
rect 1204 236 1234 330
rect 1340 299 1374 300
rect 1340 298 1341 299
rect 1264 268 1341 298
rect 1340 267 1341 268
rect 1373 298 1374 299
rect 1410 299 1444 300
rect 1410 298 1411 299
rect 1373 268 1376 298
rect 1408 268 1411 298
rect 1373 267 1374 268
rect 1340 266 1374 267
rect 1410 267 1411 268
rect 1443 298 1444 299
rect 1443 268 1522 298
rect 1443 267 1444 268
rect 1410 266 1444 267
rect 1552 236 1582 330
rect 1688 299 1722 300
rect 1688 298 1689 299
rect 1612 268 1689 298
rect 1688 267 1689 268
rect 1721 298 1722 299
rect 1758 299 1792 300
rect 1758 298 1759 299
rect 1721 268 1724 298
rect 1756 268 1759 298
rect 1721 267 1722 268
rect 1688 266 1722 267
rect 1758 267 1759 268
rect 1791 298 1792 299
rect 1791 268 1870 298
rect 1791 267 1792 268
rect 1758 266 1792 267
rect 1900 236 1930 330
rect 2036 299 2070 300
rect 2036 298 2037 299
rect 1960 268 2037 298
rect 2036 267 2037 268
rect 2069 298 2070 299
rect 2106 299 2140 300
rect 2106 298 2107 299
rect 2069 268 2072 298
rect 2104 268 2107 298
rect 2069 267 2070 268
rect 2036 266 2070 267
rect 2106 267 2107 268
rect 2139 298 2140 299
rect 2139 268 2218 298
rect 2139 267 2140 268
rect 2106 266 2140 267
rect 2248 236 2278 330
rect 2384 299 2418 300
rect 2384 298 2385 299
rect 2308 268 2385 298
rect 2384 267 2385 268
rect 2417 298 2418 299
rect 2454 299 2488 300
rect 2454 298 2455 299
rect 2417 268 2420 298
rect 2452 268 2455 298
rect 2417 267 2418 268
rect 2384 266 2418 267
rect 2454 267 2455 268
rect 2487 298 2488 299
rect 2487 268 2566 298
rect 2596 284 2626 330
rect 2732 299 2766 300
rect 2732 298 2733 299
rect 2656 268 2733 298
rect 2487 267 2488 268
rect 2454 266 2488 267
rect 2732 267 2733 268
rect 2765 298 2766 299
rect 2802 299 2836 300
rect 2802 298 2803 299
rect 2765 268 2768 298
rect 2800 268 2803 298
rect 2765 267 2766 268
rect 2732 266 2766 267
rect 2802 267 2803 268
rect 2835 298 2836 299
rect 2835 268 2914 298
rect 2835 267 2836 268
rect 2802 266 2836 267
rect 2944 236 2974 330
rect 3080 299 3114 300
rect 3080 298 3081 299
rect 3004 268 3081 298
rect 3080 267 3081 268
rect 3113 298 3114 299
rect 3150 299 3184 300
rect 3150 298 3151 299
rect 3113 268 3116 298
rect 3148 268 3151 298
rect 3113 267 3114 268
rect 3080 266 3114 267
rect 3150 267 3151 268
rect 3183 298 3184 299
rect 3183 268 3262 298
rect 3183 267 3184 268
rect 3150 266 3184 267
rect 3292 236 3322 330
rect 3428 299 3462 300
rect 3428 298 3429 299
rect 3352 268 3429 298
rect 3428 267 3429 268
rect 3461 298 3462 299
rect 3498 299 3532 300
rect 3498 298 3499 299
rect 3461 268 3464 298
rect 3496 268 3499 298
rect 3461 267 3462 268
rect 3428 266 3462 267
rect 3498 267 3499 268
rect 3531 298 3532 299
rect 3531 268 3610 298
rect 3531 267 3532 268
rect 3498 266 3532 267
rect 3640 236 3670 330
rect 3776 299 3810 300
rect 3776 298 3777 299
rect 3700 268 3777 298
rect 3776 267 3777 268
rect 3809 298 3810 299
rect 3846 299 3880 300
rect 3846 298 3847 299
rect 3809 268 3812 298
rect 3844 268 3847 298
rect 3809 267 3810 268
rect 3776 266 3810 267
rect 3846 267 3847 268
rect 3879 298 3880 299
rect 3879 268 3958 298
rect 3879 267 3880 268
rect 3846 266 3880 267
rect 3988 236 4018 330
rect 4124 299 4158 300
rect 4124 298 4125 299
rect 4048 268 4125 298
rect 4124 267 4125 268
rect 4157 298 4158 299
rect 4194 299 4228 300
rect 4194 298 4195 299
rect 4157 268 4160 298
rect 4192 268 4195 298
rect 4157 267 4158 268
rect 4124 266 4158 267
rect 4194 267 4195 268
rect 4227 298 4228 299
rect 4227 268 4306 298
rect 4227 267 4228 268
rect 4194 266 4228 267
rect 4336 236 4366 330
rect 4472 299 4506 300
rect 4472 298 4473 299
rect 4396 268 4473 298
rect 4472 267 4473 268
rect 4505 298 4506 299
rect 4542 299 4576 300
rect 4542 298 4543 299
rect 4505 268 4508 298
rect 4540 268 4543 298
rect 4505 267 4506 268
rect 4472 266 4506 267
rect 4542 267 4543 268
rect 4575 298 4576 299
rect 4575 268 4654 298
rect 4575 267 4576 268
rect 4542 266 4576 267
rect 4684 236 4714 330
rect 4820 299 4854 300
rect 4820 298 4821 299
rect 4744 268 4821 298
rect 4820 267 4821 268
rect 4853 298 4854 299
rect 4890 299 4924 300
rect 4890 298 4891 299
rect 4853 268 4856 298
rect 4888 268 4891 298
rect 4853 267 4854 268
rect 4820 266 4854 267
rect 4890 267 4891 268
rect 4923 298 4924 299
rect 4923 268 5002 298
rect 4923 267 4924 268
rect 4890 266 4924 267
rect 5032 236 5062 330
rect 5168 299 5202 300
rect 5168 298 5169 299
rect 5092 268 5169 298
rect 5168 267 5169 268
rect 5201 298 5202 299
rect 5238 299 5272 300
rect 5238 298 5239 299
rect 5201 268 5204 298
rect 5236 268 5239 298
rect 5201 267 5202 268
rect 5168 266 5202 267
rect 5238 267 5239 268
rect 5271 298 5272 299
rect 5271 268 5350 298
rect 5271 267 5272 268
rect 5238 266 5272 267
rect 5380 236 5410 330
rect 5516 299 5550 300
rect 5516 298 5517 299
rect 5440 268 5517 298
rect 5516 267 5517 268
rect 5549 298 5550 299
rect 5586 299 5620 300
rect 5586 298 5587 299
rect 5549 268 5552 298
rect 5584 268 5587 298
rect 5549 267 5550 268
rect 5516 266 5550 267
rect 5586 267 5587 268
rect 5619 298 5620 299
rect 5619 268 5698 298
rect 5619 267 5620 268
rect 5586 266 5620 267
rect 5728 236 5758 330
rect 5864 299 5898 300
rect 5864 298 5865 299
rect 5788 268 5865 298
rect 5864 267 5865 268
rect 5897 298 5898 299
rect 5934 299 5968 300
rect 5934 298 5935 299
rect 5897 268 5900 298
rect 5932 268 5935 298
rect 5897 267 5898 268
rect 5864 266 5898 267
rect 5934 267 5935 268
rect 5967 298 5968 299
rect 5967 268 6046 298
rect 5967 267 5968 268
rect 5934 266 5968 267
rect 6076 236 6106 330
rect 6212 299 6246 300
rect 6212 298 6213 299
rect 6136 268 6213 298
rect 6212 267 6213 268
rect 6245 298 6246 299
rect 6282 299 6316 300
rect 6282 298 6283 299
rect 6245 268 6248 298
rect 6280 268 6283 298
rect 6245 267 6246 268
rect 6212 266 6246 267
rect 6282 267 6283 268
rect 6315 298 6316 299
rect 6315 268 6394 298
rect 6315 267 6316 268
rect 6282 266 6316 267
rect 6424 236 6454 330
rect 6560 299 6594 300
rect 6560 298 6561 299
rect 6484 268 6561 298
rect 6560 267 6561 268
rect 6593 298 6594 299
rect 6630 299 6664 300
rect 6630 298 6631 299
rect 6593 268 6596 298
rect 6628 268 6631 298
rect 6593 267 6594 268
rect 6560 266 6594 267
rect 6630 267 6631 268
rect 6663 298 6664 299
rect 6663 268 6742 298
rect 6663 267 6664 268
rect 6630 266 6664 267
rect 6772 236 6802 330
rect 6908 299 6942 300
rect 6908 298 6909 299
rect 6832 268 6909 298
rect 6908 267 6909 268
rect 6941 298 6942 299
rect 6978 299 7012 300
rect 6978 298 6979 299
rect 6941 268 6944 298
rect 6976 268 6979 298
rect 6941 267 6942 268
rect 6908 266 6942 267
rect 6978 267 6979 268
rect 7011 298 7012 299
rect 7011 268 7090 298
rect 7011 267 7012 268
rect 6978 266 7012 267
rect 7120 236 7150 330
rect 7256 299 7290 300
rect 7256 298 7257 299
rect 7180 268 7257 298
rect 7256 267 7257 268
rect 7289 298 7290 299
rect 7289 268 7292 298
rect 7289 267 7290 268
rect 7256 266 7290 267
rect 0 206 2406 236
rect 2436 206 2784 236
rect 2814 206 4146 236
rect 4176 206 4524 236
rect 4554 206 5886 236
rect 5916 206 6264 236
rect 6294 206 7307 236
rect 18 175 52 176
rect 18 174 19 175
rect 16 144 19 174
rect 18 143 19 144
rect 51 174 52 175
rect 51 144 130 174
rect 51 143 52 144
rect 18 142 52 143
rect 160 112 190 206
rect 296 175 330 176
rect 296 174 297 175
rect 220 144 297 174
rect 296 143 297 144
rect 329 174 330 175
rect 366 175 400 176
rect 366 174 367 175
rect 329 144 332 174
rect 364 144 367 174
rect 329 143 330 144
rect 296 142 330 143
rect 366 143 367 144
rect 399 174 400 175
rect 399 144 478 174
rect 399 143 400 144
rect 366 142 400 143
rect 508 112 538 206
rect 644 175 678 176
rect 644 174 645 175
rect 568 144 645 174
rect 644 143 645 144
rect 677 174 678 175
rect 714 175 748 176
rect 714 174 715 175
rect 677 144 680 174
rect 712 144 715 174
rect 677 143 678 144
rect 644 142 678 143
rect 714 143 715 144
rect 747 174 748 175
rect 747 144 826 174
rect 747 143 748 144
rect 714 142 748 143
rect 856 112 886 206
rect 992 175 1026 176
rect 992 174 993 175
rect 916 144 993 174
rect 992 143 993 144
rect 1025 174 1026 175
rect 1062 175 1096 176
rect 1062 174 1063 175
rect 1025 144 1028 174
rect 1060 144 1063 174
rect 1025 143 1026 144
rect 992 142 1026 143
rect 1062 143 1063 144
rect 1095 174 1096 175
rect 1095 144 1174 174
rect 1095 143 1096 144
rect 1062 142 1096 143
rect 1204 112 1234 206
rect 1340 175 1374 176
rect 1340 174 1341 175
rect 1264 144 1341 174
rect 1340 143 1341 144
rect 1373 174 1374 175
rect 1410 175 1444 176
rect 1410 174 1411 175
rect 1373 144 1376 174
rect 1408 144 1411 174
rect 1373 143 1374 144
rect 1340 142 1374 143
rect 1410 143 1411 144
rect 1443 174 1444 175
rect 1443 144 1522 174
rect 1443 143 1444 144
rect 1410 142 1444 143
rect 1552 112 1582 206
rect 1688 175 1722 176
rect 1688 174 1689 175
rect 1612 144 1689 174
rect 1688 143 1689 144
rect 1721 174 1722 175
rect 1758 175 1792 176
rect 1758 174 1759 175
rect 1721 144 1724 174
rect 1756 144 1759 174
rect 1721 143 1722 144
rect 1688 142 1722 143
rect 1758 143 1759 144
rect 1791 174 1792 175
rect 1791 144 1870 174
rect 1791 143 1792 144
rect 1758 142 1792 143
rect 1900 112 1930 206
rect 2036 175 2070 176
rect 2036 174 2037 175
rect 1960 144 2037 174
rect 2036 143 2037 144
rect 2069 174 2070 175
rect 2106 175 2140 176
rect 2106 174 2107 175
rect 2069 144 2072 174
rect 2104 144 2107 174
rect 2069 143 2070 144
rect 2036 142 2070 143
rect 2106 143 2107 144
rect 2139 174 2140 175
rect 2139 144 2218 174
rect 2139 143 2140 144
rect 2106 142 2140 143
rect 2248 112 2278 206
rect 2384 175 2418 176
rect 2384 174 2385 175
rect 2308 144 2385 174
rect 2384 143 2385 144
rect 2417 174 2418 175
rect 2454 175 2488 176
rect 2454 174 2455 175
rect 2417 144 2420 174
rect 2452 144 2455 174
rect 2417 143 2418 144
rect 2384 142 2418 143
rect 2454 143 2455 144
rect 2487 174 2488 175
rect 2487 144 2566 174
rect 2487 143 2488 144
rect 2454 142 2488 143
rect 2596 112 2626 206
rect 2732 175 2766 176
rect 2732 174 2733 175
rect 2656 144 2733 174
rect 2732 143 2733 144
rect 2765 174 2766 175
rect 2802 175 2836 176
rect 2802 174 2803 175
rect 2765 144 2768 174
rect 2800 144 2803 174
rect 2765 143 2766 144
rect 2732 142 2766 143
rect 2802 143 2803 144
rect 2835 174 2836 175
rect 2835 144 2914 174
rect 2835 143 2836 144
rect 2802 142 2836 143
rect 2944 112 2974 206
rect 3080 175 3114 176
rect 3080 174 3081 175
rect 3004 144 3081 174
rect 3080 143 3081 144
rect 3113 174 3114 175
rect 3150 175 3184 176
rect 3150 174 3151 175
rect 3113 144 3116 174
rect 3148 144 3151 174
rect 3113 143 3114 144
rect 3080 142 3114 143
rect 3150 143 3151 144
rect 3183 174 3184 175
rect 3183 144 3262 174
rect 3183 143 3184 144
rect 3150 142 3184 143
rect 3292 112 3322 206
rect 3428 175 3462 176
rect 3428 174 3429 175
rect 3352 144 3429 174
rect 3428 143 3429 144
rect 3461 174 3462 175
rect 3498 175 3532 176
rect 3498 174 3499 175
rect 3461 144 3464 174
rect 3496 144 3499 174
rect 3461 143 3462 144
rect 3428 142 3462 143
rect 3498 143 3499 144
rect 3531 174 3532 175
rect 3531 144 3610 174
rect 3531 143 3532 144
rect 3498 142 3532 143
rect 3640 112 3670 206
rect 3776 175 3810 176
rect 3776 174 3777 175
rect 3700 144 3777 174
rect 3776 143 3777 144
rect 3809 174 3810 175
rect 3846 175 3880 176
rect 3846 174 3847 175
rect 3809 144 3812 174
rect 3844 144 3847 174
rect 3809 143 3810 144
rect 3776 142 3810 143
rect 3846 143 3847 144
rect 3879 174 3880 175
rect 3879 144 3958 174
rect 3879 143 3880 144
rect 3846 142 3880 143
rect 3988 112 4018 206
rect 4124 175 4158 176
rect 4124 174 4125 175
rect 4048 144 4125 174
rect 4124 143 4125 144
rect 4157 174 4158 175
rect 4194 175 4228 176
rect 4194 174 4195 175
rect 4157 144 4160 174
rect 4192 144 4195 174
rect 4157 143 4158 144
rect 4124 142 4158 143
rect 4194 143 4195 144
rect 4227 174 4228 175
rect 4227 144 4306 174
rect 4227 143 4228 144
rect 4194 142 4228 143
rect 4336 112 4366 206
rect 4472 175 4506 176
rect 4472 174 4473 175
rect 4396 144 4473 174
rect 4472 143 4473 144
rect 4505 174 4506 175
rect 4542 175 4576 176
rect 4542 174 4543 175
rect 4505 144 4508 174
rect 4540 144 4543 174
rect 4505 143 4506 144
rect 4472 142 4506 143
rect 4542 143 4543 144
rect 4575 174 4576 175
rect 4575 144 4654 174
rect 4575 143 4576 144
rect 4542 142 4576 143
rect 4684 112 4714 206
rect 4820 175 4854 176
rect 4820 174 4821 175
rect 4744 144 4821 174
rect 4820 143 4821 144
rect 4853 174 4854 175
rect 4890 175 4924 176
rect 4890 174 4891 175
rect 4853 144 4856 174
rect 4888 144 4891 174
rect 4853 143 4854 144
rect 4820 142 4854 143
rect 4890 143 4891 144
rect 4923 174 4924 175
rect 4923 144 5002 174
rect 4923 143 4924 144
rect 4890 142 4924 143
rect 5032 112 5062 206
rect 5168 175 5202 176
rect 5168 174 5169 175
rect 5092 144 5169 174
rect 5168 143 5169 144
rect 5201 174 5202 175
rect 5238 175 5272 176
rect 5238 174 5239 175
rect 5201 144 5204 174
rect 5236 144 5239 174
rect 5201 143 5202 144
rect 5168 142 5202 143
rect 5238 143 5239 144
rect 5271 174 5272 175
rect 5271 144 5350 174
rect 5271 143 5272 144
rect 5238 142 5272 143
rect 5380 112 5410 206
rect 5516 175 5550 176
rect 5516 174 5517 175
rect 5440 144 5517 174
rect 5516 143 5517 144
rect 5549 174 5550 175
rect 5586 175 5620 176
rect 5586 174 5587 175
rect 5549 144 5552 174
rect 5584 144 5587 174
rect 5549 143 5550 144
rect 5516 142 5550 143
rect 5586 143 5587 144
rect 5619 174 5620 175
rect 5619 144 5698 174
rect 5619 143 5620 144
rect 5586 142 5620 143
rect 5728 112 5758 206
rect 5864 175 5898 176
rect 5864 174 5865 175
rect 5788 144 5865 174
rect 5864 143 5865 144
rect 5897 174 5898 175
rect 5934 175 5968 176
rect 5934 174 5935 175
rect 5897 144 5900 174
rect 5932 144 5935 174
rect 5897 143 5898 144
rect 5864 142 5898 143
rect 5934 143 5935 144
rect 5967 174 5968 175
rect 5967 144 6046 174
rect 5967 143 5968 144
rect 5934 142 5968 143
rect 6076 112 6106 206
rect 6212 175 6246 176
rect 6212 174 6213 175
rect 6136 144 6213 174
rect 6212 143 6213 144
rect 6245 174 6246 175
rect 6282 175 6316 176
rect 6282 174 6283 175
rect 6245 144 6248 174
rect 6280 144 6283 174
rect 6245 143 6246 144
rect 6212 142 6246 143
rect 6282 143 6283 144
rect 6315 174 6316 175
rect 6315 144 6394 174
rect 6315 143 6316 144
rect 6282 142 6316 143
rect 6424 112 6454 206
rect 6560 175 6594 176
rect 6560 174 6561 175
rect 6484 144 6561 174
rect 6560 143 6561 144
rect 6593 174 6594 175
rect 6630 175 6664 176
rect 6630 174 6631 175
rect 6593 144 6596 174
rect 6628 144 6631 174
rect 6593 143 6594 144
rect 6560 142 6594 143
rect 6630 143 6631 144
rect 6663 174 6664 175
rect 6663 144 6742 174
rect 6663 143 6664 144
rect 6630 142 6664 143
rect 6772 112 6802 206
rect 6908 175 6942 176
rect 6908 174 6909 175
rect 6832 144 6909 174
rect 6908 143 6909 144
rect 6941 174 6942 175
rect 6978 175 7012 176
rect 6978 174 6979 175
rect 6941 144 6944 174
rect 6976 144 6979 174
rect 6941 143 6942 144
rect 6908 142 6942 143
rect 6978 143 6979 144
rect 7011 174 7012 175
rect 7011 144 7090 174
rect 7011 143 7012 144
rect 6978 142 7012 143
rect 7120 112 7150 206
rect 7256 175 7290 176
rect 7256 174 7257 175
rect 7180 144 7257 174
rect 7256 143 7257 144
rect 7289 174 7290 175
rect 7289 144 7292 174
rect 7289 143 7290 144
rect 7256 142 7290 143
rect 0 82 2406 112
rect 2436 82 2785 112
rect 2815 82 4146 112
rect 4176 82 4524 112
rect 4554 82 5886 112
rect 5916 82 6264 112
rect 6294 82 7307 112
rect 18 51 52 52
rect 18 50 19 51
rect 16 20 19 50
rect 18 19 19 20
rect 51 50 52 51
rect 51 20 130 50
rect 51 19 52 20
rect 18 18 52 19
rect 160 0 190 82
rect 296 51 330 52
rect 296 50 297 51
rect 220 20 297 50
rect 296 19 297 20
rect 329 50 330 51
rect 366 51 400 52
rect 366 50 367 51
rect 329 20 332 50
rect 364 20 367 50
rect 329 19 330 20
rect 296 18 330 19
rect 366 19 367 20
rect 399 50 400 51
rect 399 20 478 50
rect 399 19 400 20
rect 366 18 400 19
rect 508 0 538 82
rect 644 51 678 52
rect 644 50 645 51
rect 568 20 645 50
rect 644 19 645 20
rect 677 50 678 51
rect 714 51 748 52
rect 714 50 715 51
rect 677 20 680 50
rect 712 20 715 50
rect 677 19 678 20
rect 644 18 678 19
rect 714 19 715 20
rect 747 50 748 51
rect 747 20 826 50
rect 747 19 748 20
rect 714 18 748 19
rect 856 0 886 82
rect 992 51 1026 52
rect 992 50 993 51
rect 916 20 993 50
rect 992 19 993 20
rect 1025 50 1026 51
rect 1062 51 1096 52
rect 1062 50 1063 51
rect 1025 20 1028 50
rect 1060 20 1063 50
rect 1025 19 1026 20
rect 992 18 1026 19
rect 1062 19 1063 20
rect 1095 50 1096 51
rect 1095 20 1174 50
rect 1095 19 1096 20
rect 1062 18 1096 19
rect 1204 0 1234 82
rect 1340 51 1374 52
rect 1340 50 1341 51
rect 1264 20 1341 50
rect 1340 19 1341 20
rect 1373 50 1374 51
rect 1410 51 1444 52
rect 1410 50 1411 51
rect 1373 20 1376 50
rect 1408 20 1411 50
rect 1373 19 1374 20
rect 1340 18 1374 19
rect 1410 19 1411 20
rect 1443 50 1444 51
rect 1443 20 1522 50
rect 1443 19 1444 20
rect 1410 18 1444 19
rect 1552 0 1582 82
rect 1688 51 1722 52
rect 1688 50 1689 51
rect 1612 20 1689 50
rect 1688 19 1689 20
rect 1721 50 1722 51
rect 1758 51 1792 52
rect 1758 50 1759 51
rect 1721 20 1724 50
rect 1756 20 1759 50
rect 1721 19 1722 20
rect 1688 18 1722 19
rect 1758 19 1759 20
rect 1791 50 1792 51
rect 1791 20 1870 50
rect 1791 19 1792 20
rect 1758 18 1792 19
rect 1900 0 1930 82
rect 2036 51 2070 52
rect 2036 50 2037 51
rect 1960 20 2037 50
rect 2036 19 2037 20
rect 2069 50 2070 51
rect 2106 51 2140 52
rect 2106 50 2107 51
rect 2069 20 2072 50
rect 2104 20 2107 50
rect 2069 19 2070 20
rect 2036 18 2070 19
rect 2106 19 2107 20
rect 2139 50 2140 51
rect 2139 20 2218 50
rect 2139 19 2140 20
rect 2106 18 2140 19
rect 2248 0 2278 82
rect 2384 51 2418 52
rect 2384 50 2385 51
rect 2308 20 2385 50
rect 2384 19 2385 20
rect 2417 50 2418 51
rect 2454 51 2488 52
rect 2454 50 2455 51
rect 2417 20 2420 50
rect 2452 20 2455 50
rect 2417 19 2418 20
rect 2384 18 2418 19
rect 2454 19 2455 20
rect 2487 50 2488 51
rect 2487 20 2566 50
rect 2487 19 2488 20
rect 2454 18 2488 19
rect 2596 0 2626 82
rect 2732 51 2766 52
rect 2732 50 2733 51
rect 2656 20 2733 50
rect 2732 19 2733 20
rect 2765 50 2766 51
rect 2802 51 2836 52
rect 2802 50 2803 51
rect 2765 20 2768 50
rect 2800 20 2803 50
rect 2765 19 2766 20
rect 2732 18 2766 19
rect 2802 19 2803 20
rect 2835 50 2836 51
rect 2835 20 2914 50
rect 2835 19 2836 20
rect 2802 18 2836 19
rect 2944 0 2974 82
rect 3080 51 3114 52
rect 3080 50 3081 51
rect 3004 20 3081 50
rect 3080 19 3081 20
rect 3113 50 3114 51
rect 3150 51 3184 52
rect 3150 50 3151 51
rect 3113 20 3116 50
rect 3148 20 3151 50
rect 3113 19 3114 20
rect 3080 18 3114 19
rect 3150 19 3151 20
rect 3183 50 3184 51
rect 3183 20 3262 50
rect 3183 19 3184 20
rect 3150 18 3184 19
rect 3292 0 3322 82
rect 3428 51 3462 52
rect 3428 50 3429 51
rect 3352 20 3429 50
rect 3428 19 3429 20
rect 3461 50 3462 51
rect 3498 51 3532 52
rect 3498 50 3499 51
rect 3461 20 3464 50
rect 3496 20 3499 50
rect 3461 19 3462 20
rect 3428 18 3462 19
rect 3498 19 3499 20
rect 3531 50 3532 51
rect 3531 20 3610 50
rect 3531 19 3532 20
rect 3498 18 3532 19
rect 3640 0 3670 82
rect 3776 51 3810 52
rect 3776 50 3777 51
rect 3700 20 3777 50
rect 3776 19 3777 20
rect 3809 50 3810 51
rect 3846 51 3880 52
rect 3846 50 3847 51
rect 3809 20 3812 50
rect 3844 20 3847 50
rect 3809 19 3810 20
rect 3776 18 3810 19
rect 3846 19 3847 20
rect 3879 50 3880 51
rect 3879 20 3958 50
rect 3879 19 3880 20
rect 3846 18 3880 19
rect 3988 0 4018 82
rect 4124 51 4158 52
rect 4124 50 4125 51
rect 4048 20 4125 50
rect 4124 19 4125 20
rect 4157 50 4158 51
rect 4194 51 4228 52
rect 4194 50 4195 51
rect 4157 20 4160 50
rect 4192 20 4195 50
rect 4157 19 4158 20
rect 4124 18 4158 19
rect 4194 19 4195 20
rect 4227 50 4228 51
rect 4227 20 4306 50
rect 4227 19 4228 20
rect 4194 18 4228 19
rect 4336 0 4366 82
rect 4472 51 4506 52
rect 4472 50 4473 51
rect 4396 20 4473 50
rect 4472 19 4473 20
rect 4505 50 4506 51
rect 4542 51 4576 52
rect 4542 50 4543 51
rect 4505 20 4508 50
rect 4540 20 4543 50
rect 4505 19 4506 20
rect 4472 18 4506 19
rect 4542 19 4543 20
rect 4575 50 4576 51
rect 4575 20 4654 50
rect 4575 19 4576 20
rect 4542 18 4576 19
rect 4684 0 4714 82
rect 4820 51 4854 52
rect 4820 50 4821 51
rect 4744 20 4821 50
rect 4820 19 4821 20
rect 4853 50 4854 51
rect 4890 51 4924 52
rect 4890 50 4891 51
rect 4853 20 4856 50
rect 4888 20 4891 50
rect 4853 19 4854 20
rect 4820 18 4854 19
rect 4890 19 4891 20
rect 4923 50 4924 51
rect 4923 20 5002 50
rect 4923 19 4924 20
rect 4890 18 4924 19
rect 5032 0 5062 82
rect 5168 51 5202 52
rect 5168 50 5169 51
rect 5092 20 5169 50
rect 5168 19 5169 20
rect 5201 50 5202 51
rect 5238 51 5272 52
rect 5238 50 5239 51
rect 5201 20 5204 50
rect 5236 20 5239 50
rect 5201 19 5202 20
rect 5168 18 5202 19
rect 5238 19 5239 20
rect 5271 50 5272 51
rect 5271 20 5350 50
rect 5271 19 5272 20
rect 5238 18 5272 19
rect 5380 0 5410 82
rect 5516 51 5550 52
rect 5516 50 5517 51
rect 5440 20 5517 50
rect 5516 19 5517 20
rect 5549 50 5550 51
rect 5586 51 5620 52
rect 5586 50 5587 51
rect 5549 20 5552 50
rect 5584 20 5587 50
rect 5549 19 5550 20
rect 5516 18 5550 19
rect 5586 19 5587 20
rect 5619 50 5620 51
rect 5619 20 5698 50
rect 5619 19 5620 20
rect 5586 18 5620 19
rect 5728 0 5758 82
rect 5864 51 5898 52
rect 5864 50 5865 51
rect 5788 20 5865 50
rect 5864 19 5865 20
rect 5897 50 5898 51
rect 5934 51 5968 52
rect 5934 50 5935 51
rect 5897 20 5900 50
rect 5932 20 5935 50
rect 5897 19 5898 20
rect 5864 18 5898 19
rect 5934 19 5935 20
rect 5967 50 5968 51
rect 5967 20 6046 50
rect 5967 19 5968 20
rect 5934 18 5968 19
rect 6076 0 6106 82
rect 6212 51 6246 52
rect 6212 50 6213 51
rect 6136 20 6213 50
rect 6212 19 6213 20
rect 6245 50 6246 51
rect 6282 51 6316 52
rect 6282 50 6283 51
rect 6245 20 6248 50
rect 6280 20 6283 50
rect 6245 19 6246 20
rect 6212 18 6246 19
rect 6282 19 6283 20
rect 6315 50 6316 51
rect 6315 20 6394 50
rect 6315 19 6316 20
rect 6282 18 6316 19
rect 6424 0 6454 82
rect 6560 51 6594 52
rect 6560 50 6561 51
rect 6484 20 6561 50
rect 6560 19 6561 20
rect 6593 50 6594 51
rect 6630 51 6664 52
rect 6630 50 6631 51
rect 6593 20 6596 50
rect 6628 20 6631 50
rect 6593 19 6594 20
rect 6560 18 6594 19
rect 6630 19 6631 20
rect 6663 50 6664 51
rect 6663 20 6742 50
rect 6663 19 6664 20
rect 6630 18 6664 19
rect 6772 0 6802 82
rect 6908 51 6942 52
rect 6908 50 6909 51
rect 6832 20 6909 50
rect 6908 19 6909 20
rect 6941 50 6942 51
rect 6978 51 7012 52
rect 6978 50 6979 51
rect 6941 20 6944 50
rect 6976 20 6979 50
rect 6941 19 6942 20
rect 6908 18 6942 19
rect 6978 19 6979 20
rect 7011 50 7012 51
rect 7011 20 7090 50
rect 7011 19 7012 20
rect 6978 18 7012 19
rect 7120 0 7150 82
rect 7256 51 7290 52
rect 7256 50 7257 51
rect 7180 20 7257 50
rect 7256 19 7257 20
rect 7289 50 7290 51
rect 7289 20 7292 50
rect 7289 19 7290 20
rect 7256 18 7290 19
<< comment >>
rect 382 637 1325 1639
rect 2119 651 3062 1653
rect 3840 644 4783 1646
rect 5606 651 6549 1653
<< labels >>
rlabel metal4 0 206 0 236 7 dummy_top
rlabel metal2 14 142 14 172 7 dummy_bot
rlabel metal4 348 648 348 678 7 top_8
rlabel metal2 362 601 362 631 7 bot_8
rlabel metal4 2088 648 2088 678 7 top_4
rlabel metal2 2102 592 2102 622 7 bot_4
rlabel metal4 3828 648 3828 678 7 top_2
rlabel metal2 3842 605 3842 635 7 bot_2
rlabel metal4 5568 648 5568 678 7 top_1
rlabel metal2 5582 608 5582 638 7 bot_1
<< end >>
