magic
tech sky130A
magscale 1 2
timestamp 1658921500
<< nwell >>
rect 234 1182 1042 1322
rect 234 1152 742 1182
rect 818 1174 852 1182
rect 234 1144 404 1152
rect 464 1144 742 1152
rect 234 1130 742 1144
rect 234 1094 418 1130
rect 452 1094 742 1130
rect 234 984 742 1094
rect 908 1068 954 1154
rect 964 984 1042 1182
rect 234 978 1042 984
rect 468 950 532 978
<< pdiff >>
rect 406 1130 464 1144
rect 406 1094 418 1130
rect 452 1094 464 1130
rect 406 1010 464 1094
rect 908 1068 954 1154
<< psubdiff >>
rect 322 590 370 624
rect 404 590 466 624
rect 500 590 570 624
rect 604 590 674 624
rect 708 590 768 624
rect 802 590 866 624
rect 900 590 932 624
<< nsubdiff >>
rect 442 1280 946 1286
rect 442 1246 466 1280
rect 500 1246 570 1280
rect 604 1246 674 1280
rect 708 1246 770 1280
rect 804 1246 864 1280
rect 898 1246 946 1280
rect 442 1240 946 1246
<< psubdiffcont >>
rect 370 590 404 624
rect 466 590 500 624
rect 570 590 604 624
rect 674 590 708 624
rect 768 590 802 624
rect 866 590 900 624
<< nsubdiffcont >>
rect 466 1246 500 1280
rect 570 1246 604 1280
rect 674 1246 708 1280
rect 770 1246 804 1280
rect 864 1246 898 1280
<< poly >>
rect 352 1260 420 1270
rect 352 1224 368 1260
rect 404 1224 420 1260
rect 352 1160 420 1224
rect 372 804 402 1160
rect 868 1000 898 1004
rect 468 950 498 990
rect 676 978 706 998
rect 634 958 706 978
rect 468 930 536 950
rect 468 892 486 930
rect 520 892 536 930
rect 468 794 536 892
rect 634 924 650 958
rect 684 924 706 958
rect 634 890 706 924
rect 748 968 816 990
rect 868 970 974 1000
rect 748 934 764 968
rect 800 934 816 968
rect 748 922 816 934
rect 906 962 974 970
rect 906 928 922 962
rect 958 928 974 962
rect 906 918 974 928
rect 634 856 650 890
rect 684 856 706 890
rect 784 868 816 872
rect 634 840 706 856
rect 676 776 706 840
rect 748 852 816 868
rect 748 818 764 852
rect 800 818 816 852
rect 748 804 816 818
rect 868 662 1028 678
rect 868 648 984 662
rect 974 628 984 648
rect 1018 628 1028 662
rect 974 612 1028 628
<< polycont >>
rect 368 1224 404 1260
rect 486 892 520 930
rect 650 924 684 958
rect 764 934 800 968
rect 922 928 958 962
rect 650 856 684 890
rect 764 818 800 852
rect 984 628 1018 662
<< locali >>
rect 254 1148 288 1328
rect 442 1280 946 1286
rect 368 1260 404 1276
rect 442 1246 466 1280
rect 500 1246 570 1280
rect 604 1246 674 1280
rect 708 1246 770 1280
rect 804 1246 864 1280
rect 898 1246 946 1280
rect 442 1240 946 1246
rect 368 1214 404 1224
rect 368 1180 370 1214
rect 514 1154 626 1180
rect 722 1164 756 1240
rect 818 1174 852 1204
rect 514 1148 660 1154
rect 254 982 322 1148
rect 548 1142 660 1148
rect 548 1106 572 1142
rect 606 1106 638 1142
rect 548 1064 660 1106
rect 548 1028 572 1064
rect 606 1028 638 1064
rect 548 1012 660 1028
rect 254 708 288 982
rect 418 782 452 994
rect 548 980 588 1012
rect 818 1002 852 1026
rect 486 930 520 946
rect 486 856 520 892
rect 486 816 520 822
rect 554 850 588 980
rect 748 934 764 968
rect 800 934 884 968
rect 650 890 684 924
rect 554 816 616 850
rect 650 840 684 856
rect 748 852 784 866
rect 748 818 764 852
rect 800 818 816 852
rect 850 850 884 934
rect 922 962 958 978
rect 922 918 958 928
rect 994 850 1028 1328
rect 850 816 1028 850
rect 582 782 616 816
rect 322 778 368 782
rect 322 744 334 778
rect 322 734 368 744
rect 582 778 660 782
rect 582 744 598 778
rect 632 744 660 778
rect 582 742 660 744
rect 722 766 756 782
rect 332 690 356 734
rect 514 702 548 740
rect 254 570 288 674
rect 514 662 548 668
rect 818 624 852 782
rect 914 766 948 782
rect 994 678 1028 816
rect 980 662 1028 678
rect 980 628 984 662
rect 1018 628 1028 662
rect 322 590 370 624
rect 404 590 466 624
rect 500 590 570 624
rect 604 590 674 624
rect 708 590 768 624
rect 802 590 866 624
rect 900 590 932 624
rect 980 612 1028 628
rect 994 570 1028 612
<< viali >>
rect 466 1246 500 1280
rect 570 1246 604 1280
rect 674 1246 708 1280
rect 770 1246 804 1280
rect 864 1246 898 1280
rect 370 1180 404 1214
rect 418 1094 452 1130
rect 572 1106 606 1142
rect 914 1106 948 1142
rect 418 1016 452 1052
rect 572 1028 606 1064
rect 914 1028 948 1064
rect 486 822 520 856
rect 650 958 684 974
rect 650 940 684 958
rect 748 866 784 900
rect 922 884 958 918
rect 334 744 368 778
rect 598 744 632 778
rect 254 674 288 708
rect 722 732 756 766
rect 514 668 548 702
rect 914 732 948 766
rect 370 590 404 624
rect 466 590 500 624
rect 570 590 604 624
rect 674 590 708 624
rect 768 590 802 624
rect 866 590 900 624
<< metal1 >>
rect 234 1280 1042 1296
rect 234 1248 466 1280
rect 234 1240 336 1248
rect 438 1246 466 1248
rect 500 1246 570 1280
rect 604 1246 674 1280
rect 708 1246 770 1280
rect 804 1246 864 1280
rect 898 1246 1042 1280
rect 438 1240 1042 1246
rect 358 1214 416 1220
rect 358 1212 370 1214
rect 234 1182 370 1212
rect 358 1180 370 1182
rect 404 1212 416 1214
rect 404 1182 1042 1212
rect 404 1180 416 1182
rect 358 1174 416 1180
rect 406 1140 464 1144
rect 566 1142 612 1154
rect 404 1088 410 1140
rect 462 1088 468 1140
rect 404 1062 468 1088
rect 404 1010 410 1062
rect 462 1010 468 1062
rect 566 1106 572 1142
rect 606 1108 612 1142
rect 908 1142 954 1154
rect 908 1108 914 1142
rect 606 1106 914 1108
rect 948 1106 954 1142
rect 566 1080 954 1106
rect 566 1064 612 1080
rect 566 1028 572 1064
rect 606 1028 612 1064
rect 566 1016 612 1028
rect 908 1064 954 1080
rect 908 1028 914 1064
rect 948 1028 954 1064
rect 908 1016 954 1028
rect 914 1010 948 1016
rect 234 974 1042 982
rect 234 954 650 974
rect 636 940 650 954
rect 684 954 1042 974
rect 684 940 694 954
rect 636 928 694 940
rect 306 900 590 920
rect 910 918 970 926
rect 734 900 796 906
rect 910 900 922 918
rect 234 890 748 900
rect 234 872 334 890
rect 562 872 748 890
rect 734 866 748 872
rect 784 884 922 900
rect 958 900 970 918
rect 958 884 1042 900
rect 784 872 1042 884
rect 784 866 796 872
rect 474 856 532 862
rect 734 860 796 866
rect 474 844 486 856
rect 234 822 486 844
rect 520 844 532 856
rect 520 832 706 844
rect 876 832 1042 844
rect 520 822 1042 832
rect 234 816 1042 822
rect 474 810 532 816
rect 670 804 956 816
rect 322 778 380 788
rect 322 744 334 778
rect 368 770 380 778
rect 586 778 644 788
rect 586 770 598 778
rect 368 744 598 770
rect 632 744 644 778
rect 322 742 644 744
rect 322 734 380 742
rect 586 734 644 742
rect 710 766 960 774
rect 710 732 722 766
rect 756 732 914 766
rect 948 732 960 766
rect 710 726 960 732
rect 248 708 294 720
rect 248 690 254 708
rect 234 674 254 690
rect 288 690 294 708
rect 508 702 556 714
rect 508 690 514 702
rect 288 674 514 690
rect 234 668 514 674
rect 548 690 556 702
rect 548 668 1042 690
rect 234 662 1042 668
rect 234 624 1042 634
rect 234 590 370 624
rect 404 590 466 624
rect 500 590 570 624
rect 604 590 674 624
rect 708 590 768 624
rect 802 590 866 624
rect 900 590 1042 624
rect 234 578 1042 590
<< via1 >>
rect 410 1130 462 1140
rect 410 1094 418 1130
rect 418 1094 452 1130
rect 452 1094 462 1130
rect 410 1088 462 1094
rect 410 1052 462 1062
rect 410 1016 418 1052
rect 418 1016 452 1052
rect 452 1016 462 1052
rect 410 1010 462 1016
<< metal2 >>
rect 404 1140 468 1144
rect 404 1088 410 1140
rect 462 1088 468 1140
rect 404 1062 468 1088
rect 404 1010 410 1062
rect 462 1010 468 1062
rect 404 1000 468 1010
use sky130_fd_pr__nfet_01v8_J7MSU8  sky130_fd_pr__nfet_01v8_J7MSU8_0
timestamp 1658837386
transform 1 0 787 0 1 736
box -173 -68 173 68
use sky130_fd_pr__nfet_01v8_MJPTSJ  sky130_fd_pr__nfet_01v8_MJPTSJ_0
timestamp 1658840561
transform 1 0 435 0 1 736
box -125 -68 125 68
use sky130_fd_pr__pfet_01v8_5CE3MA  sky130_fd_pr__pfet_01v8_5CE3MA_0
timestamp 1658837386
transform 1 0 787 0 1 1096
box -209 -116 209 116
use sky130_fd_pr__pfet_01v8_5CSGFE  sky130_fd_pr__pfet_01v8_5CSGFE_0
timestamp 1658918966
transform 1 0 435 0 1 1064
box -161 -116 161 116
<< labels >>
rlabel metal1 234 872 234 900 7 col_n
rlabel metal1 234 954 234 982 7 colon_n
rlabel metal1 234 662 234 690 7 vcom
rlabel metal1 234 1182 234 1212 7 sample_n
rlabel metal1 234 816 234 844 7 sample
rlabel metal1 234 578 234 634 7 VSS
rlabel metal1 234 1240 234 1296 7 VDD
rlabel locali 818 1002 852 1002 5 vint1
rlabel locali 994 574 1028 574 5 row_n
<< end >>
