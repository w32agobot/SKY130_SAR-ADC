* SPICE3 file created from adc_array_wafflecap_16_6420x6420nm.ext - technology: sky130A

.subckt adc_array_wafflecap_16_6420x6420nm ctop cbot
C0 cbot ctop 8.71fF
C1 cbot VSUBS 2.76fF
.ends
