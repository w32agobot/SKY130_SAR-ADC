* NGSPICE file created from adc_array_matrix_12bit.ext - technology: sky130A

.subckt adc_array_wafflecap_dummy vcom ctop col col_n row_n rowon_n sample sample_n
+ off_n cbot VDD VSS
X0 VDD rowon_n a_170_212# VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1 a_662_574# col_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2 a_170_212# row_n a_662_574# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3 a_566_252# rowon_n a_170_212# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4 VSS row_n a_566_252# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5 a_566_252# col_n VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_262_212# sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=2.48e+11p ps=2.22e+06u w=800000u l=150000u
X7 a_170_212# sample a_262_212# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8 a_262_212# sample_n a_170_212# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X9 vcom sample a_262_212# VSS sky130_fd_pr__nfet_01v8 ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
.ends

.subckt adc_array_wafflecap_1 vcom ctop col col_n row_n rowon_n sample sample_n off_n
+ a_482_57# cbot VDD VSS
X0 VDD a_482_57# a_170_212# VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1 a_662_574# a_482_57# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2 a_170_212# a_482_57# a_662_574# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3 a_566_252# a_482_57# a_170_212# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4 VSS a_482_57# a_566_252# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5 a_566_252# a_482_57# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 cbot sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=2.48e+11p ps=2.22e+06u w=800000u l=150000u
X7 a_170_212# sample cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8 cbot sample_n a_170_212# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X9 vcom sample cbot VSS sky130_fd_pr__nfet_01v8 ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
C6 ctop cbot 0.36fF
.ends

.subckt adc_array_wafflecap_drv vcom ctop col col_n row_n rowon_n sample_i sample_o
+ sample_n_i sample_n_o off_n cbot VDD VSS
X0 VSS sample_i sample_n_o VSS sky130_fd_pr__nfet_01v8 ad=5.208e+11p pd=5.84e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1 sample_n_o sample_i VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VDD sample_i sample_n_o VDD sky130_fd_pr__pfet_01v8 ad=9.92e+11p pd=8.88e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3 sample_n_o sample_i VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4 sample_o sample_n_i VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5 VSS sample_n_i sample_o VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 sample_o sample_n_i VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X7 VDD sample_n_i sample_o VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
.ends

.subckt adc_array_wafflecap_8 vcom ctop col col_n row_n rowon_n sample sample_n off_n
+ VDD VSS
X0 VDD rowon_n a_170_212# VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1 a_662_574# col_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2 a_170_212# row_n a_662_574# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3 a_566_252# rowon_n a_170_212# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4 VSS row_n a_566_252# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5 a_566_252# col_n VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 cbot sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=2.48e+11p ps=2.22e+06u w=800000u l=150000u
X7 a_170_212# sample cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8 cbot sample_n a_170_212# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X9 vcom sample cbot VSS sky130_fd_pr__nfet_01v8 ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
C1 ctop cbot 2.89fF
.ends

.subckt adc_noise_decoup_cell1 nmoscap_top nmoscap_bot mimcap_top mimcap_bot pwell
X0 mimcap_top mimcap_bot sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X1 nmoscap_bot nmoscap_top nmoscap_bot pwell sky130_fd_pr__nfet_01v8 ad=2.296e+13p pd=6.84e+07u as=0p ps=0u w=1.64e+07u l=1.6e+07u
.ends

.subckt adc_array_wafflecap_4 vcom ctop col col_n row_n rowon_n sample sample_n off_n
+ a_482_57# cbot VDD VSS
X0 VDD a_482_57# a_170_212# VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1 a_662_574# a_482_57# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2 a_170_212# a_482_57# a_662_574# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3 a_566_252# a_482_57# a_170_212# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4 VSS a_482_57# a_566_252# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5 a_566_252# a_482_57# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 cbot sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=2.48e+11p ps=2.22e+06u w=800000u l=150000u
X7 a_170_212# sample cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8 cbot sample_n a_170_212# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X9 vcom sample cbot VSS sky130_fd_pr__nfet_01v8 ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
C3 ctop cbot 1.46fF
.ends

.subckt adc_array_wafflecap_2 vcom ctop col col_n row_n rowon_n sample sample_n off_n
+ a_482_57# cbot VDD VSS
X0 VDD a_482_57# a_170_212# VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1 a_662_574# a_482_57# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2 a_170_212# a_482_57# a_662_574# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3 a_566_252# a_482_57# a_170_212# VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4 VSS a_482_57# a_566_252# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5 a_566_252# a_482_57# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 cbot sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=2.48e+11p ps=2.22e+06u w=800000u l=150000u
X7 a_170_212# sample cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X8 cbot sample_n a_170_212# VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X9 vcom sample cbot VSS sky130_fd_pr__nfet_01v8 ad=1.302e+11p pd=1.46e+06u as=0p ps=0u w=420000u l=150000u
C4 ctop cbot 0.72fF
.ends

.subckt adc_array_wafflecap_gate sample_n rowon_n row_n vcom col_n analog_in sw sw_n
+ m2_32_32# m1_0_568# m1_0_374# li_856_970# a_169_51# VDD VSS li_34_0#
X0 a_169_51# sw_n analog_in VDD sky130_fd_pr__pfet_01v8 ad=2.7075e+12p pd=2.185e+07u as=1.102e+12p ps=8.76e+06u w=1.9e+06u l=220000u
X1 analog_in sw a_169_51# VSS sky130_fd_pr__nfet_01v8 ad=1.102e+12p pd=8.76e+06u as=2.7645e+12p ps=2.191e+07u w=1.9e+06u l=220000u
X2 analog_in sw_n a_169_51# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.9e+06u l=220000u
X3 a_169_51# sw_n analog_in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.9e+06u l=220000u
X4 a_169_51# sw_n a_169_51# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.9e+06u l=220000u
X5 a_169_51# sw analog_in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.9e+06u l=220000u
X6 a_169_51# sw analog_in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.9e+06u l=220000u
X7 a_169_51# sw a_169_51# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.9e+06u l=220000u
X8 analog_in sw a_169_51# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.9e+06u l=220000u
X9 a_169_51# sw a_169_51# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.9e+06u l=220000u
X10 a_169_51# sw_n a_169_51# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.9e+06u l=220000u
X11 analog_in sw_n a_169_51# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.9e+06u l=220000u
.ends

.subckt adc_array_matrix_12bit VDD VSS vcm sample sample_n row_n[0] row_n[1] row_n[2] row_n[3]
+ row_n[4] row_n[5] row_n[6] row_n[7] row_n[8] row_n[9] row_n[10] row_n[11] row_n[12] row_n[13] row_n[14]
+ row_n[15] rowon_n[0] rowon_n[1] rowon_n[2] rowon_n[3] rowon_n[4] rowon_n[5] rowon_n[6] rowon_n[7] rowon_n[8]
+ rowon_n[9] rowon_n[10] rowon_n[11] rowon_n[12] rowon_n[13] rowon_n[14] rowon_n[15] col_n[0] col_n[1] col_n[2]
+ col_n[3] col_n[4] col_n[5] col_n[6] col_n[7] col_n[8] col_n[9] col_n[10] col_n[11] col_n[12] col_n[13]
+ col_n[14] col_n[15] col_n[16] col_n[17] col_n[18] col_n[19] col_n[20] col_n[21] col_n[22] col_n[23] col_n[24]
+ col_n[25] col_n[26] col_n[27] col_n[28] col_n[29] col_n[30] col_n[31] en_bit_n[0] en_bit_n[1] en_bit_n[2] en_C0_n sw sw_n analog_in ctop col[0] col[1] col[2] col[3] col[4] col[5] col[6] col[7] col[8] col[9]
+ col[10] col[11] col[12] col[13] col[14] col[15] col[16] col[17] col[18] col[19] col[20] col[21] col[22]
+ col[23] col[24] col[25] col[26] col[27] col[28] col[29] col[30] col[31] rowoff_n[0] rowoff_n[1] rowoff_n[2]
+ rowoff_n[3] rowoff_n[4] rowoff_n[5] rowoff_n[6] rowoff_n[7] rowoff_n[8] rowoff_n[9] rowoff_n[10] rowoff_n[11]
+ rowoff_n[12] rowoff_n[13] rowoff_n[14] rowoff_n[15]
Xadc_array_wafflecap_dummy_5[0] vcm adc_array_wafflecap_dummy_5[0]/ctop VSS VDD row_n[0]
+ rowon_n[0] adc_array_wafflecap_8_1[9]/sample adc_array_wafflecap_8_1[9]/sample_n
+ rowoff_n[0] adc_array_wafflecap_dummy_5[0]/cbot VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_5[1] vcm adc_array_wafflecap_dummy_5[1]/ctop VSS VDD row_n[1]
+ rowon_n[1] adc_array_wafflecap_8_0[0|9]/sample adc_array_wafflecap_8_0[0|9]/sample_n
+ rowoff_n[1] adc_array_wafflecap_dummy_5[1]/cbot VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_5[2] vcm adc_array_wafflecap_dummy_5[2]/ctop VSS VDD row_n[2]
+ rowon_n[2] adc_array_wafflecap_8_0[1|9]/sample adc_array_wafflecap_8_0[1|9]/sample_n
+ rowoff_n[2] adc_array_wafflecap_dummy_5[2]/cbot VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_5[3] vcm adc_array_wafflecap_dummy_5[3]/ctop VSS VDD row_n[3]
+ rowon_n[3] adc_array_wafflecap_8_0[2|9]/sample adc_array_wafflecap_8_0[2|9]/sample_n
+ rowoff_n[3] adc_array_wafflecap_dummy_5[3]/cbot VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_5[4] vcm adc_array_wafflecap_dummy_5[4]/ctop VSS VDD row_n[4]
+ rowon_n[4] adc_array_wafflecap_8_0[3|9]/sample adc_array_wafflecap_8_0[3|9]/sample_n
+ rowoff_n[4] adc_array_wafflecap_dummy_5[4]/cbot VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_5[5] vcm adc_array_wafflecap_dummy_5[5]/ctop VSS VDD row_n[5]
+ rowon_n[5] adc_array_wafflecap_8_0[4|9]/sample adc_array_wafflecap_8_0[4|9]/sample_n
+ rowoff_n[5] adc_array_wafflecap_dummy_5[5]/cbot VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_5[6] vcm adc_array_wafflecap_dummy_5[6]/ctop VSS VDD row_n[6]
+ rowon_n[6] adc_array_wafflecap_8_0[5|9]/sample adc_array_wafflecap_8_0[5|9]/sample_n
+ rowoff_n[6] adc_array_wafflecap_dummy_5[6]/cbot VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_5[7] vcm adc_array_wafflecap_dummy_5[7]/ctop VSS VDD row_n[7]
+ rowon_n[7] adc_array_wafflecap_8_0[6|9]/sample adc_array_wafflecap_8_0[6|9]/sample_n
+ rowoff_n[7] adc_array_wafflecap_dummy_5[7]/cbot VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_5[8] vcm adc_array_wafflecap_dummy_5[8]/ctop VSS VDD row_n[8]
+ rowon_n[8] adc_array_wafflecap_8_0[7|9]/sample adc_array_wafflecap_8_0[7|9]/sample_n
+ rowoff_n[8] adc_array_wafflecap_dummy_5[8]/cbot VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_5[9] vcm adc_array_wafflecap_dummy_5[9]/ctop VSS VDD row_n[9]
+ rowon_n[9] adc_array_wafflecap_8_0[8|9]/sample adc_array_wafflecap_8_0[8|9]/sample_n
+ rowoff_n[9] adc_array_wafflecap_dummy_5[9]/cbot VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_5[10] vcm adc_array_wafflecap_dummy_5[10]/ctop VSS VDD
+ row_n[10] rowon_n[10] adc_array_wafflecap_8_0[9|9]/sample adc_array_wafflecap_8_0[9|9]/sample_n
+ rowoff_n[10] adc_array_wafflecap_dummy_5[10]/cbot VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_5[11] vcm adc_array_wafflecap_dummy_5[11]/ctop VSS VDD
+ row_n[11] rowon_n[11] adc_array_wafflecap_8_0[10|9]/sample adc_array_wafflecap_8_0[10|9]/sample_n
+ rowoff_n[11] adc_array_wafflecap_dummy_5[11]/cbot VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_5[12] vcm adc_array_wafflecap_dummy_5[12]/ctop VSS VDD
+ row_n[12] rowon_n[12] adc_array_wafflecap_8_0[11|9]/sample adc_array_wafflecap_8_0[11|9]/sample_n
+ rowoff_n[12] adc_array_wafflecap_dummy_5[12]/cbot VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_5[13] vcm adc_array_wafflecap_dummy_5[13]/ctop VSS VDD
+ row_n[13] rowon_n[13] adc_array_wafflecap_8_0[12|9]/sample adc_array_wafflecap_8_0[12|9]/sample_n
+ rowoff_n[13] adc_array_wafflecap_dummy_5[13]/cbot VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_5[14] vcm adc_array_wafflecap_dummy_5[14]/ctop VSS VDD
+ row_n[14] rowon_n[14] adc_array_wafflecap_8_0[13|9]/sample adc_array_wafflecap_8_0[13|9]/sample_n
+ rowoff_n[14] adc_array_wafflecap_dummy_5[14]/cbot VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_5[15] vcm adc_array_wafflecap_dummy_5[15]/ctop VSS VDD
+ row_n[15] rowon_n[15] adc_array_wafflecap_8_0[14|9]/sample adc_array_wafflecap_8_0[14|9]/sample_n
+ rowoff_n[15] adc_array_wafflecap_dummy_5[15]/cbot VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_6 vcm adc_array_wafflecap_dummy_6/ctop VSS VDD VDD VSS
+ adc_array_wafflecap_4_0/sample adc_array_wafflecap_4_0/sample_n VDD adc_array_wafflecap_dummy_6/cbot
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_7 vcm adc_array_wafflecap_dummy_7/ctop col[0] col_n[0]
+ row_n[0] rowon_n[0] adc_array_wafflecap_8_1[9]/sample adc_array_wafflecap_8_1[9]/sample_n
+ rowoff_n[0] adc_array_wafflecap_dummy_7/cbot VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_1_0 vcm ctop col[17] col_n[17] VDD VSS adc_array_wafflecap_4_0/sample
+ adc_array_wafflecap_4_0/sample_n VDD en_bit_n[0] adc_array_wafflecap_1_0/cbot VDD
+ VSS adc_array_wafflecap_1
Xadc_array_wafflecap_drv_0[0] vcm adc_array_wafflecap_drv_0[0]/ctop adc_array_wafflecap_drv_2/col
+ VDD row_n[0] rowon_n[0] sample adc_array_wafflecap_8_1[9]/sample sample_n adc_array_wafflecap_8_1[9]/sample_n
+ rowoff_n[0] adc_array_wafflecap_drv_0[0]/cbot VDD VSS adc_array_wafflecap_drv
Xadc_array_wafflecap_drv_0[1] vcm adc_array_wafflecap_drv_0[1]/ctop adc_array_wafflecap_drv_2/col
+ VDD row_n[1] rowon_n[1] sample adc_array_wafflecap_8_0[0|9]/sample sample_n adc_array_wafflecap_8_0[0|9]/sample_n
+ rowoff_n[1] adc_array_wafflecap_drv_0[1]/cbot VDD VSS adc_array_wafflecap_drv
Xadc_array_wafflecap_drv_0[2] vcm adc_array_wafflecap_drv_0[2]/ctop adc_array_wafflecap_drv_2/col
+ VDD row_n[2] rowon_n[2] sample adc_array_wafflecap_8_0[1|9]/sample sample_n adc_array_wafflecap_8_0[1|9]/sample_n
+ rowoff_n[2] adc_array_wafflecap_drv_0[2]/cbot VDD VSS adc_array_wafflecap_drv
Xadc_array_wafflecap_drv_0[3] vcm adc_array_wafflecap_drv_0[3]/ctop adc_array_wafflecap_drv_2/col
+ VDD row_n[3] rowon_n[3] sample adc_array_wafflecap_8_0[2|9]/sample sample_n adc_array_wafflecap_8_0[2|9]/sample_n
+ rowoff_n[3] adc_array_wafflecap_drv_0[3]/cbot VDD VSS adc_array_wafflecap_drv
Xadc_array_wafflecap_drv_0[4] vcm adc_array_wafflecap_drv_0[4]/ctop adc_array_wafflecap_drv_2/col
+ VDD row_n[4] rowon_n[4] sample adc_array_wafflecap_8_0[3|9]/sample sample_n adc_array_wafflecap_8_0[3|9]/sample_n
+ rowoff_n[4] adc_array_wafflecap_drv_0[4]/cbot VDD VSS adc_array_wafflecap_drv
Xadc_array_wafflecap_drv_0[5] vcm adc_array_wafflecap_drv_0[5]/ctop adc_array_wafflecap_drv_2/col
+ VDD row_n[5] rowon_n[5] sample adc_array_wafflecap_8_0[4|9]/sample sample_n adc_array_wafflecap_8_0[4|9]/sample_n
+ rowoff_n[5] adc_array_wafflecap_drv_0[5]/cbot VDD VSS adc_array_wafflecap_drv
Xadc_array_wafflecap_drv_0[6] vcm adc_array_wafflecap_drv_0[6]/ctop adc_array_wafflecap_drv_2/col
+ VDD row_n[6] rowon_n[6] sample adc_array_wafflecap_8_0[5|9]/sample sample_n adc_array_wafflecap_8_0[5|9]/sample_n
+ rowoff_n[6] adc_array_wafflecap_drv_0[6]/cbot VDD VSS adc_array_wafflecap_drv
Xadc_array_wafflecap_drv_0[7] vcm adc_array_wafflecap_drv_0[7]/ctop adc_array_wafflecap_drv_2/col
+ VDD row_n[7] rowon_n[7] sample adc_array_wafflecap_8_0[6|9]/sample sample_n adc_array_wafflecap_8_0[6|9]/sample_n
+ rowoff_n[7] adc_array_wafflecap_drv_0[7]/cbot VDD VSS adc_array_wafflecap_drv
Xadc_array_wafflecap_drv_0[8] vcm adc_array_wafflecap_drv_0[8]/ctop adc_array_wafflecap_drv_2/col
+ VDD row_n[8] rowon_n[8] sample adc_array_wafflecap_8_0[7|9]/sample sample_n adc_array_wafflecap_8_0[7|9]/sample_n
+ rowoff_n[8] adc_array_wafflecap_drv_0[8]/cbot VDD VSS adc_array_wafflecap_drv
Xadc_array_wafflecap_drv_0[9] vcm adc_array_wafflecap_drv_0[9]/ctop adc_array_wafflecap_drv_2/col
+ VDD row_n[9] rowon_n[9] sample adc_array_wafflecap_8_0[8|9]/sample sample_n adc_array_wafflecap_8_0[8|9]/sample_n
+ rowoff_n[9] adc_array_wafflecap_drv_0[9]/cbot VDD VSS adc_array_wafflecap_drv
Xadc_array_wafflecap_drv_0[10] vcm adc_array_wafflecap_drv_0[10]/ctop adc_array_wafflecap_drv_2/col
+ VDD row_n[10] rowon_n[10] sample adc_array_wafflecap_8_0[9|9]/sample sample_n adc_array_wafflecap_8_0[9|9]/sample_n
+ rowoff_n[10] adc_array_wafflecap_drv_0[10]/cbot VDD VSS adc_array_wafflecap_drv
Xadc_array_wafflecap_drv_0[11] vcm adc_array_wafflecap_drv_0[11]/ctop adc_array_wafflecap_drv_2/col
+ VDD row_n[11] rowon_n[11] sample adc_array_wafflecap_8_0[10|9]/sample sample_n adc_array_wafflecap_8_0[10|9]/sample_n
+ rowoff_n[11] adc_array_wafflecap_drv_0[11]/cbot VDD VSS adc_array_wafflecap_drv
Xadc_array_wafflecap_drv_0[12] vcm adc_array_wafflecap_drv_0[12]/ctop adc_array_wafflecap_drv_2/col
+ VDD row_n[12] rowon_n[12] sample adc_array_wafflecap_8_0[11|9]/sample sample_n adc_array_wafflecap_8_0[11|9]/sample_n
+ rowoff_n[12] adc_array_wafflecap_drv_0[12]/cbot VDD VSS adc_array_wafflecap_drv
Xadc_array_wafflecap_drv_0[13] vcm adc_array_wafflecap_drv_0[13]/ctop adc_array_wafflecap_drv_2/col
+ VDD row_n[13] rowon_n[13] sample adc_array_wafflecap_8_0[12|9]/sample sample_n adc_array_wafflecap_8_0[12|9]/sample_n
+ rowoff_n[13] adc_array_wafflecap_drv_0[13]/cbot VDD VSS adc_array_wafflecap_drv
Xadc_array_wafflecap_drv_0[14] vcm adc_array_wafflecap_drv_0[14]/ctop adc_array_wafflecap_drv_2/col
+ VDD row_n[14] rowon_n[14] sample adc_array_wafflecap_8_0[13|9]/sample sample_n adc_array_wafflecap_8_0[13|9]/sample_n
+ rowoff_n[14] adc_array_wafflecap_drv_0[14]/cbot VDD VSS adc_array_wafflecap_drv
Xadc_array_wafflecap_drv_0[15] vcm adc_array_wafflecap_drv_0[15]/ctop adc_array_wafflecap_drv_2/col
+ VDD row_n[15] rowon_n[15] sample adc_array_wafflecap_8_0[14|9]/sample sample_n adc_array_wafflecap_8_0[14|9]/sample_n
+ rowoff_n[15] adc_array_wafflecap_drv_0[15]/cbot VDD VSS adc_array_wafflecap_drv
Xadc_array_wafflecap_1_1 vcm ctop col[1] col_n[1] VDD VSS adc_array_wafflecap_4_0/sample
+ adc_array_wafflecap_4_0/sample_n VDD en_C0_n adc_array_wafflecap_1_1/cbot VDD VSS
+ adc_array_wafflecap_1
Xadc_array_wafflecap_drv_1 vcm adc_array_wafflecap_drv_1/ctop adc_array_wafflecap_drv_2/col
+ VDD VDD VSS sample adc_array_wafflecap_4_0/sample sample_n adc_array_wafflecap_4_0/sample_n
+ VDD adc_array_wafflecap_drv_1/cbot VDD VSS adc_array_wafflecap_drv
Xadc_array_wafflecap_drv_2 vcm adc_array_wafflecap_drv_2/ctop adc_array_wafflecap_drv_2/col
+ VDD VDD VDD sample adc_array_wafflecap_drv_2/sample_o sample_n adc_array_wafflecap_drv_2/sample_n_o
+ VSS adc_array_wafflecap_drv_2/cbot VDD VSS adc_array_wafflecap_drv
Xadc_array_wafflecap_8_0[0|0] vcm ctop col[0] col_n[0] row_n[1] rowon_n[1] adc_array_wafflecap_8_0[0|9]/sample
+ adc_array_wafflecap_8_0[0|9]/sample_n rowoff_n[1] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|0] vcm ctop col[0] col_n[0] row_n[2] rowon_n[2] adc_array_wafflecap_8_0[1|9]/sample
+ adc_array_wafflecap_8_0[1|9]/sample_n rowoff_n[2] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|0] vcm ctop col[0] col_n[0] row_n[3] rowon_n[3] adc_array_wafflecap_8_0[2|9]/sample
+ adc_array_wafflecap_8_0[2|9]/sample_n rowoff_n[3] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|0] vcm ctop col[0] col_n[0] row_n[4] rowon_n[4] adc_array_wafflecap_8_0[3|9]/sample
+ adc_array_wafflecap_8_0[3|9]/sample_n rowoff_n[4] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|0] vcm ctop col[0] col_n[0] row_n[5] rowon_n[5] adc_array_wafflecap_8_0[4|9]/sample
+ adc_array_wafflecap_8_0[4|9]/sample_n rowoff_n[5] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|0] vcm ctop col[0] col_n[0] row_n[6] rowon_n[6] adc_array_wafflecap_8_0[5|9]/sample
+ adc_array_wafflecap_8_0[5|9]/sample_n rowoff_n[6] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|0] vcm ctop col[0] col_n[0] row_n[7] rowon_n[7] adc_array_wafflecap_8_0[6|9]/sample
+ adc_array_wafflecap_8_0[6|9]/sample_n rowoff_n[7] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|0] vcm ctop col[0] col_n[0] row_n[8] rowon_n[8] adc_array_wafflecap_8_0[7|9]/sample
+ adc_array_wafflecap_8_0[7|9]/sample_n rowoff_n[8] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|0] vcm ctop col[0] col_n[0] row_n[9] rowon_n[9] adc_array_wafflecap_8_0[8|9]/sample
+ adc_array_wafflecap_8_0[8|9]/sample_n rowoff_n[9] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|0] vcm ctop col[0] col_n[0] row_n[10] rowon_n[10] adc_array_wafflecap_8_0[9|9]/sample
+ adc_array_wafflecap_8_0[9|9]/sample_n rowoff_n[10] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|0] vcm ctop col[0] col_n[0] row_n[11] rowon_n[11] adc_array_wafflecap_8_0[10|9]/sample
+ adc_array_wafflecap_8_0[10|9]/sample_n rowoff_n[11] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|0] vcm ctop col[0] col_n[0] row_n[12] rowon_n[12] adc_array_wafflecap_8_0[11|9]/sample
+ adc_array_wafflecap_8_0[11|9]/sample_n rowoff_n[12] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|0] vcm ctop col[0] col_n[0] row_n[13] rowon_n[13] adc_array_wafflecap_8_0[12|9]/sample
+ adc_array_wafflecap_8_0[12|9]/sample_n rowoff_n[13] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|0] vcm ctop col[0] col_n[0] row_n[14] rowon_n[14] adc_array_wafflecap_8_0[13|9]/sample
+ adc_array_wafflecap_8_0[13|9]/sample_n rowoff_n[14] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|0] vcm ctop col[0] col_n[0] row_n[15] rowon_n[15] adc_array_wafflecap_8_0[14|9]/sample
+ adc_array_wafflecap_8_0[14|9]/sample_n rowoff_n[15] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|1] vcm ctop col[1] col_n[1] row_n[1] rowon_n[1] adc_array_wafflecap_8_0[0|9]/sample
+ adc_array_wafflecap_8_0[0|9]/sample_n rowoff_n[1] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|1] vcm ctop col[1] col_n[1] row_n[2] rowon_n[2] adc_array_wafflecap_8_0[1|9]/sample
+ adc_array_wafflecap_8_0[1|9]/sample_n rowoff_n[2] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|1] vcm ctop col[1] col_n[1] row_n[3] rowon_n[3] adc_array_wafflecap_8_0[2|9]/sample
+ adc_array_wafflecap_8_0[2|9]/sample_n rowoff_n[3] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|1] vcm ctop col[1] col_n[1] row_n[4] rowon_n[4] adc_array_wafflecap_8_0[3|9]/sample
+ adc_array_wafflecap_8_0[3|9]/sample_n rowoff_n[4] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|1] vcm ctop col[1] col_n[1] row_n[5] rowon_n[5] adc_array_wafflecap_8_0[4|9]/sample
+ adc_array_wafflecap_8_0[4|9]/sample_n rowoff_n[5] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|1] vcm ctop col[1] col_n[1] row_n[6] rowon_n[6] adc_array_wafflecap_8_0[5|9]/sample
+ adc_array_wafflecap_8_0[5|9]/sample_n rowoff_n[6] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|1] vcm ctop col[1] col_n[1] row_n[7] rowon_n[7] adc_array_wafflecap_8_0[6|9]/sample
+ adc_array_wafflecap_8_0[6|9]/sample_n rowoff_n[7] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|1] vcm ctop col[1] col_n[1] row_n[8] rowon_n[8] adc_array_wafflecap_8_0[7|9]/sample
+ adc_array_wafflecap_8_0[7|9]/sample_n rowoff_n[8] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|1] vcm ctop col[1] col_n[1] row_n[9] rowon_n[9] adc_array_wafflecap_8_0[8|9]/sample
+ adc_array_wafflecap_8_0[8|9]/sample_n rowoff_n[9] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|1] vcm ctop col[1] col_n[1] row_n[10] rowon_n[10] adc_array_wafflecap_8_0[9|9]/sample
+ adc_array_wafflecap_8_0[9|9]/sample_n rowoff_n[10] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|1] vcm ctop col[1] col_n[1] row_n[11] rowon_n[11] adc_array_wafflecap_8_0[10|9]/sample
+ adc_array_wafflecap_8_0[10|9]/sample_n rowoff_n[11] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|1] vcm ctop col[1] col_n[1] row_n[12] rowon_n[12] adc_array_wafflecap_8_0[11|9]/sample
+ adc_array_wafflecap_8_0[11|9]/sample_n rowoff_n[12] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|1] vcm ctop col[1] col_n[1] row_n[13] rowon_n[13] adc_array_wafflecap_8_0[12|9]/sample
+ adc_array_wafflecap_8_0[12|9]/sample_n rowoff_n[13] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|1] vcm ctop col[1] col_n[1] row_n[14] rowon_n[14] adc_array_wafflecap_8_0[13|9]/sample
+ adc_array_wafflecap_8_0[13|9]/sample_n rowoff_n[14] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|1] vcm ctop col[1] col_n[1] row_n[15] rowon_n[15] adc_array_wafflecap_8_0[14|9]/sample
+ adc_array_wafflecap_8_0[14|9]/sample_n rowoff_n[15] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|2] vcm ctop col[2] col_n[2] row_n[1] rowon_n[1] adc_array_wafflecap_8_0[0|9]/sample
+ adc_array_wafflecap_8_0[0|9]/sample_n rowoff_n[1] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|2] vcm ctop col[2] col_n[2] row_n[2] rowon_n[2] adc_array_wafflecap_8_0[1|9]/sample
+ adc_array_wafflecap_8_0[1|9]/sample_n rowoff_n[2] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|2] vcm ctop col[2] col_n[2] row_n[3] rowon_n[3] adc_array_wafflecap_8_0[2|9]/sample
+ adc_array_wafflecap_8_0[2|9]/sample_n rowoff_n[3] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|2] vcm ctop col[2] col_n[2] row_n[4] rowon_n[4] adc_array_wafflecap_8_0[3|9]/sample
+ adc_array_wafflecap_8_0[3|9]/sample_n rowoff_n[4] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|2] vcm ctop col[2] col_n[2] row_n[5] rowon_n[5] adc_array_wafflecap_8_0[4|9]/sample
+ adc_array_wafflecap_8_0[4|9]/sample_n rowoff_n[5] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|2] vcm ctop col[2] col_n[2] row_n[6] rowon_n[6] adc_array_wafflecap_8_0[5|9]/sample
+ adc_array_wafflecap_8_0[5|9]/sample_n rowoff_n[6] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|2] vcm ctop col[2] col_n[2] row_n[7] rowon_n[7] adc_array_wafflecap_8_0[6|9]/sample
+ adc_array_wafflecap_8_0[6|9]/sample_n rowoff_n[7] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|2] vcm ctop col[2] col_n[2] row_n[8] rowon_n[8] adc_array_wafflecap_8_0[7|9]/sample
+ adc_array_wafflecap_8_0[7|9]/sample_n rowoff_n[8] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|2] vcm ctop col[2] col_n[2] row_n[9] rowon_n[9] adc_array_wafflecap_8_0[8|9]/sample
+ adc_array_wafflecap_8_0[8|9]/sample_n rowoff_n[9] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|2] vcm ctop col[2] col_n[2] row_n[10] rowon_n[10] adc_array_wafflecap_8_0[9|9]/sample
+ adc_array_wafflecap_8_0[9|9]/sample_n rowoff_n[10] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|2] vcm ctop col[2] col_n[2] row_n[11] rowon_n[11] adc_array_wafflecap_8_0[10|9]/sample
+ adc_array_wafflecap_8_0[10|9]/sample_n rowoff_n[11] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|2] vcm ctop col[2] col_n[2] row_n[12] rowon_n[12] adc_array_wafflecap_8_0[11|9]/sample
+ adc_array_wafflecap_8_0[11|9]/sample_n rowoff_n[12] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|2] vcm ctop col[2] col_n[2] row_n[13] rowon_n[13] adc_array_wafflecap_8_0[12|9]/sample
+ adc_array_wafflecap_8_0[12|9]/sample_n rowoff_n[13] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|2] vcm ctop col[2] col_n[2] row_n[14] rowon_n[14] adc_array_wafflecap_8_0[13|9]/sample
+ adc_array_wafflecap_8_0[13|9]/sample_n rowoff_n[14] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|2] vcm ctop col[2] col_n[2] row_n[15] rowon_n[15] adc_array_wafflecap_8_0[14|9]/sample
+ adc_array_wafflecap_8_0[14|9]/sample_n rowoff_n[15] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|3] vcm ctop col[3] col_n[3] row_n[1] rowon_n[1] adc_array_wafflecap_8_0[0|9]/sample
+ adc_array_wafflecap_8_0[0|9]/sample_n rowoff_n[1] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|3] vcm ctop col[3] col_n[3] row_n[2] rowon_n[2] adc_array_wafflecap_8_0[1|9]/sample
+ adc_array_wafflecap_8_0[1|9]/sample_n rowoff_n[2] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|3] vcm ctop col[3] col_n[3] row_n[3] rowon_n[3] adc_array_wafflecap_8_0[2|9]/sample
+ adc_array_wafflecap_8_0[2|9]/sample_n rowoff_n[3] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|3] vcm ctop col[3] col_n[3] row_n[4] rowon_n[4] adc_array_wafflecap_8_0[3|9]/sample
+ adc_array_wafflecap_8_0[3|9]/sample_n rowoff_n[4] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|3] vcm ctop col[3] col_n[3] row_n[5] rowon_n[5] adc_array_wafflecap_8_0[4|9]/sample
+ adc_array_wafflecap_8_0[4|9]/sample_n rowoff_n[5] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|3] vcm ctop col[3] col_n[3] row_n[6] rowon_n[6] adc_array_wafflecap_8_0[5|9]/sample
+ adc_array_wafflecap_8_0[5|9]/sample_n rowoff_n[6] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|3] vcm ctop col[3] col_n[3] row_n[7] rowon_n[7] adc_array_wafflecap_8_0[6|9]/sample
+ adc_array_wafflecap_8_0[6|9]/sample_n rowoff_n[7] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|3] vcm ctop col[3] col_n[3] row_n[8] rowon_n[8] adc_array_wafflecap_8_0[7|9]/sample
+ adc_array_wafflecap_8_0[7|9]/sample_n rowoff_n[8] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|3] vcm ctop col[3] col_n[3] row_n[9] rowon_n[9] adc_array_wafflecap_8_0[8|9]/sample
+ adc_array_wafflecap_8_0[8|9]/sample_n rowoff_n[9] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|3] vcm ctop col[3] col_n[3] row_n[10] rowon_n[10] adc_array_wafflecap_8_0[9|9]/sample
+ adc_array_wafflecap_8_0[9|9]/sample_n rowoff_n[10] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|3] vcm ctop col[3] col_n[3] row_n[11] rowon_n[11] adc_array_wafflecap_8_0[10|9]/sample
+ adc_array_wafflecap_8_0[10|9]/sample_n rowoff_n[11] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|3] vcm ctop col[3] col_n[3] row_n[12] rowon_n[12] adc_array_wafflecap_8_0[11|9]/sample
+ adc_array_wafflecap_8_0[11|9]/sample_n rowoff_n[12] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|3] vcm ctop col[3] col_n[3] row_n[13] rowon_n[13] adc_array_wafflecap_8_0[12|9]/sample
+ adc_array_wafflecap_8_0[12|9]/sample_n rowoff_n[13] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|3] vcm ctop col[3] col_n[3] row_n[14] rowon_n[14] adc_array_wafflecap_8_0[13|9]/sample
+ adc_array_wafflecap_8_0[13|9]/sample_n rowoff_n[14] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|3] vcm ctop col[3] col_n[3] row_n[15] rowon_n[15] adc_array_wafflecap_8_0[14|9]/sample
+ adc_array_wafflecap_8_0[14|9]/sample_n rowoff_n[15] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|4] vcm ctop col[4] col_n[4] row_n[1] rowon_n[1] adc_array_wafflecap_8_0[0|9]/sample
+ adc_array_wafflecap_8_0[0|9]/sample_n rowoff_n[1] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|4] vcm ctop col[4] col_n[4] row_n[2] rowon_n[2] adc_array_wafflecap_8_0[1|9]/sample
+ adc_array_wafflecap_8_0[1|9]/sample_n rowoff_n[2] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|4] vcm ctop col[4] col_n[4] row_n[3] rowon_n[3] adc_array_wafflecap_8_0[2|9]/sample
+ adc_array_wafflecap_8_0[2|9]/sample_n rowoff_n[3] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|4] vcm ctop col[4] col_n[4] row_n[4] rowon_n[4] adc_array_wafflecap_8_0[3|9]/sample
+ adc_array_wafflecap_8_0[3|9]/sample_n rowoff_n[4] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|4] vcm ctop col[4] col_n[4] row_n[5] rowon_n[5] adc_array_wafflecap_8_0[4|9]/sample
+ adc_array_wafflecap_8_0[4|9]/sample_n rowoff_n[5] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|4] vcm ctop col[4] col_n[4] row_n[6] rowon_n[6] adc_array_wafflecap_8_0[5|9]/sample
+ adc_array_wafflecap_8_0[5|9]/sample_n rowoff_n[6] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|4] vcm ctop col[4] col_n[4] row_n[7] rowon_n[7] adc_array_wafflecap_8_0[6|9]/sample
+ adc_array_wafflecap_8_0[6|9]/sample_n rowoff_n[7] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|4] vcm ctop col[4] col_n[4] row_n[8] rowon_n[8] adc_array_wafflecap_8_0[7|9]/sample
+ adc_array_wafflecap_8_0[7|9]/sample_n rowoff_n[8] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|4] vcm ctop col[4] col_n[4] row_n[9] rowon_n[9] adc_array_wafflecap_8_0[8|9]/sample
+ adc_array_wafflecap_8_0[8|9]/sample_n rowoff_n[9] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|4] vcm ctop col[4] col_n[4] row_n[10] rowon_n[10] adc_array_wafflecap_8_0[9|9]/sample
+ adc_array_wafflecap_8_0[9|9]/sample_n rowoff_n[10] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|4] vcm ctop col[4] col_n[4] row_n[11] rowon_n[11] adc_array_wafflecap_8_0[10|9]/sample
+ adc_array_wafflecap_8_0[10|9]/sample_n rowoff_n[11] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|4] vcm ctop col[4] col_n[4] row_n[12] rowon_n[12] adc_array_wafflecap_8_0[11|9]/sample
+ adc_array_wafflecap_8_0[11|9]/sample_n rowoff_n[12] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|4] vcm ctop col[4] col_n[4] row_n[13] rowon_n[13] adc_array_wafflecap_8_0[12|9]/sample
+ adc_array_wafflecap_8_0[12|9]/sample_n rowoff_n[13] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|4] vcm ctop col[4] col_n[4] row_n[14] rowon_n[14] adc_array_wafflecap_8_0[13|9]/sample
+ adc_array_wafflecap_8_0[13|9]/sample_n rowoff_n[14] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|4] vcm ctop col[4] col_n[4] row_n[15] rowon_n[15] adc_array_wafflecap_8_0[14|9]/sample
+ adc_array_wafflecap_8_0[14|9]/sample_n rowoff_n[15] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|5] vcm ctop col[5] col_n[5] row_n[1] rowon_n[1] adc_array_wafflecap_8_0[0|9]/sample
+ adc_array_wafflecap_8_0[0|9]/sample_n rowoff_n[1] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|5] vcm ctop col[5] col_n[5] row_n[2] rowon_n[2] adc_array_wafflecap_8_0[1|9]/sample
+ adc_array_wafflecap_8_0[1|9]/sample_n rowoff_n[2] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|5] vcm ctop col[5] col_n[5] row_n[3] rowon_n[3] adc_array_wafflecap_8_0[2|9]/sample
+ adc_array_wafflecap_8_0[2|9]/sample_n rowoff_n[3] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|5] vcm ctop col[5] col_n[5] row_n[4] rowon_n[4] adc_array_wafflecap_8_0[3|9]/sample
+ adc_array_wafflecap_8_0[3|9]/sample_n rowoff_n[4] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|5] vcm ctop col[5] col_n[5] row_n[5] rowon_n[5] adc_array_wafflecap_8_0[4|9]/sample
+ adc_array_wafflecap_8_0[4|9]/sample_n rowoff_n[5] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|5] vcm ctop col[5] col_n[5] row_n[6] rowon_n[6] adc_array_wafflecap_8_0[5|9]/sample
+ adc_array_wafflecap_8_0[5|9]/sample_n rowoff_n[6] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|5] vcm ctop col[5] col_n[5] row_n[7] rowon_n[7] adc_array_wafflecap_8_0[6|9]/sample
+ adc_array_wafflecap_8_0[6|9]/sample_n rowoff_n[7] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|5] vcm ctop col[5] col_n[5] row_n[8] rowon_n[8] adc_array_wafflecap_8_0[7|9]/sample
+ adc_array_wafflecap_8_0[7|9]/sample_n rowoff_n[8] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|5] vcm ctop col[5] col_n[5] row_n[9] rowon_n[9] adc_array_wafflecap_8_0[8|9]/sample
+ adc_array_wafflecap_8_0[8|9]/sample_n rowoff_n[9] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|5] vcm ctop col[5] col_n[5] row_n[10] rowon_n[10] adc_array_wafflecap_8_0[9|9]/sample
+ adc_array_wafflecap_8_0[9|9]/sample_n rowoff_n[10] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|5] vcm ctop col[5] col_n[5] row_n[11] rowon_n[11] adc_array_wafflecap_8_0[10|9]/sample
+ adc_array_wafflecap_8_0[10|9]/sample_n rowoff_n[11] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|5] vcm ctop col[5] col_n[5] row_n[12] rowon_n[12] adc_array_wafflecap_8_0[11|9]/sample
+ adc_array_wafflecap_8_0[11|9]/sample_n rowoff_n[12] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|5] vcm ctop col[5] col_n[5] row_n[13] rowon_n[13] adc_array_wafflecap_8_0[12|9]/sample
+ adc_array_wafflecap_8_0[12|9]/sample_n rowoff_n[13] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|5] vcm ctop col[5] col_n[5] row_n[14] rowon_n[14] adc_array_wafflecap_8_0[13|9]/sample
+ adc_array_wafflecap_8_0[13|9]/sample_n rowoff_n[14] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|5] vcm ctop col[5] col_n[5] row_n[15] rowon_n[15] adc_array_wafflecap_8_0[14|9]/sample
+ adc_array_wafflecap_8_0[14|9]/sample_n rowoff_n[15] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|6] vcm ctop col[6] col_n[6] row_n[1] rowon_n[1] adc_array_wafflecap_8_0[0|9]/sample
+ adc_array_wafflecap_8_0[0|9]/sample_n rowoff_n[1] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|6] vcm ctop col[6] col_n[6] row_n[2] rowon_n[2] adc_array_wafflecap_8_0[1|9]/sample
+ adc_array_wafflecap_8_0[1|9]/sample_n rowoff_n[2] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|6] vcm ctop col[6] col_n[6] row_n[3] rowon_n[3] adc_array_wafflecap_8_0[2|9]/sample
+ adc_array_wafflecap_8_0[2|9]/sample_n rowoff_n[3] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|6] vcm ctop col[6] col_n[6] row_n[4] rowon_n[4] adc_array_wafflecap_8_0[3|9]/sample
+ adc_array_wafflecap_8_0[3|9]/sample_n rowoff_n[4] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|6] vcm ctop col[6] col_n[6] row_n[5] rowon_n[5] adc_array_wafflecap_8_0[4|9]/sample
+ adc_array_wafflecap_8_0[4|9]/sample_n rowoff_n[5] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|6] vcm ctop col[6] col_n[6] row_n[6] rowon_n[6] adc_array_wafflecap_8_0[5|9]/sample
+ adc_array_wafflecap_8_0[5|9]/sample_n rowoff_n[6] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|6] vcm ctop col[6] col_n[6] row_n[7] rowon_n[7] adc_array_wafflecap_8_0[6|9]/sample
+ adc_array_wafflecap_8_0[6|9]/sample_n rowoff_n[7] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|6] vcm ctop col[6] col_n[6] row_n[8] rowon_n[8] adc_array_wafflecap_8_0[7|9]/sample
+ adc_array_wafflecap_8_0[7|9]/sample_n rowoff_n[8] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|6] vcm ctop col[6] col_n[6] row_n[9] rowon_n[9] adc_array_wafflecap_8_0[8|9]/sample
+ adc_array_wafflecap_8_0[8|9]/sample_n rowoff_n[9] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|6] vcm ctop col[6] col_n[6] row_n[10] rowon_n[10] adc_array_wafflecap_8_0[9|9]/sample
+ adc_array_wafflecap_8_0[9|9]/sample_n rowoff_n[10] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|6] vcm ctop col[6] col_n[6] row_n[11] rowon_n[11] adc_array_wafflecap_8_0[10|9]/sample
+ adc_array_wafflecap_8_0[10|9]/sample_n rowoff_n[11] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|6] vcm ctop col[6] col_n[6] row_n[12] rowon_n[12] adc_array_wafflecap_8_0[11|9]/sample
+ adc_array_wafflecap_8_0[11|9]/sample_n rowoff_n[12] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|6] vcm ctop col[6] col_n[6] row_n[13] rowon_n[13] adc_array_wafflecap_8_0[12|9]/sample
+ adc_array_wafflecap_8_0[12|9]/sample_n rowoff_n[13] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|6] vcm ctop col[6] col_n[6] row_n[14] rowon_n[14] adc_array_wafflecap_8_0[13|9]/sample
+ adc_array_wafflecap_8_0[13|9]/sample_n rowoff_n[14] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|6] vcm ctop col[6] col_n[6] row_n[15] rowon_n[15] adc_array_wafflecap_8_0[14|9]/sample
+ adc_array_wafflecap_8_0[14|9]/sample_n rowoff_n[15] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|7] vcm ctop col[7] col_n[7] row_n[1] rowon_n[1] adc_array_wafflecap_8_0[0|9]/sample
+ adc_array_wafflecap_8_0[0|9]/sample_n rowoff_n[1] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|7] vcm ctop col[7] col_n[7] row_n[2] rowon_n[2] adc_array_wafflecap_8_0[1|9]/sample
+ adc_array_wafflecap_8_0[1|9]/sample_n rowoff_n[2] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|7] vcm ctop col[7] col_n[7] row_n[3] rowon_n[3] adc_array_wafflecap_8_0[2|9]/sample
+ adc_array_wafflecap_8_0[2|9]/sample_n rowoff_n[3] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|7] vcm ctop col[7] col_n[7] row_n[4] rowon_n[4] adc_array_wafflecap_8_0[3|9]/sample
+ adc_array_wafflecap_8_0[3|9]/sample_n rowoff_n[4] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|7] vcm ctop col[7] col_n[7] row_n[5] rowon_n[5] adc_array_wafflecap_8_0[4|9]/sample
+ adc_array_wafflecap_8_0[4|9]/sample_n rowoff_n[5] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|7] vcm ctop col[7] col_n[7] row_n[6] rowon_n[6] adc_array_wafflecap_8_0[5|9]/sample
+ adc_array_wafflecap_8_0[5|9]/sample_n rowoff_n[6] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|7] vcm ctop col[7] col_n[7] row_n[7] rowon_n[7] adc_array_wafflecap_8_0[6|9]/sample
+ adc_array_wafflecap_8_0[6|9]/sample_n rowoff_n[7] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|7] vcm ctop col[7] col_n[7] row_n[8] rowon_n[8] adc_array_wafflecap_8_0[7|9]/sample
+ adc_array_wafflecap_8_0[7|9]/sample_n rowoff_n[8] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|7] vcm ctop col[7] col_n[7] row_n[9] rowon_n[9] adc_array_wafflecap_8_0[8|9]/sample
+ adc_array_wafflecap_8_0[8|9]/sample_n rowoff_n[9] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|7] vcm ctop col[7] col_n[7] row_n[10] rowon_n[10] adc_array_wafflecap_8_0[9|9]/sample
+ adc_array_wafflecap_8_0[9|9]/sample_n rowoff_n[10] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|7] vcm ctop col[7] col_n[7] row_n[11] rowon_n[11] adc_array_wafflecap_8_0[10|9]/sample
+ adc_array_wafflecap_8_0[10|9]/sample_n rowoff_n[11] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|7] vcm ctop col[7] col_n[7] row_n[12] rowon_n[12] adc_array_wafflecap_8_0[11|9]/sample
+ adc_array_wafflecap_8_0[11|9]/sample_n rowoff_n[12] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|7] vcm ctop col[7] col_n[7] row_n[13] rowon_n[13] adc_array_wafflecap_8_0[12|9]/sample
+ adc_array_wafflecap_8_0[12|9]/sample_n rowoff_n[13] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|7] vcm ctop col[7] col_n[7] row_n[14] rowon_n[14] adc_array_wafflecap_8_0[13|9]/sample
+ adc_array_wafflecap_8_0[13|9]/sample_n rowoff_n[14] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|7] vcm ctop col[7] col_n[7] row_n[15] rowon_n[15] adc_array_wafflecap_8_0[14|9]/sample
+ adc_array_wafflecap_8_0[14|9]/sample_n rowoff_n[15] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|8] vcm ctop col[8] col_n[8] row_n[1] rowon_n[1] adc_array_wafflecap_8_0[0|9]/sample
+ adc_array_wafflecap_8_0[0|9]/sample_n rowoff_n[1] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|8] vcm ctop col[8] col_n[8] row_n[2] rowon_n[2] adc_array_wafflecap_8_0[1|9]/sample
+ adc_array_wafflecap_8_0[1|9]/sample_n rowoff_n[2] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|8] vcm ctop col[8] col_n[8] row_n[3] rowon_n[3] adc_array_wafflecap_8_0[2|9]/sample
+ adc_array_wafflecap_8_0[2|9]/sample_n rowoff_n[3] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|8] vcm ctop col[8] col_n[8] row_n[4] rowon_n[4] adc_array_wafflecap_8_0[3|9]/sample
+ adc_array_wafflecap_8_0[3|9]/sample_n rowoff_n[4] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|8] vcm ctop col[8] col_n[8] row_n[5] rowon_n[5] adc_array_wafflecap_8_0[4|9]/sample
+ adc_array_wafflecap_8_0[4|9]/sample_n rowoff_n[5] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|8] vcm ctop col[8] col_n[8] row_n[6] rowon_n[6] adc_array_wafflecap_8_0[5|9]/sample
+ adc_array_wafflecap_8_0[5|9]/sample_n rowoff_n[6] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|8] vcm ctop col[8] col_n[8] row_n[7] rowon_n[7] adc_array_wafflecap_8_0[6|9]/sample
+ adc_array_wafflecap_8_0[6|9]/sample_n rowoff_n[7] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|8] vcm ctop col[8] col_n[8] row_n[8] rowon_n[8] adc_array_wafflecap_8_0[7|9]/sample
+ adc_array_wafflecap_8_0[7|9]/sample_n rowoff_n[8] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|8] vcm ctop col[8] col_n[8] row_n[9] rowon_n[9] adc_array_wafflecap_8_0[8|9]/sample
+ adc_array_wafflecap_8_0[8|9]/sample_n rowoff_n[9] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|8] vcm ctop col[8] col_n[8] row_n[10] rowon_n[10] adc_array_wafflecap_8_0[9|9]/sample
+ adc_array_wafflecap_8_0[9|9]/sample_n rowoff_n[10] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|8] vcm ctop col[8] col_n[8] row_n[11] rowon_n[11] adc_array_wafflecap_8_0[10|9]/sample
+ adc_array_wafflecap_8_0[10|9]/sample_n rowoff_n[11] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|8] vcm ctop col[8] col_n[8] row_n[12] rowon_n[12] adc_array_wafflecap_8_0[11|9]/sample
+ adc_array_wafflecap_8_0[11|9]/sample_n rowoff_n[12] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|8] vcm ctop col[8] col_n[8] row_n[13] rowon_n[13] adc_array_wafflecap_8_0[12|9]/sample
+ adc_array_wafflecap_8_0[12|9]/sample_n rowoff_n[13] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|8] vcm ctop col[8] col_n[8] row_n[14] rowon_n[14] adc_array_wafflecap_8_0[13|9]/sample
+ adc_array_wafflecap_8_0[13|9]/sample_n rowoff_n[14] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|8] vcm ctop col[8] col_n[8] row_n[15] rowon_n[15] adc_array_wafflecap_8_0[14|9]/sample
+ adc_array_wafflecap_8_0[14|9]/sample_n rowoff_n[15] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|9] vcm ctop col[9] col_n[9] row_n[1] rowon_n[1] adc_array_wafflecap_8_0[0|9]/sample
+ adc_array_wafflecap_8_0[0|9]/sample_n rowoff_n[1] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|9] vcm ctop col[9] col_n[9] row_n[2] rowon_n[2] adc_array_wafflecap_8_0[1|9]/sample
+ adc_array_wafflecap_8_0[1|9]/sample_n rowoff_n[2] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|9] vcm ctop col[9] col_n[9] row_n[3] rowon_n[3] adc_array_wafflecap_8_0[2|9]/sample
+ adc_array_wafflecap_8_0[2|9]/sample_n rowoff_n[3] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|9] vcm ctop col[9] col_n[9] row_n[4] rowon_n[4] adc_array_wafflecap_8_0[3|9]/sample
+ adc_array_wafflecap_8_0[3|9]/sample_n rowoff_n[4] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|9] vcm ctop col[9] col_n[9] row_n[5] rowon_n[5] adc_array_wafflecap_8_0[4|9]/sample
+ adc_array_wafflecap_8_0[4|9]/sample_n rowoff_n[5] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|9] vcm ctop col[9] col_n[9] row_n[6] rowon_n[6] adc_array_wafflecap_8_0[5|9]/sample
+ adc_array_wafflecap_8_0[5|9]/sample_n rowoff_n[6] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|9] vcm ctop col[9] col_n[9] row_n[7] rowon_n[7] adc_array_wafflecap_8_0[6|9]/sample
+ adc_array_wafflecap_8_0[6|9]/sample_n rowoff_n[7] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|9] vcm ctop col[9] col_n[9] row_n[8] rowon_n[8] adc_array_wafflecap_8_0[7|9]/sample
+ adc_array_wafflecap_8_0[7|9]/sample_n rowoff_n[8] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|9] vcm ctop col[9] col_n[9] row_n[9] rowon_n[9] adc_array_wafflecap_8_0[8|9]/sample
+ adc_array_wafflecap_8_0[8|9]/sample_n rowoff_n[9] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|9] vcm ctop col[9] col_n[9] row_n[10] rowon_n[10] adc_array_wafflecap_8_0[9|9]/sample
+ adc_array_wafflecap_8_0[9|9]/sample_n rowoff_n[10] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|9] vcm ctop col[9] col_n[9] row_n[11] rowon_n[11] adc_array_wafflecap_8_0[10|9]/sample
+ adc_array_wafflecap_8_0[10|9]/sample_n rowoff_n[11] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|9] vcm ctop col[9] col_n[9] row_n[12] rowon_n[12] adc_array_wafflecap_8_0[11|9]/sample
+ adc_array_wafflecap_8_0[11|9]/sample_n rowoff_n[12] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|9] vcm ctop col[9] col_n[9] row_n[13] rowon_n[13] adc_array_wafflecap_8_0[12|9]/sample
+ adc_array_wafflecap_8_0[12|9]/sample_n rowoff_n[13] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|9] vcm ctop col[9] col_n[9] row_n[14] rowon_n[14] adc_array_wafflecap_8_0[13|9]/sample
+ adc_array_wafflecap_8_0[13|9]/sample_n rowoff_n[14] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|9] vcm ctop col[9] col_n[9] row_n[15] rowon_n[15] adc_array_wafflecap_8_0[14|9]/sample
+ adc_array_wafflecap_8_0[14|9]/sample_n rowoff_n[15] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|10] vcm ctop col[10] col_n[10] row_n[1] rowon_n[1] adc_array_wafflecap_8_0[0|9]/sample
+ adc_array_wafflecap_8_0[0|9]/sample_n rowoff_n[1] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|10] vcm ctop col[10] col_n[10] row_n[2] rowon_n[2] adc_array_wafflecap_8_0[1|9]/sample
+ adc_array_wafflecap_8_0[1|9]/sample_n rowoff_n[2] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|10] vcm ctop col[10] col_n[10] row_n[3] rowon_n[3] adc_array_wafflecap_8_0[2|9]/sample
+ adc_array_wafflecap_8_0[2|9]/sample_n rowoff_n[3] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|10] vcm ctop col[10] col_n[10] row_n[4] rowon_n[4] adc_array_wafflecap_8_0[3|9]/sample
+ adc_array_wafflecap_8_0[3|9]/sample_n rowoff_n[4] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|10] vcm ctop col[10] col_n[10] row_n[5] rowon_n[5] adc_array_wafflecap_8_0[4|9]/sample
+ adc_array_wafflecap_8_0[4|9]/sample_n rowoff_n[5] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|10] vcm ctop col[10] col_n[10] row_n[6] rowon_n[6] adc_array_wafflecap_8_0[5|9]/sample
+ adc_array_wafflecap_8_0[5|9]/sample_n rowoff_n[6] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|10] vcm ctop col[10] col_n[10] row_n[7] rowon_n[7] adc_array_wafflecap_8_0[6|9]/sample
+ adc_array_wafflecap_8_0[6|9]/sample_n rowoff_n[7] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|10] vcm ctop col[10] col_n[10] row_n[8] rowon_n[8] adc_array_wafflecap_8_0[7|9]/sample
+ adc_array_wafflecap_8_0[7|9]/sample_n rowoff_n[8] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|10] vcm ctop col[10] col_n[10] row_n[9] rowon_n[9] adc_array_wafflecap_8_0[8|9]/sample
+ adc_array_wafflecap_8_0[8|9]/sample_n rowoff_n[9] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|10] vcm ctop col[10] col_n[10] row_n[10] rowon_n[10] adc_array_wafflecap_8_0[9|9]/sample
+ adc_array_wafflecap_8_0[9|9]/sample_n rowoff_n[10] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|10] vcm ctop col[10] col_n[10] row_n[11] rowon_n[11] adc_array_wafflecap_8_0[10|9]/sample
+ adc_array_wafflecap_8_0[10|9]/sample_n rowoff_n[11] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|10] vcm ctop col[10] col_n[10] row_n[12] rowon_n[12] adc_array_wafflecap_8_0[11|9]/sample
+ adc_array_wafflecap_8_0[11|9]/sample_n rowoff_n[12] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|10] vcm ctop col[10] col_n[10] row_n[13] rowon_n[13] adc_array_wafflecap_8_0[12|9]/sample
+ adc_array_wafflecap_8_0[12|9]/sample_n rowoff_n[13] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|10] vcm ctop col[10] col_n[10] row_n[14] rowon_n[14] adc_array_wafflecap_8_0[13|9]/sample
+ adc_array_wafflecap_8_0[13|9]/sample_n rowoff_n[14] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|10] vcm ctop col[10] col_n[10] row_n[15] rowon_n[15] adc_array_wafflecap_8_0[14|9]/sample
+ adc_array_wafflecap_8_0[14|9]/sample_n rowoff_n[15] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|11] vcm ctop col[11] col_n[11] row_n[1] rowon_n[1] adc_array_wafflecap_8_0[0|9]/sample
+ adc_array_wafflecap_8_0[0|9]/sample_n rowoff_n[1] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|11] vcm ctop col[11] col_n[11] row_n[2] rowon_n[2] adc_array_wafflecap_8_0[1|9]/sample
+ adc_array_wafflecap_8_0[1|9]/sample_n rowoff_n[2] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|11] vcm ctop col[11] col_n[11] row_n[3] rowon_n[3] adc_array_wafflecap_8_0[2|9]/sample
+ adc_array_wafflecap_8_0[2|9]/sample_n rowoff_n[3] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|11] vcm ctop col[11] col_n[11] row_n[4] rowon_n[4] adc_array_wafflecap_8_0[3|9]/sample
+ adc_array_wafflecap_8_0[3|9]/sample_n rowoff_n[4] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|11] vcm ctop col[11] col_n[11] row_n[5] rowon_n[5] adc_array_wafflecap_8_0[4|9]/sample
+ adc_array_wafflecap_8_0[4|9]/sample_n rowoff_n[5] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|11] vcm ctop col[11] col_n[11] row_n[6] rowon_n[6] adc_array_wafflecap_8_0[5|9]/sample
+ adc_array_wafflecap_8_0[5|9]/sample_n rowoff_n[6] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|11] vcm ctop col[11] col_n[11] row_n[7] rowon_n[7] adc_array_wafflecap_8_0[6|9]/sample
+ adc_array_wafflecap_8_0[6|9]/sample_n rowoff_n[7] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|11] vcm ctop col[11] col_n[11] row_n[8] rowon_n[8] adc_array_wafflecap_8_0[7|9]/sample
+ adc_array_wafflecap_8_0[7|9]/sample_n rowoff_n[8] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|11] vcm ctop col[11] col_n[11] row_n[9] rowon_n[9] adc_array_wafflecap_8_0[8|9]/sample
+ adc_array_wafflecap_8_0[8|9]/sample_n rowoff_n[9] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|11] vcm ctop col[11] col_n[11] row_n[10] rowon_n[10] adc_array_wafflecap_8_0[9|9]/sample
+ adc_array_wafflecap_8_0[9|9]/sample_n rowoff_n[10] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|11] vcm ctop col[11] col_n[11] row_n[11] rowon_n[11] adc_array_wafflecap_8_0[10|9]/sample
+ adc_array_wafflecap_8_0[10|9]/sample_n rowoff_n[11] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|11] vcm ctop col[11] col_n[11] row_n[12] rowon_n[12] adc_array_wafflecap_8_0[11|9]/sample
+ adc_array_wafflecap_8_0[11|9]/sample_n rowoff_n[12] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|11] vcm ctop col[11] col_n[11] row_n[13] rowon_n[13] adc_array_wafflecap_8_0[12|9]/sample
+ adc_array_wafflecap_8_0[12|9]/sample_n rowoff_n[13] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|11] vcm ctop col[11] col_n[11] row_n[14] rowon_n[14] adc_array_wafflecap_8_0[13|9]/sample
+ adc_array_wafflecap_8_0[13|9]/sample_n rowoff_n[14] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|11] vcm ctop col[11] col_n[11] row_n[15] rowon_n[15] adc_array_wafflecap_8_0[14|9]/sample
+ adc_array_wafflecap_8_0[14|9]/sample_n rowoff_n[15] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|12] vcm ctop col[12] col_n[12] row_n[1] rowon_n[1] adc_array_wafflecap_8_0[0|9]/sample
+ adc_array_wafflecap_8_0[0|9]/sample_n rowoff_n[1] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|12] vcm ctop col[12] col_n[12] row_n[2] rowon_n[2] adc_array_wafflecap_8_0[1|9]/sample
+ adc_array_wafflecap_8_0[1|9]/sample_n rowoff_n[2] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|12] vcm ctop col[12] col_n[12] row_n[3] rowon_n[3] adc_array_wafflecap_8_0[2|9]/sample
+ adc_array_wafflecap_8_0[2|9]/sample_n rowoff_n[3] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|12] vcm ctop col[12] col_n[12] row_n[4] rowon_n[4] adc_array_wafflecap_8_0[3|9]/sample
+ adc_array_wafflecap_8_0[3|9]/sample_n rowoff_n[4] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|12] vcm ctop col[12] col_n[12] row_n[5] rowon_n[5] adc_array_wafflecap_8_0[4|9]/sample
+ adc_array_wafflecap_8_0[4|9]/sample_n rowoff_n[5] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|12] vcm ctop col[12] col_n[12] row_n[6] rowon_n[6] adc_array_wafflecap_8_0[5|9]/sample
+ adc_array_wafflecap_8_0[5|9]/sample_n rowoff_n[6] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|12] vcm ctop col[12] col_n[12] row_n[7] rowon_n[7] adc_array_wafflecap_8_0[6|9]/sample
+ adc_array_wafflecap_8_0[6|9]/sample_n rowoff_n[7] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|12] vcm ctop col[12] col_n[12] row_n[8] rowon_n[8] adc_array_wafflecap_8_0[7|9]/sample
+ adc_array_wafflecap_8_0[7|9]/sample_n rowoff_n[8] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|12] vcm ctop col[12] col_n[12] row_n[9] rowon_n[9] adc_array_wafflecap_8_0[8|9]/sample
+ adc_array_wafflecap_8_0[8|9]/sample_n rowoff_n[9] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|12] vcm ctop col[12] col_n[12] row_n[10] rowon_n[10] adc_array_wafflecap_8_0[9|9]/sample
+ adc_array_wafflecap_8_0[9|9]/sample_n rowoff_n[10] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|12] vcm ctop col[12] col_n[12] row_n[11] rowon_n[11] adc_array_wafflecap_8_0[10|9]/sample
+ adc_array_wafflecap_8_0[10|9]/sample_n rowoff_n[11] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|12] vcm ctop col[12] col_n[12] row_n[12] rowon_n[12] adc_array_wafflecap_8_0[11|9]/sample
+ adc_array_wafflecap_8_0[11|9]/sample_n rowoff_n[12] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|12] vcm ctop col[12] col_n[12] row_n[13] rowon_n[13] adc_array_wafflecap_8_0[12|9]/sample
+ adc_array_wafflecap_8_0[12|9]/sample_n rowoff_n[13] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|12] vcm ctop col[12] col_n[12] row_n[14] rowon_n[14] adc_array_wafflecap_8_0[13|9]/sample
+ adc_array_wafflecap_8_0[13|9]/sample_n rowoff_n[14] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|12] vcm ctop col[12] col_n[12] row_n[15] rowon_n[15] adc_array_wafflecap_8_0[14|9]/sample
+ adc_array_wafflecap_8_0[14|9]/sample_n rowoff_n[15] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|13] vcm ctop col[13] col_n[13] row_n[1] rowon_n[1] adc_array_wafflecap_8_0[0|9]/sample
+ adc_array_wafflecap_8_0[0|9]/sample_n rowoff_n[1] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|13] vcm ctop col[13] col_n[13] row_n[2] rowon_n[2] adc_array_wafflecap_8_0[1|9]/sample
+ adc_array_wafflecap_8_0[1|9]/sample_n rowoff_n[2] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|13] vcm ctop col[13] col_n[13] row_n[3] rowon_n[3] adc_array_wafflecap_8_0[2|9]/sample
+ adc_array_wafflecap_8_0[2|9]/sample_n rowoff_n[3] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|13] vcm ctop col[13] col_n[13] row_n[4] rowon_n[4] adc_array_wafflecap_8_0[3|9]/sample
+ adc_array_wafflecap_8_0[3|9]/sample_n rowoff_n[4] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|13] vcm ctop col[13] col_n[13] row_n[5] rowon_n[5] adc_array_wafflecap_8_0[4|9]/sample
+ adc_array_wafflecap_8_0[4|9]/sample_n rowoff_n[5] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|13] vcm ctop col[13] col_n[13] row_n[6] rowon_n[6] adc_array_wafflecap_8_0[5|9]/sample
+ adc_array_wafflecap_8_0[5|9]/sample_n rowoff_n[6] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|13] vcm ctop col[13] col_n[13] row_n[7] rowon_n[7] adc_array_wafflecap_8_0[6|9]/sample
+ adc_array_wafflecap_8_0[6|9]/sample_n rowoff_n[7] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|13] vcm ctop col[13] col_n[13] row_n[8] rowon_n[8] adc_array_wafflecap_8_0[7|9]/sample
+ adc_array_wafflecap_8_0[7|9]/sample_n rowoff_n[8] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|13] vcm ctop col[13] col_n[13] row_n[9] rowon_n[9] adc_array_wafflecap_8_0[8|9]/sample
+ adc_array_wafflecap_8_0[8|9]/sample_n rowoff_n[9] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|13] vcm ctop col[13] col_n[13] row_n[10] rowon_n[10] adc_array_wafflecap_8_0[9|9]/sample
+ adc_array_wafflecap_8_0[9|9]/sample_n rowoff_n[10] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|13] vcm ctop col[13] col_n[13] row_n[11] rowon_n[11] adc_array_wafflecap_8_0[10|9]/sample
+ adc_array_wafflecap_8_0[10|9]/sample_n rowoff_n[11] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|13] vcm ctop col[13] col_n[13] row_n[12] rowon_n[12] adc_array_wafflecap_8_0[11|9]/sample
+ adc_array_wafflecap_8_0[11|9]/sample_n rowoff_n[12] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|13] vcm ctop col[13] col_n[13] row_n[13] rowon_n[13] adc_array_wafflecap_8_0[12|9]/sample
+ adc_array_wafflecap_8_0[12|9]/sample_n rowoff_n[13] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|13] vcm ctop col[13] col_n[13] row_n[14] rowon_n[14] adc_array_wafflecap_8_0[13|9]/sample
+ adc_array_wafflecap_8_0[13|9]/sample_n rowoff_n[14] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|13] vcm ctop col[13] col_n[13] row_n[15] rowon_n[15] adc_array_wafflecap_8_0[14|9]/sample
+ adc_array_wafflecap_8_0[14|9]/sample_n rowoff_n[15] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|14] vcm ctop col[14] col_n[14] row_n[1] rowon_n[1] adc_array_wafflecap_8_0[0|9]/sample
+ adc_array_wafflecap_8_0[0|9]/sample_n rowoff_n[1] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|14] vcm ctop col[14] col_n[14] row_n[2] rowon_n[2] adc_array_wafflecap_8_0[1|9]/sample
+ adc_array_wafflecap_8_0[1|9]/sample_n rowoff_n[2] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|14] vcm ctop col[14] col_n[14] row_n[3] rowon_n[3] adc_array_wafflecap_8_0[2|9]/sample
+ adc_array_wafflecap_8_0[2|9]/sample_n rowoff_n[3] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|14] vcm ctop col[14] col_n[14] row_n[4] rowon_n[4] adc_array_wafflecap_8_0[3|9]/sample
+ adc_array_wafflecap_8_0[3|9]/sample_n rowoff_n[4] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|14] vcm ctop col[14] col_n[14] row_n[5] rowon_n[5] adc_array_wafflecap_8_0[4|9]/sample
+ adc_array_wafflecap_8_0[4|9]/sample_n rowoff_n[5] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|14] vcm ctop col[14] col_n[14] row_n[6] rowon_n[6] adc_array_wafflecap_8_0[5|9]/sample
+ adc_array_wafflecap_8_0[5|9]/sample_n rowoff_n[6] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|14] vcm ctop col[14] col_n[14] row_n[7] rowon_n[7] adc_array_wafflecap_8_0[6|9]/sample
+ adc_array_wafflecap_8_0[6|9]/sample_n rowoff_n[7] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|14] vcm ctop col[14] col_n[14] row_n[8] rowon_n[8] adc_array_wafflecap_8_0[7|9]/sample
+ adc_array_wafflecap_8_0[7|9]/sample_n rowoff_n[8] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|14] vcm ctop col[14] col_n[14] row_n[9] rowon_n[9] adc_array_wafflecap_8_0[8|9]/sample
+ adc_array_wafflecap_8_0[8|9]/sample_n rowoff_n[9] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|14] vcm ctop col[14] col_n[14] row_n[10] rowon_n[10] adc_array_wafflecap_8_0[9|9]/sample
+ adc_array_wafflecap_8_0[9|9]/sample_n rowoff_n[10] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|14] vcm ctop col[14] col_n[14] row_n[11] rowon_n[11] adc_array_wafflecap_8_0[10|9]/sample
+ adc_array_wafflecap_8_0[10|9]/sample_n rowoff_n[11] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|14] vcm ctop col[14] col_n[14] row_n[12] rowon_n[12] adc_array_wafflecap_8_0[11|9]/sample
+ adc_array_wafflecap_8_0[11|9]/sample_n rowoff_n[12] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|14] vcm ctop col[14] col_n[14] row_n[13] rowon_n[13] adc_array_wafflecap_8_0[12|9]/sample
+ adc_array_wafflecap_8_0[12|9]/sample_n rowoff_n[13] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|14] vcm ctop col[14] col_n[14] row_n[14] rowon_n[14] adc_array_wafflecap_8_0[13|9]/sample
+ adc_array_wafflecap_8_0[13|9]/sample_n rowoff_n[14] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|14] vcm ctop col[14] col_n[14] row_n[15] rowon_n[15] adc_array_wafflecap_8_0[14|9]/sample
+ adc_array_wafflecap_8_0[14|9]/sample_n rowoff_n[15] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|15] vcm ctop col[15] col_n[15] row_n[1] rowon_n[1] adc_array_wafflecap_8_0[0|9]/sample
+ adc_array_wafflecap_8_0[0|9]/sample_n rowoff_n[1] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|15] vcm ctop col[15] col_n[15] row_n[2] rowon_n[2] adc_array_wafflecap_8_0[1|9]/sample
+ adc_array_wafflecap_8_0[1|9]/sample_n rowoff_n[2] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|15] vcm ctop col[15] col_n[15] row_n[3] rowon_n[3] adc_array_wafflecap_8_0[2|9]/sample
+ adc_array_wafflecap_8_0[2|9]/sample_n rowoff_n[3] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|15] vcm ctop col[15] col_n[15] row_n[4] rowon_n[4] adc_array_wafflecap_8_0[3|9]/sample
+ adc_array_wafflecap_8_0[3|9]/sample_n rowoff_n[4] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|15] vcm ctop col[15] col_n[15] row_n[5] rowon_n[5] adc_array_wafflecap_8_0[4|9]/sample
+ adc_array_wafflecap_8_0[4|9]/sample_n rowoff_n[5] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|15] vcm ctop col[15] col_n[15] row_n[6] rowon_n[6] adc_array_wafflecap_8_0[5|9]/sample
+ adc_array_wafflecap_8_0[5|9]/sample_n rowoff_n[6] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|15] vcm ctop col[15] col_n[15] row_n[7] rowon_n[7] adc_array_wafflecap_8_0[6|9]/sample
+ adc_array_wafflecap_8_0[6|9]/sample_n rowoff_n[7] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|15] vcm ctop col[15] col_n[15] row_n[8] rowon_n[8] adc_array_wafflecap_8_0[7|9]/sample
+ adc_array_wafflecap_8_0[7|9]/sample_n rowoff_n[8] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|15] vcm ctop col[15] col_n[15] row_n[9] rowon_n[9] adc_array_wafflecap_8_0[8|9]/sample
+ adc_array_wafflecap_8_0[8|9]/sample_n rowoff_n[9] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|15] vcm ctop col[15] col_n[15] row_n[10] rowon_n[10] adc_array_wafflecap_8_0[9|9]/sample
+ adc_array_wafflecap_8_0[9|9]/sample_n rowoff_n[10] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|15] vcm ctop col[15] col_n[15] row_n[11] rowon_n[11] adc_array_wafflecap_8_0[10|9]/sample
+ adc_array_wafflecap_8_0[10|9]/sample_n rowoff_n[11] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|15] vcm ctop col[15] col_n[15] row_n[12] rowon_n[12] adc_array_wafflecap_8_0[11|9]/sample
+ adc_array_wafflecap_8_0[11|9]/sample_n rowoff_n[12] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|15] vcm ctop col[15] col_n[15] row_n[13] rowon_n[13] adc_array_wafflecap_8_0[12|9]/sample
+ adc_array_wafflecap_8_0[12|9]/sample_n rowoff_n[13] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|15] vcm ctop col[15] col_n[15] row_n[14] rowon_n[14] adc_array_wafflecap_8_0[13|9]/sample
+ adc_array_wafflecap_8_0[13|9]/sample_n rowoff_n[14] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|15] vcm ctop col[15] col_n[15] row_n[15] rowon_n[15] adc_array_wafflecap_8_0[14|9]/sample
+ adc_array_wafflecap_8_0[14|9]/sample_n rowoff_n[15] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|16] vcm ctop col[16] col_n[16] row_n[1] rowon_n[1] adc_array_wafflecap_8_0[0|9]/sample
+ adc_array_wafflecap_8_0[0|9]/sample_n rowoff_n[1] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|16] vcm ctop col[16] col_n[16] row_n[2] rowon_n[2] adc_array_wafflecap_8_0[1|9]/sample
+ adc_array_wafflecap_8_0[1|9]/sample_n rowoff_n[2] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|16] vcm ctop col[16] col_n[16] row_n[3] rowon_n[3] adc_array_wafflecap_8_0[2|9]/sample
+ adc_array_wafflecap_8_0[2|9]/sample_n rowoff_n[3] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|16] vcm ctop col[16] col_n[16] row_n[4] rowon_n[4] adc_array_wafflecap_8_0[3|9]/sample
+ adc_array_wafflecap_8_0[3|9]/sample_n rowoff_n[4] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|16] vcm ctop col[16] col_n[16] row_n[5] rowon_n[5] adc_array_wafflecap_8_0[4|9]/sample
+ adc_array_wafflecap_8_0[4|9]/sample_n rowoff_n[5] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|16] vcm ctop col[16] col_n[16] row_n[6] rowon_n[6] adc_array_wafflecap_8_0[5|9]/sample
+ adc_array_wafflecap_8_0[5|9]/sample_n rowoff_n[6] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|16] vcm ctop col[16] col_n[16] row_n[7] rowon_n[7] adc_array_wafflecap_8_0[6|9]/sample
+ adc_array_wafflecap_8_0[6|9]/sample_n rowoff_n[7] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|16] vcm ctop col[16] col_n[16] row_n[8] rowon_n[8] adc_array_wafflecap_8_0[7|9]/sample
+ adc_array_wafflecap_8_0[7|9]/sample_n rowoff_n[8] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|16] vcm ctop col[16] col_n[16] row_n[9] rowon_n[9] adc_array_wafflecap_8_0[8|9]/sample
+ adc_array_wafflecap_8_0[8|9]/sample_n rowoff_n[9] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|16] vcm ctop col[16] col_n[16] row_n[10] rowon_n[10] adc_array_wafflecap_8_0[9|9]/sample
+ adc_array_wafflecap_8_0[9|9]/sample_n rowoff_n[10] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|16] vcm ctop col[16] col_n[16] row_n[11] rowon_n[11] adc_array_wafflecap_8_0[10|9]/sample
+ adc_array_wafflecap_8_0[10|9]/sample_n rowoff_n[11] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|16] vcm ctop col[16] col_n[16] row_n[12] rowon_n[12] adc_array_wafflecap_8_0[11|9]/sample
+ adc_array_wafflecap_8_0[11|9]/sample_n rowoff_n[12] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|16] vcm ctop col[16] col_n[16] row_n[13] rowon_n[13] adc_array_wafflecap_8_0[12|9]/sample
+ adc_array_wafflecap_8_0[12|9]/sample_n rowoff_n[13] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|16] vcm ctop col[16] col_n[16] row_n[14] rowon_n[14] adc_array_wafflecap_8_0[13|9]/sample
+ adc_array_wafflecap_8_0[13|9]/sample_n rowoff_n[14] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|16] vcm ctop col[16] col_n[16] row_n[15] rowon_n[15] adc_array_wafflecap_8_0[14|9]/sample
+ adc_array_wafflecap_8_0[14|9]/sample_n rowoff_n[15] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|17] vcm ctop col[17] col_n[17] row_n[1] rowon_n[1] adc_array_wafflecap_8_0[0|9]/sample
+ adc_array_wafflecap_8_0[0|9]/sample_n rowoff_n[1] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|17] vcm ctop col[17] col_n[17] row_n[2] rowon_n[2] adc_array_wafflecap_8_0[1|9]/sample
+ adc_array_wafflecap_8_0[1|9]/sample_n rowoff_n[2] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|17] vcm ctop col[17] col_n[17] row_n[3] rowon_n[3] adc_array_wafflecap_8_0[2|9]/sample
+ adc_array_wafflecap_8_0[2|9]/sample_n rowoff_n[3] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|17] vcm ctop col[17] col_n[17] row_n[4] rowon_n[4] adc_array_wafflecap_8_0[3|9]/sample
+ adc_array_wafflecap_8_0[3|9]/sample_n rowoff_n[4] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|17] vcm ctop col[17] col_n[17] row_n[5] rowon_n[5] adc_array_wafflecap_8_0[4|9]/sample
+ adc_array_wafflecap_8_0[4|9]/sample_n rowoff_n[5] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|17] vcm ctop col[17] col_n[17] row_n[6] rowon_n[6] adc_array_wafflecap_8_0[5|9]/sample
+ adc_array_wafflecap_8_0[5|9]/sample_n rowoff_n[6] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|17] vcm ctop col[17] col_n[17] row_n[7] rowon_n[7] adc_array_wafflecap_8_0[6|9]/sample
+ adc_array_wafflecap_8_0[6|9]/sample_n rowoff_n[7] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|17] vcm ctop col[17] col_n[17] row_n[8] rowon_n[8] adc_array_wafflecap_8_0[7|9]/sample
+ adc_array_wafflecap_8_0[7|9]/sample_n rowoff_n[8] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|17] vcm ctop col[17] col_n[17] row_n[9] rowon_n[9] adc_array_wafflecap_8_0[8|9]/sample
+ adc_array_wafflecap_8_0[8|9]/sample_n rowoff_n[9] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|17] vcm ctop col[17] col_n[17] row_n[10] rowon_n[10] adc_array_wafflecap_8_0[9|9]/sample
+ adc_array_wafflecap_8_0[9|9]/sample_n rowoff_n[10] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|17] vcm ctop col[17] col_n[17] row_n[11] rowon_n[11] adc_array_wafflecap_8_0[10|9]/sample
+ adc_array_wafflecap_8_0[10|9]/sample_n rowoff_n[11] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|17] vcm ctop col[17] col_n[17] row_n[12] rowon_n[12] adc_array_wafflecap_8_0[11|9]/sample
+ adc_array_wafflecap_8_0[11|9]/sample_n rowoff_n[12] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|17] vcm ctop col[17] col_n[17] row_n[13] rowon_n[13] adc_array_wafflecap_8_0[12|9]/sample
+ adc_array_wafflecap_8_0[12|9]/sample_n rowoff_n[13] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|17] vcm ctop col[17] col_n[17] row_n[14] rowon_n[14] adc_array_wafflecap_8_0[13|9]/sample
+ adc_array_wafflecap_8_0[13|9]/sample_n rowoff_n[14] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|17] vcm ctop col[17] col_n[17] row_n[15] rowon_n[15] adc_array_wafflecap_8_0[14|9]/sample
+ adc_array_wafflecap_8_0[14|9]/sample_n rowoff_n[15] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|18] vcm ctop col[18] col_n[18] row_n[1] rowon_n[1] adc_array_wafflecap_8_0[0|9]/sample
+ adc_array_wafflecap_8_0[0|9]/sample_n rowoff_n[1] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|18] vcm ctop col[18] col_n[18] row_n[2] rowon_n[2] adc_array_wafflecap_8_0[1|9]/sample
+ adc_array_wafflecap_8_0[1|9]/sample_n rowoff_n[2] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|18] vcm ctop col[18] col_n[18] row_n[3] rowon_n[3] adc_array_wafflecap_8_0[2|9]/sample
+ adc_array_wafflecap_8_0[2|9]/sample_n rowoff_n[3] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|18] vcm ctop col[18] col_n[18] row_n[4] rowon_n[4] adc_array_wafflecap_8_0[3|9]/sample
+ adc_array_wafflecap_8_0[3|9]/sample_n rowoff_n[4] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|18] vcm ctop col[18] col_n[18] row_n[5] rowon_n[5] adc_array_wafflecap_8_0[4|9]/sample
+ adc_array_wafflecap_8_0[4|9]/sample_n rowoff_n[5] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|18] vcm ctop col[18] col_n[18] row_n[6] rowon_n[6] adc_array_wafflecap_8_0[5|9]/sample
+ adc_array_wafflecap_8_0[5|9]/sample_n rowoff_n[6] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|18] vcm ctop col[18] col_n[18] row_n[7] rowon_n[7] adc_array_wafflecap_8_0[6|9]/sample
+ adc_array_wafflecap_8_0[6|9]/sample_n rowoff_n[7] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|18] vcm ctop col[18] col_n[18] row_n[8] rowon_n[8] adc_array_wafflecap_8_0[7|9]/sample
+ adc_array_wafflecap_8_0[7|9]/sample_n rowoff_n[8] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|18] vcm ctop col[18] col_n[18] row_n[9] rowon_n[9] adc_array_wafflecap_8_0[8|9]/sample
+ adc_array_wafflecap_8_0[8|9]/sample_n rowoff_n[9] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|18] vcm ctop col[18] col_n[18] row_n[10] rowon_n[10] adc_array_wafflecap_8_0[9|9]/sample
+ adc_array_wafflecap_8_0[9|9]/sample_n rowoff_n[10] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|18] vcm ctop col[18] col_n[18] row_n[11] rowon_n[11] adc_array_wafflecap_8_0[10|9]/sample
+ adc_array_wafflecap_8_0[10|9]/sample_n rowoff_n[11] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|18] vcm ctop col[18] col_n[18] row_n[12] rowon_n[12] adc_array_wafflecap_8_0[11|9]/sample
+ adc_array_wafflecap_8_0[11|9]/sample_n rowoff_n[12] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|18] vcm ctop col[18] col_n[18] row_n[13] rowon_n[13] adc_array_wafflecap_8_0[12|9]/sample
+ adc_array_wafflecap_8_0[12|9]/sample_n rowoff_n[13] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|18] vcm ctop col[18] col_n[18] row_n[14] rowon_n[14] adc_array_wafflecap_8_0[13|9]/sample
+ adc_array_wafflecap_8_0[13|9]/sample_n rowoff_n[14] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|18] vcm ctop col[18] col_n[18] row_n[15] rowon_n[15] adc_array_wafflecap_8_0[14|9]/sample
+ adc_array_wafflecap_8_0[14|9]/sample_n rowoff_n[15] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|19] vcm ctop col[19] col_n[19] row_n[1] rowon_n[1] adc_array_wafflecap_8_0[0|9]/sample
+ adc_array_wafflecap_8_0[0|9]/sample_n rowoff_n[1] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|19] vcm ctop col[19] col_n[19] row_n[2] rowon_n[2] adc_array_wafflecap_8_0[1|9]/sample
+ adc_array_wafflecap_8_0[1|9]/sample_n rowoff_n[2] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|19] vcm ctop col[19] col_n[19] row_n[3] rowon_n[3] adc_array_wafflecap_8_0[2|9]/sample
+ adc_array_wafflecap_8_0[2|9]/sample_n rowoff_n[3] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|19] vcm ctop col[19] col_n[19] row_n[4] rowon_n[4] adc_array_wafflecap_8_0[3|9]/sample
+ adc_array_wafflecap_8_0[3|9]/sample_n rowoff_n[4] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|19] vcm ctop col[19] col_n[19] row_n[5] rowon_n[5] adc_array_wafflecap_8_0[4|9]/sample
+ adc_array_wafflecap_8_0[4|9]/sample_n rowoff_n[5] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|19] vcm ctop col[19] col_n[19] row_n[6] rowon_n[6] adc_array_wafflecap_8_0[5|9]/sample
+ adc_array_wafflecap_8_0[5|9]/sample_n rowoff_n[6] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|19] vcm ctop col[19] col_n[19] row_n[7] rowon_n[7] adc_array_wafflecap_8_0[6|9]/sample
+ adc_array_wafflecap_8_0[6|9]/sample_n rowoff_n[7] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|19] vcm ctop col[19] col_n[19] row_n[8] rowon_n[8] adc_array_wafflecap_8_0[7|9]/sample
+ adc_array_wafflecap_8_0[7|9]/sample_n rowoff_n[8] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|19] vcm ctop col[19] col_n[19] row_n[9] rowon_n[9] adc_array_wafflecap_8_0[8|9]/sample
+ adc_array_wafflecap_8_0[8|9]/sample_n rowoff_n[9] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|19] vcm ctop col[19] col_n[19] row_n[10] rowon_n[10] adc_array_wafflecap_8_0[9|9]/sample
+ adc_array_wafflecap_8_0[9|9]/sample_n rowoff_n[10] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|19] vcm ctop col[19] col_n[19] row_n[11] rowon_n[11] adc_array_wafflecap_8_0[10|9]/sample
+ adc_array_wafflecap_8_0[10|9]/sample_n rowoff_n[11] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|19] vcm ctop col[19] col_n[19] row_n[12] rowon_n[12] adc_array_wafflecap_8_0[11|9]/sample
+ adc_array_wafflecap_8_0[11|9]/sample_n rowoff_n[12] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|19] vcm ctop col[19] col_n[19] row_n[13] rowon_n[13] adc_array_wafflecap_8_0[12|9]/sample
+ adc_array_wafflecap_8_0[12|9]/sample_n rowoff_n[13] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|19] vcm ctop col[19] col_n[19] row_n[14] rowon_n[14] adc_array_wafflecap_8_0[13|9]/sample
+ adc_array_wafflecap_8_0[13|9]/sample_n rowoff_n[14] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|19] vcm ctop col[19] col_n[19] row_n[15] rowon_n[15] adc_array_wafflecap_8_0[14|9]/sample
+ adc_array_wafflecap_8_0[14|9]/sample_n rowoff_n[15] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|20] vcm ctop col[20] col_n[20] row_n[1] rowon_n[1] adc_array_wafflecap_8_0[0|9]/sample
+ adc_array_wafflecap_8_0[0|9]/sample_n rowoff_n[1] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|20] vcm ctop col[20] col_n[20] row_n[2] rowon_n[2] adc_array_wafflecap_8_0[1|9]/sample
+ adc_array_wafflecap_8_0[1|9]/sample_n rowoff_n[2] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|20] vcm ctop col[20] col_n[20] row_n[3] rowon_n[3] adc_array_wafflecap_8_0[2|9]/sample
+ adc_array_wafflecap_8_0[2|9]/sample_n rowoff_n[3] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|20] vcm ctop col[20] col_n[20] row_n[4] rowon_n[4] adc_array_wafflecap_8_0[3|9]/sample
+ adc_array_wafflecap_8_0[3|9]/sample_n rowoff_n[4] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|20] vcm ctop col[20] col_n[20] row_n[5] rowon_n[5] adc_array_wafflecap_8_0[4|9]/sample
+ adc_array_wafflecap_8_0[4|9]/sample_n rowoff_n[5] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|20] vcm ctop col[20] col_n[20] row_n[6] rowon_n[6] adc_array_wafflecap_8_0[5|9]/sample
+ adc_array_wafflecap_8_0[5|9]/sample_n rowoff_n[6] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|20] vcm ctop col[20] col_n[20] row_n[7] rowon_n[7] adc_array_wafflecap_8_0[6|9]/sample
+ adc_array_wafflecap_8_0[6|9]/sample_n rowoff_n[7] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|20] vcm ctop col[20] col_n[20] row_n[8] rowon_n[8] adc_array_wafflecap_8_0[7|9]/sample
+ adc_array_wafflecap_8_0[7|9]/sample_n rowoff_n[8] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|20] vcm ctop col[20] col_n[20] row_n[9] rowon_n[9] adc_array_wafflecap_8_0[8|9]/sample
+ adc_array_wafflecap_8_0[8|9]/sample_n rowoff_n[9] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|20] vcm ctop col[20] col_n[20] row_n[10] rowon_n[10] adc_array_wafflecap_8_0[9|9]/sample
+ adc_array_wafflecap_8_0[9|9]/sample_n rowoff_n[10] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|20] vcm ctop col[20] col_n[20] row_n[11] rowon_n[11] adc_array_wafflecap_8_0[10|9]/sample
+ adc_array_wafflecap_8_0[10|9]/sample_n rowoff_n[11] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|20] vcm ctop col[20] col_n[20] row_n[12] rowon_n[12] adc_array_wafflecap_8_0[11|9]/sample
+ adc_array_wafflecap_8_0[11|9]/sample_n rowoff_n[12] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|20] vcm ctop col[20] col_n[20] row_n[13] rowon_n[13] adc_array_wafflecap_8_0[12|9]/sample
+ adc_array_wafflecap_8_0[12|9]/sample_n rowoff_n[13] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|20] vcm ctop col[20] col_n[20] row_n[14] rowon_n[14] adc_array_wafflecap_8_0[13|9]/sample
+ adc_array_wafflecap_8_0[13|9]/sample_n rowoff_n[14] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|20] vcm ctop col[20] col_n[20] row_n[15] rowon_n[15] adc_array_wafflecap_8_0[14|9]/sample
+ adc_array_wafflecap_8_0[14|9]/sample_n rowoff_n[15] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|21] vcm ctop col[21] col_n[21] row_n[1] rowon_n[1] adc_array_wafflecap_8_0[0|9]/sample
+ adc_array_wafflecap_8_0[0|9]/sample_n rowoff_n[1] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|21] vcm ctop col[21] col_n[21] row_n[2] rowon_n[2] adc_array_wafflecap_8_0[1|9]/sample
+ adc_array_wafflecap_8_0[1|9]/sample_n rowoff_n[2] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|21] vcm ctop col[21] col_n[21] row_n[3] rowon_n[3] adc_array_wafflecap_8_0[2|9]/sample
+ adc_array_wafflecap_8_0[2|9]/sample_n rowoff_n[3] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|21] vcm ctop col[21] col_n[21] row_n[4] rowon_n[4] adc_array_wafflecap_8_0[3|9]/sample
+ adc_array_wafflecap_8_0[3|9]/sample_n rowoff_n[4] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|21] vcm ctop col[21] col_n[21] row_n[5] rowon_n[5] adc_array_wafflecap_8_0[4|9]/sample
+ adc_array_wafflecap_8_0[4|9]/sample_n rowoff_n[5] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|21] vcm ctop col[21] col_n[21] row_n[6] rowon_n[6] adc_array_wafflecap_8_0[5|9]/sample
+ adc_array_wafflecap_8_0[5|9]/sample_n rowoff_n[6] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|21] vcm ctop col[21] col_n[21] row_n[7] rowon_n[7] adc_array_wafflecap_8_0[6|9]/sample
+ adc_array_wafflecap_8_0[6|9]/sample_n rowoff_n[7] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|21] vcm ctop col[21] col_n[21] row_n[8] rowon_n[8] adc_array_wafflecap_8_0[7|9]/sample
+ adc_array_wafflecap_8_0[7|9]/sample_n rowoff_n[8] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|21] vcm ctop col[21] col_n[21] row_n[9] rowon_n[9] adc_array_wafflecap_8_0[8|9]/sample
+ adc_array_wafflecap_8_0[8|9]/sample_n rowoff_n[9] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|21] vcm ctop col[21] col_n[21] row_n[10] rowon_n[10] adc_array_wafflecap_8_0[9|9]/sample
+ adc_array_wafflecap_8_0[9|9]/sample_n rowoff_n[10] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|21] vcm ctop col[21] col_n[21] row_n[11] rowon_n[11] adc_array_wafflecap_8_0[10|9]/sample
+ adc_array_wafflecap_8_0[10|9]/sample_n rowoff_n[11] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|21] vcm ctop col[21] col_n[21] row_n[12] rowon_n[12] adc_array_wafflecap_8_0[11|9]/sample
+ adc_array_wafflecap_8_0[11|9]/sample_n rowoff_n[12] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|21] vcm ctop col[21] col_n[21] row_n[13] rowon_n[13] adc_array_wafflecap_8_0[12|9]/sample
+ adc_array_wafflecap_8_0[12|9]/sample_n rowoff_n[13] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|21] vcm ctop col[21] col_n[21] row_n[14] rowon_n[14] adc_array_wafflecap_8_0[13|9]/sample
+ adc_array_wafflecap_8_0[13|9]/sample_n rowoff_n[14] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|21] vcm ctop col[21] col_n[21] row_n[15] rowon_n[15] adc_array_wafflecap_8_0[14|9]/sample
+ adc_array_wafflecap_8_0[14|9]/sample_n rowoff_n[15] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|22] vcm ctop col[22] col_n[22] row_n[1] rowon_n[1] adc_array_wafflecap_8_0[0|9]/sample
+ adc_array_wafflecap_8_0[0|9]/sample_n rowoff_n[1] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|22] vcm ctop col[22] col_n[22] row_n[2] rowon_n[2] adc_array_wafflecap_8_0[1|9]/sample
+ adc_array_wafflecap_8_0[1|9]/sample_n rowoff_n[2] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|22] vcm ctop col[22] col_n[22] row_n[3] rowon_n[3] adc_array_wafflecap_8_0[2|9]/sample
+ adc_array_wafflecap_8_0[2|9]/sample_n rowoff_n[3] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|22] vcm ctop col[22] col_n[22] row_n[4] rowon_n[4] adc_array_wafflecap_8_0[3|9]/sample
+ adc_array_wafflecap_8_0[3|9]/sample_n rowoff_n[4] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|22] vcm ctop col[22] col_n[22] row_n[5] rowon_n[5] adc_array_wafflecap_8_0[4|9]/sample
+ adc_array_wafflecap_8_0[4|9]/sample_n rowoff_n[5] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|22] vcm ctop col[22] col_n[22] row_n[6] rowon_n[6] adc_array_wafflecap_8_0[5|9]/sample
+ adc_array_wafflecap_8_0[5|9]/sample_n rowoff_n[6] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|22] vcm ctop col[22] col_n[22] row_n[7] rowon_n[7] adc_array_wafflecap_8_0[6|9]/sample
+ adc_array_wafflecap_8_0[6|9]/sample_n rowoff_n[7] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|22] vcm ctop col[22] col_n[22] row_n[8] rowon_n[8] adc_array_wafflecap_8_0[7|9]/sample
+ adc_array_wafflecap_8_0[7|9]/sample_n rowoff_n[8] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|22] vcm ctop col[22] col_n[22] row_n[9] rowon_n[9] adc_array_wafflecap_8_0[8|9]/sample
+ adc_array_wafflecap_8_0[8|9]/sample_n rowoff_n[9] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|22] vcm ctop col[22] col_n[22] row_n[10] rowon_n[10] adc_array_wafflecap_8_0[9|9]/sample
+ adc_array_wafflecap_8_0[9|9]/sample_n rowoff_n[10] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|22] vcm ctop col[22] col_n[22] row_n[11] rowon_n[11] adc_array_wafflecap_8_0[10|9]/sample
+ adc_array_wafflecap_8_0[10|9]/sample_n rowoff_n[11] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|22] vcm ctop col[22] col_n[22] row_n[12] rowon_n[12] adc_array_wafflecap_8_0[11|9]/sample
+ adc_array_wafflecap_8_0[11|9]/sample_n rowoff_n[12] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|22] vcm ctop col[22] col_n[22] row_n[13] rowon_n[13] adc_array_wafflecap_8_0[12|9]/sample
+ adc_array_wafflecap_8_0[12|9]/sample_n rowoff_n[13] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|22] vcm ctop col[22] col_n[22] row_n[14] rowon_n[14] adc_array_wafflecap_8_0[13|9]/sample
+ adc_array_wafflecap_8_0[13|9]/sample_n rowoff_n[14] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|22] vcm ctop col[22] col_n[22] row_n[15] rowon_n[15] adc_array_wafflecap_8_0[14|9]/sample
+ adc_array_wafflecap_8_0[14|9]/sample_n rowoff_n[15] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|23] vcm ctop col[23] col_n[23] row_n[1] rowon_n[1] adc_array_wafflecap_8_0[0|9]/sample
+ adc_array_wafflecap_8_0[0|9]/sample_n rowoff_n[1] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|23] vcm ctop col[23] col_n[23] row_n[2] rowon_n[2] adc_array_wafflecap_8_0[1|9]/sample
+ adc_array_wafflecap_8_0[1|9]/sample_n rowoff_n[2] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|23] vcm ctop col[23] col_n[23] row_n[3] rowon_n[3] adc_array_wafflecap_8_0[2|9]/sample
+ adc_array_wafflecap_8_0[2|9]/sample_n rowoff_n[3] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|23] vcm ctop col[23] col_n[23] row_n[4] rowon_n[4] adc_array_wafflecap_8_0[3|9]/sample
+ adc_array_wafflecap_8_0[3|9]/sample_n rowoff_n[4] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|23] vcm ctop col[23] col_n[23] row_n[5] rowon_n[5] adc_array_wafflecap_8_0[4|9]/sample
+ adc_array_wafflecap_8_0[4|9]/sample_n rowoff_n[5] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|23] vcm ctop col[23] col_n[23] row_n[6] rowon_n[6] adc_array_wafflecap_8_0[5|9]/sample
+ adc_array_wafflecap_8_0[5|9]/sample_n rowoff_n[6] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|23] vcm ctop col[23] col_n[23] row_n[7] rowon_n[7] adc_array_wafflecap_8_0[6|9]/sample
+ adc_array_wafflecap_8_0[6|9]/sample_n rowoff_n[7] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|23] vcm ctop col[23] col_n[23] row_n[8] rowon_n[8] adc_array_wafflecap_8_0[7|9]/sample
+ adc_array_wafflecap_8_0[7|9]/sample_n rowoff_n[8] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|23] vcm ctop col[23] col_n[23] row_n[9] rowon_n[9] adc_array_wafflecap_8_0[8|9]/sample
+ adc_array_wafflecap_8_0[8|9]/sample_n rowoff_n[9] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|23] vcm ctop col[23] col_n[23] row_n[10] rowon_n[10] adc_array_wafflecap_8_0[9|9]/sample
+ adc_array_wafflecap_8_0[9|9]/sample_n rowoff_n[10] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|23] vcm ctop col[23] col_n[23] row_n[11] rowon_n[11] adc_array_wafflecap_8_0[10|9]/sample
+ adc_array_wafflecap_8_0[10|9]/sample_n rowoff_n[11] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|23] vcm ctop col[23] col_n[23] row_n[12] rowon_n[12] adc_array_wafflecap_8_0[11|9]/sample
+ adc_array_wafflecap_8_0[11|9]/sample_n rowoff_n[12] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|23] vcm ctop col[23] col_n[23] row_n[13] rowon_n[13] adc_array_wafflecap_8_0[12|9]/sample
+ adc_array_wafflecap_8_0[12|9]/sample_n rowoff_n[13] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|23] vcm ctop col[23] col_n[23] row_n[14] rowon_n[14] adc_array_wafflecap_8_0[13|9]/sample
+ adc_array_wafflecap_8_0[13|9]/sample_n rowoff_n[14] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|23] vcm ctop col[23] col_n[23] row_n[15] rowon_n[15] adc_array_wafflecap_8_0[14|9]/sample
+ adc_array_wafflecap_8_0[14|9]/sample_n rowoff_n[15] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|24] vcm ctop col[24] col_n[24] row_n[1] rowon_n[1] adc_array_wafflecap_8_0[0|9]/sample
+ adc_array_wafflecap_8_0[0|9]/sample_n rowoff_n[1] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|24] vcm ctop col[24] col_n[24] row_n[2] rowon_n[2] adc_array_wafflecap_8_0[1|9]/sample
+ adc_array_wafflecap_8_0[1|9]/sample_n rowoff_n[2] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|24] vcm ctop col[24] col_n[24] row_n[3] rowon_n[3] adc_array_wafflecap_8_0[2|9]/sample
+ adc_array_wafflecap_8_0[2|9]/sample_n rowoff_n[3] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|24] vcm ctop col[24] col_n[24] row_n[4] rowon_n[4] adc_array_wafflecap_8_0[3|9]/sample
+ adc_array_wafflecap_8_0[3|9]/sample_n rowoff_n[4] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|24] vcm ctop col[24] col_n[24] row_n[5] rowon_n[5] adc_array_wafflecap_8_0[4|9]/sample
+ adc_array_wafflecap_8_0[4|9]/sample_n rowoff_n[5] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|24] vcm ctop col[24] col_n[24] row_n[6] rowon_n[6] adc_array_wafflecap_8_0[5|9]/sample
+ adc_array_wafflecap_8_0[5|9]/sample_n rowoff_n[6] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|24] vcm ctop col[24] col_n[24] row_n[7] rowon_n[7] adc_array_wafflecap_8_0[6|9]/sample
+ adc_array_wafflecap_8_0[6|9]/sample_n rowoff_n[7] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|24] vcm ctop col[24] col_n[24] row_n[8] rowon_n[8] adc_array_wafflecap_8_0[7|9]/sample
+ adc_array_wafflecap_8_0[7|9]/sample_n rowoff_n[8] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|24] vcm ctop col[24] col_n[24] row_n[9] rowon_n[9] adc_array_wafflecap_8_0[8|9]/sample
+ adc_array_wafflecap_8_0[8|9]/sample_n rowoff_n[9] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|24] vcm ctop col[24] col_n[24] row_n[10] rowon_n[10] adc_array_wafflecap_8_0[9|9]/sample
+ adc_array_wafflecap_8_0[9|9]/sample_n rowoff_n[10] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|24] vcm ctop col[24] col_n[24] row_n[11] rowon_n[11] adc_array_wafflecap_8_0[10|9]/sample
+ adc_array_wafflecap_8_0[10|9]/sample_n rowoff_n[11] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|24] vcm ctop col[24] col_n[24] row_n[12] rowon_n[12] adc_array_wafflecap_8_0[11|9]/sample
+ adc_array_wafflecap_8_0[11|9]/sample_n rowoff_n[12] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|24] vcm ctop col[24] col_n[24] row_n[13] rowon_n[13] adc_array_wafflecap_8_0[12|9]/sample
+ adc_array_wafflecap_8_0[12|9]/sample_n rowoff_n[13] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|24] vcm ctop col[24] col_n[24] row_n[14] rowon_n[14] adc_array_wafflecap_8_0[13|9]/sample
+ adc_array_wafflecap_8_0[13|9]/sample_n rowoff_n[14] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|24] vcm ctop col[24] col_n[24] row_n[15] rowon_n[15] adc_array_wafflecap_8_0[14|9]/sample
+ adc_array_wafflecap_8_0[14|9]/sample_n rowoff_n[15] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|25] vcm ctop col[25] col_n[25] row_n[1] rowon_n[1] adc_array_wafflecap_8_0[0|9]/sample
+ adc_array_wafflecap_8_0[0|9]/sample_n rowoff_n[1] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|25] vcm ctop col[25] col_n[25] row_n[2] rowon_n[2] adc_array_wafflecap_8_0[1|9]/sample
+ adc_array_wafflecap_8_0[1|9]/sample_n rowoff_n[2] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|25] vcm ctop col[25] col_n[25] row_n[3] rowon_n[3] adc_array_wafflecap_8_0[2|9]/sample
+ adc_array_wafflecap_8_0[2|9]/sample_n rowoff_n[3] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|25] vcm ctop col[25] col_n[25] row_n[4] rowon_n[4] adc_array_wafflecap_8_0[3|9]/sample
+ adc_array_wafflecap_8_0[3|9]/sample_n rowoff_n[4] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|25] vcm ctop col[25] col_n[25] row_n[5] rowon_n[5] adc_array_wafflecap_8_0[4|9]/sample
+ adc_array_wafflecap_8_0[4|9]/sample_n rowoff_n[5] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|25] vcm ctop col[25] col_n[25] row_n[6] rowon_n[6] adc_array_wafflecap_8_0[5|9]/sample
+ adc_array_wafflecap_8_0[5|9]/sample_n rowoff_n[6] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|25] vcm ctop col[25] col_n[25] row_n[7] rowon_n[7] adc_array_wafflecap_8_0[6|9]/sample
+ adc_array_wafflecap_8_0[6|9]/sample_n rowoff_n[7] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|25] vcm ctop col[25] col_n[25] row_n[8] rowon_n[8] adc_array_wafflecap_8_0[7|9]/sample
+ adc_array_wafflecap_8_0[7|9]/sample_n rowoff_n[8] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|25] vcm ctop col[25] col_n[25] row_n[9] rowon_n[9] adc_array_wafflecap_8_0[8|9]/sample
+ adc_array_wafflecap_8_0[8|9]/sample_n rowoff_n[9] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|25] vcm ctop col[25] col_n[25] row_n[10] rowon_n[10] adc_array_wafflecap_8_0[9|9]/sample
+ adc_array_wafflecap_8_0[9|9]/sample_n rowoff_n[10] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|25] vcm ctop col[25] col_n[25] row_n[11] rowon_n[11] adc_array_wafflecap_8_0[10|9]/sample
+ adc_array_wafflecap_8_0[10|9]/sample_n rowoff_n[11] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|25] vcm ctop col[25] col_n[25] row_n[12] rowon_n[12] adc_array_wafflecap_8_0[11|9]/sample
+ adc_array_wafflecap_8_0[11|9]/sample_n rowoff_n[12] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|25] vcm ctop col[25] col_n[25] row_n[13] rowon_n[13] adc_array_wafflecap_8_0[12|9]/sample
+ adc_array_wafflecap_8_0[12|9]/sample_n rowoff_n[13] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|25] vcm ctop col[25] col_n[25] row_n[14] rowon_n[14] adc_array_wafflecap_8_0[13|9]/sample
+ adc_array_wafflecap_8_0[13|9]/sample_n rowoff_n[14] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|25] vcm ctop col[25] col_n[25] row_n[15] rowon_n[15] adc_array_wafflecap_8_0[14|9]/sample
+ adc_array_wafflecap_8_0[14|9]/sample_n rowoff_n[15] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|26] vcm ctop col[26] col_n[26] row_n[1] rowon_n[1] adc_array_wafflecap_8_0[0|9]/sample
+ adc_array_wafflecap_8_0[0|9]/sample_n rowoff_n[1] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|26] vcm ctop col[26] col_n[26] row_n[2] rowon_n[2] adc_array_wafflecap_8_0[1|9]/sample
+ adc_array_wafflecap_8_0[1|9]/sample_n rowoff_n[2] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|26] vcm ctop col[26] col_n[26] row_n[3] rowon_n[3] adc_array_wafflecap_8_0[2|9]/sample
+ adc_array_wafflecap_8_0[2|9]/sample_n rowoff_n[3] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|26] vcm ctop col[26] col_n[26] row_n[4] rowon_n[4] adc_array_wafflecap_8_0[3|9]/sample
+ adc_array_wafflecap_8_0[3|9]/sample_n rowoff_n[4] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|26] vcm ctop col[26] col_n[26] row_n[5] rowon_n[5] adc_array_wafflecap_8_0[4|9]/sample
+ adc_array_wafflecap_8_0[4|9]/sample_n rowoff_n[5] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|26] vcm ctop col[26] col_n[26] row_n[6] rowon_n[6] adc_array_wafflecap_8_0[5|9]/sample
+ adc_array_wafflecap_8_0[5|9]/sample_n rowoff_n[6] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|26] vcm ctop col[26] col_n[26] row_n[7] rowon_n[7] adc_array_wafflecap_8_0[6|9]/sample
+ adc_array_wafflecap_8_0[6|9]/sample_n rowoff_n[7] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|26] vcm ctop col[26] col_n[26] row_n[8] rowon_n[8] adc_array_wafflecap_8_0[7|9]/sample
+ adc_array_wafflecap_8_0[7|9]/sample_n rowoff_n[8] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|26] vcm ctop col[26] col_n[26] row_n[9] rowon_n[9] adc_array_wafflecap_8_0[8|9]/sample
+ adc_array_wafflecap_8_0[8|9]/sample_n rowoff_n[9] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|26] vcm ctop col[26] col_n[26] row_n[10] rowon_n[10] adc_array_wafflecap_8_0[9|9]/sample
+ adc_array_wafflecap_8_0[9|9]/sample_n rowoff_n[10] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|26] vcm ctop col[26] col_n[26] row_n[11] rowon_n[11] adc_array_wafflecap_8_0[10|9]/sample
+ adc_array_wafflecap_8_0[10|9]/sample_n rowoff_n[11] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|26] vcm ctop col[26] col_n[26] row_n[12] rowon_n[12] adc_array_wafflecap_8_0[11|9]/sample
+ adc_array_wafflecap_8_0[11|9]/sample_n rowoff_n[12] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|26] vcm ctop col[26] col_n[26] row_n[13] rowon_n[13] adc_array_wafflecap_8_0[12|9]/sample
+ adc_array_wafflecap_8_0[12|9]/sample_n rowoff_n[13] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|26] vcm ctop col[26] col_n[26] row_n[14] rowon_n[14] adc_array_wafflecap_8_0[13|9]/sample
+ adc_array_wafflecap_8_0[13|9]/sample_n rowoff_n[14] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|26] vcm ctop col[26] col_n[26] row_n[15] rowon_n[15] adc_array_wafflecap_8_0[14|9]/sample
+ adc_array_wafflecap_8_0[14|9]/sample_n rowoff_n[15] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|27] vcm ctop col[27] col_n[27] row_n[1] rowon_n[1] adc_array_wafflecap_8_0[0|9]/sample
+ adc_array_wafflecap_8_0[0|9]/sample_n rowoff_n[1] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|27] vcm ctop col[27] col_n[27] row_n[2] rowon_n[2] adc_array_wafflecap_8_0[1|9]/sample
+ adc_array_wafflecap_8_0[1|9]/sample_n rowoff_n[2] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|27] vcm ctop col[27] col_n[27] row_n[3] rowon_n[3] adc_array_wafflecap_8_0[2|9]/sample
+ adc_array_wafflecap_8_0[2|9]/sample_n rowoff_n[3] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|27] vcm ctop col[27] col_n[27] row_n[4] rowon_n[4] adc_array_wafflecap_8_0[3|9]/sample
+ adc_array_wafflecap_8_0[3|9]/sample_n rowoff_n[4] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|27] vcm ctop col[27] col_n[27] row_n[5] rowon_n[5] adc_array_wafflecap_8_0[4|9]/sample
+ adc_array_wafflecap_8_0[4|9]/sample_n rowoff_n[5] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|27] vcm ctop col[27] col_n[27] row_n[6] rowon_n[6] adc_array_wafflecap_8_0[5|9]/sample
+ adc_array_wafflecap_8_0[5|9]/sample_n rowoff_n[6] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|27] vcm ctop col[27] col_n[27] row_n[7] rowon_n[7] adc_array_wafflecap_8_0[6|9]/sample
+ adc_array_wafflecap_8_0[6|9]/sample_n rowoff_n[7] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|27] vcm ctop col[27] col_n[27] row_n[8] rowon_n[8] adc_array_wafflecap_8_0[7|9]/sample
+ adc_array_wafflecap_8_0[7|9]/sample_n rowoff_n[8] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|27] vcm ctop col[27] col_n[27] row_n[9] rowon_n[9] adc_array_wafflecap_8_0[8|9]/sample
+ adc_array_wafflecap_8_0[8|9]/sample_n rowoff_n[9] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|27] vcm ctop col[27] col_n[27] row_n[10] rowon_n[10] adc_array_wafflecap_8_0[9|9]/sample
+ adc_array_wafflecap_8_0[9|9]/sample_n rowoff_n[10] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|27] vcm ctop col[27] col_n[27] row_n[11] rowon_n[11] adc_array_wafflecap_8_0[10|9]/sample
+ adc_array_wafflecap_8_0[10|9]/sample_n rowoff_n[11] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|27] vcm ctop col[27] col_n[27] row_n[12] rowon_n[12] adc_array_wafflecap_8_0[11|9]/sample
+ adc_array_wafflecap_8_0[11|9]/sample_n rowoff_n[12] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|27] vcm ctop col[27] col_n[27] row_n[13] rowon_n[13] adc_array_wafflecap_8_0[12|9]/sample
+ adc_array_wafflecap_8_0[12|9]/sample_n rowoff_n[13] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|27] vcm ctop col[27] col_n[27] row_n[14] rowon_n[14] adc_array_wafflecap_8_0[13|9]/sample
+ adc_array_wafflecap_8_0[13|9]/sample_n rowoff_n[14] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|27] vcm ctop col[27] col_n[27] row_n[15] rowon_n[15] adc_array_wafflecap_8_0[14|9]/sample
+ adc_array_wafflecap_8_0[14|9]/sample_n rowoff_n[15] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|28] vcm ctop col[28] col_n[28] row_n[1] rowon_n[1] adc_array_wafflecap_8_0[0|9]/sample
+ adc_array_wafflecap_8_0[0|9]/sample_n rowoff_n[1] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|28] vcm ctop col[28] col_n[28] row_n[2] rowon_n[2] adc_array_wafflecap_8_0[1|9]/sample
+ adc_array_wafflecap_8_0[1|9]/sample_n rowoff_n[2] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|28] vcm ctop col[28] col_n[28] row_n[3] rowon_n[3] adc_array_wafflecap_8_0[2|9]/sample
+ adc_array_wafflecap_8_0[2|9]/sample_n rowoff_n[3] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|28] vcm ctop col[28] col_n[28] row_n[4] rowon_n[4] adc_array_wafflecap_8_0[3|9]/sample
+ adc_array_wafflecap_8_0[3|9]/sample_n rowoff_n[4] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|28] vcm ctop col[28] col_n[28] row_n[5] rowon_n[5] adc_array_wafflecap_8_0[4|9]/sample
+ adc_array_wafflecap_8_0[4|9]/sample_n rowoff_n[5] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|28] vcm ctop col[28] col_n[28] row_n[6] rowon_n[6] adc_array_wafflecap_8_0[5|9]/sample
+ adc_array_wafflecap_8_0[5|9]/sample_n rowoff_n[6] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|28] vcm ctop col[28] col_n[28] row_n[7] rowon_n[7] adc_array_wafflecap_8_0[6|9]/sample
+ adc_array_wafflecap_8_0[6|9]/sample_n rowoff_n[7] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|28] vcm ctop col[28] col_n[28] row_n[8] rowon_n[8] adc_array_wafflecap_8_0[7|9]/sample
+ adc_array_wafflecap_8_0[7|9]/sample_n rowoff_n[8] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|28] vcm ctop col[28] col_n[28] row_n[9] rowon_n[9] adc_array_wafflecap_8_0[8|9]/sample
+ adc_array_wafflecap_8_0[8|9]/sample_n rowoff_n[9] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|28] vcm ctop col[28] col_n[28] row_n[10] rowon_n[10] adc_array_wafflecap_8_0[9|9]/sample
+ adc_array_wafflecap_8_0[9|9]/sample_n rowoff_n[10] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|28] vcm ctop col[28] col_n[28] row_n[11] rowon_n[11] adc_array_wafflecap_8_0[10|9]/sample
+ adc_array_wafflecap_8_0[10|9]/sample_n rowoff_n[11] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|28] vcm ctop col[28] col_n[28] row_n[12] rowon_n[12] adc_array_wafflecap_8_0[11|9]/sample
+ adc_array_wafflecap_8_0[11|9]/sample_n rowoff_n[12] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|28] vcm ctop col[28] col_n[28] row_n[13] rowon_n[13] adc_array_wafflecap_8_0[12|9]/sample
+ adc_array_wafflecap_8_0[12|9]/sample_n rowoff_n[13] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|28] vcm ctop col[28] col_n[28] row_n[14] rowon_n[14] adc_array_wafflecap_8_0[13|9]/sample
+ adc_array_wafflecap_8_0[13|9]/sample_n rowoff_n[14] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|28] vcm ctop col[28] col_n[28] row_n[15] rowon_n[15] adc_array_wafflecap_8_0[14|9]/sample
+ adc_array_wafflecap_8_0[14|9]/sample_n rowoff_n[15] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|29] vcm ctop col[29] col_n[29] row_n[1] rowon_n[1] adc_array_wafflecap_8_0[0|9]/sample
+ adc_array_wafflecap_8_0[0|9]/sample_n rowoff_n[1] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|29] vcm ctop col[29] col_n[29] row_n[2] rowon_n[2] adc_array_wafflecap_8_0[1|9]/sample
+ adc_array_wafflecap_8_0[1|9]/sample_n rowoff_n[2] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|29] vcm ctop col[29] col_n[29] row_n[3] rowon_n[3] adc_array_wafflecap_8_0[2|9]/sample
+ adc_array_wafflecap_8_0[2|9]/sample_n rowoff_n[3] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|29] vcm ctop col[29] col_n[29] row_n[4] rowon_n[4] adc_array_wafflecap_8_0[3|9]/sample
+ adc_array_wafflecap_8_0[3|9]/sample_n rowoff_n[4] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|29] vcm ctop col[29] col_n[29] row_n[5] rowon_n[5] adc_array_wafflecap_8_0[4|9]/sample
+ adc_array_wafflecap_8_0[4|9]/sample_n rowoff_n[5] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|29] vcm ctop col[29] col_n[29] row_n[6] rowon_n[6] adc_array_wafflecap_8_0[5|9]/sample
+ adc_array_wafflecap_8_0[5|9]/sample_n rowoff_n[6] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|29] vcm ctop col[29] col_n[29] row_n[7] rowon_n[7] adc_array_wafflecap_8_0[6|9]/sample
+ adc_array_wafflecap_8_0[6|9]/sample_n rowoff_n[7] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|29] vcm ctop col[29] col_n[29] row_n[8] rowon_n[8] adc_array_wafflecap_8_0[7|9]/sample
+ adc_array_wafflecap_8_0[7|9]/sample_n rowoff_n[8] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|29] vcm ctop col[29] col_n[29] row_n[9] rowon_n[9] adc_array_wafflecap_8_0[8|9]/sample
+ adc_array_wafflecap_8_0[8|9]/sample_n rowoff_n[9] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|29] vcm ctop col[29] col_n[29] row_n[10] rowon_n[10] adc_array_wafflecap_8_0[9|9]/sample
+ adc_array_wafflecap_8_0[9|9]/sample_n rowoff_n[10] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|29] vcm ctop col[29] col_n[29] row_n[11] rowon_n[11] adc_array_wafflecap_8_0[10|9]/sample
+ adc_array_wafflecap_8_0[10|9]/sample_n rowoff_n[11] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|29] vcm ctop col[29] col_n[29] row_n[12] rowon_n[12] adc_array_wafflecap_8_0[11|9]/sample
+ adc_array_wafflecap_8_0[11|9]/sample_n rowoff_n[12] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|29] vcm ctop col[29] col_n[29] row_n[13] rowon_n[13] adc_array_wafflecap_8_0[12|9]/sample
+ adc_array_wafflecap_8_0[12|9]/sample_n rowoff_n[13] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|29] vcm ctop col[29] col_n[29] row_n[14] rowon_n[14] adc_array_wafflecap_8_0[13|9]/sample
+ adc_array_wafflecap_8_0[13|9]/sample_n rowoff_n[14] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|29] vcm ctop col[29] col_n[29] row_n[15] rowon_n[15] adc_array_wafflecap_8_0[14|9]/sample
+ adc_array_wafflecap_8_0[14|9]/sample_n rowoff_n[15] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|30] vcm ctop col[30] col_n[30] row_n[1] rowon_n[1] adc_array_wafflecap_8_0[0|9]/sample
+ adc_array_wafflecap_8_0[0|9]/sample_n rowoff_n[1] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|30] vcm ctop col[30] col_n[30] row_n[2] rowon_n[2] adc_array_wafflecap_8_0[1|9]/sample
+ adc_array_wafflecap_8_0[1|9]/sample_n rowoff_n[2] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|30] vcm ctop col[30] col_n[30] row_n[3] rowon_n[3] adc_array_wafflecap_8_0[2|9]/sample
+ adc_array_wafflecap_8_0[2|9]/sample_n rowoff_n[3] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|30] vcm ctop col[30] col_n[30] row_n[4] rowon_n[4] adc_array_wafflecap_8_0[3|9]/sample
+ adc_array_wafflecap_8_0[3|9]/sample_n rowoff_n[4] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|30] vcm ctop col[30] col_n[30] row_n[5] rowon_n[5] adc_array_wafflecap_8_0[4|9]/sample
+ adc_array_wafflecap_8_0[4|9]/sample_n rowoff_n[5] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|30] vcm ctop col[30] col_n[30] row_n[6] rowon_n[6] adc_array_wafflecap_8_0[5|9]/sample
+ adc_array_wafflecap_8_0[5|9]/sample_n rowoff_n[6] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|30] vcm ctop col[30] col_n[30] row_n[7] rowon_n[7] adc_array_wafflecap_8_0[6|9]/sample
+ adc_array_wafflecap_8_0[6|9]/sample_n rowoff_n[7] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|30] vcm ctop col[30] col_n[30] row_n[8] rowon_n[8] adc_array_wafflecap_8_0[7|9]/sample
+ adc_array_wafflecap_8_0[7|9]/sample_n rowoff_n[8] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|30] vcm ctop col[30] col_n[30] row_n[9] rowon_n[9] adc_array_wafflecap_8_0[8|9]/sample
+ adc_array_wafflecap_8_0[8|9]/sample_n rowoff_n[9] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|30] vcm ctop col[30] col_n[30] row_n[10] rowon_n[10] adc_array_wafflecap_8_0[9|9]/sample
+ adc_array_wafflecap_8_0[9|9]/sample_n rowoff_n[10] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|30] vcm ctop col[30] col_n[30] row_n[11] rowon_n[11] adc_array_wafflecap_8_0[10|9]/sample
+ adc_array_wafflecap_8_0[10|9]/sample_n rowoff_n[11] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|30] vcm ctop col[30] col_n[30] row_n[12] rowon_n[12] adc_array_wafflecap_8_0[11|9]/sample
+ adc_array_wafflecap_8_0[11|9]/sample_n rowoff_n[12] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|30] vcm ctop col[30] col_n[30] row_n[13] rowon_n[13] adc_array_wafflecap_8_0[12|9]/sample
+ adc_array_wafflecap_8_0[12|9]/sample_n rowoff_n[13] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|30] vcm ctop col[30] col_n[30] row_n[14] rowon_n[14] adc_array_wafflecap_8_0[13|9]/sample
+ adc_array_wafflecap_8_0[13|9]/sample_n rowoff_n[14] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|30] vcm ctop col[30] col_n[30] row_n[15] rowon_n[15] adc_array_wafflecap_8_0[14|9]/sample
+ adc_array_wafflecap_8_0[14|9]/sample_n rowoff_n[15] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[0|31] vcm ctop col[31] col_n[31] row_n[1] rowon_n[1] adc_array_wafflecap_8_0[0|9]/sample
+ adc_array_wafflecap_8_0[0|9]/sample_n rowoff_n[1] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[1|31] vcm ctop col[31] col_n[31] row_n[2] rowon_n[2] adc_array_wafflecap_8_0[1|9]/sample
+ adc_array_wafflecap_8_0[1|9]/sample_n rowoff_n[2] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[2|31] vcm ctop col[31] col_n[31] row_n[3] rowon_n[3] adc_array_wafflecap_8_0[2|9]/sample
+ adc_array_wafflecap_8_0[2|9]/sample_n rowoff_n[3] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[3|31] vcm ctop col[31] col_n[31] row_n[4] rowon_n[4] adc_array_wafflecap_8_0[3|9]/sample
+ adc_array_wafflecap_8_0[3|9]/sample_n rowoff_n[4] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[4|31] vcm ctop col[31] col_n[31] row_n[5] rowon_n[5] adc_array_wafflecap_8_0[4|9]/sample
+ adc_array_wafflecap_8_0[4|9]/sample_n rowoff_n[5] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[5|31] vcm ctop col[31] col_n[31] row_n[6] rowon_n[6] adc_array_wafflecap_8_0[5|9]/sample
+ adc_array_wafflecap_8_0[5|9]/sample_n rowoff_n[6] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[6|31] vcm ctop col[31] col_n[31] row_n[7] rowon_n[7] adc_array_wafflecap_8_0[6|9]/sample
+ adc_array_wafflecap_8_0[6|9]/sample_n rowoff_n[7] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[7|31] vcm ctop col[31] col_n[31] row_n[8] rowon_n[8] adc_array_wafflecap_8_0[7|9]/sample
+ adc_array_wafflecap_8_0[7|9]/sample_n rowoff_n[8] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[8|31] vcm ctop col[31] col_n[31] row_n[9] rowon_n[9] adc_array_wafflecap_8_0[8|9]/sample
+ adc_array_wafflecap_8_0[8|9]/sample_n rowoff_n[9] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[9|31] vcm ctop col[31] col_n[31] row_n[10] rowon_n[10] adc_array_wafflecap_8_0[9|9]/sample
+ adc_array_wafflecap_8_0[9|9]/sample_n rowoff_n[10] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[10|31] vcm ctop col[31] col_n[31] row_n[11] rowon_n[11] adc_array_wafflecap_8_0[10|9]/sample
+ adc_array_wafflecap_8_0[10|9]/sample_n rowoff_n[11] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[11|31] vcm ctop col[31] col_n[31] row_n[12] rowon_n[12] adc_array_wafflecap_8_0[11|9]/sample
+ adc_array_wafflecap_8_0[11|9]/sample_n rowoff_n[12] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[12|31] vcm ctop col[31] col_n[31] row_n[13] rowon_n[13] adc_array_wafflecap_8_0[12|9]/sample
+ adc_array_wafflecap_8_0[12|9]/sample_n rowoff_n[13] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[13|31] vcm ctop col[31] col_n[31] row_n[14] rowon_n[14] adc_array_wafflecap_8_0[13|9]/sample
+ adc_array_wafflecap_8_0[13|9]/sample_n rowoff_n[14] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_0[14|31] vcm ctop col[31] col_n[31] row_n[15] rowon_n[15] adc_array_wafflecap_8_0[14|9]/sample
+ adc_array_wafflecap_8_0[14|9]/sample_n rowoff_n[15] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[0] vcm ctop col[1] col_n[1] row_n[0] rowon_n[0] adc_array_wafflecap_8_1[9]/sample
+ adc_array_wafflecap_8_1[9]/sample_n rowoff_n[0] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[1] vcm ctop col[2] col_n[2] row_n[0] rowon_n[0] adc_array_wafflecap_8_1[9]/sample
+ adc_array_wafflecap_8_1[9]/sample_n rowoff_n[0] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[2] vcm ctop col[3] col_n[3] row_n[0] rowon_n[0] adc_array_wafflecap_8_1[9]/sample
+ adc_array_wafflecap_8_1[9]/sample_n rowoff_n[0] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[3] vcm ctop col[4] col_n[4] row_n[0] rowon_n[0] adc_array_wafflecap_8_1[9]/sample
+ adc_array_wafflecap_8_1[9]/sample_n rowoff_n[0] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[4] vcm ctop col[5] col_n[5] row_n[0] rowon_n[0] adc_array_wafflecap_8_1[9]/sample
+ adc_array_wafflecap_8_1[9]/sample_n rowoff_n[0] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[5] vcm ctop col[6] col_n[6] row_n[0] rowon_n[0] adc_array_wafflecap_8_1[9]/sample
+ adc_array_wafflecap_8_1[9]/sample_n rowoff_n[0] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[6] vcm ctop col[7] col_n[7] row_n[0] rowon_n[0] adc_array_wafflecap_8_1[9]/sample
+ adc_array_wafflecap_8_1[9]/sample_n rowoff_n[0] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[7] vcm ctop col[8] col_n[8] row_n[0] rowon_n[0] adc_array_wafflecap_8_1[9]/sample
+ adc_array_wafflecap_8_1[9]/sample_n rowoff_n[0] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[8] vcm ctop col[9] col_n[9] row_n[0] rowon_n[0] adc_array_wafflecap_8_1[9]/sample
+ adc_array_wafflecap_8_1[9]/sample_n rowoff_n[0] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[9] vcm ctop col[10] col_n[10] row_n[0] rowon_n[0] adc_array_wafflecap_8_1[9]/sample
+ adc_array_wafflecap_8_1[9]/sample_n rowoff_n[0] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[10] vcm ctop col[11] col_n[11] row_n[0] rowon_n[0] adc_array_wafflecap_8_1[9]/sample
+ adc_array_wafflecap_8_1[9]/sample_n rowoff_n[0] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[11] vcm ctop col[12] col_n[12] row_n[0] rowon_n[0] adc_array_wafflecap_8_1[9]/sample
+ adc_array_wafflecap_8_1[9]/sample_n rowoff_n[0] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[12] vcm ctop col[13] col_n[13] row_n[0] rowon_n[0] adc_array_wafflecap_8_1[9]/sample
+ adc_array_wafflecap_8_1[9]/sample_n rowoff_n[0] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[13] vcm ctop col[14] col_n[14] row_n[0] rowon_n[0] adc_array_wafflecap_8_1[9]/sample
+ adc_array_wafflecap_8_1[9]/sample_n rowoff_n[0] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[14] vcm ctop col[15] col_n[15] row_n[0] rowon_n[0] adc_array_wafflecap_8_1[9]/sample
+ adc_array_wafflecap_8_1[9]/sample_n rowoff_n[0] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[15] vcm ctop col[16] col_n[16] row_n[0] rowon_n[0] adc_array_wafflecap_8_1[9]/sample
+ adc_array_wafflecap_8_1[9]/sample_n rowoff_n[0] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[16] vcm ctop col[17] col_n[17] row_n[0] rowon_n[0] adc_array_wafflecap_8_1[9]/sample
+ adc_array_wafflecap_8_1[9]/sample_n rowoff_n[0] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[17] vcm ctop col[18] col_n[18] row_n[0] rowon_n[0] adc_array_wafflecap_8_1[9]/sample
+ adc_array_wafflecap_8_1[9]/sample_n rowoff_n[0] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[18] vcm ctop col[19] col_n[19] row_n[0] rowon_n[0] adc_array_wafflecap_8_1[9]/sample
+ adc_array_wafflecap_8_1[9]/sample_n rowoff_n[0] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[19] vcm ctop col[20] col_n[20] row_n[0] rowon_n[0] adc_array_wafflecap_8_1[9]/sample
+ adc_array_wafflecap_8_1[9]/sample_n rowoff_n[0] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[20] vcm ctop col[21] col_n[21] row_n[0] rowon_n[0] adc_array_wafflecap_8_1[9]/sample
+ adc_array_wafflecap_8_1[9]/sample_n rowoff_n[0] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[21] vcm ctop col[22] col_n[22] row_n[0] rowon_n[0] adc_array_wafflecap_8_1[9]/sample
+ adc_array_wafflecap_8_1[9]/sample_n rowoff_n[0] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[22] vcm ctop col[23] col_n[23] row_n[0] rowon_n[0] adc_array_wafflecap_8_1[9]/sample
+ adc_array_wafflecap_8_1[9]/sample_n rowoff_n[0] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[23] vcm ctop col[24] col_n[24] row_n[0] rowon_n[0] adc_array_wafflecap_8_1[9]/sample
+ adc_array_wafflecap_8_1[9]/sample_n rowoff_n[0] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[24] vcm ctop col[25] col_n[25] row_n[0] rowon_n[0] adc_array_wafflecap_8_1[9]/sample
+ adc_array_wafflecap_8_1[9]/sample_n rowoff_n[0] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[25] vcm ctop col[26] col_n[26] row_n[0] rowon_n[0] adc_array_wafflecap_8_1[9]/sample
+ adc_array_wafflecap_8_1[9]/sample_n rowoff_n[0] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[26] vcm ctop col[27] col_n[27] row_n[0] rowon_n[0] adc_array_wafflecap_8_1[9]/sample
+ adc_array_wafflecap_8_1[9]/sample_n rowoff_n[0] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[27] vcm ctop col[28] col_n[28] row_n[0] rowon_n[0] adc_array_wafflecap_8_1[9]/sample
+ adc_array_wafflecap_8_1[9]/sample_n rowoff_n[0] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[28] vcm ctop col[29] col_n[29] row_n[0] rowon_n[0] adc_array_wafflecap_8_1[9]/sample
+ adc_array_wafflecap_8_1[9]/sample_n rowoff_n[0] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[29] vcm ctop col[30] col_n[30] row_n[0] rowon_n[0] adc_array_wafflecap_8_1[9]/sample
+ adc_array_wafflecap_8_1[9]/sample_n rowoff_n[0] VDD VSS adc_array_wafflecap_8
Xadc_array_wafflecap_8_1[30] vcm ctop col[31] col_n[31] row_n[0] rowon_n[0] adc_array_wafflecap_8_1[9]/sample
+ adc_array_wafflecap_8_1[9]/sample_n rowoff_n[0] VDD VSS adc_array_wafflecap_8
Xadc_noise_decoup_cell1_0[0] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[1] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[2] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[3] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[4] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_0[5] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[0] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[1] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[2] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[3] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[4] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[5] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[6] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[7] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_noise_decoup_cell1_1[8] VDD VSS VDD VSS VSS adc_noise_decoup_cell1
Xadc_array_wafflecap_4_0 vcm ctop col[16] col_n[16] VDD VSS adc_array_wafflecap_4_0/sample
+ adc_array_wafflecap_4_0/sample_n VDD en_bit_n[2] adc_array_wafflecap_4_0/cbot VDD
+ VSS adc_array_wafflecap_4
Xadc_array_wafflecap_2_0 vcm ctop col[15] col_n[15] VDD VSS adc_array_wafflecap_4_0/sample
+ adc_array_wafflecap_4_0/sample_n VDD en_bit_n[1] adc_array_wafflecap_2_0/cbot VDD
+ VSS adc_array_wafflecap_2
Xadc_array_wafflecap_dummy_0 vcm adc_array_wafflecap_dummy_0/ctop col[0] col_n[0]
+ VDD VSS adc_array_wafflecap_4_0/sample adc_array_wafflecap_4_0/sample_n VDD adc_array_wafflecap_dummy_0/cbot
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_1[0] vcm adc_array_wafflecap_dummy_1[0]/ctop col[2] col_n[2]
+ VDD VSS adc_array_wafflecap_4_0/sample adc_array_wafflecap_4_0/sample_n VDD adc_array_wafflecap_dummy_1[0]/cbot
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_1[1] vcm adc_array_wafflecap_dummy_1[1]/ctop col[3] col_n[3]
+ VDD VSS adc_array_wafflecap_4_0/sample adc_array_wafflecap_4_0/sample_n VDD adc_array_wafflecap_dummy_1[1]/cbot
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_1[2] vcm adc_array_wafflecap_dummy_1[2]/ctop col[4] col_n[4]
+ VDD VSS adc_array_wafflecap_4_0/sample adc_array_wafflecap_4_0/sample_n VDD adc_array_wafflecap_dummy_1[2]/cbot
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_1[3] vcm adc_array_wafflecap_dummy_1[3]/ctop col[5] col_n[5]
+ VDD VSS adc_array_wafflecap_4_0/sample adc_array_wafflecap_4_0/sample_n VDD adc_array_wafflecap_dummy_1[3]/cbot
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_1[4] vcm adc_array_wafflecap_dummy_1[4]/ctop col[6] col_n[6]
+ VDD VSS adc_array_wafflecap_4_0/sample adc_array_wafflecap_4_0/sample_n VDD adc_array_wafflecap_dummy_1[4]/cbot
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_1[5] vcm adc_array_wafflecap_dummy_1[5]/ctop col[7] col_n[7]
+ VDD VSS adc_array_wafflecap_4_0/sample adc_array_wafflecap_4_0/sample_n VDD adc_array_wafflecap_dummy_1[5]/cbot
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_1[6] vcm adc_array_wafflecap_dummy_1[6]/ctop col[8] col_n[8]
+ VDD VSS adc_array_wafflecap_4_0/sample adc_array_wafflecap_4_0/sample_n VDD adc_array_wafflecap_dummy_1[6]/cbot
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_1[7] vcm adc_array_wafflecap_dummy_1[7]/ctop col[9] col_n[9]
+ VDD VSS adc_array_wafflecap_4_0/sample adc_array_wafflecap_4_0/sample_n VDD adc_array_wafflecap_dummy_1[7]/cbot
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_1[8] vcm adc_array_wafflecap_dummy_1[8]/ctop col[10] col_n[10]
+ VDD VSS adc_array_wafflecap_4_0/sample adc_array_wafflecap_4_0/sample_n VDD adc_array_wafflecap_dummy_1[8]/cbot
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_1[9] vcm adc_array_wafflecap_dummy_1[9]/ctop col[11] col_n[11]
+ VDD VSS adc_array_wafflecap_4_0/sample adc_array_wafflecap_4_0/sample_n VDD adc_array_wafflecap_dummy_1[9]/cbot
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_1[10] vcm adc_array_wafflecap_dummy_1[10]/ctop col[12]
+ col_n[12] VDD VSS adc_array_wafflecap_4_0/sample adc_array_wafflecap_4_0/sample_n
+ VDD adc_array_wafflecap_dummy_1[10]/cbot VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_1[11] vcm adc_array_wafflecap_dummy_1[11]/ctop col[13]
+ col_n[13] VDD VSS adc_array_wafflecap_4_0/sample adc_array_wafflecap_4_0/sample_n
+ VDD adc_array_wafflecap_dummy_1[11]/cbot VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_1[12] vcm adc_array_wafflecap_dummy_1[12]/ctop col[14]
+ col_n[14] VDD VSS adc_array_wafflecap_4_0/sample adc_array_wafflecap_4_0/sample_n
+ VDD adc_array_wafflecap_dummy_1[12]/cbot VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_3[0] vcm adc_array_wafflecap_dummy_3[0]/ctop col[18] col_n[18]
+ VDD VSS adc_array_wafflecap_4_0/sample adc_array_wafflecap_4_0/sample_n VDD adc_array_wafflecap_dummy_3[0]/cbot
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_3[1] vcm adc_array_wafflecap_dummy_3[1]/ctop col[19] col_n[19]
+ VDD VSS adc_array_wafflecap_4_0/sample adc_array_wafflecap_4_0/sample_n VDD adc_array_wafflecap_dummy_3[1]/cbot
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_3[2] vcm adc_array_wafflecap_dummy_3[2]/ctop col[20] col_n[20]
+ VDD VSS adc_array_wafflecap_4_0/sample adc_array_wafflecap_4_0/sample_n VDD adc_array_wafflecap_dummy_3[2]/cbot
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_3[3] vcm adc_array_wafflecap_dummy_3[3]/ctop col[21] col_n[21]
+ VDD VSS adc_array_wafflecap_4_0/sample adc_array_wafflecap_4_0/sample_n VDD adc_array_wafflecap_dummy_3[3]/cbot
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_3[4] vcm adc_array_wafflecap_dummy_3[4]/ctop col[22] col_n[22]
+ VDD VSS adc_array_wafflecap_4_0/sample adc_array_wafflecap_4_0/sample_n VDD adc_array_wafflecap_dummy_3[4]/cbot
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_3[5] vcm adc_array_wafflecap_dummy_3[5]/ctop col[23] col_n[23]
+ VDD VSS adc_array_wafflecap_4_0/sample adc_array_wafflecap_4_0/sample_n VDD adc_array_wafflecap_dummy_3[5]/cbot
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_3[6] vcm adc_array_wafflecap_dummy_3[6]/ctop col[24] col_n[24]
+ VDD VSS adc_array_wafflecap_4_0/sample adc_array_wafflecap_4_0/sample_n VDD adc_array_wafflecap_dummy_3[6]/cbot
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_3[7] vcm adc_array_wafflecap_dummy_3[7]/ctop col[25] col_n[25]
+ VDD VSS adc_array_wafflecap_4_0/sample adc_array_wafflecap_4_0/sample_n VDD adc_array_wafflecap_dummy_3[7]/cbot
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_3[8] vcm adc_array_wafflecap_dummy_3[8]/ctop col[26] col_n[26]
+ VDD VSS adc_array_wafflecap_4_0/sample adc_array_wafflecap_4_0/sample_n VDD adc_array_wafflecap_dummy_3[8]/cbot
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_3[9] vcm adc_array_wafflecap_dummy_3[9]/ctop col[27] col_n[27]
+ VDD VSS adc_array_wafflecap_4_0/sample adc_array_wafflecap_4_0/sample_n VDD adc_array_wafflecap_dummy_3[9]/cbot
+ VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_3[10] vcm adc_array_wafflecap_dummy_3[10]/ctop col[28]
+ col_n[28] VDD VSS adc_array_wafflecap_4_0/sample adc_array_wafflecap_4_0/sample_n
+ VDD adc_array_wafflecap_dummy_3[10]/cbot VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_3[11] vcm adc_array_wafflecap_dummy_3[11]/ctop col[29]
+ col_n[29] VDD VSS adc_array_wafflecap_4_0/sample adc_array_wafflecap_4_0/sample_n
+ VDD adc_array_wafflecap_dummy_3[11]/cbot VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_3[12] vcm adc_array_wafflecap_dummy_3[12]/ctop col[30]
+ col_n[30] VDD VSS adc_array_wafflecap_4_0/sample adc_array_wafflecap_4_0/sample_n
+ VDD adc_array_wafflecap_dummy_3[12]/cbot VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[0] vcm adc_array_wafflecap_dummy_4[0]/ctop col[0] col_n[0]
+ VDD VDD adc_array_wafflecap_drv_2/sample_o adc_array_wafflecap_drv_2/sample_n_o
+ VSS adc_array_wafflecap_dummy_4[0]/cbot VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[1] vcm adc_array_wafflecap_dummy_4[1]/ctop col[1] col_n[1]
+ VDD VDD adc_array_wafflecap_drv_2/sample_o adc_array_wafflecap_drv_2/sample_n_o
+ VSS adc_array_wafflecap_dummy_4[1]/cbot VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[2] vcm adc_array_wafflecap_dummy_4[2]/ctop col[2] col_n[2]
+ VDD VDD adc_array_wafflecap_drv_2/sample_o adc_array_wafflecap_drv_2/sample_n_o
+ VSS adc_array_wafflecap_dummy_4[2]/cbot VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[3] vcm adc_array_wafflecap_dummy_4[3]/ctop col[3] col_n[3]
+ VDD VDD adc_array_wafflecap_drv_2/sample_o adc_array_wafflecap_drv_2/sample_n_o
+ VSS adc_array_wafflecap_dummy_4[3]/cbot VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[4] vcm adc_array_wafflecap_dummy_4[4]/ctop col[4] col_n[4]
+ VDD VDD adc_array_wafflecap_drv_2/sample_o adc_array_wafflecap_drv_2/sample_n_o
+ VSS adc_array_wafflecap_dummy_4[4]/cbot VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[5] vcm adc_array_wafflecap_dummy_4[5]/ctop col[5] col_n[5]
+ VDD VDD adc_array_wafflecap_drv_2/sample_o adc_array_wafflecap_drv_2/sample_n_o
+ VSS adc_array_wafflecap_dummy_4[5]/cbot VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[6] vcm adc_array_wafflecap_dummy_4[6]/ctop col[6] col_n[6]
+ VDD VDD adc_array_wafflecap_drv_2/sample_o adc_array_wafflecap_drv_2/sample_n_o
+ VSS adc_array_wafflecap_dummy_4[6]/cbot VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[7] vcm adc_array_wafflecap_dummy_4[7]/ctop col[7] col_n[7]
+ VDD VDD adc_array_wafflecap_drv_2/sample_o adc_array_wafflecap_drv_2/sample_n_o
+ VSS adc_array_wafflecap_dummy_4[7]/cbot VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[8] vcm adc_array_wafflecap_dummy_4[8]/ctop col[8] col_n[8]
+ VDD VDD adc_array_wafflecap_drv_2/sample_o adc_array_wafflecap_drv_2/sample_n_o
+ VSS adc_array_wafflecap_dummy_4[8]/cbot VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[9] vcm adc_array_wafflecap_dummy_4[9]/ctop col[9] col_n[9]
+ VDD VDD adc_array_wafflecap_drv_2/sample_o adc_array_wafflecap_drv_2/sample_n_o
+ VSS adc_array_wafflecap_dummy_4[9]/cbot VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[10] vcm adc_array_wafflecap_dummy_4[10]/ctop col[10]
+ col_n[10] VDD VDD adc_array_wafflecap_drv_2/sample_o adc_array_wafflecap_drv_2/sample_n_o
+ VSS adc_array_wafflecap_dummy_4[10]/cbot VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[11] vcm adc_array_wafflecap_dummy_4[11]/ctop col[11]
+ col_n[11] VDD VDD adc_array_wafflecap_drv_2/sample_o adc_array_wafflecap_drv_2/sample_n_o
+ VSS adc_array_wafflecap_dummy_4[11]/cbot VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[12] vcm adc_array_wafflecap_dummy_4[12]/ctop col[12]
+ col_n[12] VDD VDD adc_array_wafflecap_drv_2/sample_o adc_array_wafflecap_drv_2/sample_n_o
+ VSS adc_array_wafflecap_dummy_4[12]/cbot VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[13] vcm adc_array_wafflecap_dummy_4[13]/ctop col[13]
+ col_n[13] VDD VDD adc_array_wafflecap_drv_2/sample_o adc_array_wafflecap_drv_2/sample_n_o
+ VSS adc_array_wafflecap_dummy_4[13]/cbot VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[14] vcm adc_array_wafflecap_dummy_4[14]/ctop col[14]
+ col_n[14] VDD VDD adc_array_wafflecap_drv_2/sample_o adc_array_wafflecap_drv_2/sample_n_o
+ VSS adc_array_wafflecap_dummy_4[14]/cbot VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[15] vcm adc_array_wafflecap_dummy_4[15]/ctop col[15]
+ col_n[15] VDD VDD adc_array_wafflecap_drv_2/sample_o adc_array_wafflecap_drv_2/sample_n_o
+ VSS adc_array_wafflecap_dummy_4[15]/cbot VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[16] vcm adc_array_wafflecap_dummy_4[16]/ctop col[16]
+ col_n[16] VDD VDD adc_array_wafflecap_drv_2/sample_o adc_array_wafflecap_drv_2/sample_n_o
+ VSS adc_array_wafflecap_dummy_4[16]/cbot VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[17] vcm adc_array_wafflecap_dummy_4[17]/ctop col[17]
+ col_n[17] VDD VDD adc_array_wafflecap_drv_2/sample_o adc_array_wafflecap_drv_2/sample_n_o
+ VSS adc_array_wafflecap_dummy_4[17]/cbot VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[18] vcm adc_array_wafflecap_dummy_4[18]/ctop col[18]
+ col_n[18] VDD VDD adc_array_wafflecap_drv_2/sample_o adc_array_wafflecap_drv_2/sample_n_o
+ VSS adc_array_wafflecap_dummy_4[18]/cbot VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[19] vcm adc_array_wafflecap_dummy_4[19]/ctop col[19]
+ col_n[19] VDD VDD adc_array_wafflecap_drv_2/sample_o adc_array_wafflecap_drv_2/sample_n_o
+ VSS adc_array_wafflecap_dummy_4[19]/cbot VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[20] vcm adc_array_wafflecap_dummy_4[20]/ctop col[20]
+ col_n[20] VDD VDD adc_array_wafflecap_drv_2/sample_o adc_array_wafflecap_drv_2/sample_n_o
+ VSS adc_array_wafflecap_dummy_4[20]/cbot VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[21] vcm adc_array_wafflecap_dummy_4[21]/ctop col[21]
+ col_n[21] VDD VDD adc_array_wafflecap_drv_2/sample_o adc_array_wafflecap_drv_2/sample_n_o
+ VSS adc_array_wafflecap_dummy_4[21]/cbot VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[22] vcm adc_array_wafflecap_dummy_4[22]/ctop col[22]
+ col_n[22] VDD VDD adc_array_wafflecap_drv_2/sample_o adc_array_wafflecap_drv_2/sample_n_o
+ VSS adc_array_wafflecap_dummy_4[22]/cbot VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[23] vcm adc_array_wafflecap_dummy_4[23]/ctop col[23]
+ col_n[23] VDD VDD adc_array_wafflecap_drv_2/sample_o adc_array_wafflecap_drv_2/sample_n_o
+ VSS adc_array_wafflecap_dummy_4[23]/cbot VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[24] vcm adc_array_wafflecap_dummy_4[24]/ctop col[24]
+ col_n[24] VDD VDD adc_array_wafflecap_drv_2/sample_o adc_array_wafflecap_drv_2/sample_n_o
+ VSS adc_array_wafflecap_dummy_4[24]/cbot VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[25] vcm adc_array_wafflecap_dummy_4[25]/ctop col[25]
+ col_n[25] VDD VDD adc_array_wafflecap_drv_2/sample_o adc_array_wafflecap_drv_2/sample_n_o
+ VSS adc_array_wafflecap_dummy_4[25]/cbot VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[26] vcm adc_array_wafflecap_dummy_4[26]/ctop col[26]
+ col_n[26] VDD VDD adc_array_wafflecap_drv_2/sample_o adc_array_wafflecap_drv_2/sample_n_o
+ VSS adc_array_wafflecap_dummy_4[26]/cbot VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[27] vcm adc_array_wafflecap_dummy_4[27]/ctop col[27]
+ col_n[27] VDD VDD adc_array_wafflecap_drv_2/sample_o adc_array_wafflecap_drv_2/sample_n_o
+ VSS adc_array_wafflecap_dummy_4[27]/cbot VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[28] vcm adc_array_wafflecap_dummy_4[28]/ctop col[28]
+ col_n[28] VDD VDD adc_array_wafflecap_drv_2/sample_o adc_array_wafflecap_drv_2/sample_n_o
+ VSS adc_array_wafflecap_dummy_4[28]/cbot VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[29] vcm adc_array_wafflecap_dummy_4[29]/ctop col[29]
+ col_n[29] VDD VDD adc_array_wafflecap_drv_2/sample_o adc_array_wafflecap_drv_2/sample_n_o
+ VSS adc_array_wafflecap_dummy_4[29]/cbot VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[30] vcm adc_array_wafflecap_dummy_4[30]/ctop col[30]
+ col_n[30] VDD VDD adc_array_wafflecap_drv_2/sample_o adc_array_wafflecap_drv_2/sample_n_o
+ VSS adc_array_wafflecap_dummy_4[30]/cbot VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[31] vcm adc_array_wafflecap_dummy_4[31]/ctop col[31]
+ col_n[31] VDD VDD adc_array_wafflecap_drv_2/sample_o adc_array_wafflecap_drv_2/sample_n_o
+ VSS adc_array_wafflecap_dummy_4[31]/cbot VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_dummy_4[32] vcm adc_array_wafflecap_dummy_4[32]/ctop VSS VDD
+ VDD VDD adc_array_wafflecap_drv_2/sample_o adc_array_wafflecap_drv_2/sample_n_o
+ VSS adc_array_wafflecap_dummy_4[32]/cbot VDD VSS adc_array_wafflecap_dummy
Xadc_array_wafflecap_gate_0 adc_array_wafflecap_4_0/sample_n VSS VDD vcm col_n[31]
+ analog_in sw sw_n adc_array_wafflecap_gate_0/m2_32_32# VDD adc_array_wafflecap_4_0/sample
+ col_n[31] ctop VDD VSS col[31] adc_array_wafflecap_gate
.ends

