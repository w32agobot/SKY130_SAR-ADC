magic
tech sky130A
timestamp 1666978453
<< metal1 >>
rect 0 0 1000 3000
<< properties >>
string FIXED_BBOX 0 0 1000 3000
string LEFclass BLOCK
string LEForigin 0 0
string LEFsource USER
<< end >>
