magic
tech sky130A
timestamp 1662997094
<< metal2 >>
rect 16 16 198 486
rect 304 16 486 486
<< metal4 >>
rect 236 0 266 467
<< comment >>
rect 0 486 16 502
rect 486 486 502 502
rect 0 0 16 16
rect 486 0 502 16
<< end >>
