magic
tech sky130A
timestamp 1665394094
<< nwell >>
rect 2065 1600 2124 1804
rect 446 1361 628 1406
rect 423 1349 628 1361
rect 423 1220 451 1349
rect 506 1294 628 1349
rect 500 1275 628 1294
rect 506 1220 628 1275
rect 423 1207 628 1220
rect 2064 1028 2204 1230
<< poly >>
rect 2119 1556 2135 1570
rect 2119 1474 2134 1556
rect 2119 1465 2156 1474
rect 2119 1448 2134 1465
rect 2151 1448 2156 1465
rect 2119 1440 2156 1448
rect 1318 1062 1357 1067
rect 1318 1045 1326 1062
rect 1343 1045 1357 1062
rect 1318 1040 1357 1045
<< polycont >>
rect 2134 1448 2151 1465
rect 418 1187 435 1204
rect 1326 1045 1343 1062
<< locali >>
rect 570 1740 678 1743
rect 570 1722 576 1740
rect 593 1722 615 1740
rect 632 1722 651 1740
rect 668 1722 678 1740
rect 570 1719 678 1722
rect 570 1406 613 1719
rect 2550 1570 2617 1573
rect 2550 1552 2556 1570
rect 2574 1552 2593 1570
rect 2611 1552 2617 1570
rect 2550 1549 2617 1552
rect 454 1386 613 1406
rect 2130 1465 2154 1473
rect 2130 1448 2134 1465
rect 2151 1448 2154 1465
rect 2183 1448 2733 1474
rect 523 1294 545 1386
rect 523 1275 569 1294
rect 2130 1282 2154 1448
rect 2130 1264 2133 1282
rect 2151 1264 2154 1282
rect 410 1204 437 1212
rect 410 1187 418 1204
rect 435 1187 437 1204
rect 410 1179 437 1187
rect 527 1204 554 1212
rect 527 1187 535 1204
rect 552 1187 554 1204
rect 527 1179 554 1187
rect 2130 1106 2154 1264
rect 2171 1420 2195 1426
rect 2171 1402 2174 1420
rect 2192 1402 2195 1420
rect 2171 1252 2195 1402
rect 2264 1365 2307 1448
rect 2437 1275 2537 1278
rect 2437 1259 2475 1275
rect 2469 1257 2475 1259
rect 2493 1257 2513 1275
rect 2531 1257 2537 1275
rect 2469 1254 2537 1257
rect 2171 1234 2174 1252
rect 2192 1234 2195 1252
rect 2171 1228 2195 1234
rect 2130 1080 2259 1106
rect 1318 1062 1357 1067
rect 1318 1045 1326 1062
rect 1343 1045 1357 1062
rect 2081 1046 2249 1063
rect 1318 1040 1357 1045
<< viali >>
rect 576 1722 593 1740
rect 615 1722 632 1740
rect 651 1722 668 1740
rect 2556 1552 2574 1570
rect 2593 1552 2611 1570
rect 2133 1264 2151 1282
rect 418 1187 435 1204
rect 535 1187 552 1204
rect 2174 1402 2192 1420
rect 2475 1257 2493 1275
rect 2513 1257 2531 1275
rect 2174 1234 2192 1252
rect 1326 1045 1343 1062
rect 1365 1045 1382 1062
<< metal1 >>
rect 0 1770 14 1885
rect 570 1740 678 1770
rect 570 1722 576 1740
rect 593 1722 615 1740
rect 632 1722 651 1740
rect 668 1722 678 1740
rect 570 1719 678 1722
rect 2060 1738 2121 1755
rect 0 1541 7 1555
rect 0 1513 7 1527
rect 2060 1426 2078 1738
rect 2607 1588 3005 1602
rect 2550 1570 2617 1573
rect 2550 1552 2556 1570
rect 2574 1552 2593 1570
rect 2611 1568 2617 1570
rect 2611 1554 3005 1568
rect 2611 1552 2617 1554
rect 2550 1549 2617 1552
rect 2060 1420 2195 1426
rect 2060 1407 2174 1420
rect 2171 1402 2174 1407
rect 2192 1402 2195 1420
rect 2171 1396 2195 1402
rect 2130 1282 2154 1288
rect 2130 1277 2133 1282
rect 2032 1264 2133 1277
rect 2151 1264 2154 1282
rect 2032 1258 2154 1264
rect 2469 1275 2537 1278
rect 2171 1252 2195 1258
rect 2469 1257 2475 1275
rect 2493 1257 2513 1275
rect 2531 1273 2537 1275
rect 2531 1259 2664 1273
rect 2531 1257 2537 1259
rect 2469 1254 2537 1257
rect 2171 1234 2174 1252
rect 2192 1245 2195 1252
rect 2192 1234 2220 1245
rect 2171 1226 2220 1234
rect 407 1204 438 1212
rect 407 1203 418 1204
rect 336 1189 418 1203
rect 407 1187 418 1189
rect 435 1187 438 1204
rect 407 1179 438 1187
rect 527 1204 555 1212
rect 527 1187 535 1204
rect 552 1195 555 1204
rect 552 1187 657 1195
rect 527 1179 657 1187
rect 0 910 11 1026
rect 393 1025 621 1078
rect 636 1067 657 1179
rect 636 1062 1390 1067
rect 636 1045 1326 1062
rect 1343 1045 1365 1062
rect 1382 1045 1390 1062
rect 636 1040 1390 1045
use adc_comp_circuit  adc_comp_circuit_0
timestamp 1665394094
transform 1 0 637 0 1 1689
box -637 -1689 2355 1109
use adc_inverter  adc_inverter_0
timestamp 1664803391
transform 1 0 423 0 1 1118
box -13 -65 104 291
use adc_inverter  adc_inverter_1
timestamp 1664803391
transform 1 0 540 0 1 1118
box -13 -65 104 291
use adc_nor  adc_nor_0
timestamp 1661513809
transform 1 0 2208 0 -1 1258
box -4 -118 253 230
use adc_nor_latch  adc_nor_latch_0
timestamp 1661515501
transform 1 0 2124 0 1 1456
box -3 0 505 348
<< labels >>
flabel metal1 s 0 1513 7 1527 7 FreeSans 80 0 0 0 inn
port 30 w analog input
flabel metal1 s 0 1541 7 1555 7 FreeSans 80 0 0 0 inp
port 31 w analog input
flabel metal1 s 0 1770 14 1885 7 FreeSans 80 0 0 0 VDD
port 27 w power bidirectional
flabel metal1 s 0 910 11 1026 7 FreeSans 80 0 0 0 VSS
port 26 w power bidirectional
flabel metal1 s 2924 1588 3005 1602 3 FreeSans 80 0 0 0 latch_q
port 21 e signal output
flabel metal1 s 2924 1554 3005 1568 3 FreeSans 80 0 0 0 latch_qn
port 22 e signal output
flabel metal1 s 2583 1259 2664 1273 3 FreeSans 80 0 0 0 comp_trig
port 23 e signal output
flabel metal1 s 336 1189 343 1203 7 FreeSans 80 0 0 0 clk
port 32 w signal input
<< properties >>
string LEFclass CORE
string LEForigin 0 0
string LEFsource USER
<< end >>
