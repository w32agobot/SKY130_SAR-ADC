* SPICE3 file created from adc_array_fingercap_8(2)x360aF_topB_22um2.ext - technology: sky130A

C0 VSS cbot 3.09fF
C1 VSS ctop 0.34fF
C2 VSS floatingmetal 0.69fF
C3 cbot ctop 0.72fF
C4 cbot floatingmetal 2.02fF
C5 floatingmetal ctop 0.28fF
C6 floatingmetal VSUBS 0.61fF
C7 ctop VSUBS 0.35fF
C8 cbot VSUBS 0.43fF
C9 VSS VSUBS 1.80fF
