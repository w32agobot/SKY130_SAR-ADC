magic
tech sky130A
magscale 1 2
timestamp 1661518684
<< metal3 >>
rect -2149 50 -10 1530
rect 72 50 2210 1530
rect -1206 -50 -1052 50
rect 1110 -50 1264 50
rect -2149 -1530 -10 -50
rect 72 -1530 2210 -50
<< mimcap >>
rect -2049 1390 -209 1430
rect -2049 190 -2009 1390
rect -249 190 -209 1390
rect -2049 150 -209 190
rect 270 1390 2110 1430
rect 270 190 310 1390
rect 2070 190 2110 1390
rect 270 150 2110 190
rect -2049 -190 -209 -150
rect -2049 -1390 -2009 -190
rect -249 -1390 -209 -190
rect -2049 -1430 -209 -1390
rect 270 -190 2110 -150
rect 270 -1390 310 -190
rect 2070 -1390 2110 -190
rect 270 -1430 2110 -1390
<< mimcapcontact >>
rect -2009 190 -249 1390
rect 310 190 2070 1390
rect -2009 -1390 -249 -190
rect 310 -1390 2070 -190
<< metal4 >>
rect -1181 1391 -1077 1580
rect 1138 1391 1242 1580
rect -2010 1390 -248 1391
rect -2010 190 -2009 1390
rect -249 190 -248 1390
rect -2010 189 -248 190
rect 309 1390 2071 1391
rect 309 190 310 1390
rect 2070 190 2071 1390
rect 309 189 2071 190
rect -1181 -189 -1077 189
rect 1138 -189 1242 189
rect -2010 -190 -248 -189
rect -2010 -1390 -2009 -190
rect -249 -1390 -248 -190
rect -2010 -1391 -248 -1390
rect 309 -190 2071 -189
rect 309 -1390 310 -190
rect 2070 -1390 2071 -190
rect 309 -1391 2071 -1390
rect -1181 -1580 -1077 -1391
rect 1138 -1534 1242 -1391
<< end >>
