magic
tech sky130A
timestamp 1663934390
<< psubdiff >>
rect 238 9567 445 9731
rect 238 9550 252 9567
rect 427 9550 445 9567
rect 238 9527 445 9550
rect 238 9510 252 9527
rect 427 9510 445 9527
rect 238 9487 445 9510
rect 238 9470 252 9487
rect 427 9470 445 9487
rect 238 9447 445 9470
rect 238 9430 252 9447
rect 427 9430 445 9447
rect 238 9407 445 9430
rect 238 9390 252 9407
rect 427 9390 445 9407
rect 238 9367 445 9390
rect 238 9350 252 9367
rect 427 9350 445 9367
rect 238 9327 445 9350
rect 238 9310 252 9327
rect 427 9310 445 9327
rect 238 9287 445 9310
rect 238 9270 252 9287
rect 427 9270 445 9287
rect 238 9247 445 9270
rect 238 9230 252 9247
rect 427 9230 445 9247
rect 238 9207 445 9230
rect 238 9190 252 9207
rect 427 9190 445 9207
rect 238 9167 445 9190
rect 238 9150 252 9167
rect 427 9150 445 9167
rect 238 9127 445 9150
rect 238 9110 252 9127
rect 427 9110 445 9127
rect 238 9087 445 9110
rect 238 9070 252 9087
rect 427 9070 445 9087
rect 238 9047 445 9070
rect 238 9030 252 9047
rect 427 9030 445 9047
rect 238 9007 445 9030
rect 238 8990 252 9007
rect 427 8990 445 9007
rect 238 8967 445 8990
rect 238 8950 252 8967
rect 427 8950 445 8967
rect 238 8927 445 8950
rect 238 8910 252 8927
rect 427 8910 445 8927
rect 238 8887 445 8910
rect 238 8870 252 8887
rect 427 8870 445 8887
rect 238 8847 445 8870
rect 238 8830 252 8847
rect 427 8830 445 8847
rect 238 8807 445 8830
rect 238 8790 252 8807
rect 427 8790 445 8807
rect 238 8767 445 8790
rect 238 8750 252 8767
rect 427 8750 445 8767
rect 238 8727 445 8750
rect 238 8710 252 8727
rect 427 8710 445 8727
rect 238 8687 445 8710
rect 238 8670 252 8687
rect 427 8670 445 8687
rect 238 8647 445 8670
rect 238 8630 252 8647
rect 427 8630 445 8647
rect 238 8607 445 8630
rect 238 8590 252 8607
rect 427 8590 445 8607
rect 238 8567 445 8590
rect 238 8550 252 8567
rect 427 8550 445 8567
rect 238 8527 445 8550
rect 238 8510 252 8527
rect 427 8510 445 8527
rect 238 8487 445 8510
rect 238 8470 252 8487
rect 427 8470 445 8487
rect 238 8447 445 8470
rect 238 8430 252 8447
rect 427 8430 445 8447
rect 238 8407 445 8430
rect 238 8390 252 8407
rect 427 8390 445 8407
rect 238 8367 445 8390
rect 238 8350 252 8367
rect 427 8350 445 8367
rect 238 8327 445 8350
rect 238 8310 252 8327
rect 427 8310 445 8327
rect 238 8287 445 8310
rect 238 8270 252 8287
rect 427 8270 445 8287
rect 238 8247 445 8270
rect 238 8230 252 8247
rect 427 8230 445 8247
rect 238 8207 445 8230
rect 238 8190 252 8207
rect 427 8190 445 8207
rect 238 8167 445 8190
rect 238 8150 252 8167
rect 427 8150 445 8167
rect 238 8127 445 8150
rect 238 8110 252 8127
rect 427 8110 445 8127
rect 238 8087 445 8110
rect 238 8070 252 8087
rect 427 8070 445 8087
rect 238 8047 445 8070
rect 238 8030 252 8047
rect 427 8030 445 8047
rect 238 8007 445 8030
rect 238 7990 252 8007
rect 427 7990 445 8007
rect 238 7967 445 7990
rect 238 7950 252 7967
rect 427 7950 445 7967
rect 238 7927 445 7950
rect 238 7910 252 7927
rect 427 7910 445 7927
rect 238 7887 445 7910
rect 238 7870 252 7887
rect 427 7870 445 7887
rect 238 7847 445 7870
rect 238 7830 252 7847
rect 427 7830 445 7847
rect 238 7807 445 7830
rect 238 7790 252 7807
rect 427 7790 445 7807
rect 238 7767 445 7790
rect 238 7750 252 7767
rect 427 7750 445 7767
rect 238 7727 445 7750
rect 238 7710 252 7727
rect 427 7710 445 7727
rect 238 7687 445 7710
rect 238 7670 252 7687
rect 427 7670 445 7687
rect 238 7647 445 7670
rect 238 7630 252 7647
rect 427 7630 445 7647
rect 238 7607 445 7630
rect 238 7590 252 7607
rect 427 7590 445 7607
rect 238 7567 445 7590
rect 238 7550 252 7567
rect 427 7550 445 7567
rect 238 7527 445 7550
rect 238 7510 252 7527
rect 427 7510 445 7527
rect 238 7487 445 7510
rect 238 7470 252 7487
rect 427 7470 445 7487
rect 238 7447 445 7470
rect 238 7430 252 7447
rect 427 7430 445 7447
rect 238 7407 445 7430
rect 238 7390 252 7407
rect 427 7390 445 7407
rect 238 7367 445 7390
rect 238 7350 252 7367
rect 427 7350 445 7367
rect 238 7327 445 7350
rect 238 7310 252 7327
rect 427 7310 445 7327
rect 238 7287 445 7310
rect 238 7270 252 7287
rect 427 7270 445 7287
rect 238 7247 445 7270
rect 238 7230 252 7247
rect 427 7230 445 7247
rect 238 7207 445 7230
rect 238 7190 252 7207
rect 427 7190 445 7207
rect 238 7167 445 7190
rect 238 7150 252 7167
rect 427 7150 445 7167
rect 238 7127 445 7150
rect 238 7110 252 7127
rect 427 7110 445 7127
rect 238 7087 445 7110
rect 238 7070 252 7087
rect 427 7070 445 7087
rect 238 7047 445 7070
rect 238 7030 252 7047
rect 427 7030 445 7047
rect 238 7007 445 7030
rect 238 6990 252 7007
rect 427 6990 445 7007
rect 238 6967 445 6990
rect 238 6950 252 6967
rect 427 6950 445 6967
rect 238 6927 445 6950
rect 238 6910 252 6927
rect 427 6910 445 6927
rect 238 6887 445 6910
rect 238 6870 252 6887
rect 427 6870 445 6887
rect 238 6847 445 6870
rect 238 6830 252 6847
rect 427 6830 445 6847
rect 238 6807 445 6830
rect 238 6790 252 6807
rect 427 6790 445 6807
rect 238 6767 445 6790
rect 238 6750 252 6767
rect 427 6750 445 6767
rect 238 6727 445 6750
rect 238 6710 252 6727
rect 427 6710 445 6727
rect 238 6687 445 6710
rect 238 6670 252 6687
rect 427 6670 445 6687
rect 238 6647 445 6670
rect 238 6630 252 6647
rect 427 6630 445 6647
rect 238 6607 445 6630
rect 238 6590 252 6607
rect 427 6590 445 6607
rect 238 6567 445 6590
rect 238 6550 252 6567
rect 427 6550 445 6567
rect 238 6527 445 6550
rect 238 6510 252 6527
rect 427 6510 445 6527
rect 238 6487 445 6510
rect 238 6470 252 6487
rect 427 6470 445 6487
rect 238 6447 445 6470
rect 238 6430 252 6447
rect 427 6430 445 6447
rect 238 6407 445 6430
rect 238 6390 252 6407
rect 427 6390 445 6407
rect 238 6367 445 6390
rect 238 6350 252 6367
rect 427 6350 445 6367
rect 238 6327 445 6350
rect 238 6310 252 6327
rect 427 6310 445 6327
rect 238 6287 445 6310
rect 238 6270 252 6287
rect 427 6270 445 6287
rect 238 6247 445 6270
rect 238 6230 252 6247
rect 427 6230 445 6247
rect 238 6207 445 6230
rect 238 6190 252 6207
rect 427 6190 445 6207
rect 238 6167 445 6190
rect 238 6150 252 6167
rect 427 6150 445 6167
rect 238 6127 445 6150
rect 238 6110 252 6127
rect 427 6110 445 6127
rect 238 6087 445 6110
rect 238 6070 252 6087
rect 427 6070 445 6087
rect 238 6047 445 6070
rect 238 6030 252 6047
rect 427 6030 445 6047
rect 238 6007 445 6030
rect 238 5990 252 6007
rect 427 5990 445 6007
rect 238 5967 445 5990
rect 238 5950 252 5967
rect 427 5950 445 5967
rect 238 5927 445 5950
rect 238 5910 252 5927
rect 427 5910 445 5927
rect 238 5887 445 5910
rect 238 5870 252 5887
rect 427 5870 445 5887
rect 238 5847 445 5870
rect 238 5830 252 5847
rect 427 5830 445 5847
rect 238 5807 445 5830
rect 238 5790 252 5807
rect 427 5790 445 5807
rect 238 5767 445 5790
rect 238 5750 252 5767
rect 427 5750 445 5767
rect 238 5727 445 5750
rect 238 5710 252 5727
rect 427 5710 445 5727
rect 238 5687 445 5710
rect 238 5670 252 5687
rect 427 5670 445 5687
rect 238 5647 445 5670
rect 238 5630 252 5647
rect 427 5630 445 5647
rect 238 5607 445 5630
rect 238 5590 252 5607
rect 427 5590 445 5607
rect 238 5567 445 5590
rect 238 5550 252 5567
rect 427 5550 445 5567
rect 238 5527 445 5550
rect 238 5510 252 5527
rect 427 5510 445 5527
rect 238 5487 445 5510
rect 238 5470 252 5487
rect 427 5470 445 5487
rect 238 5447 445 5470
rect 238 5430 252 5447
rect 427 5430 445 5447
rect 238 5407 445 5430
rect 238 5390 252 5407
rect 427 5390 445 5407
rect 238 5367 445 5390
rect 238 5350 252 5367
rect 427 5350 445 5367
rect 238 5327 445 5350
rect 238 5310 252 5327
rect 427 5310 445 5327
rect 238 5287 445 5310
rect 238 5270 252 5287
rect 427 5270 445 5287
rect 238 5247 445 5270
rect 238 5230 252 5247
rect 427 5230 445 5247
rect 238 5207 445 5230
rect 238 5190 252 5207
rect 427 5190 445 5207
rect 238 5167 445 5190
rect 238 5150 252 5167
rect 427 5150 445 5167
rect 238 5127 445 5150
rect 238 5110 252 5127
rect 427 5110 445 5127
rect 238 5087 445 5110
rect 238 5070 252 5087
rect 427 5070 445 5087
rect 238 5047 445 5070
rect 238 5030 252 5047
rect 427 5030 445 5047
rect 238 5007 445 5030
rect 238 4990 252 5007
rect 427 4990 445 5007
rect 238 4967 445 4990
rect 238 4950 252 4967
rect 427 4950 445 4967
rect 238 4927 445 4950
rect 238 4910 252 4927
rect 427 4910 445 4927
rect 238 4887 445 4910
rect 238 4870 252 4887
rect 427 4870 445 4887
rect 238 4847 445 4870
rect 238 4830 252 4847
rect 427 4830 445 4847
rect 238 4807 445 4830
rect 238 4790 252 4807
rect 427 4790 445 4807
rect 238 4767 445 4790
rect 238 4750 252 4767
rect 427 4750 445 4767
rect 238 4727 445 4750
rect 238 4710 252 4727
rect 427 4710 445 4727
rect 238 4687 445 4710
rect 238 4670 252 4687
rect 427 4670 445 4687
rect 238 4647 445 4670
rect 238 4630 252 4647
rect 427 4630 445 4647
rect 238 4607 445 4630
rect 238 4590 252 4607
rect 427 4590 445 4607
rect 238 4567 445 4590
rect 238 4550 252 4567
rect 427 4550 445 4567
rect 238 4527 445 4550
rect 238 4510 252 4527
rect 427 4510 445 4527
rect 238 4487 445 4510
rect 238 4470 252 4487
rect 427 4470 445 4487
rect 238 4447 445 4470
rect 238 4430 252 4447
rect 427 4430 445 4447
rect 238 4407 445 4430
rect 238 4390 252 4407
rect 427 4390 445 4407
rect 238 4367 445 4390
rect 238 4350 252 4367
rect 427 4350 445 4367
rect 238 4327 445 4350
rect 238 4310 252 4327
rect 427 4310 445 4327
rect 238 4287 445 4310
rect 238 4270 252 4287
rect 427 4270 445 4287
rect 238 4247 445 4270
rect 238 4230 252 4247
rect 427 4230 445 4247
rect 238 4207 445 4230
rect 238 4190 252 4207
rect 427 4190 445 4207
rect 238 4167 445 4190
rect 238 4150 252 4167
rect 427 4150 445 4167
rect 238 4127 445 4150
rect 238 4110 252 4127
rect 427 4110 445 4127
rect 238 4087 445 4110
rect 238 4070 252 4087
rect 427 4070 445 4087
rect 238 4047 445 4070
rect 238 4030 252 4047
rect 427 4030 445 4047
rect 238 4007 445 4030
rect 238 3990 252 4007
rect 427 3990 445 4007
rect 238 3967 445 3990
rect 238 3950 252 3967
rect 427 3950 445 3967
rect 238 3927 445 3950
rect 238 3910 252 3927
rect 427 3910 445 3927
rect 238 3887 445 3910
rect 238 3870 252 3887
rect 427 3870 445 3887
rect 238 3847 445 3870
rect 238 3830 252 3847
rect 427 3830 445 3847
rect 238 3807 445 3830
rect 238 3790 252 3807
rect 427 3790 445 3807
rect 238 3767 445 3790
rect 238 3750 252 3767
rect 427 3750 445 3767
rect 238 3727 445 3750
rect 238 3710 252 3727
rect 427 3710 445 3727
rect 238 3687 445 3710
rect 238 3670 252 3687
rect 427 3670 445 3687
rect 238 3647 445 3670
rect 238 3630 252 3647
rect 427 3630 445 3647
rect 238 3607 445 3630
rect 238 3590 252 3607
rect 427 3590 445 3607
rect 238 3567 445 3590
rect 238 3550 252 3567
rect 427 3550 445 3567
rect 238 3527 445 3550
rect 238 3510 252 3527
rect 427 3510 445 3527
rect 238 3487 445 3510
rect 238 3470 252 3487
rect 427 3470 445 3487
rect 238 3447 445 3470
rect 238 3430 252 3447
rect 427 3430 445 3447
rect 238 3407 445 3430
rect 238 3390 252 3407
rect 427 3390 445 3407
rect 238 3367 445 3390
rect 238 3350 252 3367
rect 427 3350 445 3367
rect 238 3327 445 3350
rect 238 3310 252 3327
rect 427 3310 445 3327
rect 238 3287 445 3310
rect 238 3270 252 3287
rect 427 3270 445 3287
rect 238 3247 445 3270
rect 238 3230 252 3247
rect 427 3230 445 3247
rect 238 3207 445 3230
rect 238 3190 252 3207
rect 427 3190 445 3207
rect 238 3167 445 3190
rect 238 3150 252 3167
rect 427 3150 445 3167
rect 238 3127 445 3150
rect 238 3110 252 3127
rect 427 3110 445 3127
rect 238 3087 445 3110
rect 238 3070 252 3087
rect 427 3070 445 3087
rect 238 3047 445 3070
rect 238 3030 252 3047
rect 427 3030 445 3047
rect 238 3007 445 3030
rect 238 2990 252 3007
rect 427 2990 445 3007
rect 238 2967 445 2990
rect 238 2950 252 2967
rect 427 2950 445 2967
rect 238 2927 445 2950
rect 238 2910 252 2927
rect 427 2910 445 2927
rect 238 2887 445 2910
rect 238 2870 252 2887
rect 427 2870 445 2887
rect 238 2847 445 2870
rect 238 2830 252 2847
rect 427 2830 445 2847
rect 238 2807 445 2830
rect 238 2790 252 2807
rect 427 2790 445 2807
rect 238 2767 445 2790
rect 238 2750 252 2767
rect 427 2750 445 2767
rect 238 2727 445 2750
rect 238 2710 252 2727
rect 427 2710 445 2727
rect 238 2687 445 2710
rect 238 2670 252 2687
rect 427 2670 445 2687
rect 238 2647 445 2670
rect 238 2630 252 2647
rect 427 2630 445 2647
rect 238 2607 445 2630
rect 238 2590 252 2607
rect 427 2590 445 2607
rect 238 2567 445 2590
rect 238 2550 252 2567
rect 427 2550 445 2567
rect 238 2527 445 2550
rect 238 2510 252 2527
rect 427 2510 445 2527
rect 238 2487 445 2510
rect 238 2470 252 2487
rect 427 2470 445 2487
rect 238 2447 445 2470
rect 238 2430 252 2447
rect 427 2430 445 2447
rect 238 2407 445 2430
rect 238 2390 252 2407
rect 427 2390 445 2407
rect 238 2367 445 2390
rect 238 2350 252 2367
rect 427 2350 445 2367
rect 238 2327 445 2350
rect 238 2310 252 2327
rect 427 2310 445 2327
rect 238 2287 445 2310
rect 238 2270 252 2287
rect 427 2270 445 2287
rect 238 2247 445 2270
rect 238 2230 252 2247
rect 427 2230 445 2247
rect 238 2207 445 2230
rect 238 2190 252 2207
rect 427 2190 445 2207
rect 238 2167 445 2190
rect 238 2150 252 2167
rect 427 2150 445 2167
rect 238 2127 445 2150
rect 238 2110 252 2127
rect 427 2110 445 2127
rect 238 2087 445 2110
rect 238 2070 252 2087
rect 427 2070 445 2087
rect 238 2047 445 2070
rect 238 2030 252 2047
rect 427 2030 445 2047
rect 238 2007 445 2030
rect 238 1990 252 2007
rect 427 1990 445 2007
rect 238 1967 445 1990
rect 238 1950 252 1967
rect 427 1950 445 1967
rect 238 1927 445 1950
rect 238 1910 252 1927
rect 427 1910 445 1927
rect 238 1887 445 1910
rect 238 1870 252 1887
rect 427 1870 445 1887
rect 238 1847 445 1870
rect 238 1830 252 1847
rect 427 1830 445 1847
rect 238 1807 445 1830
rect 238 1790 252 1807
rect 427 1790 445 1807
rect 238 1767 445 1790
rect 238 1750 252 1767
rect 427 1750 445 1767
rect 238 1727 445 1750
rect 238 1710 252 1727
rect 427 1710 445 1727
rect 238 1687 445 1710
rect 238 1670 252 1687
rect 427 1670 445 1687
rect 238 1647 445 1670
rect 238 1630 252 1647
rect 427 1630 445 1647
rect 238 1607 445 1630
rect 238 1590 252 1607
rect 427 1590 445 1607
rect 238 1567 445 1590
rect 238 1550 252 1567
rect 427 1550 445 1567
rect 238 1527 445 1550
rect 238 1510 252 1527
rect 427 1510 445 1527
rect 238 1487 445 1510
rect 238 1470 252 1487
rect 427 1470 445 1487
rect 238 1447 445 1470
rect 238 1430 252 1447
rect 427 1430 445 1447
rect 238 1407 445 1430
rect 238 1390 252 1407
rect 427 1390 445 1407
rect 238 1367 445 1390
rect 238 1350 252 1367
rect 427 1350 445 1367
rect 238 1327 445 1350
rect 238 1310 252 1327
rect 427 1310 445 1327
rect 238 1287 445 1310
rect 18827 9567 19034 9731
rect 18827 9550 18845 9567
rect 19020 9550 19034 9567
rect 18827 9527 19034 9550
rect 18827 9510 18845 9527
rect 19020 9510 19034 9527
rect 18827 9487 19034 9510
rect 18827 9470 18845 9487
rect 19020 9470 19034 9487
rect 18827 9447 19034 9470
rect 18827 9430 18845 9447
rect 19020 9430 19034 9447
rect 18827 9407 19034 9430
rect 18827 9390 18845 9407
rect 19020 9390 19034 9407
rect 18827 9367 19034 9390
rect 18827 9350 18845 9367
rect 19020 9350 19034 9367
rect 18827 9331 19034 9350
rect 18827 9327 19035 9331
rect 18827 9310 18845 9327
rect 19020 9310 19035 9327
rect 18827 9287 19035 9310
rect 18827 9270 18845 9287
rect 19020 9270 19035 9287
rect 18827 9247 19035 9270
rect 18827 9230 18845 9247
rect 19020 9230 19035 9247
rect 18827 9207 19035 9230
rect 18827 9190 18845 9207
rect 19020 9190 19035 9207
rect 18827 9167 19034 9190
rect 18827 9150 18845 9167
rect 19020 9150 19034 9167
rect 18827 9127 19034 9150
rect 18827 9110 18845 9127
rect 19020 9110 19034 9127
rect 18827 9087 19034 9110
rect 18827 9070 18845 9087
rect 19020 9070 19034 9087
rect 18827 9047 19034 9070
rect 18827 9030 18845 9047
rect 19020 9030 19034 9047
rect 18827 9007 19034 9030
rect 18827 8990 18845 9007
rect 19020 8990 19034 9007
rect 18827 8967 19034 8990
rect 18827 8950 18845 8967
rect 19020 8950 19034 8967
rect 18827 8927 19034 8950
rect 18827 8910 18845 8927
rect 19020 8910 19034 8927
rect 18827 8887 19034 8910
rect 18827 8870 18845 8887
rect 19020 8870 19034 8887
rect 18827 8847 19034 8870
rect 18827 8830 18845 8847
rect 19020 8830 19034 8847
rect 18827 8807 19034 8830
rect 18827 8790 18845 8807
rect 19020 8790 19034 8807
rect 18827 8767 19034 8790
rect 18827 8750 18845 8767
rect 19020 8750 19034 8767
rect 18827 8727 19034 8750
rect 18827 8710 18845 8727
rect 19020 8710 19034 8727
rect 18827 8687 19034 8710
rect 18827 8670 18845 8687
rect 19020 8670 19034 8687
rect 18827 8647 19034 8670
rect 18827 8630 18845 8647
rect 19020 8630 19034 8647
rect 18827 8607 19034 8630
rect 18827 8590 18845 8607
rect 19020 8590 19034 8607
rect 18827 8567 19034 8590
rect 18827 8550 18845 8567
rect 19020 8550 19034 8567
rect 18827 8527 19034 8550
rect 18827 8510 18845 8527
rect 19020 8510 19034 8527
rect 18827 8487 19034 8510
rect 18827 8470 18845 8487
rect 19020 8470 19034 8487
rect 18827 8447 19034 8470
rect 18827 8430 18845 8447
rect 19020 8430 19034 8447
rect 18827 8407 19034 8430
rect 18827 8390 18845 8407
rect 19020 8390 19034 8407
rect 18827 8367 19034 8390
rect 18827 8350 18845 8367
rect 19020 8350 19034 8367
rect 18827 8327 19034 8350
rect 18827 8310 18845 8327
rect 19020 8310 19034 8327
rect 18827 8287 19034 8310
rect 18827 8270 18845 8287
rect 19020 8270 19034 8287
rect 18827 8247 19034 8270
rect 18827 8230 18845 8247
rect 19020 8230 19034 8247
rect 18827 8207 19034 8230
rect 18827 8190 18845 8207
rect 19020 8190 19034 8207
rect 18827 8167 19034 8190
rect 18827 8150 18845 8167
rect 19020 8150 19034 8167
rect 18827 8127 19034 8150
rect 18827 8110 18845 8127
rect 19020 8110 19034 8127
rect 18827 8087 19034 8110
rect 18827 8070 18845 8087
rect 19020 8070 19034 8087
rect 18827 8047 19034 8070
rect 18827 8030 18845 8047
rect 19020 8030 19034 8047
rect 18827 8007 19034 8030
rect 18827 7990 18845 8007
rect 19020 7990 19034 8007
rect 18827 7967 19034 7990
rect 18827 7950 18845 7967
rect 19020 7950 19034 7967
rect 18827 7927 19034 7950
rect 18827 7910 18845 7927
rect 19020 7910 19034 7927
rect 18827 7887 19034 7910
rect 18827 7870 18845 7887
rect 19020 7870 19034 7887
rect 18827 7847 19034 7870
rect 18827 7830 18845 7847
rect 19020 7830 19034 7847
rect 18827 7807 19034 7830
rect 18827 7790 18845 7807
rect 19020 7790 19034 7807
rect 18827 7767 19034 7790
rect 18827 7750 18845 7767
rect 19020 7750 19034 7767
rect 18827 7727 19034 7750
rect 18827 7710 18845 7727
rect 19020 7710 19034 7727
rect 18827 7687 19034 7710
rect 18827 7670 18845 7687
rect 19020 7670 19034 7687
rect 18827 7647 19034 7670
rect 18827 7630 18845 7647
rect 19020 7630 19034 7647
rect 18827 7607 19034 7630
rect 18827 7590 18845 7607
rect 19020 7590 19034 7607
rect 18827 7567 19034 7590
rect 18827 7550 18845 7567
rect 19020 7550 19034 7567
rect 18827 7527 19034 7550
rect 18827 7510 18845 7527
rect 19020 7510 19034 7527
rect 18827 7487 19034 7510
rect 18827 7470 18845 7487
rect 19020 7470 19034 7487
rect 18827 7447 19034 7470
rect 18827 7430 18845 7447
rect 19020 7430 19034 7447
rect 18827 7407 19034 7430
rect 18827 7390 18845 7407
rect 19020 7390 19034 7407
rect 18827 7367 19034 7390
rect 18827 7350 18845 7367
rect 19020 7350 19034 7367
rect 18827 7327 19034 7350
rect 18827 7310 18845 7327
rect 19020 7310 19034 7327
rect 18827 7287 19034 7310
rect 18827 7270 18845 7287
rect 19020 7270 19034 7287
rect 18827 7247 19034 7270
rect 18827 7230 18845 7247
rect 19020 7230 19034 7247
rect 18827 7207 19034 7230
rect 18827 7190 18845 7207
rect 19020 7190 19034 7207
rect 18827 7167 19034 7190
rect 18827 7150 18845 7167
rect 19020 7150 19034 7167
rect 18827 7127 19034 7150
rect 18827 7110 18845 7127
rect 19020 7110 19034 7127
rect 18827 7087 19034 7110
rect 18827 7070 18845 7087
rect 19020 7070 19034 7087
rect 18827 7047 19034 7070
rect 18827 7030 18845 7047
rect 19020 7030 19034 7047
rect 18827 7007 19034 7030
rect 18827 6990 18845 7007
rect 19020 6990 19034 7007
rect 18827 6967 19034 6990
rect 18827 6950 18845 6967
rect 19020 6950 19034 6967
rect 18827 6927 19034 6950
rect 18827 6910 18845 6927
rect 19020 6910 19034 6927
rect 18827 6887 19034 6910
rect 18827 6870 18845 6887
rect 19020 6870 19034 6887
rect 18827 6847 19034 6870
rect 18827 6830 18845 6847
rect 19020 6830 19034 6847
rect 18827 6807 19034 6830
rect 18827 6790 18845 6807
rect 19020 6790 19034 6807
rect 18827 6767 19034 6790
rect 18827 6750 18845 6767
rect 19020 6750 19034 6767
rect 18827 6727 19034 6750
rect 18827 6710 18845 6727
rect 19020 6710 19034 6727
rect 18827 6686 19034 6710
rect 18827 6669 18846 6686
rect 19021 6669 19034 6686
rect 18827 6647 19034 6669
rect 18827 6630 18845 6647
rect 19020 6630 19034 6647
rect 18827 6607 19034 6630
rect 18827 6590 18845 6607
rect 19020 6590 19034 6607
rect 18827 6567 19034 6590
rect 18827 6550 18845 6567
rect 19020 6550 19034 6567
rect 18827 6527 19034 6550
rect 18827 6510 18845 6527
rect 19020 6510 19034 6527
rect 18827 6487 19034 6510
rect 18827 6470 18845 6487
rect 19020 6470 19034 6487
rect 18827 6447 19034 6470
rect 18827 6430 18845 6447
rect 19020 6430 19034 6447
rect 18827 6407 19034 6430
rect 18827 6390 18845 6407
rect 19020 6390 19034 6407
rect 18827 6367 19034 6390
rect 18827 6350 18845 6367
rect 19020 6361 19034 6367
rect 19020 6350 19035 6361
rect 18827 6327 19035 6350
rect 18827 6310 18845 6327
rect 19020 6310 19035 6327
rect 18827 6287 19035 6310
rect 18827 6270 18845 6287
rect 19020 6270 19035 6287
rect 18827 6247 19035 6270
rect 18827 6230 18845 6247
rect 19020 6230 19035 6247
rect 18827 6220 19035 6230
rect 18827 6207 19034 6220
rect 18827 6190 18845 6207
rect 19020 6190 19034 6207
rect 18827 6167 19034 6190
rect 18827 6150 18845 6167
rect 19020 6150 19034 6167
rect 18827 6127 19034 6150
rect 18827 6110 18845 6127
rect 19020 6110 19034 6127
rect 18827 6087 19034 6110
rect 18827 6070 18845 6087
rect 19020 6070 19034 6087
rect 18827 6047 19034 6070
rect 18827 6030 18845 6047
rect 19020 6030 19034 6047
rect 18827 6007 19034 6030
rect 18827 5990 18845 6007
rect 19020 5990 19034 6007
rect 18827 5967 19034 5990
rect 18827 5950 18845 5967
rect 19020 5950 19034 5967
rect 18827 5927 19034 5950
rect 18827 5910 18845 5927
rect 19020 5910 19034 5927
rect 18827 5887 19034 5910
rect 18827 5870 18845 5887
rect 19020 5870 19034 5887
rect 18827 5847 19034 5870
rect 18827 5830 18845 5847
rect 19020 5830 19034 5847
rect 18827 5806 19034 5830
rect 18827 5789 18844 5806
rect 19019 5789 19034 5806
rect 18827 5767 19034 5789
rect 18827 5750 18845 5767
rect 19020 5750 19034 5767
rect 18827 5727 19034 5750
rect 18827 5710 18845 5727
rect 19020 5710 19034 5727
rect 18827 5687 19034 5710
rect 18827 5670 18845 5687
rect 19020 5670 19034 5687
rect 18827 5647 19034 5670
rect 18827 5630 18845 5647
rect 19020 5630 19034 5647
rect 18827 5607 19034 5630
rect 18827 5590 18845 5607
rect 19020 5590 19034 5607
rect 18827 5567 19034 5590
rect 18827 5550 18845 5567
rect 19020 5550 19034 5567
rect 18827 5527 19034 5550
rect 18827 5510 18845 5527
rect 19020 5510 19034 5527
rect 18827 5487 19034 5510
rect 18827 5470 18845 5487
rect 19020 5470 19034 5487
rect 18827 5447 19034 5470
rect 18827 5430 18845 5447
rect 19020 5430 19034 5447
rect 18827 5407 19034 5430
rect 18827 5390 18845 5407
rect 19020 5390 19034 5407
rect 18827 5367 19034 5390
rect 18827 5350 18845 5367
rect 19020 5350 19034 5367
rect 18827 5327 19034 5350
rect 18827 5310 18845 5327
rect 19020 5310 19034 5327
rect 18827 5287 19034 5310
rect 18827 5270 18845 5287
rect 19020 5270 19034 5287
rect 18827 5247 19034 5270
rect 18827 5230 18845 5247
rect 19020 5230 19034 5247
rect 18827 5207 19034 5230
rect 18827 5190 18845 5207
rect 19020 5190 19034 5207
rect 18827 5167 19034 5190
rect 18827 5150 18845 5167
rect 19020 5150 19034 5167
rect 18827 5127 19034 5150
rect 18827 5110 18845 5127
rect 19020 5110 19034 5127
rect 18827 5087 19034 5110
rect 18827 5070 18845 5087
rect 19020 5070 19034 5087
rect 18827 5047 19034 5070
rect 18827 5030 18845 5047
rect 19020 5030 19034 5047
rect 18827 5007 19034 5030
rect 18827 4990 18845 5007
rect 19020 4990 19034 5007
rect 18827 4967 19034 4990
rect 18827 4950 18845 4967
rect 19020 4950 19034 4967
rect 18827 4927 19034 4950
rect 18827 4910 18845 4927
rect 19020 4910 19034 4927
rect 18827 4887 19034 4910
rect 18827 4870 18845 4887
rect 19020 4870 19034 4887
rect 18827 4847 19034 4870
rect 18827 4830 18845 4847
rect 19020 4830 19034 4847
rect 18827 4807 19034 4830
rect 18827 4790 18845 4807
rect 19020 4790 19034 4807
rect 18827 4767 19034 4790
rect 18827 4750 18845 4767
rect 19020 4750 19034 4767
rect 18827 4727 19034 4750
rect 18827 4710 18845 4727
rect 19020 4710 19034 4727
rect 18827 4687 19034 4710
rect 18827 4670 18845 4687
rect 19020 4670 19034 4687
rect 18827 4647 19034 4670
rect 18827 4630 18845 4647
rect 19020 4630 19034 4647
rect 18827 4607 19034 4630
rect 18827 4590 18845 4607
rect 19020 4590 19034 4607
rect 18827 4567 19034 4590
rect 18827 4550 18845 4567
rect 19020 4550 19034 4567
rect 18827 4527 19034 4550
rect 18827 4510 18845 4527
rect 19020 4510 19034 4527
rect 18827 4487 19034 4510
rect 18827 4470 18845 4487
rect 19020 4470 19034 4487
rect 18827 4447 19034 4470
rect 18827 4430 18845 4447
rect 19020 4430 19034 4447
rect 18827 4407 19034 4430
rect 18827 4390 18845 4407
rect 19020 4390 19034 4407
rect 18827 4367 19034 4390
rect 18827 4350 18845 4367
rect 19020 4350 19034 4367
rect 18827 4327 19034 4350
rect 18827 4310 18845 4327
rect 19020 4310 19034 4327
rect 18827 4287 19035 4310
rect 18827 4270 18845 4287
rect 19020 4270 19035 4287
rect 18827 4247 19035 4270
rect 18827 4230 18845 4247
rect 19020 4230 19035 4247
rect 18827 4207 19035 4230
rect 18827 4190 18845 4207
rect 19020 4190 19035 4207
rect 18827 4169 19035 4190
rect 18827 4167 19034 4169
rect 18827 4150 18845 4167
rect 19020 4150 19034 4167
rect 18827 4127 19034 4150
rect 18827 4110 18845 4127
rect 19020 4110 19034 4127
rect 18827 4087 19034 4110
rect 18827 4070 18845 4087
rect 19020 4070 19034 4087
rect 18827 4047 19034 4070
rect 18827 4030 18845 4047
rect 19020 4030 19034 4047
rect 18827 4007 19034 4030
rect 18827 3990 18845 4007
rect 19020 3990 19034 4007
rect 18827 3967 19034 3990
rect 18827 3950 18845 3967
rect 19020 3950 19034 3967
rect 18827 3927 19034 3950
rect 18827 3910 18845 3927
rect 19020 3910 19034 3927
rect 18827 3887 19034 3910
rect 18827 3870 18845 3887
rect 19020 3870 19034 3887
rect 18827 3847 19034 3870
rect 18827 3830 18845 3847
rect 19020 3830 19034 3847
rect 18827 3807 19034 3830
rect 18827 3790 18845 3807
rect 19020 3790 19034 3807
rect 18827 3767 19034 3790
rect 18827 3750 18845 3767
rect 19020 3750 19034 3767
rect 18827 3727 19034 3750
rect 18827 3710 18845 3727
rect 19020 3710 19034 3727
rect 18827 3687 19034 3710
rect 18827 3670 18845 3687
rect 19020 3670 19034 3687
rect 18827 3647 19034 3670
rect 18827 3630 18845 3647
rect 19020 3630 19034 3647
rect 18827 3607 19034 3630
rect 18827 3590 18845 3607
rect 19020 3590 19034 3607
rect 18827 3567 19034 3590
rect 18827 3550 18845 3567
rect 19020 3550 19034 3567
rect 18827 3527 19034 3550
rect 18827 3510 18845 3527
rect 19020 3510 19034 3527
rect 18827 3487 19034 3510
rect 18827 3470 18845 3487
rect 19020 3470 19034 3487
rect 18827 3447 19034 3470
rect 18827 3430 18845 3447
rect 19020 3430 19034 3447
rect 18827 3407 19034 3430
rect 18827 3390 18845 3407
rect 19020 3390 19034 3407
rect 18827 3367 19034 3390
rect 18827 3350 18845 3367
rect 19020 3350 19034 3367
rect 18827 3327 19034 3350
rect 18827 3310 18845 3327
rect 19020 3310 19034 3327
rect 18827 3288 19034 3310
rect 18827 3287 19035 3288
rect 18827 3270 18845 3287
rect 19020 3270 19035 3287
rect 18827 3247 19035 3270
rect 18827 3230 18845 3247
rect 19020 3230 19035 3247
rect 18827 3207 19035 3230
rect 18827 3190 18845 3207
rect 19020 3190 19035 3207
rect 18827 3167 19035 3190
rect 18827 3150 18845 3167
rect 19020 3150 19035 3167
rect 18827 3147 19035 3150
rect 18827 3127 19034 3147
rect 18827 3110 18845 3127
rect 19020 3110 19034 3127
rect 18827 3087 19034 3110
rect 18827 3070 18845 3087
rect 19020 3070 19034 3087
rect 18827 3047 19034 3070
rect 18827 3030 18845 3047
rect 19020 3030 19034 3047
rect 18827 3007 19034 3030
rect 18827 2990 18845 3007
rect 19020 2990 19034 3007
rect 18827 2967 19034 2990
rect 18827 2950 18845 2967
rect 19020 2950 19034 2967
rect 18827 2927 19034 2950
rect 18827 2910 18845 2927
rect 19020 2910 19034 2927
rect 18827 2887 19034 2910
rect 18827 2870 18845 2887
rect 19020 2870 19034 2887
rect 18827 2847 19034 2870
rect 18827 2830 18845 2847
rect 19020 2830 19034 2847
rect 18827 2807 19034 2830
rect 18827 2790 18845 2807
rect 19020 2790 19034 2807
rect 18827 2767 19034 2790
rect 18827 2750 18845 2767
rect 19020 2750 19034 2767
rect 18827 2724 19034 2750
rect 18827 2707 18845 2724
rect 19020 2707 19034 2724
rect 18827 2687 19034 2707
rect 18827 2670 18845 2687
rect 19020 2670 19034 2687
rect 18827 2647 19034 2670
rect 18827 2630 18845 2647
rect 19020 2630 19034 2647
rect 18827 2607 19034 2630
rect 18827 2590 18845 2607
rect 19020 2590 19034 2607
rect 18827 2567 19034 2590
rect 18827 2550 18845 2567
rect 19020 2550 19034 2567
rect 18827 2527 19034 2550
rect 18827 2510 18845 2527
rect 19020 2510 19034 2527
rect 18827 2487 19034 2510
rect 18827 2470 18845 2487
rect 19020 2470 19034 2487
rect 18827 2447 19034 2470
rect 18827 2430 18845 2447
rect 19020 2430 19034 2447
rect 18827 2407 19034 2430
rect 18827 2390 18845 2407
rect 19020 2390 19034 2407
rect 18827 2367 19034 2390
rect 18827 2350 18845 2367
rect 19020 2350 19034 2367
rect 18827 2327 19034 2350
rect 18827 2310 18845 2327
rect 19020 2310 19034 2327
rect 18827 2287 19034 2310
rect 18827 2270 18845 2287
rect 19020 2270 19034 2287
rect 18827 2247 19034 2270
rect 18827 2230 18845 2247
rect 19020 2230 19034 2247
rect 18827 2207 19034 2230
rect 18827 2190 18845 2207
rect 19020 2190 19034 2207
rect 18827 2167 19034 2190
rect 18827 2150 18845 2167
rect 19020 2150 19034 2167
rect 18827 2127 19034 2150
rect 18827 2110 18845 2127
rect 19020 2110 19034 2127
rect 18827 2087 19034 2110
rect 18827 2070 18845 2087
rect 19020 2070 19034 2087
rect 18827 2047 19034 2070
rect 18827 2030 18845 2047
rect 19020 2030 19034 2047
rect 18827 2007 19034 2030
rect 18827 1990 18845 2007
rect 19020 1990 19034 2007
rect 18827 1967 19034 1990
rect 18827 1950 18845 1967
rect 19020 1950 19034 1967
rect 18827 1927 19034 1950
rect 18827 1910 18845 1927
rect 19020 1910 19034 1927
rect 18827 1887 19034 1910
rect 18827 1870 18845 1887
rect 19020 1870 19034 1887
rect 18827 1847 19034 1870
rect 18827 1830 18845 1847
rect 19020 1830 19034 1847
rect 18827 1807 19034 1830
rect 18827 1790 18845 1807
rect 19020 1790 19034 1807
rect 18827 1767 19034 1790
rect 18827 1750 18845 1767
rect 19020 1750 19034 1767
rect 18827 1727 19034 1750
rect 18827 1710 18845 1727
rect 19020 1710 19034 1727
rect 18827 1687 19034 1710
rect 18827 1670 18845 1687
rect 19020 1670 19034 1687
rect 18827 1647 19034 1670
rect 18827 1630 18845 1647
rect 19020 1630 19034 1647
rect 18827 1607 19034 1630
rect 18827 1590 18845 1607
rect 19020 1590 19034 1607
rect 18827 1567 19034 1590
rect 18827 1550 18845 1567
rect 19020 1550 19034 1567
rect 18827 1527 19034 1550
rect 18827 1510 18845 1527
rect 19020 1510 19034 1527
rect 18827 1487 19034 1510
rect 18827 1470 18845 1487
rect 19020 1470 19034 1487
rect 18827 1447 19034 1470
rect 18827 1430 18845 1447
rect 19020 1430 19034 1447
rect 18827 1407 19034 1430
rect 18827 1390 18845 1407
rect 19020 1390 19034 1407
rect 18827 1367 19034 1390
rect 18827 1350 18845 1367
rect 19020 1350 19034 1367
rect 18827 1327 19034 1350
rect 18827 1310 18845 1327
rect 19020 1310 19034 1327
rect 18827 1291 19034 1310
rect 238 1270 252 1287
rect 427 1270 445 1287
rect 238 1247 445 1270
rect 238 1230 252 1247
rect 427 1230 445 1247
rect 238 1207 445 1230
rect 238 1190 252 1207
rect 427 1190 445 1207
rect 238 1167 445 1190
rect 238 1150 252 1167
rect 427 1150 445 1167
rect 18826 1287 19034 1291
rect 18826 1270 18845 1287
rect 19020 1270 19034 1287
rect 18826 1247 19034 1270
rect 18826 1230 18845 1247
rect 19020 1230 19034 1247
rect 18826 1207 19034 1230
rect 18826 1190 18845 1207
rect 19020 1190 19034 1207
rect 18826 1167 19034 1190
rect 18826 1150 18845 1167
rect 19020 1150 19034 1167
rect 238 1127 445 1150
rect 238 1110 252 1127
rect 427 1110 445 1127
rect 238 1087 445 1110
rect 238 1070 252 1087
rect 427 1070 445 1087
rect 238 1047 445 1070
rect 238 1030 252 1047
rect 427 1030 445 1047
rect 238 1007 445 1030
rect 238 990 252 1007
rect 427 990 445 1007
rect 238 967 445 990
rect 238 950 252 967
rect 427 950 445 967
rect 238 927 445 950
rect 238 910 252 927
rect 427 910 445 927
rect 238 887 445 910
rect 238 870 252 887
rect 427 870 445 887
rect 238 847 445 870
rect 238 830 252 847
rect 427 830 445 847
rect 238 807 445 830
rect 238 790 252 807
rect 427 790 445 807
rect 238 767 445 790
rect 238 750 252 767
rect 427 750 445 767
rect 238 727 445 750
rect 238 710 252 727
rect 427 710 445 727
rect 238 687 445 710
rect 238 670 252 687
rect 427 670 445 687
rect 238 647 445 670
rect 238 630 252 647
rect 427 630 445 647
rect 238 607 445 630
rect 238 590 252 607
rect 427 590 445 607
rect 238 567 445 590
rect 238 550 252 567
rect 427 550 445 567
rect 238 527 445 550
rect 238 510 252 527
rect 427 510 445 527
rect 238 487 445 510
rect 238 470 252 487
rect 427 470 445 487
rect 238 240 445 470
rect 18827 1127 19034 1150
rect 18827 1110 18845 1127
rect 19020 1110 19034 1127
rect 18827 1087 19034 1110
rect 18827 1070 18845 1087
rect 19020 1070 19034 1087
rect 18827 1047 19034 1070
rect 18827 1030 18845 1047
rect 19020 1030 19034 1047
rect 18827 1007 19034 1030
rect 18827 990 18845 1007
rect 19020 990 19034 1007
rect 18827 967 19034 990
rect 18827 950 18845 967
rect 19020 950 19034 967
rect 18827 927 19034 950
rect 18827 910 18845 927
rect 19020 910 19034 927
rect 18827 887 19034 910
rect 18827 870 18845 887
rect 19020 870 19034 887
rect 18827 847 19034 870
rect 18827 830 18845 847
rect 19020 830 19034 847
rect 18827 807 19034 830
rect 18827 790 18845 807
rect 19020 790 19034 807
rect 18827 767 19034 790
rect 18827 750 18845 767
rect 19020 750 19034 767
rect 18827 727 19034 750
rect 18827 710 18845 727
rect 19020 710 19034 727
rect 18827 687 19034 710
rect 18827 670 18845 687
rect 19020 670 19034 687
rect 18827 647 19034 670
rect 18827 630 18845 647
rect 19020 630 19034 647
rect 18827 607 19034 630
rect 18827 590 18845 607
rect 19020 590 19034 607
rect 18827 567 19034 590
rect 18827 550 18845 567
rect 19020 550 19034 567
rect 18827 527 19034 550
rect 18827 510 18845 527
rect 19020 510 19034 527
rect 18827 487 19034 510
rect 18827 470 18845 487
rect 19020 470 19034 487
rect 18827 305 19034 470
<< psubdiffcont >>
rect 252 9550 427 9567
rect 252 9510 427 9527
rect 252 9470 427 9487
rect 252 9430 427 9447
rect 252 9390 427 9407
rect 252 9350 427 9367
rect 252 9310 427 9327
rect 252 9270 427 9287
rect 252 9230 427 9247
rect 252 9190 427 9207
rect 252 9150 427 9167
rect 252 9110 427 9127
rect 252 9070 427 9087
rect 252 9030 427 9047
rect 252 8990 427 9007
rect 252 8950 427 8967
rect 252 8910 427 8927
rect 252 8870 427 8887
rect 252 8830 427 8847
rect 252 8790 427 8807
rect 252 8750 427 8767
rect 252 8710 427 8727
rect 252 8670 427 8687
rect 252 8630 427 8647
rect 252 8590 427 8607
rect 252 8550 427 8567
rect 252 8510 427 8527
rect 252 8470 427 8487
rect 252 8430 427 8447
rect 252 8390 427 8407
rect 252 8350 427 8367
rect 252 8310 427 8327
rect 252 8270 427 8287
rect 252 8230 427 8247
rect 252 8190 427 8207
rect 252 8150 427 8167
rect 252 8110 427 8127
rect 252 8070 427 8087
rect 252 8030 427 8047
rect 252 7990 427 8007
rect 252 7950 427 7967
rect 252 7910 427 7927
rect 252 7870 427 7887
rect 252 7830 427 7847
rect 252 7790 427 7807
rect 252 7750 427 7767
rect 252 7710 427 7727
rect 252 7670 427 7687
rect 252 7630 427 7647
rect 252 7590 427 7607
rect 252 7550 427 7567
rect 252 7510 427 7527
rect 252 7470 427 7487
rect 252 7430 427 7447
rect 252 7390 427 7407
rect 252 7350 427 7367
rect 252 7310 427 7327
rect 252 7270 427 7287
rect 252 7230 427 7247
rect 252 7190 427 7207
rect 252 7150 427 7167
rect 252 7110 427 7127
rect 252 7070 427 7087
rect 252 7030 427 7047
rect 252 6990 427 7007
rect 252 6950 427 6967
rect 252 6910 427 6927
rect 252 6870 427 6887
rect 252 6830 427 6847
rect 252 6790 427 6807
rect 252 6750 427 6767
rect 252 6710 427 6727
rect 252 6670 427 6687
rect 252 6630 427 6647
rect 252 6590 427 6607
rect 252 6550 427 6567
rect 252 6510 427 6527
rect 252 6470 427 6487
rect 252 6430 427 6447
rect 252 6390 427 6407
rect 252 6350 427 6367
rect 252 6310 427 6327
rect 252 6270 427 6287
rect 252 6230 427 6247
rect 252 6190 427 6207
rect 252 6150 427 6167
rect 252 6110 427 6127
rect 252 6070 427 6087
rect 252 6030 427 6047
rect 252 5990 427 6007
rect 252 5950 427 5967
rect 252 5910 427 5927
rect 252 5870 427 5887
rect 252 5830 427 5847
rect 252 5790 427 5807
rect 252 5750 427 5767
rect 252 5710 427 5727
rect 252 5670 427 5687
rect 252 5630 427 5647
rect 252 5590 427 5607
rect 252 5550 427 5567
rect 252 5510 427 5527
rect 252 5470 427 5487
rect 252 5430 427 5447
rect 252 5390 427 5407
rect 252 5350 427 5367
rect 252 5310 427 5327
rect 252 5270 427 5287
rect 252 5230 427 5247
rect 252 5190 427 5207
rect 252 5150 427 5167
rect 252 5110 427 5127
rect 252 5070 427 5087
rect 252 5030 427 5047
rect 252 4990 427 5007
rect 252 4950 427 4967
rect 252 4910 427 4927
rect 252 4870 427 4887
rect 252 4830 427 4847
rect 252 4790 427 4807
rect 252 4750 427 4767
rect 252 4710 427 4727
rect 252 4670 427 4687
rect 252 4630 427 4647
rect 252 4590 427 4607
rect 252 4550 427 4567
rect 252 4510 427 4527
rect 252 4470 427 4487
rect 252 4430 427 4447
rect 252 4390 427 4407
rect 252 4350 427 4367
rect 252 4310 427 4327
rect 252 4270 427 4287
rect 252 4230 427 4247
rect 252 4190 427 4207
rect 252 4150 427 4167
rect 252 4110 427 4127
rect 252 4070 427 4087
rect 252 4030 427 4047
rect 252 3990 427 4007
rect 252 3950 427 3967
rect 252 3910 427 3927
rect 252 3870 427 3887
rect 252 3830 427 3847
rect 252 3790 427 3807
rect 252 3750 427 3767
rect 252 3710 427 3727
rect 252 3670 427 3687
rect 252 3630 427 3647
rect 252 3590 427 3607
rect 252 3550 427 3567
rect 252 3510 427 3527
rect 252 3470 427 3487
rect 252 3430 427 3447
rect 252 3390 427 3407
rect 252 3350 427 3367
rect 252 3310 427 3327
rect 252 3270 427 3287
rect 252 3230 427 3247
rect 252 3190 427 3207
rect 252 3150 427 3167
rect 252 3110 427 3127
rect 252 3070 427 3087
rect 252 3030 427 3047
rect 252 2990 427 3007
rect 252 2950 427 2967
rect 252 2910 427 2927
rect 252 2870 427 2887
rect 252 2830 427 2847
rect 252 2790 427 2807
rect 252 2750 427 2767
rect 252 2710 427 2727
rect 252 2670 427 2687
rect 252 2630 427 2647
rect 252 2590 427 2607
rect 252 2550 427 2567
rect 252 2510 427 2527
rect 252 2470 427 2487
rect 252 2430 427 2447
rect 252 2390 427 2407
rect 252 2350 427 2367
rect 252 2310 427 2327
rect 252 2270 427 2287
rect 252 2230 427 2247
rect 252 2190 427 2207
rect 252 2150 427 2167
rect 252 2110 427 2127
rect 252 2070 427 2087
rect 252 2030 427 2047
rect 252 1990 427 2007
rect 252 1950 427 1967
rect 252 1910 427 1927
rect 252 1870 427 1887
rect 252 1830 427 1847
rect 252 1790 427 1807
rect 252 1750 427 1767
rect 252 1710 427 1727
rect 252 1670 427 1687
rect 252 1630 427 1647
rect 252 1590 427 1607
rect 252 1550 427 1567
rect 252 1510 427 1527
rect 252 1470 427 1487
rect 252 1430 427 1447
rect 252 1390 427 1407
rect 252 1350 427 1367
rect 252 1310 427 1327
rect 18845 9550 19020 9567
rect 18845 9510 19020 9527
rect 18845 9470 19020 9487
rect 18845 9430 19020 9447
rect 18845 9390 19020 9407
rect 18845 9350 19020 9367
rect 18845 9310 19020 9327
rect 18845 9270 19020 9287
rect 18845 9230 19020 9247
rect 18845 9190 19020 9207
rect 18845 9150 19020 9167
rect 18845 9110 19020 9127
rect 18845 9070 19020 9087
rect 18845 9030 19020 9047
rect 18845 8990 19020 9007
rect 18845 8950 19020 8967
rect 18845 8910 19020 8927
rect 18845 8870 19020 8887
rect 18845 8830 19020 8847
rect 18845 8790 19020 8807
rect 18845 8750 19020 8767
rect 18845 8710 19020 8727
rect 18845 8670 19020 8687
rect 18845 8630 19020 8647
rect 18845 8590 19020 8607
rect 18845 8550 19020 8567
rect 18845 8510 19020 8527
rect 18845 8470 19020 8487
rect 18845 8430 19020 8447
rect 18845 8390 19020 8407
rect 18845 8350 19020 8367
rect 18845 8310 19020 8327
rect 18845 8270 19020 8287
rect 18845 8230 19020 8247
rect 18845 8190 19020 8207
rect 18845 8150 19020 8167
rect 18845 8110 19020 8127
rect 18845 8070 19020 8087
rect 18845 8030 19020 8047
rect 18845 7990 19020 8007
rect 18845 7950 19020 7967
rect 18845 7910 19020 7927
rect 18845 7870 19020 7887
rect 18845 7830 19020 7847
rect 18845 7790 19020 7807
rect 18845 7750 19020 7767
rect 18845 7710 19020 7727
rect 18845 7670 19020 7687
rect 18845 7630 19020 7647
rect 18845 7590 19020 7607
rect 18845 7550 19020 7567
rect 18845 7510 19020 7527
rect 18845 7470 19020 7487
rect 18845 7430 19020 7447
rect 18845 7390 19020 7407
rect 18845 7350 19020 7367
rect 18845 7310 19020 7327
rect 18845 7270 19020 7287
rect 18845 7230 19020 7247
rect 18845 7190 19020 7207
rect 18845 7150 19020 7167
rect 18845 7110 19020 7127
rect 18845 7070 19020 7087
rect 18845 7030 19020 7047
rect 18845 6990 19020 7007
rect 18845 6950 19020 6967
rect 18845 6910 19020 6927
rect 18845 6870 19020 6887
rect 18845 6830 19020 6847
rect 18845 6790 19020 6807
rect 18845 6750 19020 6767
rect 18845 6710 19020 6727
rect 18846 6669 19021 6686
rect 18845 6630 19020 6647
rect 18845 6590 19020 6607
rect 18845 6550 19020 6567
rect 18845 6510 19020 6527
rect 18845 6470 19020 6487
rect 18845 6430 19020 6447
rect 18845 6390 19020 6407
rect 18845 6350 19020 6367
rect 18845 6310 19020 6327
rect 18845 6270 19020 6287
rect 18845 6230 19020 6247
rect 18845 6190 19020 6207
rect 18845 6150 19020 6167
rect 18845 6110 19020 6127
rect 18845 6070 19020 6087
rect 18845 6030 19020 6047
rect 18845 5990 19020 6007
rect 18845 5950 19020 5967
rect 18845 5910 19020 5927
rect 18845 5870 19020 5887
rect 18845 5830 19020 5847
rect 18844 5789 19019 5806
rect 18845 5750 19020 5767
rect 18845 5710 19020 5727
rect 18845 5670 19020 5687
rect 18845 5630 19020 5647
rect 18845 5590 19020 5607
rect 18845 5550 19020 5567
rect 18845 5510 19020 5527
rect 18845 5470 19020 5487
rect 18845 5430 19020 5447
rect 18845 5390 19020 5407
rect 18845 5350 19020 5367
rect 18845 5310 19020 5327
rect 18845 5270 19020 5287
rect 18845 5230 19020 5247
rect 18845 5190 19020 5207
rect 18845 5150 19020 5167
rect 18845 5110 19020 5127
rect 18845 5070 19020 5087
rect 18845 5030 19020 5047
rect 18845 4990 19020 5007
rect 18845 4950 19020 4967
rect 18845 4910 19020 4927
rect 18845 4870 19020 4887
rect 18845 4830 19020 4847
rect 18845 4790 19020 4807
rect 18845 4750 19020 4767
rect 18845 4710 19020 4727
rect 18845 4670 19020 4687
rect 18845 4630 19020 4647
rect 18845 4590 19020 4607
rect 18845 4550 19020 4567
rect 18845 4510 19020 4527
rect 18845 4470 19020 4487
rect 18845 4430 19020 4447
rect 18845 4390 19020 4407
rect 18845 4350 19020 4367
rect 18845 4310 19020 4327
rect 18845 4270 19020 4287
rect 18845 4230 19020 4247
rect 18845 4190 19020 4207
rect 18845 4150 19020 4167
rect 18845 4110 19020 4127
rect 18845 4070 19020 4087
rect 18845 4030 19020 4047
rect 18845 3990 19020 4007
rect 18845 3950 19020 3967
rect 18845 3910 19020 3927
rect 18845 3870 19020 3887
rect 18845 3830 19020 3847
rect 18845 3790 19020 3807
rect 18845 3750 19020 3767
rect 18845 3710 19020 3727
rect 18845 3670 19020 3687
rect 18845 3630 19020 3647
rect 18845 3590 19020 3607
rect 18845 3550 19020 3567
rect 18845 3510 19020 3527
rect 18845 3470 19020 3487
rect 18845 3430 19020 3447
rect 18845 3390 19020 3407
rect 18845 3350 19020 3367
rect 18845 3310 19020 3327
rect 18845 3270 19020 3287
rect 18845 3230 19020 3247
rect 18845 3190 19020 3207
rect 18845 3150 19020 3167
rect 18845 3110 19020 3127
rect 18845 3070 19020 3087
rect 18845 3030 19020 3047
rect 18845 2990 19020 3007
rect 18845 2950 19020 2967
rect 18845 2910 19020 2927
rect 18845 2870 19020 2887
rect 18845 2830 19020 2847
rect 18845 2790 19020 2807
rect 18845 2750 19020 2767
rect 18845 2707 19020 2724
rect 18845 2670 19020 2687
rect 18845 2630 19020 2647
rect 18845 2590 19020 2607
rect 18845 2550 19020 2567
rect 18845 2510 19020 2527
rect 18845 2470 19020 2487
rect 18845 2430 19020 2447
rect 18845 2390 19020 2407
rect 18845 2350 19020 2367
rect 18845 2310 19020 2327
rect 18845 2270 19020 2287
rect 18845 2230 19020 2247
rect 18845 2190 19020 2207
rect 18845 2150 19020 2167
rect 18845 2110 19020 2127
rect 18845 2070 19020 2087
rect 18845 2030 19020 2047
rect 18845 1990 19020 2007
rect 18845 1950 19020 1967
rect 18845 1910 19020 1927
rect 18845 1870 19020 1887
rect 18845 1830 19020 1847
rect 18845 1790 19020 1807
rect 18845 1750 19020 1767
rect 18845 1710 19020 1727
rect 18845 1670 19020 1687
rect 18845 1630 19020 1647
rect 18845 1590 19020 1607
rect 18845 1550 19020 1567
rect 18845 1510 19020 1527
rect 18845 1470 19020 1487
rect 18845 1430 19020 1447
rect 18845 1390 19020 1407
rect 18845 1350 19020 1367
rect 18845 1310 19020 1327
rect 252 1270 427 1287
rect 252 1230 427 1247
rect 252 1190 427 1207
rect 252 1150 427 1167
rect 18845 1270 19020 1287
rect 18845 1230 19020 1247
rect 18845 1190 19020 1207
rect 18845 1150 19020 1167
rect 252 1110 427 1127
rect 252 1070 427 1087
rect 252 1030 427 1047
rect 252 990 427 1007
rect 252 950 427 967
rect 252 910 427 927
rect 252 870 427 887
rect 252 830 427 847
rect 252 790 427 807
rect 252 750 427 767
rect 252 710 427 727
rect 252 670 427 687
rect 252 630 427 647
rect 252 590 427 607
rect 252 550 427 567
rect 252 510 427 527
rect 252 470 427 487
rect 18845 1110 19020 1127
rect 18845 1070 19020 1087
rect 18845 1030 19020 1047
rect 18845 990 19020 1007
rect 18845 950 19020 967
rect 18845 910 19020 927
rect 18845 870 19020 887
rect 18845 830 19020 847
rect 18845 790 19020 807
rect 18845 750 19020 767
rect 18845 710 19020 727
rect 18845 670 19020 687
rect 18845 630 19020 647
rect 18845 590 19020 607
rect 18845 550 19020 567
rect 18845 510 19020 527
rect 18845 470 19020 487
<< locali >>
rect 21346 11625 21762 11638
rect 21346 11419 21643 11625
rect 21749 11419 21762 11625
rect 21346 11407 21762 11419
rect 21346 10746 21762 10759
rect 21346 10540 21643 10746
rect 21749 10540 21762 10746
rect 21346 10528 21762 10540
rect 1487 10052 1633 10060
rect 1487 9973 1494 10052
rect 1625 9973 1633 10052
rect 0 21 207 9950
rect 755 9940 901 9971
rect 755 9912 765 9940
rect 793 9912 812 9940
rect 840 9912 859 9940
rect 887 9912 901 9940
rect 755 9893 901 9912
rect 755 9865 765 9893
rect 793 9865 812 9893
rect 840 9865 859 9893
rect 887 9865 901 9893
rect 755 9846 901 9865
rect 755 9818 765 9846
rect 793 9818 812 9846
rect 840 9818 859 9846
rect 887 9818 901 9846
rect 238 9567 445 9731
rect 238 9550 252 9567
rect 427 9550 445 9567
rect 238 9527 445 9550
rect 238 9510 252 9527
rect 427 9510 445 9527
rect 238 9487 445 9510
rect 238 9470 252 9487
rect 427 9470 445 9487
rect 238 9447 445 9470
rect 238 9430 252 9447
rect 427 9430 445 9447
rect 238 9407 445 9430
rect 238 9390 252 9407
rect 427 9390 445 9407
rect 238 9367 445 9390
rect 238 9350 252 9367
rect 427 9350 445 9367
rect 238 9327 445 9350
rect 238 9310 252 9327
rect 427 9310 445 9327
rect 238 9287 445 9310
rect 238 9270 252 9287
rect 427 9270 445 9287
rect 238 9247 445 9270
rect 238 9230 252 9247
rect 427 9230 445 9247
rect 238 9207 445 9230
rect 238 9190 252 9207
rect 427 9190 445 9207
rect 238 9167 445 9190
rect 238 9150 252 9167
rect 427 9150 445 9167
rect 238 9127 445 9150
rect 238 9110 252 9127
rect 427 9110 445 9127
rect 238 9087 445 9110
rect 238 9070 252 9087
rect 427 9070 445 9087
rect 238 9047 445 9070
rect 238 9030 252 9047
rect 427 9030 445 9047
rect 238 9007 445 9030
rect 238 8990 252 9007
rect 427 8990 445 9007
rect 238 8967 445 8990
rect 238 8950 252 8967
rect 427 8950 445 8967
rect 238 8927 445 8950
rect 238 8910 252 8927
rect 427 8910 445 8927
rect 238 8887 445 8910
rect 238 8870 252 8887
rect 427 8870 445 8887
rect 238 8847 445 8870
rect 238 8830 252 8847
rect 427 8830 445 8847
rect 238 8807 445 8830
rect 238 8790 252 8807
rect 427 8790 445 8807
rect 238 8767 445 8790
rect 238 8750 252 8767
rect 427 8750 445 8767
rect 238 8727 445 8750
rect 238 8710 252 8727
rect 427 8710 445 8727
rect 238 8687 445 8710
rect 238 8670 252 8687
rect 427 8670 445 8687
rect 238 8647 445 8670
rect 238 8630 252 8647
rect 427 8630 445 8647
rect 238 8607 445 8630
rect 238 8590 252 8607
rect 427 8590 445 8607
rect 238 8567 445 8590
rect 238 8550 252 8567
rect 427 8550 445 8567
rect 238 8527 445 8550
rect 238 8510 252 8527
rect 427 8510 445 8527
rect 238 8487 445 8510
rect 238 8470 252 8487
rect 427 8470 445 8487
rect 238 8447 445 8470
rect 238 8430 252 8447
rect 427 8430 445 8447
rect 238 8407 445 8430
rect 238 8390 252 8407
rect 427 8390 445 8407
rect 238 8367 445 8390
rect 238 8350 252 8367
rect 427 8350 445 8367
rect 238 8327 445 8350
rect 238 8310 252 8327
rect 427 8310 445 8327
rect 238 8287 445 8310
rect 238 8270 252 8287
rect 427 8270 445 8287
rect 238 8247 445 8270
rect 238 8230 252 8247
rect 427 8230 445 8247
rect 238 8207 445 8230
rect 238 8190 252 8207
rect 427 8190 445 8207
rect 238 8167 445 8190
rect 238 8150 252 8167
rect 427 8150 445 8167
rect 238 8127 445 8150
rect 238 8110 252 8127
rect 427 8110 445 8127
rect 238 8087 445 8110
rect 238 8070 252 8087
rect 427 8070 445 8087
rect 238 8047 445 8070
rect 238 8030 252 8047
rect 427 8030 445 8047
rect 238 8007 445 8030
rect 238 7990 252 8007
rect 427 7990 445 8007
rect 238 7967 445 7990
rect 238 7950 252 7967
rect 427 7950 445 7967
rect 238 7927 445 7950
rect 238 7910 252 7927
rect 427 7910 445 7927
rect 238 7887 445 7910
rect 238 7870 252 7887
rect 427 7870 445 7887
rect 238 7847 445 7870
rect 238 7830 252 7847
rect 427 7830 445 7847
rect 238 7807 445 7830
rect 238 7790 252 7807
rect 427 7790 445 7807
rect 238 7767 445 7790
rect 238 7750 252 7767
rect 427 7750 445 7767
rect 238 7727 445 7750
rect 238 7710 252 7727
rect 427 7710 445 7727
rect 238 7687 445 7710
rect 238 7670 252 7687
rect 427 7670 445 7687
rect 238 7647 445 7670
rect 238 7630 252 7647
rect 427 7630 445 7647
rect 238 7607 445 7630
rect 238 7590 252 7607
rect 427 7590 445 7607
rect 238 7567 445 7590
rect 238 7550 252 7567
rect 427 7550 445 7567
rect 238 7527 445 7550
rect 238 7510 252 7527
rect 427 7510 445 7527
rect 238 7487 445 7510
rect 238 7470 252 7487
rect 427 7470 445 7487
rect 238 7447 445 7470
rect 238 7430 252 7447
rect 427 7430 445 7447
rect 238 7407 445 7430
rect 238 7390 252 7407
rect 427 7390 445 7407
rect 238 7367 445 7390
rect 238 7350 252 7367
rect 427 7350 445 7367
rect 238 7327 445 7350
rect 238 7310 252 7327
rect 427 7310 445 7327
rect 238 7287 445 7310
rect 238 7270 252 7287
rect 427 7270 445 7287
rect 238 7247 445 7270
rect 238 7230 252 7247
rect 427 7230 445 7247
rect 238 7207 445 7230
rect 238 7190 252 7207
rect 427 7190 445 7207
rect 238 7167 445 7190
rect 238 7150 252 7167
rect 427 7150 445 7167
rect 238 7127 445 7150
rect 238 7110 252 7127
rect 427 7110 445 7127
rect 238 7087 445 7110
rect 238 7070 252 7087
rect 427 7070 445 7087
rect 238 7047 445 7070
rect 238 7030 252 7047
rect 427 7030 445 7047
rect 238 7007 445 7030
rect 238 6990 252 7007
rect 427 6990 445 7007
rect 238 6967 445 6990
rect 238 6950 252 6967
rect 427 6950 445 6967
rect 238 6927 445 6950
rect 238 6910 252 6927
rect 427 6910 445 6927
rect 238 6887 445 6910
rect 238 6870 252 6887
rect 427 6870 445 6887
rect 238 6847 445 6870
rect 238 6830 252 6847
rect 427 6830 445 6847
rect 238 6807 445 6830
rect 238 6790 252 6807
rect 427 6790 445 6807
rect 238 6767 445 6790
rect 238 6750 252 6767
rect 427 6750 445 6767
rect 238 6727 445 6750
rect 238 6710 252 6727
rect 427 6710 445 6727
rect 238 6687 445 6710
rect 238 6670 252 6687
rect 427 6670 445 6687
rect 238 6647 445 6670
rect 238 6630 252 6647
rect 427 6630 445 6647
rect 238 6607 445 6630
rect 238 6590 252 6607
rect 427 6590 445 6607
rect 238 6567 445 6590
rect 238 6550 252 6567
rect 427 6550 445 6567
rect 238 6527 445 6550
rect 238 6510 252 6527
rect 427 6510 445 6527
rect 238 6487 445 6510
rect 238 6470 252 6487
rect 427 6470 445 6487
rect 238 6447 445 6470
rect 238 6430 252 6447
rect 427 6430 445 6447
rect 238 6407 445 6430
rect 238 6390 252 6407
rect 427 6390 445 6407
rect 238 6367 445 6390
rect 238 6350 252 6367
rect 427 6350 445 6367
rect 238 6327 445 6350
rect 238 6310 252 6327
rect 427 6310 445 6327
rect 238 6287 445 6310
rect 238 6270 252 6287
rect 427 6270 445 6287
rect 238 6247 445 6270
rect 238 6230 252 6247
rect 427 6230 445 6247
rect 238 6207 445 6230
rect 238 6190 252 6207
rect 427 6190 445 6207
rect 238 6167 445 6190
rect 238 6150 252 6167
rect 427 6150 445 6167
rect 238 6127 445 6150
rect 238 6110 252 6127
rect 427 6110 445 6127
rect 238 6087 445 6110
rect 238 6070 252 6087
rect 427 6070 445 6087
rect 238 6047 445 6070
rect 238 6030 252 6047
rect 427 6030 445 6047
rect 238 6007 445 6030
rect 238 5990 252 6007
rect 427 5990 445 6007
rect 238 5967 445 5990
rect 238 5950 252 5967
rect 427 5950 445 5967
rect 238 5927 445 5950
rect 238 5910 252 5927
rect 427 5910 445 5927
rect 238 5887 445 5910
rect 238 5870 252 5887
rect 427 5870 445 5887
rect 238 5847 445 5870
rect 238 5830 252 5847
rect 427 5830 445 5847
rect 238 5807 445 5830
rect 238 5790 252 5807
rect 427 5790 445 5807
rect 238 5767 445 5790
rect 238 5750 252 5767
rect 427 5750 445 5767
rect 238 5727 445 5750
rect 238 5710 252 5727
rect 427 5710 445 5727
rect 238 5687 445 5710
rect 238 5670 252 5687
rect 427 5670 445 5687
rect 238 5647 445 5670
rect 238 5630 252 5647
rect 427 5630 445 5647
rect 238 5607 445 5630
rect 238 5590 252 5607
rect 427 5590 445 5607
rect 238 5567 445 5590
rect 238 5550 252 5567
rect 427 5550 445 5567
rect 238 5527 445 5550
rect 238 5510 252 5527
rect 427 5510 445 5527
rect 238 5487 445 5510
rect 238 5470 252 5487
rect 427 5470 445 5487
rect 238 5447 445 5470
rect 238 5430 252 5447
rect 427 5430 445 5447
rect 238 5407 445 5430
rect 238 5390 252 5407
rect 427 5390 445 5407
rect 238 5367 445 5390
rect 238 5350 252 5367
rect 427 5350 445 5367
rect 238 5327 445 5350
rect 238 5310 252 5327
rect 427 5310 445 5327
rect 238 5287 445 5310
rect 238 5270 252 5287
rect 427 5270 445 5287
rect 238 5247 445 5270
rect 238 5230 252 5247
rect 427 5230 445 5247
rect 238 5207 445 5230
rect 238 5190 252 5207
rect 427 5190 445 5207
rect 238 5167 445 5190
rect 238 5150 252 5167
rect 427 5150 445 5167
rect 238 5127 445 5150
rect 238 5110 252 5127
rect 427 5110 445 5127
rect 238 5087 445 5110
rect 238 5070 252 5087
rect 427 5070 445 5087
rect 238 5047 445 5070
rect 238 5030 252 5047
rect 427 5030 445 5047
rect 238 5007 445 5030
rect 238 4990 252 5007
rect 427 4990 445 5007
rect 238 4967 445 4990
rect 238 4950 252 4967
rect 427 4950 445 4967
rect 238 4927 445 4950
rect 238 4910 252 4927
rect 427 4910 445 4927
rect 238 4887 445 4910
rect 238 4870 252 4887
rect 427 4870 445 4887
rect 238 4847 445 4870
rect 238 4830 252 4847
rect 427 4830 445 4847
rect 238 4807 445 4830
rect 238 4790 252 4807
rect 427 4790 445 4807
rect 238 4767 445 4790
rect 238 4750 252 4767
rect 427 4750 445 4767
rect 238 4727 445 4750
rect 238 4710 252 4727
rect 427 4710 445 4727
rect 238 4687 445 4710
rect 238 4670 252 4687
rect 427 4670 445 4687
rect 238 4647 445 4670
rect 238 4630 252 4647
rect 427 4630 445 4647
rect 238 4607 445 4630
rect 238 4590 252 4607
rect 427 4590 445 4607
rect 238 4567 445 4590
rect 238 4550 252 4567
rect 427 4550 445 4567
rect 238 4527 445 4550
rect 238 4510 252 4527
rect 427 4510 445 4527
rect 238 4487 445 4510
rect 238 4470 252 4487
rect 427 4470 445 4487
rect 238 4447 445 4470
rect 238 4430 252 4447
rect 427 4430 445 4447
rect 238 4407 445 4430
rect 238 4390 252 4407
rect 427 4390 445 4407
rect 238 4367 445 4390
rect 238 4350 252 4367
rect 427 4350 445 4367
rect 238 4327 445 4350
rect 238 4310 252 4327
rect 427 4310 445 4327
rect 238 4287 445 4310
rect 238 4270 252 4287
rect 427 4270 445 4287
rect 238 4247 445 4270
rect 238 4230 252 4247
rect 427 4230 445 4247
rect 238 4207 445 4230
rect 238 4190 252 4207
rect 427 4190 445 4207
rect 238 4167 445 4190
rect 238 4150 252 4167
rect 427 4150 445 4167
rect 238 4127 445 4150
rect 238 4110 252 4127
rect 427 4110 445 4127
rect 238 4087 445 4110
rect 238 4070 252 4087
rect 427 4070 445 4087
rect 238 4047 445 4070
rect 238 4030 252 4047
rect 427 4030 445 4047
rect 238 4007 445 4030
rect 238 3990 252 4007
rect 427 3990 445 4007
rect 238 3967 445 3990
rect 238 3950 252 3967
rect 427 3950 445 3967
rect 238 3927 445 3950
rect 238 3910 252 3927
rect 427 3910 445 3927
rect 238 3887 445 3910
rect 238 3870 252 3887
rect 427 3870 445 3887
rect 238 3847 445 3870
rect 238 3830 252 3847
rect 427 3830 445 3847
rect 238 3807 445 3830
rect 238 3790 252 3807
rect 427 3790 445 3807
rect 238 3767 445 3790
rect 238 3750 252 3767
rect 427 3750 445 3767
rect 238 3727 445 3750
rect 238 3710 252 3727
rect 427 3710 445 3727
rect 238 3687 445 3710
rect 238 3670 252 3687
rect 427 3670 445 3687
rect 238 3647 445 3670
rect 238 3630 252 3647
rect 427 3630 445 3647
rect 238 3607 445 3630
rect 238 3590 252 3607
rect 427 3590 445 3607
rect 238 3567 445 3590
rect 238 3550 252 3567
rect 427 3550 445 3567
rect 238 3527 445 3550
rect 238 3510 252 3527
rect 427 3510 445 3527
rect 238 3487 445 3510
rect 238 3470 252 3487
rect 427 3470 445 3487
rect 238 3447 445 3470
rect 238 3430 252 3447
rect 427 3430 445 3447
rect 238 3407 445 3430
rect 238 3390 252 3407
rect 427 3390 445 3407
rect 238 3367 445 3390
rect 238 3350 252 3367
rect 427 3350 445 3367
rect 238 3327 445 3350
rect 238 3310 252 3327
rect 427 3310 445 3327
rect 238 3287 445 3310
rect 238 3270 252 3287
rect 427 3270 445 3287
rect 238 3247 445 3270
rect 238 3230 252 3247
rect 427 3230 445 3247
rect 238 3207 445 3230
rect 238 3190 252 3207
rect 427 3190 445 3207
rect 238 3167 445 3190
rect 238 3150 252 3167
rect 427 3150 445 3167
rect 238 3127 445 3150
rect 238 3110 252 3127
rect 427 3110 445 3127
rect 238 3087 445 3110
rect 238 3070 252 3087
rect 427 3070 445 3087
rect 238 3047 445 3070
rect 238 3030 252 3047
rect 427 3030 445 3047
rect 238 3007 445 3030
rect 238 2990 252 3007
rect 427 2990 445 3007
rect 238 2967 445 2990
rect 238 2950 252 2967
rect 427 2950 445 2967
rect 238 2927 445 2950
rect 238 2910 252 2927
rect 427 2910 445 2927
rect 238 2887 445 2910
rect 238 2870 252 2887
rect 427 2870 445 2887
rect 238 2847 445 2870
rect 238 2830 252 2847
rect 427 2830 445 2847
rect 238 2807 445 2830
rect 238 2790 252 2807
rect 427 2790 445 2807
rect 238 2767 445 2790
rect 238 2750 252 2767
rect 427 2750 445 2767
rect 238 2727 445 2750
rect 238 2710 252 2727
rect 427 2710 445 2727
rect 238 2687 445 2710
rect 238 2670 252 2687
rect 427 2670 445 2687
rect 238 2647 445 2670
rect 238 2630 252 2647
rect 427 2630 445 2647
rect 238 2607 445 2630
rect 238 2590 252 2607
rect 427 2590 445 2607
rect 238 2567 445 2590
rect 238 2550 252 2567
rect 427 2550 445 2567
rect 238 2527 445 2550
rect 238 2510 252 2527
rect 427 2510 445 2527
rect 238 2487 445 2510
rect 238 2470 252 2487
rect 427 2470 445 2487
rect 238 2447 445 2470
rect 238 2430 252 2447
rect 427 2430 445 2447
rect 238 2407 445 2430
rect 238 2390 252 2407
rect 427 2390 445 2407
rect 238 2367 445 2390
rect 238 2350 252 2367
rect 427 2350 445 2367
rect 238 2327 445 2350
rect 238 2310 252 2327
rect 427 2310 445 2327
rect 238 2287 445 2310
rect 238 2270 252 2287
rect 427 2270 445 2287
rect 238 2247 445 2270
rect 238 2230 252 2247
rect 427 2230 445 2247
rect 238 2207 445 2230
rect 238 2190 252 2207
rect 427 2190 445 2207
rect 238 2167 445 2190
rect 238 2150 252 2167
rect 427 2150 445 2167
rect 238 2127 445 2150
rect 238 2110 252 2127
rect 427 2110 445 2127
rect 238 2087 445 2110
rect 238 2070 252 2087
rect 427 2070 445 2087
rect 238 2047 445 2070
rect 238 2030 252 2047
rect 427 2030 445 2047
rect 238 2007 445 2030
rect 238 1990 252 2007
rect 427 1990 445 2007
rect 238 1967 445 1990
rect 238 1950 252 1967
rect 427 1950 445 1967
rect 238 1927 445 1950
rect 238 1910 252 1927
rect 427 1910 445 1927
rect 238 1887 445 1910
rect 238 1870 252 1887
rect 427 1870 445 1887
rect 238 1847 445 1870
rect 238 1830 252 1847
rect 427 1830 445 1847
rect 238 1807 445 1830
rect 238 1790 252 1807
rect 427 1790 445 1807
rect 238 1767 445 1790
rect 238 1750 252 1767
rect 427 1750 445 1767
rect 238 1727 445 1750
rect 238 1710 252 1727
rect 427 1710 445 1727
rect 238 1687 445 1710
rect 238 1670 252 1687
rect 427 1670 445 1687
rect 238 1647 445 1670
rect 238 1630 252 1647
rect 427 1630 445 1647
rect 238 1607 445 1630
rect 238 1590 252 1607
rect 427 1590 445 1607
rect 238 1567 445 1590
rect 238 1550 252 1567
rect 427 1550 445 1567
rect 238 1527 445 1550
rect 238 1510 252 1527
rect 427 1510 445 1527
rect 238 1487 445 1510
rect 238 1470 252 1487
rect 427 1470 445 1487
rect 238 1447 445 1470
rect 238 1430 252 1447
rect 427 1430 445 1447
rect 238 1407 445 1430
rect 238 1390 252 1407
rect 427 1390 445 1407
rect 238 1367 445 1390
rect 238 1350 252 1367
rect 427 1350 445 1367
rect 238 1327 445 1350
rect 238 1310 252 1327
rect 427 1310 445 1327
rect 238 1287 445 1310
rect 238 1270 252 1287
rect 427 1270 445 1287
rect 238 1247 445 1270
rect 238 1230 252 1247
rect 427 1230 445 1247
rect 238 1207 445 1230
rect 238 1190 252 1207
rect 427 1190 445 1207
rect 238 1167 445 1190
rect 238 1150 252 1167
rect 427 1150 445 1167
rect 238 1127 445 1150
rect 238 1110 252 1127
rect 427 1110 445 1127
rect 238 1087 445 1110
rect 238 1070 252 1087
rect 427 1070 445 1087
rect 238 1047 445 1070
rect 238 1030 252 1047
rect 427 1030 445 1047
rect 238 1007 445 1030
rect 238 990 252 1007
rect 427 990 445 1007
rect 238 967 445 990
rect 238 950 252 967
rect 427 950 445 967
rect 238 927 445 950
rect 238 910 252 927
rect 427 910 445 927
rect 238 887 445 910
rect 238 870 252 887
rect 427 870 445 887
rect 238 847 445 870
rect 238 830 252 847
rect 427 830 445 847
rect 238 807 445 830
rect 238 790 252 807
rect 427 790 445 807
rect 238 767 445 790
rect 238 750 252 767
rect 427 750 445 767
rect 238 727 445 750
rect 238 710 252 727
rect 427 710 445 727
rect 238 687 445 710
rect 238 670 252 687
rect 427 670 445 687
rect 238 647 445 670
rect 238 630 252 647
rect 427 630 445 647
rect 238 607 445 630
rect 238 590 252 607
rect 427 590 445 607
rect 238 567 445 590
rect 238 550 252 567
rect 427 550 445 567
rect 238 527 445 550
rect 238 510 252 527
rect 427 510 445 527
rect 238 487 445 510
rect 238 470 252 487
rect 427 470 445 487
rect 238 240 445 470
rect 536 8881 570 9493
rect 536 8864 544 8881
rect 561 8864 570 8881
rect 536 8379 570 8864
rect 536 8362 544 8379
rect 561 8362 570 8379
rect 536 7877 570 8362
rect 536 7860 544 7877
rect 561 7860 570 7877
rect 536 7375 570 7860
rect 536 7358 544 7375
rect 561 7358 570 7375
rect 536 6873 570 7358
rect 536 6856 544 6873
rect 561 6856 570 6873
rect 536 6371 570 6856
rect 536 6354 544 6371
rect 561 6354 570 6371
rect 536 5869 570 6354
rect 536 5852 544 5869
rect 561 5852 570 5869
rect 536 5367 570 5852
rect 536 5350 544 5367
rect 561 5350 570 5367
rect 536 4865 570 5350
rect 536 4848 544 4865
rect 561 4848 570 4865
rect 536 4363 570 4848
rect 536 4346 544 4363
rect 561 4346 570 4363
rect 536 3861 570 4346
rect 536 3844 544 3861
rect 561 3844 570 3861
rect 536 3359 570 3844
rect 536 3342 544 3359
rect 561 3342 570 3359
rect 536 2857 570 3342
rect 536 2840 544 2857
rect 561 2840 570 2857
rect 536 2355 570 2840
rect 536 2338 544 2355
rect 561 2338 570 2355
rect 536 1853 570 2338
rect 536 1836 544 1853
rect 561 1836 570 1853
rect 536 1351 570 1836
rect 536 1334 544 1351
rect 561 1334 570 1351
rect 536 0 570 1334
rect 590 8687 624 9493
rect 590 8670 598 8687
rect 615 8670 624 8687
rect 590 8185 624 8670
rect 590 8168 598 8185
rect 615 8168 624 8185
rect 590 7683 624 8168
rect 590 7666 598 7683
rect 615 7666 624 7683
rect 590 7181 624 7666
rect 590 7164 598 7181
rect 615 7164 624 7181
rect 590 6679 624 7164
rect 590 6662 598 6679
rect 615 6662 624 6679
rect 590 6177 624 6662
rect 590 6160 598 6177
rect 615 6160 624 6177
rect 590 5675 624 6160
rect 590 5658 598 5675
rect 615 5658 624 5675
rect 590 5173 624 5658
rect 590 5156 598 5173
rect 615 5156 624 5173
rect 590 4671 624 5156
rect 590 4654 598 4671
rect 615 4654 624 4671
rect 590 4169 624 4654
rect 590 4152 598 4169
rect 615 4152 624 4169
rect 590 3667 624 4152
rect 590 3650 598 3667
rect 615 3650 624 3667
rect 590 3165 624 3650
rect 590 3148 598 3165
rect 615 3148 624 3165
rect 590 2663 624 3148
rect 590 2646 598 2663
rect 615 2646 624 2663
rect 590 2161 624 2646
rect 590 2144 598 2161
rect 615 2144 624 2161
rect 590 1659 624 2144
rect 590 1642 598 1659
rect 615 1642 624 1659
rect 590 1157 624 1642
rect 590 1140 598 1157
rect 615 1140 624 1157
rect 590 0 624 1140
rect 644 9118 712 9493
rect 644 9098 650 9118
rect 670 9098 689 9118
rect 709 9098 712 9118
rect 644 8616 712 9098
rect 644 8596 650 8616
rect 670 8596 689 8616
rect 709 8596 712 8616
rect 644 8114 712 8596
rect 644 8094 650 8114
rect 670 8094 689 8114
rect 709 8094 712 8114
rect 644 7612 712 8094
rect 644 7592 650 7612
rect 670 7592 689 7612
rect 709 7592 712 7612
rect 644 7110 712 7592
rect 644 7090 650 7110
rect 670 7090 689 7110
rect 709 7090 712 7110
rect 644 6608 712 7090
rect 644 6588 650 6608
rect 670 6588 689 6608
rect 709 6588 712 6608
rect 644 6106 712 6588
rect 644 6086 650 6106
rect 670 6086 689 6106
rect 709 6086 712 6106
rect 644 5604 712 6086
rect 644 5584 650 5604
rect 670 5584 689 5604
rect 709 5584 712 5604
rect 644 5102 712 5584
rect 644 5082 650 5102
rect 670 5082 689 5102
rect 709 5082 712 5102
rect 644 4600 712 5082
rect 644 4580 650 4600
rect 670 4580 689 4600
rect 709 4580 712 4600
rect 644 4098 712 4580
rect 644 4078 650 4098
rect 670 4078 689 4098
rect 709 4078 712 4098
rect 644 3596 712 4078
rect 644 3576 650 3596
rect 670 3576 689 3596
rect 709 3576 712 3596
rect 644 3094 712 3576
rect 644 3074 650 3094
rect 670 3074 689 3094
rect 709 3074 712 3094
rect 644 2592 712 3074
rect 644 2572 650 2592
rect 670 2572 689 2592
rect 709 2572 712 2592
rect 644 2090 712 2572
rect 644 2070 650 2090
rect 670 2070 689 2090
rect 709 2070 712 2090
rect 644 1588 712 2070
rect 644 1568 650 1588
rect 670 1568 689 1588
rect 709 1568 712 1588
rect 644 1086 712 1568
rect 644 1066 650 1086
rect 670 1066 689 1086
rect 709 1066 712 1086
rect 644 584 712 1066
rect 644 564 650 584
rect 670 564 689 584
rect 709 564 712 584
rect 644 0 712 564
rect 755 9414 901 9818
rect 755 9394 761 9414
rect 781 9394 800 9414
rect 820 9394 839 9414
rect 859 9394 878 9414
rect 898 9394 901 9414
rect 755 9372 901 9394
rect 755 9352 761 9372
rect 781 9352 800 9372
rect 820 9352 839 9372
rect 859 9352 878 9372
rect 898 9352 901 9372
rect 755 9244 901 9352
rect 755 9224 761 9244
rect 781 9224 800 9244
rect 820 9224 839 9244
rect 859 9224 878 9244
rect 898 9224 901 9244
rect 755 8912 901 9224
rect 755 8892 761 8912
rect 781 8892 800 8912
rect 820 8892 839 8912
rect 859 8892 878 8912
rect 898 8892 901 8912
rect 755 8410 901 8892
rect 755 8390 761 8410
rect 781 8390 800 8410
rect 820 8390 839 8410
rect 859 8390 878 8410
rect 898 8390 901 8410
rect 755 7908 901 8390
rect 755 7888 761 7908
rect 781 7888 800 7908
rect 820 7888 839 7908
rect 859 7888 878 7908
rect 898 7888 901 7908
rect 755 7406 901 7888
rect 755 7386 761 7406
rect 781 7386 800 7406
rect 820 7386 839 7406
rect 859 7386 878 7406
rect 898 7386 901 7406
rect 755 6904 901 7386
rect 755 6884 761 6904
rect 781 6884 800 6904
rect 820 6884 839 6904
rect 859 6884 878 6904
rect 898 6884 901 6904
rect 755 6402 901 6884
rect 755 6382 761 6402
rect 781 6382 800 6402
rect 820 6382 839 6402
rect 859 6382 878 6402
rect 898 6382 901 6402
rect 755 5900 901 6382
rect 755 5880 761 5900
rect 781 5880 800 5900
rect 820 5880 839 5900
rect 859 5880 878 5900
rect 898 5880 901 5900
rect 755 5398 901 5880
rect 755 5378 761 5398
rect 781 5378 800 5398
rect 820 5378 839 5398
rect 859 5378 878 5398
rect 898 5378 901 5398
rect 755 4896 901 5378
rect 755 4876 761 4896
rect 781 4876 800 4896
rect 820 4876 839 4896
rect 859 4876 878 4896
rect 898 4876 901 4896
rect 755 4394 901 4876
rect 755 4374 761 4394
rect 781 4374 800 4394
rect 820 4374 839 4394
rect 859 4374 878 4394
rect 898 4374 901 4394
rect 755 3892 901 4374
rect 755 3872 761 3892
rect 781 3872 800 3892
rect 820 3872 839 3892
rect 859 3872 878 3892
rect 898 3872 901 3892
rect 755 3390 901 3872
rect 755 3370 761 3390
rect 781 3370 800 3390
rect 820 3370 839 3390
rect 859 3370 878 3390
rect 898 3370 901 3390
rect 755 2888 901 3370
rect 755 2868 761 2888
rect 781 2868 800 2888
rect 820 2868 839 2888
rect 859 2868 878 2888
rect 898 2868 901 2888
rect 755 2386 901 2868
rect 755 2366 761 2386
rect 781 2366 800 2386
rect 820 2366 839 2386
rect 859 2366 878 2386
rect 898 2366 901 2386
rect 755 1884 901 2366
rect 755 1864 761 1884
rect 781 1864 800 1884
rect 820 1864 839 1884
rect 859 1864 878 1884
rect 898 1864 901 1884
rect 755 1382 901 1864
rect 755 1362 761 1382
rect 781 1362 800 1382
rect 820 1362 839 1382
rect 859 1362 878 1382
rect 898 1362 901 1382
rect 755 880 901 1362
rect 755 860 761 880
rect 781 860 800 880
rect 820 860 839 880
rect 859 860 878 880
rect 898 860 901 880
rect 755 838 901 860
rect 755 818 761 838
rect 781 818 800 838
rect 820 818 839 838
rect 859 818 878 838
rect 898 818 901 838
rect 755 153 901 818
rect 755 125 765 153
rect 793 125 812 153
rect 840 125 859 153
rect 887 125 901 153
rect 755 106 901 125
rect 755 78 765 106
rect 793 78 812 106
rect 840 78 859 106
rect 887 78 901 106
rect 755 59 901 78
rect 755 31 765 59
rect 793 31 812 59
rect 840 31 859 59
rect 887 31 901 59
rect 755 0 901 31
rect 944 9721 1090 9971
rect 944 9693 954 9721
rect 982 9693 1001 9721
rect 1029 9693 1048 9721
rect 1076 9693 1090 9721
rect 944 9674 1090 9693
rect 944 9646 954 9674
rect 982 9646 1001 9674
rect 1029 9646 1048 9674
rect 1076 9646 1090 9674
rect 944 9627 1090 9646
rect 944 9599 954 9627
rect 982 9599 1001 9627
rect 1029 9599 1048 9627
rect 1076 9599 1090 9627
rect 944 9188 1090 9599
rect 1487 9721 1633 9973
rect 1487 9693 1497 9721
rect 1525 9693 1544 9721
rect 1572 9693 1591 9721
rect 1619 9693 1633 9721
rect 1487 9674 1633 9693
rect 1487 9646 1497 9674
rect 1525 9646 1544 9674
rect 1572 9646 1591 9674
rect 1619 9646 1633 9674
rect 1487 9627 1633 9646
rect 1487 9599 1497 9627
rect 1525 9599 1544 9627
rect 1572 9599 1591 9627
rect 1619 9599 1633 9627
rect 1487 9591 1633 9599
rect 1837 9721 1983 10083
rect 1837 9693 1847 9721
rect 1875 9693 1894 9721
rect 1922 9693 1941 9721
rect 1969 9693 1983 9721
rect 1837 9674 1983 9693
rect 1837 9646 1847 9674
rect 1875 9646 1894 9674
rect 1922 9646 1941 9674
rect 1969 9646 1983 9674
rect 1837 9627 1983 9646
rect 1837 9599 1847 9627
rect 1875 9599 1894 9627
rect 1922 9599 1941 9627
rect 1969 9599 1983 9627
rect 1837 9591 1983 9599
rect 3051 10052 3197 10060
rect 3051 9973 3058 10052
rect 3189 9973 3197 10052
rect 3051 9721 3197 9973
rect 3051 9693 3061 9721
rect 3089 9693 3108 9721
rect 3136 9693 3155 9721
rect 3183 9693 3197 9721
rect 3051 9674 3197 9693
rect 3051 9646 3061 9674
rect 3089 9646 3108 9674
rect 3136 9646 3155 9674
rect 3183 9646 3197 9674
rect 3051 9627 3197 9646
rect 3051 9599 3061 9627
rect 3089 9599 3108 9627
rect 3136 9599 3155 9627
rect 3183 9599 3197 9627
rect 3051 9591 3197 9599
rect 3487 10052 3633 10060
rect 3487 9973 3494 10052
rect 3625 9973 3633 10052
rect 3487 9721 3633 9973
rect 3487 9693 3497 9721
rect 3525 9693 3544 9721
rect 3572 9693 3591 9721
rect 3619 9693 3633 9721
rect 3487 9674 3633 9693
rect 3487 9646 3497 9674
rect 3525 9646 3544 9674
rect 3572 9646 3591 9674
rect 3619 9646 3633 9674
rect 3487 9627 3633 9646
rect 3487 9599 3497 9627
rect 3525 9599 3544 9627
rect 3572 9599 3591 9627
rect 3619 9599 3633 9627
rect 3487 9591 3633 9599
rect 3837 9721 3983 10083
rect 3837 9693 3847 9721
rect 3875 9693 3894 9721
rect 3922 9693 3941 9721
rect 3969 9693 3983 9721
rect 3837 9674 3983 9693
rect 3837 9646 3847 9674
rect 3875 9646 3894 9674
rect 3922 9646 3941 9674
rect 3969 9646 3983 9674
rect 3837 9627 3983 9646
rect 3837 9599 3847 9627
rect 3875 9599 3894 9627
rect 3922 9599 3941 9627
rect 3969 9599 3983 9627
rect 3837 9591 3983 9599
rect 5051 10052 5197 10060
rect 5051 9973 5058 10052
rect 5189 9973 5197 10052
rect 5051 9721 5197 9973
rect 5051 9693 5061 9721
rect 5089 9693 5108 9721
rect 5136 9693 5155 9721
rect 5183 9693 5197 9721
rect 5051 9674 5197 9693
rect 5051 9646 5061 9674
rect 5089 9646 5108 9674
rect 5136 9646 5155 9674
rect 5183 9646 5197 9674
rect 5051 9627 5197 9646
rect 5051 9599 5061 9627
rect 5089 9599 5108 9627
rect 5136 9599 5155 9627
rect 5183 9599 5197 9627
rect 5051 9591 5197 9599
rect 5487 10052 5633 10060
rect 5487 9973 5494 10052
rect 5625 9973 5633 10052
rect 5487 9721 5633 9973
rect 5487 9693 5497 9721
rect 5525 9693 5544 9721
rect 5572 9693 5591 9721
rect 5619 9693 5633 9721
rect 5487 9674 5633 9693
rect 5487 9646 5497 9674
rect 5525 9646 5544 9674
rect 5572 9646 5591 9674
rect 5619 9646 5633 9674
rect 5487 9627 5633 9646
rect 5487 9599 5497 9627
rect 5525 9599 5544 9627
rect 5572 9599 5591 9627
rect 5619 9599 5633 9627
rect 5487 9591 5633 9599
rect 5837 9721 5983 10083
rect 5837 9693 5847 9721
rect 5875 9693 5894 9721
rect 5922 9693 5941 9721
rect 5969 9693 5983 9721
rect 5837 9674 5983 9693
rect 5837 9646 5847 9674
rect 5875 9646 5894 9674
rect 5922 9646 5941 9674
rect 5969 9646 5983 9674
rect 5837 9627 5983 9646
rect 5837 9599 5847 9627
rect 5875 9599 5894 9627
rect 5922 9599 5941 9627
rect 5969 9599 5983 9627
rect 5837 9591 5983 9599
rect 7051 10052 7197 10060
rect 7051 9973 7058 10052
rect 7189 9973 7197 10052
rect 7051 9721 7197 9973
rect 7051 9693 7061 9721
rect 7089 9693 7108 9721
rect 7136 9693 7155 9721
rect 7183 9693 7197 9721
rect 7051 9674 7197 9693
rect 7051 9646 7061 9674
rect 7089 9646 7108 9674
rect 7136 9646 7155 9674
rect 7183 9646 7197 9674
rect 7051 9627 7197 9646
rect 7051 9599 7061 9627
rect 7089 9599 7108 9627
rect 7136 9599 7155 9627
rect 7183 9599 7197 9627
rect 7051 9591 7197 9599
rect 7487 10052 7633 10060
rect 7487 9973 7494 10052
rect 7625 9973 7633 10052
rect 7487 9721 7633 9973
rect 7487 9693 7497 9721
rect 7525 9693 7544 9721
rect 7572 9693 7591 9721
rect 7619 9693 7633 9721
rect 7487 9674 7633 9693
rect 7487 9646 7497 9674
rect 7525 9646 7544 9674
rect 7572 9646 7591 9674
rect 7619 9646 7633 9674
rect 7487 9627 7633 9646
rect 7487 9599 7497 9627
rect 7525 9599 7544 9627
rect 7572 9599 7591 9627
rect 7619 9599 7633 9627
rect 7487 9591 7633 9599
rect 7837 9721 7983 10083
rect 7837 9693 7847 9721
rect 7875 9693 7894 9721
rect 7922 9693 7941 9721
rect 7969 9693 7983 9721
rect 7837 9674 7983 9693
rect 7837 9646 7847 9674
rect 7875 9646 7894 9674
rect 7922 9646 7941 9674
rect 7969 9646 7983 9674
rect 7837 9627 7983 9646
rect 7837 9599 7847 9627
rect 7875 9599 7894 9627
rect 7922 9599 7941 9627
rect 7969 9599 7983 9627
rect 7837 9591 7983 9599
rect 9051 10052 9197 10060
rect 9051 9973 9058 10052
rect 9189 9973 9197 10052
rect 9051 9721 9197 9973
rect 9051 9693 9061 9721
rect 9089 9693 9108 9721
rect 9136 9693 9155 9721
rect 9183 9693 9197 9721
rect 9051 9674 9197 9693
rect 9051 9646 9061 9674
rect 9089 9646 9108 9674
rect 9136 9646 9155 9674
rect 9183 9646 9197 9674
rect 9051 9627 9197 9646
rect 9051 9599 9061 9627
rect 9089 9599 9108 9627
rect 9136 9599 9155 9627
rect 9183 9599 9197 9627
rect 9051 9591 9197 9599
rect 9487 10052 9633 10060
rect 9487 9973 9494 10052
rect 9625 9973 9633 10052
rect 9487 9721 9633 9973
rect 9487 9693 9497 9721
rect 9525 9693 9544 9721
rect 9572 9693 9591 9721
rect 9619 9693 9633 9721
rect 9487 9674 9633 9693
rect 9487 9646 9497 9674
rect 9525 9646 9544 9674
rect 9572 9646 9591 9674
rect 9619 9646 9633 9674
rect 9487 9627 9633 9646
rect 9487 9599 9497 9627
rect 9525 9599 9544 9627
rect 9572 9599 9591 9627
rect 9619 9599 9633 9627
rect 9487 9591 9633 9599
rect 9837 9721 9983 10083
rect 9837 9693 9847 9721
rect 9875 9693 9894 9721
rect 9922 9693 9941 9721
rect 9969 9693 9983 9721
rect 9837 9674 9983 9693
rect 9837 9646 9847 9674
rect 9875 9646 9894 9674
rect 9922 9646 9941 9674
rect 9969 9646 9983 9674
rect 9837 9627 9983 9646
rect 9837 9599 9847 9627
rect 9875 9599 9894 9627
rect 9922 9599 9941 9627
rect 9969 9599 9983 9627
rect 9837 9591 9983 9599
rect 11051 10052 11197 10060
rect 11051 9973 11058 10052
rect 11189 9973 11197 10052
rect 11051 9721 11197 9973
rect 11051 9693 11061 9721
rect 11089 9693 11108 9721
rect 11136 9693 11155 9721
rect 11183 9693 11197 9721
rect 11051 9674 11197 9693
rect 11051 9646 11061 9674
rect 11089 9646 11108 9674
rect 11136 9646 11155 9674
rect 11183 9646 11197 9674
rect 11051 9627 11197 9646
rect 11051 9599 11061 9627
rect 11089 9599 11108 9627
rect 11136 9599 11155 9627
rect 11183 9599 11197 9627
rect 11051 9591 11197 9599
rect 11487 10052 11633 10060
rect 11487 9973 11494 10052
rect 11625 9973 11633 10052
rect 11487 9721 11633 9973
rect 11487 9693 11497 9721
rect 11525 9693 11544 9721
rect 11572 9693 11591 9721
rect 11619 9693 11633 9721
rect 11487 9674 11633 9693
rect 11487 9646 11497 9674
rect 11525 9646 11544 9674
rect 11572 9646 11591 9674
rect 11619 9646 11633 9674
rect 11487 9627 11633 9646
rect 11487 9599 11497 9627
rect 11525 9599 11544 9627
rect 11572 9599 11591 9627
rect 11619 9599 11633 9627
rect 11487 9591 11633 9599
rect 11837 9721 11983 10083
rect 11837 9693 11847 9721
rect 11875 9693 11894 9721
rect 11922 9693 11941 9721
rect 11969 9693 11983 9721
rect 11837 9674 11983 9693
rect 11837 9646 11847 9674
rect 11875 9646 11894 9674
rect 11922 9646 11941 9674
rect 11969 9646 11983 9674
rect 11837 9627 11983 9646
rect 11837 9599 11847 9627
rect 11875 9599 11894 9627
rect 11922 9599 11941 9627
rect 11969 9599 11983 9627
rect 11837 9591 11983 9599
rect 13051 10052 13197 10060
rect 13051 9973 13058 10052
rect 13189 9973 13197 10052
rect 13051 9721 13197 9973
rect 13051 9693 13061 9721
rect 13089 9693 13108 9721
rect 13136 9693 13155 9721
rect 13183 9693 13197 9721
rect 13051 9674 13197 9693
rect 13051 9646 13061 9674
rect 13089 9646 13108 9674
rect 13136 9646 13155 9674
rect 13183 9646 13197 9674
rect 13051 9627 13197 9646
rect 13051 9599 13061 9627
rect 13089 9599 13108 9627
rect 13136 9599 13155 9627
rect 13183 9599 13197 9627
rect 13051 9591 13197 9599
rect 13487 10052 13633 10060
rect 13487 9973 13494 10052
rect 13625 9973 13633 10052
rect 13487 9721 13633 9973
rect 13487 9693 13497 9721
rect 13525 9693 13544 9721
rect 13572 9693 13591 9721
rect 13619 9693 13633 9721
rect 13487 9674 13633 9693
rect 13487 9646 13497 9674
rect 13525 9646 13544 9674
rect 13572 9646 13591 9674
rect 13619 9646 13633 9674
rect 13487 9627 13633 9646
rect 13487 9599 13497 9627
rect 13525 9599 13544 9627
rect 13572 9599 13591 9627
rect 13619 9599 13633 9627
rect 13487 9591 13633 9599
rect 13837 9721 13983 10083
rect 13837 9693 13847 9721
rect 13875 9693 13894 9721
rect 13922 9693 13941 9721
rect 13969 9693 13983 9721
rect 13837 9674 13983 9693
rect 13837 9646 13847 9674
rect 13875 9646 13894 9674
rect 13922 9646 13941 9674
rect 13969 9646 13983 9674
rect 13837 9627 13983 9646
rect 13837 9599 13847 9627
rect 13875 9599 13894 9627
rect 13922 9599 13941 9627
rect 13969 9599 13983 9627
rect 13837 9591 13983 9599
rect 15051 10052 15197 10060
rect 15051 9973 15058 10052
rect 15189 9973 15197 10052
rect 15051 9721 15197 9973
rect 15051 9693 15061 9721
rect 15089 9693 15108 9721
rect 15136 9693 15155 9721
rect 15183 9693 15197 9721
rect 15051 9674 15197 9693
rect 15051 9646 15061 9674
rect 15089 9646 15108 9674
rect 15136 9646 15155 9674
rect 15183 9646 15197 9674
rect 15051 9627 15197 9646
rect 15051 9599 15061 9627
rect 15089 9599 15108 9627
rect 15136 9599 15155 9627
rect 15183 9599 15197 9627
rect 15051 9591 15197 9599
rect 15487 10052 15633 10060
rect 15487 9973 15494 10052
rect 15625 9973 15633 10052
rect 15487 9721 15633 9973
rect 15487 9693 15497 9721
rect 15525 9693 15544 9721
rect 15572 9693 15591 9721
rect 15619 9693 15633 9721
rect 15487 9674 15633 9693
rect 15487 9646 15497 9674
rect 15525 9646 15544 9674
rect 15572 9646 15591 9674
rect 15619 9646 15633 9674
rect 15487 9627 15633 9646
rect 15487 9599 15497 9627
rect 15525 9599 15544 9627
rect 15572 9599 15591 9627
rect 15619 9599 15633 9627
rect 15487 9591 15633 9599
rect 15837 9721 15983 10083
rect 15837 9693 15847 9721
rect 15875 9693 15894 9721
rect 15922 9693 15941 9721
rect 15969 9693 15983 9721
rect 15837 9674 15983 9693
rect 15837 9646 15847 9674
rect 15875 9646 15894 9674
rect 15922 9646 15941 9674
rect 15969 9646 15983 9674
rect 15837 9627 15983 9646
rect 15837 9599 15847 9627
rect 15875 9599 15894 9627
rect 15922 9599 15941 9627
rect 15969 9599 15983 9627
rect 15837 9591 15983 9599
rect 17051 10052 17197 10060
rect 17051 9973 17058 10052
rect 17189 9973 17197 10052
rect 17051 9721 17197 9973
rect 17051 9693 17061 9721
rect 17089 9693 17108 9721
rect 17136 9693 17155 9721
rect 17183 9693 17197 9721
rect 17051 9674 17197 9693
rect 17051 9646 17061 9674
rect 17089 9646 17108 9674
rect 17136 9646 17155 9674
rect 17183 9646 17197 9674
rect 17051 9627 17197 9646
rect 17051 9599 17061 9627
rect 17089 9599 17108 9627
rect 17136 9599 17155 9627
rect 17183 9599 17197 9627
rect 17051 9591 17197 9599
rect 17487 10052 17633 10060
rect 17487 9973 17494 10052
rect 17625 9973 17633 10052
rect 17487 9721 17633 9973
rect 17487 9693 17497 9721
rect 17525 9693 17544 9721
rect 17572 9693 17591 9721
rect 17619 9693 17633 9721
rect 17487 9674 17633 9693
rect 17487 9646 17497 9674
rect 17525 9646 17544 9674
rect 17572 9646 17591 9674
rect 17619 9646 17633 9674
rect 17487 9627 17633 9646
rect 17487 9599 17497 9627
rect 17525 9599 17544 9627
rect 17572 9599 17591 9627
rect 17619 9599 17633 9627
rect 17487 9591 17633 9599
rect 17837 9721 17983 10083
rect 19051 10052 19197 10060
rect 19051 9990 19058 10052
rect 19189 9990 19197 10052
rect 17837 9693 17847 9721
rect 17875 9693 17894 9721
rect 17922 9693 17941 9721
rect 17969 9693 17983 9721
rect 17837 9674 17983 9693
rect 17837 9646 17847 9674
rect 17875 9646 17894 9674
rect 17922 9646 17941 9674
rect 17969 9646 17983 9674
rect 17837 9627 17983 9646
rect 17837 9599 17847 9627
rect 17875 9599 17894 9627
rect 17922 9599 17941 9627
rect 17969 9599 17983 9627
rect 17837 9591 17983 9599
rect 18362 9716 18510 9966
rect 18362 9688 18376 9716
rect 18404 9688 18423 9716
rect 18451 9688 18470 9716
rect 18498 9688 18510 9716
rect 18362 9669 18510 9688
rect 18362 9641 18376 9669
rect 18404 9641 18423 9669
rect 18451 9641 18470 9669
rect 18498 9641 18510 9669
rect 18362 9622 18510 9641
rect 18362 9594 18376 9622
rect 18404 9594 18423 9622
rect 18451 9594 18470 9622
rect 18498 9594 18510 9622
rect 944 9168 950 9188
rect 970 9168 989 9188
rect 1009 9168 1028 9188
rect 1048 9168 1067 9188
rect 1087 9168 1090 9188
rect 944 9083 1090 9168
rect 944 9063 950 9083
rect 970 9063 989 9083
rect 1009 9063 1028 9083
rect 1048 9063 1067 9083
rect 1087 9063 1090 9083
rect 944 8581 1090 9063
rect 944 8561 950 8581
rect 970 8561 989 8581
rect 1009 8561 1028 8581
rect 1048 8561 1067 8581
rect 1087 8561 1090 8581
rect 944 8079 1090 8561
rect 944 8059 950 8079
rect 970 8059 989 8079
rect 1009 8059 1028 8079
rect 1048 8059 1067 8079
rect 1087 8059 1090 8079
rect 944 7577 1090 8059
rect 944 7557 950 7577
rect 970 7557 989 7577
rect 1009 7557 1028 7577
rect 1048 7557 1067 7577
rect 1087 7557 1090 7577
rect 944 7075 1090 7557
rect 944 7055 950 7075
rect 970 7055 989 7075
rect 1009 7055 1028 7075
rect 1048 7055 1067 7075
rect 1087 7055 1090 7075
rect 944 6573 1090 7055
rect 944 6553 950 6573
rect 970 6553 989 6573
rect 1009 6553 1028 6573
rect 1048 6553 1067 6573
rect 1087 6553 1090 6573
rect 944 6071 1090 6553
rect 944 6051 950 6071
rect 970 6051 989 6071
rect 1009 6051 1028 6071
rect 1048 6051 1067 6071
rect 1087 6051 1090 6071
rect 944 5569 1090 6051
rect 944 5549 950 5569
rect 970 5549 989 5569
rect 1009 5549 1028 5569
rect 1048 5549 1067 5569
rect 1087 5549 1090 5569
rect 944 5067 1090 5549
rect 944 5047 950 5067
rect 970 5047 989 5067
rect 1009 5047 1028 5067
rect 1048 5047 1067 5067
rect 1087 5047 1090 5067
rect 944 4565 1090 5047
rect 944 4545 950 4565
rect 970 4545 989 4565
rect 1009 4545 1028 4565
rect 1048 4545 1067 4565
rect 1087 4545 1090 4565
rect 944 4063 1090 4545
rect 944 4043 950 4063
rect 970 4043 989 4063
rect 1009 4043 1028 4063
rect 1048 4043 1067 4063
rect 1087 4043 1090 4063
rect 944 3561 1090 4043
rect 944 3541 950 3561
rect 970 3541 989 3561
rect 1009 3541 1028 3561
rect 1048 3541 1067 3561
rect 1087 3541 1090 3561
rect 944 3059 1090 3541
rect 944 3039 950 3059
rect 970 3039 989 3059
rect 1009 3039 1028 3059
rect 1048 3039 1067 3059
rect 1087 3039 1090 3059
rect 944 2557 1090 3039
rect 944 2537 950 2557
rect 970 2537 989 2557
rect 1009 2537 1028 2557
rect 1048 2537 1067 2557
rect 1087 2537 1090 2557
rect 944 2055 1090 2537
rect 944 2035 950 2055
rect 970 2035 989 2055
rect 1009 2035 1028 2055
rect 1048 2035 1067 2055
rect 1087 2035 1090 2055
rect 944 1553 1090 2035
rect 944 1533 950 1553
rect 970 1533 989 1553
rect 1009 1533 1028 1553
rect 1048 1533 1067 1553
rect 1087 1533 1090 1553
rect 944 1051 1090 1533
rect 18362 9322 18510 9594
rect 18362 9294 18377 9322
rect 18405 9294 18424 9322
rect 18452 9294 18471 9322
rect 18499 9294 18510 9322
rect 18362 9275 18510 9294
rect 18362 9247 18377 9275
rect 18405 9247 18424 9275
rect 18452 9247 18471 9275
rect 18499 9247 18510 9275
rect 18362 9228 18510 9247
rect 18362 9200 18377 9228
rect 18405 9200 18424 9228
rect 18452 9200 18471 9228
rect 18499 9200 18510 9228
rect 18362 9083 18510 9200
rect 18362 9063 18365 9083
rect 18385 9063 18404 9083
rect 18424 9063 18443 9083
rect 18463 9063 18482 9083
rect 18502 9063 18510 9083
rect 18362 8581 18510 9063
rect 18362 8561 18365 8581
rect 18385 8561 18404 8581
rect 18424 8561 18443 8581
rect 18463 8561 18482 8581
rect 18502 8561 18510 8581
rect 18362 8314 18510 8561
rect 18362 8286 18376 8314
rect 18404 8286 18423 8314
rect 18451 8286 18470 8314
rect 18498 8286 18510 8314
rect 18362 8267 18510 8286
rect 18362 8239 18376 8267
rect 18404 8239 18423 8267
rect 18451 8239 18470 8267
rect 18498 8239 18510 8267
rect 18362 8220 18510 8239
rect 18362 8192 18376 8220
rect 18404 8192 18423 8220
rect 18451 8192 18470 8220
rect 18498 8192 18510 8220
rect 18362 8079 18510 8192
rect 18362 8059 18365 8079
rect 18385 8059 18404 8079
rect 18424 8059 18443 8079
rect 18463 8059 18482 8079
rect 18502 8059 18510 8079
rect 18362 7577 18510 8059
rect 18362 7557 18365 7577
rect 18385 7557 18404 7577
rect 18424 7557 18443 7577
rect 18463 7557 18482 7577
rect 18502 7557 18510 7577
rect 18362 7314 18510 7557
rect 18362 7286 18376 7314
rect 18404 7286 18423 7314
rect 18451 7286 18470 7314
rect 18498 7286 18510 7314
rect 18362 7267 18510 7286
rect 18362 7239 18376 7267
rect 18404 7239 18423 7267
rect 18451 7239 18470 7267
rect 18498 7239 18510 7267
rect 18362 7220 18510 7239
rect 18362 7192 18376 7220
rect 18404 7192 18423 7220
rect 18451 7192 18470 7220
rect 18498 7192 18510 7220
rect 18362 7075 18510 7192
rect 18362 7055 18365 7075
rect 18385 7055 18404 7075
rect 18424 7055 18443 7075
rect 18463 7055 18482 7075
rect 18502 7055 18510 7075
rect 18362 6573 18510 7055
rect 18550 9935 18697 9966
rect 18550 9907 18565 9935
rect 18593 9907 18612 9935
rect 18640 9907 18659 9935
rect 18687 9907 18697 9935
rect 18550 9888 18697 9907
rect 18550 9860 18565 9888
rect 18593 9860 18612 9888
rect 18640 9860 18659 9888
rect 18687 9860 18697 9888
rect 18550 9841 18697 9860
rect 18550 9813 18565 9841
rect 18593 9813 18612 9841
rect 18640 9813 18659 9841
rect 18687 9813 18697 9841
rect 18550 9493 18697 9813
rect 19051 9950 19197 9990
rect 18827 9567 19034 9731
rect 19051 9721 19272 9950
rect 19051 9693 19061 9721
rect 19089 9693 19108 9721
rect 19136 9693 19155 9721
rect 19183 9693 19272 9721
rect 19051 9674 19272 9693
rect 19051 9646 19061 9674
rect 19089 9646 19108 9674
rect 19136 9646 19155 9674
rect 19183 9646 19272 9674
rect 19051 9627 19272 9646
rect 19051 9599 19061 9627
rect 19089 9599 19108 9627
rect 19136 9599 19155 9627
rect 19183 9599 19272 9627
rect 19051 9591 19272 9599
rect 18827 9550 18845 9567
rect 19020 9550 19034 9567
rect 18827 9527 19034 9550
rect 18827 9510 18845 9527
rect 19020 9510 19034 9527
rect 18550 9414 18698 9493
rect 18550 9394 18554 9414
rect 18574 9394 18593 9414
rect 18613 9394 18632 9414
rect 18652 9394 18671 9414
rect 18691 9394 18698 9414
rect 18550 9331 18698 9394
rect 18550 9190 18699 9331
rect 18550 8912 18698 9190
rect 18550 8892 18554 8912
rect 18574 8892 18593 8912
rect 18613 8892 18632 8912
rect 18652 8892 18671 8912
rect 18691 8892 18698 8912
rect 18550 8830 18698 8892
rect 18550 8802 18565 8830
rect 18593 8802 18612 8830
rect 18640 8802 18659 8830
rect 18687 8802 18698 8830
rect 18550 8783 18698 8802
rect 18550 8755 18565 8783
rect 18593 8755 18612 8783
rect 18640 8755 18659 8783
rect 18687 8755 18698 8783
rect 18550 8736 18698 8755
rect 18550 8708 18565 8736
rect 18593 8708 18612 8736
rect 18640 8708 18659 8736
rect 18687 8708 18698 8736
rect 18550 8410 18698 8708
rect 18550 8390 18554 8410
rect 18574 8390 18593 8410
rect 18613 8390 18632 8410
rect 18652 8390 18671 8410
rect 18691 8390 18698 8410
rect 18550 7908 18698 8390
rect 18550 7888 18554 7908
rect 18574 7888 18593 7908
rect 18613 7888 18632 7908
rect 18652 7888 18671 7908
rect 18691 7888 18698 7908
rect 18550 7776 18698 7888
rect 18550 7748 18565 7776
rect 18593 7748 18612 7776
rect 18640 7748 18659 7776
rect 18687 7748 18698 7776
rect 18550 7729 18698 7748
rect 18550 7701 18565 7729
rect 18593 7701 18612 7729
rect 18640 7701 18659 7729
rect 18687 7701 18698 7729
rect 18550 7682 18698 7701
rect 18550 7654 18565 7682
rect 18593 7654 18612 7682
rect 18640 7654 18659 7682
rect 18687 7654 18698 7682
rect 18550 7406 18698 7654
rect 18550 7386 18554 7406
rect 18574 7386 18593 7406
rect 18613 7386 18632 7406
rect 18652 7386 18671 7406
rect 18691 7386 18698 7406
rect 18550 6904 18698 7386
rect 18550 6884 18554 6904
rect 18574 6884 18593 6904
rect 18613 6884 18632 6904
rect 18652 6884 18671 6904
rect 18691 6884 18698 6904
rect 18550 6818 18698 6884
rect 18549 6811 18698 6818
rect 18549 6783 18564 6811
rect 18592 6783 18611 6811
rect 18639 6783 18658 6811
rect 18686 6783 18698 6811
rect 18549 6764 18698 6783
rect 18549 6736 18564 6764
rect 18592 6736 18611 6764
rect 18639 6736 18658 6764
rect 18686 6736 18698 6764
rect 18549 6717 18698 6736
rect 18549 6689 18564 6717
rect 18592 6689 18611 6717
rect 18639 6689 18658 6717
rect 18686 6689 18698 6717
rect 18549 6678 18698 6689
rect 18362 6553 18365 6573
rect 18385 6553 18404 6573
rect 18424 6553 18443 6573
rect 18463 6553 18482 6573
rect 18502 6553 18510 6573
rect 18362 6352 18510 6553
rect 18362 6324 18377 6352
rect 18405 6324 18424 6352
rect 18452 6324 18471 6352
rect 18499 6324 18510 6352
rect 18362 6305 18510 6324
rect 18362 6277 18377 6305
rect 18405 6277 18424 6305
rect 18452 6277 18471 6305
rect 18499 6277 18510 6305
rect 18362 6258 18510 6277
rect 18362 6230 18377 6258
rect 18405 6230 18424 6258
rect 18452 6230 18471 6258
rect 18499 6230 18510 6258
rect 18362 6071 18510 6230
rect 18362 6051 18365 6071
rect 18385 6051 18404 6071
rect 18424 6051 18443 6071
rect 18463 6051 18482 6071
rect 18502 6051 18510 6071
rect 18362 5569 18510 6051
rect 18362 5549 18365 5569
rect 18385 5549 18404 5569
rect 18424 5549 18443 5569
rect 18463 5549 18482 5569
rect 18502 5549 18510 5569
rect 18362 5289 18510 5549
rect 18362 5261 18376 5289
rect 18404 5261 18423 5289
rect 18451 5261 18470 5289
rect 18498 5261 18510 5289
rect 18362 5242 18510 5261
rect 18362 5214 18376 5242
rect 18404 5214 18423 5242
rect 18451 5214 18470 5242
rect 18498 5214 18510 5242
rect 18362 5195 18510 5214
rect 18362 5167 18376 5195
rect 18404 5167 18423 5195
rect 18451 5167 18470 5195
rect 18498 5167 18510 5195
rect 18362 5067 18510 5167
rect 18362 5047 18365 5067
rect 18385 5047 18404 5067
rect 18424 5047 18443 5067
rect 18463 5047 18482 5067
rect 18502 5047 18510 5067
rect 18362 4565 18510 5047
rect 18362 4545 18365 4565
rect 18385 4545 18404 4565
rect 18424 4545 18443 4565
rect 18463 4545 18482 4565
rect 18502 4545 18510 4565
rect 18362 4301 18510 4545
rect 18362 4273 18377 4301
rect 18405 4273 18424 4301
rect 18452 4273 18471 4301
rect 18499 4273 18510 4301
rect 18362 4254 18510 4273
rect 18362 4226 18377 4254
rect 18405 4226 18424 4254
rect 18452 4226 18471 4254
rect 18499 4226 18510 4254
rect 18362 4207 18510 4226
rect 18362 4179 18377 4207
rect 18405 4179 18424 4207
rect 18452 4179 18471 4207
rect 18499 4179 18510 4207
rect 18362 4063 18510 4179
rect 18362 4043 18365 4063
rect 18385 4043 18404 4063
rect 18424 4043 18443 4063
rect 18463 4043 18482 4063
rect 18502 4043 18510 4063
rect 18362 3561 18510 4043
rect 18550 6402 18698 6678
rect 18550 6382 18554 6402
rect 18574 6382 18593 6402
rect 18613 6382 18632 6402
rect 18652 6382 18671 6402
rect 18691 6382 18698 6402
rect 18550 6361 18698 6382
rect 18740 9118 18808 9493
rect 18740 9098 18743 9118
rect 18763 9098 18782 9118
rect 18802 9098 18808 9118
rect 18740 8616 18808 9098
rect 18740 8596 18743 8616
rect 18763 8596 18782 8616
rect 18802 8596 18808 8616
rect 18740 8114 18808 8596
rect 18740 8094 18743 8114
rect 18763 8094 18782 8114
rect 18802 8094 18808 8114
rect 18740 7612 18808 8094
rect 18740 7592 18743 7612
rect 18763 7592 18782 7612
rect 18802 7592 18808 7612
rect 18740 7110 18808 7592
rect 18740 7090 18743 7110
rect 18763 7090 18782 7110
rect 18802 7090 18808 7110
rect 18740 6608 18808 7090
rect 18740 6588 18743 6608
rect 18763 6588 18782 6608
rect 18802 6588 18808 6608
rect 18550 6220 18699 6361
rect 18550 5900 18698 6220
rect 18550 5880 18554 5900
rect 18574 5880 18593 5900
rect 18613 5880 18632 5900
rect 18652 5880 18671 5900
rect 18691 5880 18698 5900
rect 18550 5803 18698 5880
rect 18550 5775 18565 5803
rect 18593 5775 18612 5803
rect 18640 5775 18659 5803
rect 18687 5775 18698 5803
rect 18550 5756 18698 5775
rect 18550 5728 18565 5756
rect 18593 5728 18612 5756
rect 18640 5728 18659 5756
rect 18687 5728 18698 5756
rect 18550 5709 18698 5728
rect 18550 5681 18565 5709
rect 18593 5681 18612 5709
rect 18640 5681 18659 5709
rect 18687 5681 18698 5709
rect 18550 5398 18698 5681
rect 18550 5378 18554 5398
rect 18574 5378 18593 5398
rect 18613 5378 18632 5398
rect 18652 5378 18671 5398
rect 18691 5378 18698 5398
rect 18550 4896 18698 5378
rect 18550 4876 18554 4896
rect 18574 4876 18593 4896
rect 18613 4876 18632 4896
rect 18652 4876 18671 4896
rect 18691 4876 18698 4896
rect 18550 4802 18698 4876
rect 18550 4774 18565 4802
rect 18593 4774 18612 4802
rect 18640 4774 18659 4802
rect 18687 4774 18698 4802
rect 18550 4755 18698 4774
rect 18550 4727 18565 4755
rect 18593 4727 18612 4755
rect 18640 4727 18659 4755
rect 18687 4727 18698 4755
rect 18550 4708 18698 4727
rect 18550 4680 18565 4708
rect 18593 4680 18612 4708
rect 18640 4680 18659 4708
rect 18687 4680 18698 4708
rect 18550 4394 18698 4680
rect 18550 4374 18554 4394
rect 18574 4374 18593 4394
rect 18613 4374 18632 4394
rect 18652 4374 18671 4394
rect 18691 4374 18698 4394
rect 18550 4310 18698 4374
rect 18740 6106 18808 6588
rect 18740 6086 18743 6106
rect 18763 6086 18782 6106
rect 18802 6086 18808 6106
rect 18740 5604 18808 6086
rect 18740 5584 18743 5604
rect 18763 5584 18782 5604
rect 18802 5584 18808 5604
rect 18740 5102 18808 5584
rect 18740 5082 18743 5102
rect 18763 5082 18782 5102
rect 18802 5082 18808 5102
rect 18740 4600 18808 5082
rect 18740 4580 18743 4600
rect 18763 4580 18782 4600
rect 18802 4580 18808 4600
rect 18550 4169 18699 4310
rect 18550 3892 18698 4169
rect 18550 3872 18554 3892
rect 18574 3872 18593 3892
rect 18613 3872 18632 3892
rect 18652 3872 18671 3892
rect 18691 3872 18698 3892
rect 18550 3810 18698 3872
rect 18549 3803 18698 3810
rect 18549 3775 18564 3803
rect 18592 3775 18611 3803
rect 18639 3775 18658 3803
rect 18686 3775 18698 3803
rect 18549 3756 18698 3775
rect 18549 3728 18564 3756
rect 18592 3728 18611 3756
rect 18639 3728 18658 3756
rect 18686 3728 18698 3756
rect 18549 3709 18698 3728
rect 18549 3681 18564 3709
rect 18592 3681 18611 3709
rect 18639 3681 18658 3709
rect 18686 3681 18698 3709
rect 18549 3670 18698 3681
rect 18362 3541 18365 3561
rect 18385 3541 18404 3561
rect 18424 3541 18443 3561
rect 18463 3541 18482 3561
rect 18502 3541 18510 3561
rect 18362 3279 18510 3541
rect 18362 3251 18377 3279
rect 18405 3251 18424 3279
rect 18452 3251 18471 3279
rect 18499 3251 18510 3279
rect 18362 3232 18510 3251
rect 18362 3204 18377 3232
rect 18405 3204 18424 3232
rect 18452 3204 18471 3232
rect 18499 3204 18510 3232
rect 18362 3185 18510 3204
rect 18362 3157 18377 3185
rect 18405 3157 18424 3185
rect 18452 3157 18471 3185
rect 18499 3157 18510 3185
rect 18362 3059 18510 3157
rect 18362 3039 18365 3059
rect 18385 3039 18404 3059
rect 18424 3039 18443 3059
rect 18463 3039 18482 3059
rect 18502 3039 18510 3059
rect 18362 2557 18510 3039
rect 18362 2537 18365 2557
rect 18385 2537 18404 2557
rect 18424 2537 18443 2557
rect 18463 2537 18482 2557
rect 18502 2537 18510 2557
rect 18362 2282 18510 2537
rect 18362 2254 18377 2282
rect 18405 2254 18424 2282
rect 18452 2254 18471 2282
rect 18499 2254 18510 2282
rect 18362 2235 18510 2254
rect 18362 2207 18377 2235
rect 18405 2207 18424 2235
rect 18452 2207 18471 2235
rect 18499 2207 18510 2235
rect 18362 2188 18510 2207
rect 18362 2160 18377 2188
rect 18405 2160 18424 2188
rect 18452 2160 18471 2188
rect 18499 2160 18510 2188
rect 18362 2055 18510 2160
rect 18362 2035 18365 2055
rect 18385 2035 18404 2055
rect 18424 2035 18443 2055
rect 18463 2035 18482 2055
rect 18502 2035 18510 2055
rect 18362 1553 18510 2035
rect 18362 1533 18365 1553
rect 18385 1533 18404 1553
rect 18424 1533 18443 1553
rect 18463 1533 18482 1553
rect 18502 1533 18510 1553
rect 18362 1291 18510 1533
rect 18550 3390 18698 3670
rect 18550 3370 18554 3390
rect 18574 3370 18593 3390
rect 18613 3370 18632 3390
rect 18652 3370 18671 3390
rect 18691 3370 18698 3390
rect 18550 3288 18698 3370
rect 18740 4098 18808 4580
rect 18740 4078 18743 4098
rect 18763 4078 18782 4098
rect 18802 4078 18808 4098
rect 18740 3596 18808 4078
rect 18740 3576 18743 3596
rect 18763 3576 18782 3596
rect 18802 3576 18808 3596
rect 18550 3147 18699 3288
rect 18550 2888 18698 3147
rect 18550 2868 18554 2888
rect 18574 2868 18593 2888
rect 18613 2868 18632 2888
rect 18652 2868 18671 2888
rect 18691 2868 18698 2888
rect 18550 2769 18698 2868
rect 18550 2741 18565 2769
rect 18593 2741 18612 2769
rect 18640 2741 18659 2769
rect 18687 2741 18698 2769
rect 18550 2722 18698 2741
rect 18550 2694 18565 2722
rect 18593 2694 18612 2722
rect 18640 2694 18659 2722
rect 18687 2694 18698 2722
rect 18550 2675 18698 2694
rect 18550 2647 18565 2675
rect 18593 2647 18612 2675
rect 18640 2647 18659 2675
rect 18687 2647 18698 2675
rect 18550 2386 18698 2647
rect 18550 2366 18554 2386
rect 18574 2366 18593 2386
rect 18613 2366 18632 2386
rect 18652 2366 18671 2386
rect 18691 2366 18698 2386
rect 18550 2290 18698 2366
rect 18740 3094 18808 3576
rect 18740 3074 18743 3094
rect 18763 3074 18782 3094
rect 18802 3074 18808 3094
rect 18740 2592 18808 3074
rect 18740 2572 18743 2592
rect 18763 2572 18782 2592
rect 18802 2572 18808 2592
rect 18550 2149 18699 2290
rect 18550 1884 18698 2149
rect 18550 1864 18554 1884
rect 18574 1864 18593 1884
rect 18613 1864 18632 1884
rect 18652 1864 18671 1884
rect 18691 1864 18698 1884
rect 18550 1767 18698 1864
rect 18550 1739 18565 1767
rect 18593 1739 18612 1767
rect 18640 1739 18659 1767
rect 18687 1739 18698 1767
rect 18550 1720 18698 1739
rect 18550 1692 18565 1720
rect 18593 1692 18612 1720
rect 18640 1692 18659 1720
rect 18687 1692 18698 1720
rect 18550 1673 18698 1692
rect 18550 1645 18565 1673
rect 18593 1645 18612 1673
rect 18640 1645 18659 1673
rect 18687 1645 18698 1673
rect 18550 1382 18698 1645
rect 18550 1362 18554 1382
rect 18574 1362 18593 1382
rect 18613 1362 18632 1382
rect 18652 1362 18671 1382
rect 18691 1362 18698 1382
rect 18550 1291 18698 1362
rect 18361 1282 18510 1291
rect 18361 1254 18375 1282
rect 18403 1254 18422 1282
rect 18450 1254 18469 1282
rect 18497 1254 18510 1282
rect 18361 1235 18510 1254
rect 18361 1207 18375 1235
rect 18403 1207 18422 1235
rect 18450 1207 18469 1235
rect 18497 1207 18510 1235
rect 18361 1188 18510 1207
rect 18361 1160 18375 1188
rect 18403 1160 18422 1188
rect 18450 1160 18469 1188
rect 18497 1160 18510 1188
rect 18361 1150 18510 1160
rect 18549 1150 18698 1291
rect 944 1031 950 1051
rect 970 1031 989 1051
rect 1009 1031 1028 1051
rect 1048 1031 1067 1051
rect 1087 1031 1090 1051
rect 944 710 1090 1031
rect 944 690 950 710
rect 970 690 989 710
rect 1009 690 1028 710
rect 1048 690 1067 710
rect 1087 690 1090 710
rect 944 654 1090 690
rect 944 634 950 654
rect 970 634 989 654
rect 1009 634 1028 654
rect 1048 634 1067 654
rect 1087 634 1090 654
rect 944 549 1090 634
rect 944 529 950 549
rect 970 529 989 549
rect 1009 529 1028 549
rect 1048 529 1067 549
rect 1087 529 1090 549
rect 944 372 1090 529
rect 18362 1051 18510 1150
rect 18362 1031 18365 1051
rect 18385 1031 18404 1051
rect 18424 1031 18443 1051
rect 18463 1031 18482 1051
rect 18502 1031 18510 1051
rect 18362 549 18510 1031
rect 18362 529 18365 549
rect 18385 529 18404 549
rect 18424 529 18443 549
rect 18463 529 18482 549
rect 18502 529 18510 549
rect 944 344 954 372
rect 982 344 1001 372
rect 1029 344 1048 372
rect 1076 344 1090 372
rect 944 325 1090 344
rect 944 297 954 325
rect 982 297 1001 325
rect 1029 297 1048 325
rect 1076 297 1090 325
rect 944 278 1090 297
rect 944 250 954 278
rect 982 250 1001 278
rect 1029 250 1048 278
rect 1076 250 1090 278
rect 944 0 1090 250
rect 1622 165 1639 457
rect 1617 162 1639 165
rect 1617 145 1620 162
rect 1637 145 1639 162
rect 1617 141 1639 145
rect 2124 0 2141 457
rect 2626 0 2643 457
rect 3128 0 3145 457
rect 3630 0 3647 457
rect 4132 0 4149 457
rect 4634 0 4651 457
rect 5136 0 5153 457
rect 5638 0 5655 457
rect 5974 0 5991 457
rect 6140 0 6157 457
rect 6642 0 6659 457
rect 7144 0 7161 457
rect 7646 0 7663 457
rect 8148 0 8165 457
rect 8650 0 8667 457
rect 9152 0 9169 457
rect 9654 0 9671 457
rect 9990 0 10007 457
rect 10156 0 10173 457
rect 10658 0 10675 457
rect 11160 0 11177 457
rect 11662 0 11679 457
rect 12164 0 12181 457
rect 12666 0 12683 457
rect 13168 0 13185 457
rect 13670 0 13687 457
rect 14006 0 14023 457
rect 14172 0 14189 457
rect 14674 397 14691 457
rect 14274 380 14691 397
rect 14274 0 14291 380
rect 15176 362 15193 457
rect 14376 345 15193 362
rect 14376 0 14393 345
rect 14478 321 14495 322
rect 14478 0 14495 304
rect 15678 321 15695 457
rect 15678 300 15695 304
rect 14580 282 14597 283
rect 14580 0 14597 265
rect 16180 282 16197 457
rect 16180 261 16197 265
rect 14682 244 14699 245
rect 14682 0 14699 227
rect 16682 244 16699 457
rect 16682 223 16699 227
rect 14784 206 14801 207
rect 14784 0 14801 189
rect 17184 206 17201 457
rect 17433 431 17450 457
rect 17184 185 17201 189
rect 17238 414 17450 431
rect 14886 168 14903 169
rect 14886 0 14903 151
rect 17238 1 17255 414
rect 17299 393 17316 396
rect 17299 1 17316 376
rect 17469 344 17486 457
rect 17543 393 17560 457
rect 17543 372 17560 376
rect 17469 322 17613 344
rect 17596 25 17613 322
rect 17686 168 17703 457
rect 17686 147 17703 151
rect 18188 162 18205 457
rect 18362 437 18510 529
rect 18362 409 18376 437
rect 18404 409 18423 437
rect 18451 409 18470 437
rect 18498 409 18510 437
rect 18362 390 18510 409
rect 18362 362 18376 390
rect 18404 362 18423 390
rect 18451 362 18470 390
rect 18498 362 18510 390
rect 18362 343 18510 362
rect 18362 315 18376 343
rect 18404 315 18423 343
rect 18451 315 18470 343
rect 18498 315 18510 343
rect 18188 159 18209 162
rect 18188 142 18190 159
rect 18207 142 18209 159
rect 18188 139 18209 142
rect 18362 65 18510 315
rect 18550 880 18698 1150
rect 18550 860 18554 880
rect 18574 860 18593 880
rect 18613 860 18632 880
rect 18652 860 18671 880
rect 18691 860 18698 880
rect 18550 770 18698 860
rect 18550 742 18565 770
rect 18593 742 18612 770
rect 18640 742 18659 770
rect 18687 742 18698 770
rect 18550 723 18698 742
rect 18550 695 18565 723
rect 18593 695 18612 723
rect 18640 695 18659 723
rect 18687 695 18698 723
rect 18550 676 18698 695
rect 18550 648 18565 676
rect 18593 648 18612 676
rect 18640 648 18659 676
rect 18687 648 18698 676
rect 18550 219 18698 648
rect 18740 2090 18808 2572
rect 18740 2070 18743 2090
rect 18763 2070 18782 2090
rect 18802 2070 18808 2090
rect 18740 1588 18808 2070
rect 18740 1568 18743 1588
rect 18763 1568 18782 1588
rect 18802 1568 18808 1588
rect 18740 1086 18808 1568
rect 18827 9487 19034 9510
rect 18827 9470 18845 9487
rect 19020 9470 19034 9487
rect 18827 9447 19034 9470
rect 18827 9430 18845 9447
rect 19020 9430 19034 9447
rect 18827 9407 19034 9430
rect 18827 9390 18845 9407
rect 19020 9390 19034 9407
rect 18827 9367 19034 9390
rect 18827 9350 18845 9367
rect 19020 9350 19034 9367
rect 18827 9331 19034 9350
rect 18827 9327 19035 9331
rect 18827 9310 18845 9327
rect 19020 9310 19035 9327
rect 18827 9287 19035 9310
rect 18827 9270 18845 9287
rect 19020 9270 19035 9287
rect 18827 9247 19035 9270
rect 18827 9230 18845 9247
rect 19020 9230 19035 9247
rect 18827 9207 19035 9230
rect 18827 9190 18845 9207
rect 19020 9190 19035 9207
rect 18827 9167 19034 9190
rect 18827 9150 18845 9167
rect 19020 9150 19034 9167
rect 18827 9127 19034 9150
rect 18827 9110 18845 9127
rect 19020 9110 19034 9127
rect 18827 9087 19034 9110
rect 18827 9070 18845 9087
rect 19020 9070 19034 9087
rect 18827 9047 19034 9070
rect 18827 9030 18845 9047
rect 19020 9030 19034 9047
rect 18827 9007 19034 9030
rect 18827 8990 18845 9007
rect 19020 8990 19034 9007
rect 18827 8967 19034 8990
rect 18827 8950 18845 8967
rect 19020 8950 19034 8967
rect 18827 8927 19034 8950
rect 18827 8910 18845 8927
rect 19020 8910 19034 8927
rect 18827 8887 19034 8910
rect 18827 8870 18845 8887
rect 19020 8870 19034 8887
rect 18827 8847 19034 8870
rect 18827 8830 18845 8847
rect 19020 8830 19034 8847
rect 18827 8807 19034 8830
rect 18827 8790 18845 8807
rect 19020 8790 19034 8807
rect 18827 8767 19034 8790
rect 18827 8750 18845 8767
rect 19020 8750 19034 8767
rect 18827 8727 19034 8750
rect 18827 8710 18845 8727
rect 19020 8710 19034 8727
rect 18827 8687 19034 8710
rect 18827 8670 18845 8687
rect 19020 8670 19034 8687
rect 18827 8647 19034 8670
rect 18827 8630 18845 8647
rect 19020 8630 19034 8647
rect 18827 8607 19034 8630
rect 18827 8590 18845 8607
rect 19020 8590 19034 8607
rect 18827 8567 19034 8590
rect 18827 8550 18845 8567
rect 19020 8550 19034 8567
rect 18827 8527 19034 8550
rect 18827 8510 18845 8527
rect 19020 8510 19034 8527
rect 18827 8487 19034 8510
rect 18827 8470 18845 8487
rect 19020 8470 19034 8487
rect 18827 8447 19034 8470
rect 18827 8430 18845 8447
rect 19020 8430 19034 8447
rect 18827 8407 19034 8430
rect 18827 8390 18845 8407
rect 19020 8390 19034 8407
rect 18827 8367 19034 8390
rect 18827 8350 18845 8367
rect 19020 8350 19034 8367
rect 18827 8327 19034 8350
rect 18827 8310 18845 8327
rect 19020 8310 19034 8327
rect 18827 8287 19034 8310
rect 18827 8270 18845 8287
rect 19020 8270 19034 8287
rect 18827 8247 19034 8270
rect 18827 8230 18845 8247
rect 19020 8230 19034 8247
rect 18827 8207 19034 8230
rect 18827 8190 18845 8207
rect 19020 8190 19034 8207
rect 18827 8167 19034 8190
rect 18827 8150 18845 8167
rect 19020 8150 19034 8167
rect 18827 8127 19034 8150
rect 18827 8110 18845 8127
rect 19020 8110 19034 8127
rect 18827 8087 19034 8110
rect 18827 8070 18845 8087
rect 19020 8070 19034 8087
rect 18827 8047 19034 8070
rect 18827 8030 18845 8047
rect 19020 8030 19034 8047
rect 18827 8007 19034 8030
rect 18827 7990 18845 8007
rect 19020 7990 19034 8007
rect 18827 7967 19034 7990
rect 18827 7950 18845 7967
rect 19020 7950 19034 7967
rect 18827 7927 19034 7950
rect 18827 7910 18845 7927
rect 19020 7910 19034 7927
rect 18827 7887 19034 7910
rect 18827 7870 18845 7887
rect 19020 7870 19034 7887
rect 18827 7847 19034 7870
rect 18827 7830 18845 7847
rect 19020 7830 19034 7847
rect 18827 7807 19034 7830
rect 18827 7790 18845 7807
rect 19020 7790 19034 7807
rect 18827 7767 19034 7790
rect 18827 7750 18845 7767
rect 19020 7750 19034 7767
rect 18827 7727 19034 7750
rect 18827 7710 18845 7727
rect 19020 7710 19034 7727
rect 18827 7687 19034 7710
rect 18827 7670 18845 7687
rect 19020 7670 19034 7687
rect 18827 7647 19034 7670
rect 18827 7630 18845 7647
rect 19020 7630 19034 7647
rect 18827 7607 19034 7630
rect 18827 7590 18845 7607
rect 19020 7590 19034 7607
rect 18827 7567 19034 7590
rect 18827 7550 18845 7567
rect 19020 7550 19034 7567
rect 18827 7527 19034 7550
rect 18827 7510 18845 7527
rect 19020 7510 19034 7527
rect 18827 7487 19034 7510
rect 18827 7470 18845 7487
rect 19020 7470 19034 7487
rect 18827 7447 19034 7470
rect 18827 7430 18845 7447
rect 19020 7430 19034 7447
rect 18827 7407 19034 7430
rect 18827 7390 18845 7407
rect 19020 7390 19034 7407
rect 18827 7367 19034 7390
rect 18827 7350 18845 7367
rect 19020 7350 19034 7367
rect 18827 7327 19034 7350
rect 18827 7310 18845 7327
rect 19020 7310 19034 7327
rect 18827 7287 19034 7310
rect 18827 7270 18845 7287
rect 19020 7270 19034 7287
rect 18827 7247 19034 7270
rect 18827 7230 18845 7247
rect 19020 7230 19034 7247
rect 18827 7207 19034 7230
rect 18827 7190 18845 7207
rect 19020 7190 19034 7207
rect 18827 7167 19034 7190
rect 18827 7150 18845 7167
rect 19020 7150 19034 7167
rect 18827 7127 19034 7150
rect 18827 7110 18845 7127
rect 19020 7110 19034 7127
rect 18827 7087 19034 7110
rect 18827 7070 18845 7087
rect 19020 7070 19034 7087
rect 18827 7047 19034 7070
rect 18827 7030 18845 7047
rect 19020 7030 19034 7047
rect 18827 7007 19034 7030
rect 18827 6990 18845 7007
rect 19020 6990 19034 7007
rect 18827 6967 19034 6990
rect 18827 6950 18845 6967
rect 19020 6950 19034 6967
rect 18827 6927 19034 6950
rect 18827 6910 18845 6927
rect 19020 6910 19034 6927
rect 18827 6887 19034 6910
rect 18827 6870 18845 6887
rect 19020 6870 19034 6887
rect 18827 6847 19034 6870
rect 18827 6830 18845 6847
rect 19020 6830 19034 6847
rect 18827 6807 19034 6830
rect 19065 6818 19272 9591
rect 21346 9625 21762 9638
rect 21346 9419 21643 9625
rect 21749 9419 21762 9625
rect 21346 9407 21762 9419
rect 21346 8746 21762 8759
rect 21346 8540 21643 8746
rect 21749 8540 21762 8746
rect 21346 8528 21762 8540
rect 21346 7625 21762 7638
rect 21346 7419 21643 7625
rect 21749 7419 21762 7625
rect 21346 7407 21762 7419
rect 18827 6790 18845 6807
rect 19020 6790 19034 6807
rect 18827 6767 19034 6790
rect 18827 6750 18845 6767
rect 19020 6750 19034 6767
rect 18827 6727 19034 6750
rect 18827 6710 18845 6727
rect 19020 6710 19034 6727
rect 18827 6686 19034 6710
rect 18827 6669 18846 6686
rect 19021 6669 19034 6686
rect 19064 6678 19272 6818
rect 18827 6647 19034 6669
rect 18827 6630 18845 6647
rect 19020 6630 19034 6647
rect 18827 6607 19034 6630
rect 18827 6590 18845 6607
rect 19020 6590 19034 6607
rect 18827 6567 19034 6590
rect 18827 6550 18845 6567
rect 19020 6550 19034 6567
rect 18827 6527 19034 6550
rect 18827 6510 18845 6527
rect 19020 6510 19034 6527
rect 18827 6487 19034 6510
rect 18827 6470 18845 6487
rect 19020 6470 19034 6487
rect 18827 6447 19034 6470
rect 18827 6430 18845 6447
rect 19020 6430 19034 6447
rect 18827 6407 19034 6430
rect 18827 6390 18845 6407
rect 19020 6390 19034 6407
rect 18827 6367 19034 6390
rect 18827 6350 18845 6367
rect 19020 6361 19034 6367
rect 19020 6350 19035 6361
rect 18827 6327 19035 6350
rect 18827 6310 18845 6327
rect 19020 6310 19035 6327
rect 18827 6287 19035 6310
rect 18827 6270 18845 6287
rect 19020 6270 19035 6287
rect 18827 6247 19035 6270
rect 18827 6230 18845 6247
rect 19020 6230 19035 6247
rect 18827 6220 19035 6230
rect 18827 6207 19034 6220
rect 18827 6190 18845 6207
rect 19020 6190 19034 6207
rect 18827 6167 19034 6190
rect 18827 6150 18845 6167
rect 19020 6150 19034 6167
rect 18827 6127 19034 6150
rect 18827 6110 18845 6127
rect 19020 6110 19034 6127
rect 18827 6087 19034 6110
rect 18827 6070 18845 6087
rect 19020 6070 19034 6087
rect 18827 6047 19034 6070
rect 18827 6030 18845 6047
rect 19020 6030 19034 6047
rect 18827 6007 19034 6030
rect 18827 5990 18845 6007
rect 19020 5990 19034 6007
rect 18827 5967 19034 5990
rect 18827 5950 18845 5967
rect 19020 5950 19034 5967
rect 18827 5927 19034 5950
rect 18827 5910 18845 5927
rect 19020 5910 19034 5927
rect 18827 5887 19034 5910
rect 18827 5870 18845 5887
rect 19020 5870 19034 5887
rect 18827 5847 19034 5870
rect 18827 5830 18845 5847
rect 19020 5830 19034 5847
rect 18827 5806 19034 5830
rect 18827 5789 18844 5806
rect 19019 5789 19034 5806
rect 18827 5767 19034 5789
rect 18827 5750 18845 5767
rect 19020 5750 19034 5767
rect 18827 5727 19034 5750
rect 18827 5710 18845 5727
rect 19020 5710 19034 5727
rect 18827 5687 19034 5710
rect 18827 5670 18845 5687
rect 19020 5670 19034 5687
rect 18827 5647 19034 5670
rect 18827 5630 18845 5647
rect 19020 5630 19034 5647
rect 18827 5607 19034 5630
rect 18827 5590 18845 5607
rect 19020 5590 19034 5607
rect 18827 5567 19034 5590
rect 18827 5550 18845 5567
rect 19020 5550 19034 5567
rect 18827 5527 19034 5550
rect 18827 5510 18845 5527
rect 19020 5510 19034 5527
rect 18827 5487 19034 5510
rect 18827 5470 18845 5487
rect 19020 5470 19034 5487
rect 18827 5447 19034 5470
rect 18827 5430 18845 5447
rect 19020 5430 19034 5447
rect 18827 5407 19034 5430
rect 18827 5390 18845 5407
rect 19020 5390 19034 5407
rect 18827 5367 19034 5390
rect 18827 5350 18845 5367
rect 19020 5350 19034 5367
rect 18827 5327 19034 5350
rect 18827 5310 18845 5327
rect 19020 5310 19034 5327
rect 18827 5287 19034 5310
rect 18827 5270 18845 5287
rect 19020 5270 19034 5287
rect 18827 5247 19034 5270
rect 18827 5230 18845 5247
rect 19020 5230 19034 5247
rect 18827 5207 19034 5230
rect 18827 5190 18845 5207
rect 19020 5190 19034 5207
rect 18827 5167 19034 5190
rect 18827 5150 18845 5167
rect 19020 5150 19034 5167
rect 18827 5127 19034 5150
rect 18827 5110 18845 5127
rect 19020 5110 19034 5127
rect 18827 5087 19034 5110
rect 18827 5070 18845 5087
rect 19020 5070 19034 5087
rect 18827 5047 19034 5070
rect 18827 5030 18845 5047
rect 19020 5030 19034 5047
rect 18827 5007 19034 5030
rect 18827 4990 18845 5007
rect 19020 4990 19034 5007
rect 18827 4967 19034 4990
rect 18827 4950 18845 4967
rect 19020 4950 19034 4967
rect 18827 4927 19034 4950
rect 18827 4910 18845 4927
rect 19020 4910 19034 4927
rect 18827 4887 19034 4910
rect 18827 4870 18845 4887
rect 19020 4870 19034 4887
rect 18827 4847 19034 4870
rect 18827 4830 18845 4847
rect 19020 4830 19034 4847
rect 18827 4807 19034 4830
rect 18827 4790 18845 4807
rect 19020 4790 19034 4807
rect 18827 4767 19034 4790
rect 18827 4750 18845 4767
rect 19020 4750 19034 4767
rect 18827 4727 19034 4750
rect 18827 4710 18845 4727
rect 19020 4710 19034 4727
rect 18827 4687 19034 4710
rect 18827 4670 18845 4687
rect 19020 4670 19034 4687
rect 18827 4647 19034 4670
rect 18827 4630 18845 4647
rect 19020 4630 19034 4647
rect 18827 4607 19034 4630
rect 18827 4590 18845 4607
rect 19020 4590 19034 4607
rect 18827 4567 19034 4590
rect 18827 4550 18845 4567
rect 19020 4550 19034 4567
rect 18827 4527 19034 4550
rect 18827 4510 18845 4527
rect 19020 4510 19034 4527
rect 18827 4487 19034 4510
rect 18827 4470 18845 4487
rect 19020 4470 19034 4487
rect 18827 4447 19034 4470
rect 18827 4430 18845 4447
rect 19020 4430 19034 4447
rect 18827 4407 19034 4430
rect 18827 4390 18845 4407
rect 19020 4390 19034 4407
rect 18827 4367 19034 4390
rect 18827 4350 18845 4367
rect 19020 4350 19034 4367
rect 18827 4327 19034 4350
rect 18827 4310 18845 4327
rect 19020 4310 19034 4327
rect 18827 4287 19035 4310
rect 18827 4270 18845 4287
rect 19020 4270 19035 4287
rect 18827 4247 19035 4270
rect 18827 4230 18845 4247
rect 19020 4230 19035 4247
rect 18827 4207 19035 4230
rect 18827 4190 18845 4207
rect 19020 4190 19035 4207
rect 18827 4169 19035 4190
rect 18827 4167 19034 4169
rect 18827 4150 18845 4167
rect 19020 4150 19034 4167
rect 18827 4127 19034 4150
rect 18827 4110 18845 4127
rect 19020 4110 19034 4127
rect 18827 4087 19034 4110
rect 18827 4070 18845 4087
rect 19020 4070 19034 4087
rect 18827 4047 19034 4070
rect 18827 4030 18845 4047
rect 19020 4030 19034 4047
rect 18827 4007 19034 4030
rect 18827 3990 18845 4007
rect 19020 3990 19034 4007
rect 18827 3967 19034 3990
rect 18827 3950 18845 3967
rect 19020 3950 19034 3967
rect 18827 3927 19034 3950
rect 18827 3910 18845 3927
rect 19020 3910 19034 3927
rect 18827 3887 19034 3910
rect 18827 3870 18845 3887
rect 19020 3870 19034 3887
rect 18827 3847 19034 3870
rect 18827 3830 18845 3847
rect 19020 3830 19034 3847
rect 18827 3807 19034 3830
rect 19065 3810 19272 6678
rect 21346 6746 21762 6759
rect 21346 6540 21643 6746
rect 21749 6540 21762 6746
rect 21346 6528 21762 6540
rect 21346 5625 21762 5638
rect 21346 5419 21643 5625
rect 21749 5419 21762 5625
rect 21346 5407 21762 5419
rect 21346 4746 21762 4759
rect 21346 4540 21643 4746
rect 21749 4540 21762 4746
rect 21346 4528 21762 4540
rect 18827 3790 18845 3807
rect 19020 3790 19034 3807
rect 18827 3767 19034 3790
rect 18827 3750 18845 3767
rect 19020 3750 19034 3767
rect 18827 3727 19034 3750
rect 18827 3710 18845 3727
rect 19020 3710 19034 3727
rect 18827 3687 19034 3710
rect 18827 3670 18845 3687
rect 19020 3670 19034 3687
rect 19064 3670 19272 3810
rect 18827 3647 19034 3670
rect 18827 3630 18845 3647
rect 19020 3630 19034 3647
rect 18827 3607 19034 3630
rect 18827 3590 18845 3607
rect 19020 3590 19034 3607
rect 18827 3567 19034 3590
rect 18827 3550 18845 3567
rect 19020 3550 19034 3567
rect 18827 3527 19034 3550
rect 18827 3510 18845 3527
rect 19020 3510 19034 3527
rect 18827 3487 19034 3510
rect 18827 3470 18845 3487
rect 19020 3470 19034 3487
rect 18827 3447 19034 3470
rect 18827 3430 18845 3447
rect 19020 3430 19034 3447
rect 18827 3407 19034 3430
rect 18827 3390 18845 3407
rect 19020 3390 19034 3407
rect 18827 3367 19034 3390
rect 18827 3350 18845 3367
rect 19020 3350 19034 3367
rect 18827 3327 19034 3350
rect 18827 3310 18845 3327
rect 19020 3310 19034 3327
rect 18827 3288 19034 3310
rect 18827 3287 19035 3288
rect 18827 3270 18845 3287
rect 19020 3270 19035 3287
rect 18827 3247 19035 3270
rect 18827 3230 18845 3247
rect 19020 3230 19035 3247
rect 18827 3207 19035 3230
rect 18827 3190 18845 3207
rect 19020 3190 19035 3207
rect 18827 3167 19035 3190
rect 18827 3150 18845 3167
rect 19020 3150 19035 3167
rect 18827 3147 19035 3150
rect 18827 3127 19034 3147
rect 18827 3110 18845 3127
rect 19020 3110 19034 3127
rect 18827 3087 19034 3110
rect 18827 3070 18845 3087
rect 19020 3070 19034 3087
rect 18827 3047 19034 3070
rect 18827 3030 18845 3047
rect 19020 3030 19034 3047
rect 18827 3007 19034 3030
rect 18827 2990 18845 3007
rect 19020 2990 19034 3007
rect 18827 2967 19034 2990
rect 18827 2950 18845 2967
rect 19020 2950 19034 2967
rect 18827 2927 19034 2950
rect 18827 2910 18845 2927
rect 19020 2910 19034 2927
rect 18827 2887 19034 2910
rect 18827 2870 18845 2887
rect 19020 2870 19034 2887
rect 18827 2847 19034 2870
rect 18827 2830 18845 2847
rect 19020 2830 19034 2847
rect 18827 2807 19034 2830
rect 18827 2790 18845 2807
rect 19020 2790 19034 2807
rect 18827 2767 19034 2790
rect 18827 2750 18845 2767
rect 19020 2750 19034 2767
rect 18827 2724 19034 2750
rect 18827 2707 18845 2724
rect 19020 2707 19034 2724
rect 18827 2687 19034 2707
rect 18827 2670 18845 2687
rect 19020 2670 19034 2687
rect 18827 2647 19034 2670
rect 18827 2630 18845 2647
rect 19020 2630 19034 2647
rect 18827 2607 19034 2630
rect 18827 2590 18845 2607
rect 19020 2590 19034 2607
rect 18827 2567 19034 2590
rect 18827 2550 18845 2567
rect 19020 2550 19034 2567
rect 18827 2527 19034 2550
rect 18827 2510 18845 2527
rect 19020 2510 19034 2527
rect 18827 2487 19034 2510
rect 18827 2470 18845 2487
rect 19020 2470 19034 2487
rect 18827 2447 19034 2470
rect 18827 2430 18845 2447
rect 19020 2430 19034 2447
rect 18827 2407 19034 2430
rect 18827 2390 18845 2407
rect 19020 2390 19034 2407
rect 18827 2367 19034 2390
rect 18827 2350 18845 2367
rect 19020 2350 19034 2367
rect 18827 2327 19034 2350
rect 18827 2310 18845 2327
rect 19020 2310 19034 2327
rect 18827 2287 19034 2310
rect 18827 2270 18845 2287
rect 19020 2270 19034 2287
rect 18827 2247 19034 2270
rect 18827 2230 18845 2247
rect 19020 2230 19034 2247
rect 18827 2207 19034 2230
rect 18827 2190 18845 2207
rect 19020 2190 19034 2207
rect 18827 2167 19034 2190
rect 18827 2150 18845 2167
rect 19020 2150 19034 2167
rect 18827 2127 19034 2150
rect 18827 2110 18845 2127
rect 19020 2110 19034 2127
rect 18827 2087 19034 2110
rect 18827 2070 18845 2087
rect 19020 2070 19034 2087
rect 18827 2047 19034 2070
rect 18827 2030 18845 2047
rect 19020 2030 19034 2047
rect 18827 2007 19034 2030
rect 18827 1990 18845 2007
rect 19020 1990 19034 2007
rect 18827 1967 19034 1990
rect 18827 1950 18845 1967
rect 19020 1950 19034 1967
rect 18827 1927 19034 1950
rect 18827 1910 18845 1927
rect 19020 1910 19034 1927
rect 18827 1887 19034 1910
rect 18827 1870 18845 1887
rect 19020 1870 19034 1887
rect 18827 1847 19034 1870
rect 18827 1830 18845 1847
rect 19020 1830 19034 1847
rect 18827 1807 19034 1830
rect 18827 1790 18845 1807
rect 19020 1790 19034 1807
rect 18827 1767 19034 1790
rect 18827 1750 18845 1767
rect 19020 1750 19034 1767
rect 18827 1727 19034 1750
rect 18827 1710 18845 1727
rect 19020 1710 19034 1727
rect 18827 1687 19034 1710
rect 18827 1670 18845 1687
rect 19020 1670 19034 1687
rect 18827 1647 19034 1670
rect 18827 1630 18845 1647
rect 19020 1630 19034 1647
rect 18827 1607 19034 1630
rect 18827 1590 18845 1607
rect 19020 1590 19034 1607
rect 18827 1567 19034 1590
rect 18827 1550 18845 1567
rect 19020 1550 19034 1567
rect 18827 1527 19034 1550
rect 18827 1510 18845 1527
rect 19020 1510 19034 1527
rect 18827 1487 19034 1510
rect 18827 1470 18845 1487
rect 19020 1470 19034 1487
rect 18827 1447 19034 1470
rect 18827 1430 18845 1447
rect 19020 1430 19034 1447
rect 18827 1407 19034 1430
rect 18827 1390 18845 1407
rect 19020 1390 19034 1407
rect 18827 1367 19034 1390
rect 18827 1350 18845 1367
rect 19020 1350 19034 1367
rect 18827 1327 19034 1350
rect 18827 1310 18845 1327
rect 19020 1310 19034 1327
rect 18827 1291 19034 1310
rect 18826 1287 19034 1291
rect 18826 1270 18845 1287
rect 19020 1270 19034 1287
rect 18826 1247 19034 1270
rect 18826 1230 18845 1247
rect 19020 1230 19034 1247
rect 18826 1207 19034 1230
rect 18826 1190 18845 1207
rect 19020 1190 19034 1207
rect 18826 1167 19034 1190
rect 18826 1150 18845 1167
rect 19020 1150 19034 1167
rect 18740 1066 18743 1086
rect 18763 1066 18782 1086
rect 18802 1066 18808 1086
rect 18740 584 18808 1066
rect 18740 564 18743 584
rect 18763 564 18782 584
rect 18802 564 18808 584
rect 18740 457 18808 564
rect 18827 1127 19034 1150
rect 18827 1110 18845 1127
rect 19020 1110 19034 1127
rect 18827 1087 19034 1110
rect 18827 1070 18845 1087
rect 19020 1070 19034 1087
rect 18827 1047 19034 1070
rect 18827 1030 18845 1047
rect 19020 1030 19034 1047
rect 18827 1007 19034 1030
rect 18827 990 18845 1007
rect 19020 990 19034 1007
rect 18827 967 19034 990
rect 18827 950 18845 967
rect 19020 950 19034 967
rect 18827 927 19034 950
rect 18827 910 18845 927
rect 19020 910 19034 927
rect 18827 887 19034 910
rect 18827 870 18845 887
rect 19020 870 19034 887
rect 18827 847 19034 870
rect 18827 830 18845 847
rect 19020 830 19034 847
rect 18827 807 19034 830
rect 18827 790 18845 807
rect 19020 790 19034 807
rect 18827 767 19034 790
rect 18827 750 18845 767
rect 19020 750 19034 767
rect 18827 727 19034 750
rect 18827 710 18845 727
rect 19020 710 19034 727
rect 18827 687 19034 710
rect 18827 670 18845 687
rect 19020 670 19034 687
rect 18827 647 19034 670
rect 18827 630 18845 647
rect 19020 630 19034 647
rect 18827 607 19034 630
rect 18827 590 18845 607
rect 19020 590 19034 607
rect 18827 567 19034 590
rect 18827 550 18845 567
rect 19020 550 19034 567
rect 18827 527 19034 550
rect 18827 510 18845 527
rect 19020 510 19034 527
rect 18827 487 19034 510
rect 18827 470 18845 487
rect 19020 470 19034 487
rect 18827 305 19034 470
rect 18550 191 18565 219
rect 18593 191 18612 219
rect 18640 191 18659 219
rect 18687 191 18698 219
rect 18550 172 18698 191
rect 18550 144 18565 172
rect 18593 144 18612 172
rect 18640 144 18659 172
rect 18687 144 18698 172
rect 18550 125 18698 144
rect 18550 97 18565 125
rect 18593 97 18612 125
rect 18640 97 18659 125
rect 18687 97 18698 125
rect 18550 65 18698 97
rect 19065 86 19272 3670
rect 21346 3625 21762 3638
rect 21346 3419 21643 3625
rect 21749 3419 21762 3625
rect 21346 3407 21762 3419
rect 21346 2746 21762 2759
rect 21346 2540 21643 2746
rect 21749 2540 21762 2746
rect 21346 2528 21762 2540
rect 21346 1625 21762 1638
rect 21346 1419 21643 1625
rect 21749 1419 21762 1625
rect 21346 1407 21762 1419
rect 21346 746 21762 759
rect 21346 540 21643 746
rect 21749 540 21762 746
rect 21346 528 21762 540
rect 17632 25 17649 28
rect 17590 8 17596 25
rect 17613 8 17632 25
rect 17649 8 17655 25
rect 17596 1 17613 8
rect 17632 4 17649 8
<< viali >>
rect 21643 11419 21749 11625
rect 21643 10540 21749 10746
rect 1494 9973 1625 10052
rect 765 9912 793 9940
rect 812 9912 840 9940
rect 859 9912 887 9940
rect 765 9865 793 9893
rect 812 9865 840 9893
rect 859 9865 887 9893
rect 765 9818 793 9846
rect 812 9818 840 9846
rect 859 9818 887 9846
rect 252 9310 427 9327
rect 252 8870 427 8887
rect 252 8430 427 8447
rect 252 7990 427 8007
rect 252 7550 427 7567
rect 252 7110 427 7127
rect 252 6670 427 6687
rect 252 6230 427 6247
rect 252 5790 427 5807
rect 252 5350 427 5367
rect 252 4910 427 4927
rect 252 4470 427 4487
rect 252 4030 427 4047
rect 252 3590 427 3607
rect 252 3150 427 3167
rect 252 2710 427 2727
rect 252 2270 427 2287
rect 252 1830 427 1847
rect 252 1390 427 1407
rect 252 950 427 967
rect 252 510 427 527
rect 544 8864 561 8881
rect 544 8362 561 8379
rect 544 7860 561 7877
rect 544 7358 561 7375
rect 544 6856 561 6873
rect 544 6354 561 6371
rect 544 5852 561 5869
rect 544 5350 561 5367
rect 544 4848 561 4865
rect 544 4346 561 4363
rect 544 3844 561 3861
rect 544 3342 561 3359
rect 544 2840 561 2857
rect 544 2338 561 2355
rect 544 1836 561 1853
rect 544 1334 561 1351
rect 598 8670 615 8687
rect 598 8168 615 8185
rect 598 7666 615 7683
rect 598 7164 615 7181
rect 598 6662 615 6679
rect 598 6160 615 6177
rect 598 5658 615 5675
rect 598 5156 615 5173
rect 598 4654 615 4671
rect 598 4152 615 4169
rect 598 3650 615 3667
rect 598 3148 615 3165
rect 598 2646 615 2663
rect 598 2144 615 2161
rect 598 1642 615 1659
rect 598 1140 615 1157
rect 650 9098 670 9118
rect 689 9098 709 9118
rect 650 8596 670 8616
rect 689 8596 709 8616
rect 650 8094 670 8114
rect 689 8094 709 8114
rect 650 7592 670 7612
rect 689 7592 709 7612
rect 650 7090 670 7110
rect 689 7090 709 7110
rect 650 6588 670 6608
rect 689 6588 709 6608
rect 650 6086 670 6106
rect 689 6086 709 6106
rect 650 5584 670 5604
rect 689 5584 709 5604
rect 650 5082 670 5102
rect 689 5082 709 5102
rect 650 4580 670 4600
rect 689 4580 709 4600
rect 650 4078 670 4098
rect 689 4078 709 4098
rect 650 3576 670 3596
rect 689 3576 709 3596
rect 650 3074 670 3094
rect 689 3074 709 3094
rect 650 2572 670 2592
rect 689 2572 709 2592
rect 650 2070 670 2090
rect 689 2070 709 2090
rect 650 1568 670 1588
rect 689 1568 709 1588
rect 650 1066 670 1086
rect 689 1066 709 1086
rect 650 564 670 584
rect 689 564 709 584
rect 761 9394 781 9414
rect 800 9394 820 9414
rect 839 9394 859 9414
rect 878 9394 898 9414
rect 761 9352 781 9372
rect 800 9352 820 9372
rect 839 9352 859 9372
rect 878 9352 898 9372
rect 761 9224 781 9244
rect 800 9224 820 9244
rect 839 9224 859 9244
rect 878 9224 898 9244
rect 761 8892 781 8912
rect 800 8892 820 8912
rect 839 8892 859 8912
rect 878 8892 898 8912
rect 761 8390 781 8410
rect 800 8390 820 8410
rect 839 8390 859 8410
rect 878 8390 898 8410
rect 761 7888 781 7908
rect 800 7888 820 7908
rect 839 7888 859 7908
rect 878 7888 898 7908
rect 761 7386 781 7406
rect 800 7386 820 7406
rect 839 7386 859 7406
rect 878 7386 898 7406
rect 761 6884 781 6904
rect 800 6884 820 6904
rect 839 6884 859 6904
rect 878 6884 898 6904
rect 761 6382 781 6402
rect 800 6382 820 6402
rect 839 6382 859 6402
rect 878 6382 898 6402
rect 761 5880 781 5900
rect 800 5880 820 5900
rect 839 5880 859 5900
rect 878 5880 898 5900
rect 761 5378 781 5398
rect 800 5378 820 5398
rect 839 5378 859 5398
rect 878 5378 898 5398
rect 761 4876 781 4896
rect 800 4876 820 4896
rect 839 4876 859 4896
rect 878 4876 898 4896
rect 761 4374 781 4394
rect 800 4374 820 4394
rect 839 4374 859 4394
rect 878 4374 898 4394
rect 761 3872 781 3892
rect 800 3872 820 3892
rect 839 3872 859 3892
rect 878 3872 898 3892
rect 761 3370 781 3390
rect 800 3370 820 3390
rect 839 3370 859 3390
rect 878 3370 898 3390
rect 761 2868 781 2888
rect 800 2868 820 2888
rect 839 2868 859 2888
rect 878 2868 898 2888
rect 761 2366 781 2386
rect 800 2366 820 2386
rect 839 2366 859 2386
rect 878 2366 898 2386
rect 761 1864 781 1884
rect 800 1864 820 1884
rect 839 1864 859 1884
rect 878 1864 898 1884
rect 761 1362 781 1382
rect 800 1362 820 1382
rect 839 1362 859 1382
rect 878 1362 898 1382
rect 761 860 781 880
rect 800 860 820 880
rect 839 860 859 880
rect 878 860 898 880
rect 761 818 781 838
rect 800 818 820 838
rect 839 818 859 838
rect 878 818 898 838
rect 765 125 793 153
rect 812 125 840 153
rect 859 125 887 153
rect 765 78 793 106
rect 812 78 840 106
rect 859 78 887 106
rect 765 31 793 59
rect 812 31 840 59
rect 859 31 887 59
rect 954 9693 982 9721
rect 1001 9693 1029 9721
rect 1048 9693 1076 9721
rect 954 9646 982 9674
rect 1001 9646 1029 9674
rect 1048 9646 1076 9674
rect 954 9599 982 9627
rect 1001 9599 1029 9627
rect 1048 9599 1076 9627
rect 1497 9693 1525 9721
rect 1544 9693 1572 9721
rect 1591 9693 1619 9721
rect 1497 9646 1525 9674
rect 1544 9646 1572 9674
rect 1591 9646 1619 9674
rect 1497 9599 1525 9627
rect 1544 9599 1572 9627
rect 1591 9599 1619 9627
rect 1847 9693 1875 9721
rect 1894 9693 1922 9721
rect 1941 9693 1969 9721
rect 1847 9646 1875 9674
rect 1894 9646 1922 9674
rect 1941 9646 1969 9674
rect 1847 9599 1875 9627
rect 1894 9599 1922 9627
rect 1941 9599 1969 9627
rect 3058 9973 3189 10052
rect 3061 9693 3089 9721
rect 3108 9693 3136 9721
rect 3155 9693 3183 9721
rect 3061 9646 3089 9674
rect 3108 9646 3136 9674
rect 3155 9646 3183 9674
rect 3061 9599 3089 9627
rect 3108 9599 3136 9627
rect 3155 9599 3183 9627
rect 3494 9973 3625 10052
rect 3497 9693 3525 9721
rect 3544 9693 3572 9721
rect 3591 9693 3619 9721
rect 3497 9646 3525 9674
rect 3544 9646 3572 9674
rect 3591 9646 3619 9674
rect 3497 9599 3525 9627
rect 3544 9599 3572 9627
rect 3591 9599 3619 9627
rect 3847 9693 3875 9721
rect 3894 9693 3922 9721
rect 3941 9693 3969 9721
rect 3847 9646 3875 9674
rect 3894 9646 3922 9674
rect 3941 9646 3969 9674
rect 3847 9599 3875 9627
rect 3894 9599 3922 9627
rect 3941 9599 3969 9627
rect 5058 9973 5189 10052
rect 5061 9693 5089 9721
rect 5108 9693 5136 9721
rect 5155 9693 5183 9721
rect 5061 9646 5089 9674
rect 5108 9646 5136 9674
rect 5155 9646 5183 9674
rect 5061 9599 5089 9627
rect 5108 9599 5136 9627
rect 5155 9599 5183 9627
rect 5494 9973 5625 10052
rect 5497 9693 5525 9721
rect 5544 9693 5572 9721
rect 5591 9693 5619 9721
rect 5497 9646 5525 9674
rect 5544 9646 5572 9674
rect 5591 9646 5619 9674
rect 5497 9599 5525 9627
rect 5544 9599 5572 9627
rect 5591 9599 5619 9627
rect 5847 9693 5875 9721
rect 5894 9693 5922 9721
rect 5941 9693 5969 9721
rect 5847 9646 5875 9674
rect 5894 9646 5922 9674
rect 5941 9646 5969 9674
rect 5847 9599 5875 9627
rect 5894 9599 5922 9627
rect 5941 9599 5969 9627
rect 7058 9973 7189 10052
rect 7061 9693 7089 9721
rect 7108 9693 7136 9721
rect 7155 9693 7183 9721
rect 7061 9646 7089 9674
rect 7108 9646 7136 9674
rect 7155 9646 7183 9674
rect 7061 9599 7089 9627
rect 7108 9599 7136 9627
rect 7155 9599 7183 9627
rect 7494 9973 7625 10052
rect 7497 9693 7525 9721
rect 7544 9693 7572 9721
rect 7591 9693 7619 9721
rect 7497 9646 7525 9674
rect 7544 9646 7572 9674
rect 7591 9646 7619 9674
rect 7497 9599 7525 9627
rect 7544 9599 7572 9627
rect 7591 9599 7619 9627
rect 7847 9693 7875 9721
rect 7894 9693 7922 9721
rect 7941 9693 7969 9721
rect 7847 9646 7875 9674
rect 7894 9646 7922 9674
rect 7941 9646 7969 9674
rect 7847 9599 7875 9627
rect 7894 9599 7922 9627
rect 7941 9599 7969 9627
rect 9058 9973 9189 10052
rect 9061 9693 9089 9721
rect 9108 9693 9136 9721
rect 9155 9693 9183 9721
rect 9061 9646 9089 9674
rect 9108 9646 9136 9674
rect 9155 9646 9183 9674
rect 9061 9599 9089 9627
rect 9108 9599 9136 9627
rect 9155 9599 9183 9627
rect 9494 9973 9625 10052
rect 9497 9693 9525 9721
rect 9544 9693 9572 9721
rect 9591 9693 9619 9721
rect 9497 9646 9525 9674
rect 9544 9646 9572 9674
rect 9591 9646 9619 9674
rect 9497 9599 9525 9627
rect 9544 9599 9572 9627
rect 9591 9599 9619 9627
rect 9847 9693 9875 9721
rect 9894 9693 9922 9721
rect 9941 9693 9969 9721
rect 9847 9646 9875 9674
rect 9894 9646 9922 9674
rect 9941 9646 9969 9674
rect 9847 9599 9875 9627
rect 9894 9599 9922 9627
rect 9941 9599 9969 9627
rect 11058 9973 11189 10052
rect 11061 9693 11089 9721
rect 11108 9693 11136 9721
rect 11155 9693 11183 9721
rect 11061 9646 11089 9674
rect 11108 9646 11136 9674
rect 11155 9646 11183 9674
rect 11061 9599 11089 9627
rect 11108 9599 11136 9627
rect 11155 9599 11183 9627
rect 11494 9973 11625 10052
rect 11497 9693 11525 9721
rect 11544 9693 11572 9721
rect 11591 9693 11619 9721
rect 11497 9646 11525 9674
rect 11544 9646 11572 9674
rect 11591 9646 11619 9674
rect 11497 9599 11525 9627
rect 11544 9599 11572 9627
rect 11591 9599 11619 9627
rect 11847 9693 11875 9721
rect 11894 9693 11922 9721
rect 11941 9693 11969 9721
rect 11847 9646 11875 9674
rect 11894 9646 11922 9674
rect 11941 9646 11969 9674
rect 11847 9599 11875 9627
rect 11894 9599 11922 9627
rect 11941 9599 11969 9627
rect 13058 9973 13189 10052
rect 13061 9693 13089 9721
rect 13108 9693 13136 9721
rect 13155 9693 13183 9721
rect 13061 9646 13089 9674
rect 13108 9646 13136 9674
rect 13155 9646 13183 9674
rect 13061 9599 13089 9627
rect 13108 9599 13136 9627
rect 13155 9599 13183 9627
rect 13494 9973 13625 10052
rect 13497 9693 13525 9721
rect 13544 9693 13572 9721
rect 13591 9693 13619 9721
rect 13497 9646 13525 9674
rect 13544 9646 13572 9674
rect 13591 9646 13619 9674
rect 13497 9599 13525 9627
rect 13544 9599 13572 9627
rect 13591 9599 13619 9627
rect 13847 9693 13875 9721
rect 13894 9693 13922 9721
rect 13941 9693 13969 9721
rect 13847 9646 13875 9674
rect 13894 9646 13922 9674
rect 13941 9646 13969 9674
rect 13847 9599 13875 9627
rect 13894 9599 13922 9627
rect 13941 9599 13969 9627
rect 15058 9973 15189 10052
rect 15061 9693 15089 9721
rect 15108 9693 15136 9721
rect 15155 9693 15183 9721
rect 15061 9646 15089 9674
rect 15108 9646 15136 9674
rect 15155 9646 15183 9674
rect 15061 9599 15089 9627
rect 15108 9599 15136 9627
rect 15155 9599 15183 9627
rect 15494 9973 15625 10052
rect 15497 9693 15525 9721
rect 15544 9693 15572 9721
rect 15591 9693 15619 9721
rect 15497 9646 15525 9674
rect 15544 9646 15572 9674
rect 15591 9646 15619 9674
rect 15497 9599 15525 9627
rect 15544 9599 15572 9627
rect 15591 9599 15619 9627
rect 15847 9693 15875 9721
rect 15894 9693 15922 9721
rect 15941 9693 15969 9721
rect 15847 9646 15875 9674
rect 15894 9646 15922 9674
rect 15941 9646 15969 9674
rect 15847 9599 15875 9627
rect 15894 9599 15922 9627
rect 15941 9599 15969 9627
rect 17058 9973 17189 10052
rect 17061 9693 17089 9721
rect 17108 9693 17136 9721
rect 17155 9693 17183 9721
rect 17061 9646 17089 9674
rect 17108 9646 17136 9674
rect 17155 9646 17183 9674
rect 17061 9599 17089 9627
rect 17108 9599 17136 9627
rect 17155 9599 17183 9627
rect 17494 9973 17625 10052
rect 17497 9693 17525 9721
rect 17544 9693 17572 9721
rect 17591 9693 17619 9721
rect 17497 9646 17525 9674
rect 17544 9646 17572 9674
rect 17591 9646 17619 9674
rect 17497 9599 17525 9627
rect 17544 9599 17572 9627
rect 17591 9599 17619 9627
rect 19058 9990 19189 10052
rect 17847 9693 17875 9721
rect 17894 9693 17922 9721
rect 17941 9693 17969 9721
rect 17847 9646 17875 9674
rect 17894 9646 17922 9674
rect 17941 9646 17969 9674
rect 17847 9599 17875 9627
rect 17894 9599 17922 9627
rect 17941 9599 17969 9627
rect 18376 9688 18404 9716
rect 18423 9688 18451 9716
rect 18470 9688 18498 9716
rect 18376 9641 18404 9669
rect 18423 9641 18451 9669
rect 18470 9641 18498 9669
rect 18376 9594 18404 9622
rect 18423 9594 18451 9622
rect 18470 9594 18498 9622
rect 950 9168 970 9188
rect 989 9168 1009 9188
rect 1028 9168 1048 9188
rect 1067 9168 1087 9188
rect 950 9063 970 9083
rect 989 9063 1009 9083
rect 1028 9063 1048 9083
rect 1067 9063 1087 9083
rect 950 8561 970 8581
rect 989 8561 1009 8581
rect 1028 8561 1048 8581
rect 1067 8561 1087 8581
rect 950 8059 970 8079
rect 989 8059 1009 8079
rect 1028 8059 1048 8079
rect 1067 8059 1087 8079
rect 950 7557 970 7577
rect 989 7557 1009 7577
rect 1028 7557 1048 7577
rect 1067 7557 1087 7577
rect 950 7055 970 7075
rect 989 7055 1009 7075
rect 1028 7055 1048 7075
rect 1067 7055 1087 7075
rect 950 6553 970 6573
rect 989 6553 1009 6573
rect 1028 6553 1048 6573
rect 1067 6553 1087 6573
rect 950 6051 970 6071
rect 989 6051 1009 6071
rect 1028 6051 1048 6071
rect 1067 6051 1087 6071
rect 950 5549 970 5569
rect 989 5549 1009 5569
rect 1028 5549 1048 5569
rect 1067 5549 1087 5569
rect 950 5047 970 5067
rect 989 5047 1009 5067
rect 1028 5047 1048 5067
rect 1067 5047 1087 5067
rect 950 4545 970 4565
rect 989 4545 1009 4565
rect 1028 4545 1048 4565
rect 1067 4545 1087 4565
rect 950 4043 970 4063
rect 989 4043 1009 4063
rect 1028 4043 1048 4063
rect 1067 4043 1087 4063
rect 950 3541 970 3561
rect 989 3541 1009 3561
rect 1028 3541 1048 3561
rect 1067 3541 1087 3561
rect 950 3039 970 3059
rect 989 3039 1009 3059
rect 1028 3039 1048 3059
rect 1067 3039 1087 3059
rect 950 2537 970 2557
rect 989 2537 1009 2557
rect 1028 2537 1048 2557
rect 1067 2537 1087 2557
rect 950 2035 970 2055
rect 989 2035 1009 2055
rect 1028 2035 1048 2055
rect 1067 2035 1087 2055
rect 950 1533 970 1553
rect 989 1533 1009 1553
rect 1028 1533 1048 1553
rect 1067 1533 1087 1553
rect 18377 9294 18405 9322
rect 18424 9294 18452 9322
rect 18471 9294 18499 9322
rect 18377 9247 18405 9275
rect 18424 9247 18452 9275
rect 18471 9247 18499 9275
rect 18377 9200 18405 9228
rect 18424 9200 18452 9228
rect 18471 9200 18499 9228
rect 18365 9063 18385 9083
rect 18404 9063 18424 9083
rect 18443 9063 18463 9083
rect 18482 9063 18502 9083
rect 18365 8561 18385 8581
rect 18404 8561 18424 8581
rect 18443 8561 18463 8581
rect 18482 8561 18502 8581
rect 18376 8286 18404 8314
rect 18423 8286 18451 8314
rect 18470 8286 18498 8314
rect 18376 8239 18404 8267
rect 18423 8239 18451 8267
rect 18470 8239 18498 8267
rect 18376 8192 18404 8220
rect 18423 8192 18451 8220
rect 18470 8192 18498 8220
rect 18365 8059 18385 8079
rect 18404 8059 18424 8079
rect 18443 8059 18463 8079
rect 18482 8059 18502 8079
rect 18365 7557 18385 7577
rect 18404 7557 18424 7577
rect 18443 7557 18463 7577
rect 18482 7557 18502 7577
rect 18376 7286 18404 7314
rect 18423 7286 18451 7314
rect 18470 7286 18498 7314
rect 18376 7239 18404 7267
rect 18423 7239 18451 7267
rect 18470 7239 18498 7267
rect 18376 7192 18404 7220
rect 18423 7192 18451 7220
rect 18470 7192 18498 7220
rect 18365 7055 18385 7075
rect 18404 7055 18424 7075
rect 18443 7055 18463 7075
rect 18482 7055 18502 7075
rect 18565 9907 18593 9935
rect 18612 9907 18640 9935
rect 18659 9907 18687 9935
rect 18565 9860 18593 9888
rect 18612 9860 18640 9888
rect 18659 9860 18687 9888
rect 18565 9813 18593 9841
rect 18612 9813 18640 9841
rect 18659 9813 18687 9841
rect 19061 9693 19089 9721
rect 19108 9693 19136 9721
rect 19155 9693 19183 9721
rect 19061 9646 19089 9674
rect 19108 9646 19136 9674
rect 19155 9646 19183 9674
rect 19061 9599 19089 9627
rect 19108 9599 19136 9627
rect 19155 9599 19183 9627
rect 18554 9394 18574 9414
rect 18593 9394 18613 9414
rect 18632 9394 18652 9414
rect 18671 9394 18691 9414
rect 18554 8892 18574 8912
rect 18593 8892 18613 8912
rect 18632 8892 18652 8912
rect 18671 8892 18691 8912
rect 18565 8802 18593 8830
rect 18612 8802 18640 8830
rect 18659 8802 18687 8830
rect 18565 8755 18593 8783
rect 18612 8755 18640 8783
rect 18659 8755 18687 8783
rect 18565 8708 18593 8736
rect 18612 8708 18640 8736
rect 18659 8708 18687 8736
rect 18554 8390 18574 8410
rect 18593 8390 18613 8410
rect 18632 8390 18652 8410
rect 18671 8390 18691 8410
rect 18554 7888 18574 7908
rect 18593 7888 18613 7908
rect 18632 7888 18652 7908
rect 18671 7888 18691 7908
rect 18565 7748 18593 7776
rect 18612 7748 18640 7776
rect 18659 7748 18687 7776
rect 18565 7701 18593 7729
rect 18612 7701 18640 7729
rect 18659 7701 18687 7729
rect 18565 7654 18593 7682
rect 18612 7654 18640 7682
rect 18659 7654 18687 7682
rect 18554 7386 18574 7406
rect 18593 7386 18613 7406
rect 18632 7386 18652 7406
rect 18671 7386 18691 7406
rect 18554 6884 18574 6904
rect 18593 6884 18613 6904
rect 18632 6884 18652 6904
rect 18671 6884 18691 6904
rect 18564 6783 18592 6811
rect 18611 6783 18639 6811
rect 18658 6783 18686 6811
rect 18564 6736 18592 6764
rect 18611 6736 18639 6764
rect 18658 6736 18686 6764
rect 18564 6689 18592 6717
rect 18611 6689 18639 6717
rect 18658 6689 18686 6717
rect 18365 6553 18385 6573
rect 18404 6553 18424 6573
rect 18443 6553 18463 6573
rect 18482 6553 18502 6573
rect 18377 6324 18405 6352
rect 18424 6324 18452 6352
rect 18471 6324 18499 6352
rect 18377 6277 18405 6305
rect 18424 6277 18452 6305
rect 18471 6277 18499 6305
rect 18377 6230 18405 6258
rect 18424 6230 18452 6258
rect 18471 6230 18499 6258
rect 18365 6051 18385 6071
rect 18404 6051 18424 6071
rect 18443 6051 18463 6071
rect 18482 6051 18502 6071
rect 18365 5549 18385 5569
rect 18404 5549 18424 5569
rect 18443 5549 18463 5569
rect 18482 5549 18502 5569
rect 18376 5261 18404 5289
rect 18423 5261 18451 5289
rect 18470 5261 18498 5289
rect 18376 5214 18404 5242
rect 18423 5214 18451 5242
rect 18470 5214 18498 5242
rect 18376 5167 18404 5195
rect 18423 5167 18451 5195
rect 18470 5167 18498 5195
rect 18365 5047 18385 5067
rect 18404 5047 18424 5067
rect 18443 5047 18463 5067
rect 18482 5047 18502 5067
rect 18365 4545 18385 4565
rect 18404 4545 18424 4565
rect 18443 4545 18463 4565
rect 18482 4545 18502 4565
rect 18377 4273 18405 4301
rect 18424 4273 18452 4301
rect 18471 4273 18499 4301
rect 18377 4226 18405 4254
rect 18424 4226 18452 4254
rect 18471 4226 18499 4254
rect 18377 4179 18405 4207
rect 18424 4179 18452 4207
rect 18471 4179 18499 4207
rect 18365 4043 18385 4063
rect 18404 4043 18424 4063
rect 18443 4043 18463 4063
rect 18482 4043 18502 4063
rect 18554 6382 18574 6402
rect 18593 6382 18613 6402
rect 18632 6382 18652 6402
rect 18671 6382 18691 6402
rect 18743 9098 18763 9118
rect 18782 9098 18802 9118
rect 18743 8596 18763 8616
rect 18782 8596 18802 8616
rect 18743 8094 18763 8114
rect 18782 8094 18802 8114
rect 18743 7592 18763 7612
rect 18782 7592 18802 7612
rect 18743 7090 18763 7110
rect 18782 7090 18802 7110
rect 18743 6588 18763 6608
rect 18782 6588 18802 6608
rect 18554 5880 18574 5900
rect 18593 5880 18613 5900
rect 18632 5880 18652 5900
rect 18671 5880 18691 5900
rect 18565 5775 18593 5803
rect 18612 5775 18640 5803
rect 18659 5775 18687 5803
rect 18565 5728 18593 5756
rect 18612 5728 18640 5756
rect 18659 5728 18687 5756
rect 18565 5681 18593 5709
rect 18612 5681 18640 5709
rect 18659 5681 18687 5709
rect 18554 5378 18574 5398
rect 18593 5378 18613 5398
rect 18632 5378 18652 5398
rect 18671 5378 18691 5398
rect 18554 4876 18574 4896
rect 18593 4876 18613 4896
rect 18632 4876 18652 4896
rect 18671 4876 18691 4896
rect 18565 4774 18593 4802
rect 18612 4774 18640 4802
rect 18659 4774 18687 4802
rect 18565 4727 18593 4755
rect 18612 4727 18640 4755
rect 18659 4727 18687 4755
rect 18565 4680 18593 4708
rect 18612 4680 18640 4708
rect 18659 4680 18687 4708
rect 18554 4374 18574 4394
rect 18593 4374 18613 4394
rect 18632 4374 18652 4394
rect 18671 4374 18691 4394
rect 18743 6086 18763 6106
rect 18782 6086 18802 6106
rect 18743 5584 18763 5604
rect 18782 5584 18802 5604
rect 18743 5082 18763 5102
rect 18782 5082 18802 5102
rect 18743 4580 18763 4600
rect 18782 4580 18802 4600
rect 18554 3872 18574 3892
rect 18593 3872 18613 3892
rect 18632 3872 18652 3892
rect 18671 3872 18691 3892
rect 18564 3775 18592 3803
rect 18611 3775 18639 3803
rect 18658 3775 18686 3803
rect 18564 3728 18592 3756
rect 18611 3728 18639 3756
rect 18658 3728 18686 3756
rect 18564 3681 18592 3709
rect 18611 3681 18639 3709
rect 18658 3681 18686 3709
rect 18365 3541 18385 3561
rect 18404 3541 18424 3561
rect 18443 3541 18463 3561
rect 18482 3541 18502 3561
rect 18377 3251 18405 3279
rect 18424 3251 18452 3279
rect 18471 3251 18499 3279
rect 18377 3204 18405 3232
rect 18424 3204 18452 3232
rect 18471 3204 18499 3232
rect 18377 3157 18405 3185
rect 18424 3157 18452 3185
rect 18471 3157 18499 3185
rect 18365 3039 18385 3059
rect 18404 3039 18424 3059
rect 18443 3039 18463 3059
rect 18482 3039 18502 3059
rect 18365 2537 18385 2557
rect 18404 2537 18424 2557
rect 18443 2537 18463 2557
rect 18482 2537 18502 2557
rect 18377 2254 18405 2282
rect 18424 2254 18452 2282
rect 18471 2254 18499 2282
rect 18377 2207 18405 2235
rect 18424 2207 18452 2235
rect 18471 2207 18499 2235
rect 18377 2160 18405 2188
rect 18424 2160 18452 2188
rect 18471 2160 18499 2188
rect 18365 2035 18385 2055
rect 18404 2035 18424 2055
rect 18443 2035 18463 2055
rect 18482 2035 18502 2055
rect 18365 1533 18385 1553
rect 18404 1533 18424 1553
rect 18443 1533 18463 1553
rect 18482 1533 18502 1553
rect 18554 3370 18574 3390
rect 18593 3370 18613 3390
rect 18632 3370 18652 3390
rect 18671 3370 18691 3390
rect 18743 4078 18763 4098
rect 18782 4078 18802 4098
rect 18743 3576 18763 3596
rect 18782 3576 18802 3596
rect 18554 2868 18574 2888
rect 18593 2868 18613 2888
rect 18632 2868 18652 2888
rect 18671 2868 18691 2888
rect 18565 2741 18593 2769
rect 18612 2741 18640 2769
rect 18659 2741 18687 2769
rect 18565 2694 18593 2722
rect 18612 2694 18640 2722
rect 18659 2694 18687 2722
rect 18565 2647 18593 2675
rect 18612 2647 18640 2675
rect 18659 2647 18687 2675
rect 18554 2366 18574 2386
rect 18593 2366 18613 2386
rect 18632 2366 18652 2386
rect 18671 2366 18691 2386
rect 18743 3074 18763 3094
rect 18782 3074 18802 3094
rect 18743 2572 18763 2592
rect 18782 2572 18802 2592
rect 18554 1864 18574 1884
rect 18593 1864 18613 1884
rect 18632 1864 18652 1884
rect 18671 1864 18691 1884
rect 18565 1739 18593 1767
rect 18612 1739 18640 1767
rect 18659 1739 18687 1767
rect 18565 1692 18593 1720
rect 18612 1692 18640 1720
rect 18659 1692 18687 1720
rect 18565 1645 18593 1673
rect 18612 1645 18640 1673
rect 18659 1645 18687 1673
rect 18554 1362 18574 1382
rect 18593 1362 18613 1382
rect 18632 1362 18652 1382
rect 18671 1362 18691 1382
rect 18375 1254 18403 1282
rect 18422 1254 18450 1282
rect 18469 1254 18497 1282
rect 18375 1207 18403 1235
rect 18422 1207 18450 1235
rect 18469 1207 18497 1235
rect 18375 1160 18403 1188
rect 18422 1160 18450 1188
rect 18469 1160 18497 1188
rect 950 1031 970 1051
rect 989 1031 1009 1051
rect 1028 1031 1048 1051
rect 1067 1031 1087 1051
rect 950 690 970 710
rect 989 690 1009 710
rect 1028 690 1048 710
rect 1067 690 1087 710
rect 950 634 970 654
rect 989 634 1009 654
rect 1028 634 1048 654
rect 1067 634 1087 654
rect 950 529 970 549
rect 989 529 1009 549
rect 1028 529 1048 549
rect 1067 529 1087 549
rect 18365 1031 18385 1051
rect 18404 1031 18424 1051
rect 18443 1031 18463 1051
rect 18482 1031 18502 1051
rect 18365 529 18385 549
rect 18404 529 18424 549
rect 18443 529 18463 549
rect 18482 529 18502 549
rect 954 344 982 372
rect 1001 344 1029 372
rect 1048 344 1076 372
rect 954 297 982 325
rect 1001 297 1029 325
rect 1048 297 1076 325
rect 954 250 982 278
rect 1001 250 1029 278
rect 1048 250 1076 278
rect 1620 145 1637 162
rect 14478 304 14495 321
rect 15678 304 15695 321
rect 14580 265 14597 282
rect 16180 265 16197 282
rect 14682 227 14699 244
rect 16682 227 16699 244
rect 14784 189 14801 206
rect 17184 189 17201 206
rect 14886 151 14903 168
rect 17299 376 17316 393
rect 17543 376 17560 393
rect 17686 151 17703 168
rect 18376 409 18404 437
rect 18423 409 18451 437
rect 18470 409 18498 437
rect 18376 362 18404 390
rect 18423 362 18451 390
rect 18470 362 18498 390
rect 18376 315 18404 343
rect 18423 315 18451 343
rect 18470 315 18498 343
rect 18190 142 18207 159
rect 18554 860 18574 880
rect 18593 860 18613 880
rect 18632 860 18652 880
rect 18671 860 18691 880
rect 18565 742 18593 770
rect 18612 742 18640 770
rect 18659 742 18687 770
rect 18565 695 18593 723
rect 18612 695 18640 723
rect 18659 695 18687 723
rect 18565 648 18593 676
rect 18612 648 18640 676
rect 18659 648 18687 676
rect 18743 2070 18763 2090
rect 18782 2070 18802 2090
rect 18743 1568 18763 1588
rect 18782 1568 18802 1588
rect 18845 9310 19020 9327
rect 18845 8870 19020 8887
rect 18845 8430 19020 8447
rect 18845 7990 19020 8007
rect 18845 7550 19020 7567
rect 18845 7110 19020 7127
rect 21643 9419 21749 9625
rect 21643 8540 21749 8746
rect 21643 7419 21749 7625
rect 18845 6230 19020 6247
rect 18845 5350 19020 5367
rect 18845 4910 19020 4927
rect 18845 4470 19020 4487
rect 18845 4030 19020 4047
rect 21643 6540 21749 6746
rect 21643 5419 21749 5625
rect 21643 4540 21749 4746
rect 18845 3590 19020 3607
rect 18845 3150 19020 3167
rect 18845 2270 19020 2287
rect 18845 1830 19020 1847
rect 18845 1390 19020 1407
rect 18743 1066 18763 1086
rect 18782 1066 18802 1086
rect 18743 564 18763 584
rect 18782 564 18802 584
rect 18845 950 19020 967
rect 18845 510 19020 527
rect 18565 191 18593 219
rect 18612 191 18640 219
rect 18659 191 18687 219
rect 18565 144 18593 172
rect 18612 144 18640 172
rect 18659 144 18687 172
rect 18565 97 18593 125
rect 18612 97 18640 125
rect 18659 97 18687 125
rect 21643 3419 21749 3625
rect 21643 2540 21749 2746
rect 21643 1419 21749 1625
rect 21643 540 21749 746
rect 17596 8 17613 25
rect 17632 8 17649 25
<< metal1 >>
rect 21346 11828 21762 11834
rect 21346 11747 21637 11828
rect 21756 11747 21762 11828
rect 21346 11742 21762 11747
rect 21630 11625 21762 11638
rect 21630 11419 21643 11625
rect 21749 11419 21762 11625
rect 21630 11407 21762 11419
rect 21346 11394 21514 11403
rect 21346 11319 21397 11394
rect 21503 11319 21514 11394
rect 21346 11312 21514 11319
rect 21346 11123 21514 11132
rect 21346 11048 21397 11123
rect 21503 11048 21514 11123
rect 21346 11041 21514 11048
rect 21346 10845 21514 10854
rect 21346 10770 21397 10845
rect 21503 10770 21514 10845
rect 21346 10763 21514 10770
rect 21630 10746 21762 10759
rect 21630 10540 21643 10746
rect 21749 10540 21762 10746
rect 21630 10528 21762 10540
rect 21346 10273 21762 10279
rect 21346 10192 21637 10273
rect 21756 10192 21762 10273
rect 21346 10187 21762 10192
rect 1487 10052 1633 10083
rect 1487 9973 1494 10052
rect 1625 9973 1633 10052
rect 1487 9967 1633 9973
rect 2255 9950 2440 10083
rect 3051 10052 3197 10083
rect 3051 9973 3058 10052
rect 3189 9973 3197 10052
rect 3051 9967 3197 9973
rect 3487 10052 3633 10083
rect 3487 9973 3494 10052
rect 3625 9973 3633 10052
rect 3487 9967 3633 9973
rect 4255 9950 4440 10083
rect 5051 10052 5197 10083
rect 5051 9973 5058 10052
rect 5189 9973 5197 10052
rect 5051 9967 5197 9973
rect 5487 10052 5633 10083
rect 5487 9973 5494 10052
rect 5625 9973 5633 10052
rect 5487 9967 5633 9973
rect 6255 9950 6440 10083
rect 7051 10052 7197 10083
rect 7051 9973 7058 10052
rect 7189 9973 7197 10052
rect 7051 9967 7197 9973
rect 7487 10052 7633 10083
rect 7487 9973 7494 10052
rect 7625 9973 7633 10052
rect 7487 9967 7633 9973
rect 8255 9950 8440 10083
rect 9051 10052 9197 10083
rect 9051 9973 9058 10052
rect 9189 9973 9197 10052
rect 9051 9967 9197 9973
rect 9487 10052 9633 10083
rect 9487 9973 9494 10052
rect 9625 9973 9633 10052
rect 9487 9967 9633 9973
rect 10255 9950 10440 10083
rect 11051 10052 11197 10083
rect 11051 9973 11058 10052
rect 11189 9973 11197 10052
rect 11051 9967 11197 9973
rect 11487 10052 11633 10083
rect 11487 9973 11494 10052
rect 11625 9973 11633 10052
rect 11487 9967 11633 9973
rect 12255 9950 12440 10083
rect 13051 10052 13197 10083
rect 13051 9973 13058 10052
rect 13189 9973 13197 10052
rect 13051 9967 13197 9973
rect 13487 10052 13633 10083
rect 13487 9973 13494 10052
rect 13625 9973 13633 10052
rect 13487 9967 13633 9973
rect 14255 9950 14440 10083
rect 15051 10052 15197 10083
rect 15051 9973 15058 10052
rect 15189 9973 15197 10052
rect 15051 9967 15197 9973
rect 15487 10052 15633 10083
rect 15487 9973 15494 10052
rect 15625 9973 15633 10052
rect 15487 9967 15633 9973
rect 16255 9950 16440 10083
rect 17051 10052 17197 10083
rect 17051 9973 17058 10052
rect 17189 9973 17197 10052
rect 17051 9967 17197 9973
rect 17487 10052 17633 10083
rect 17487 9973 17494 10052
rect 17625 9973 17633 10052
rect 17487 9967 17633 9973
rect 18255 9950 18440 10083
rect 19051 10052 19197 10083
rect 19051 9990 19058 10052
rect 19189 9990 19197 10052
rect 19051 9984 19197 9990
rect 0 9946 19272 9950
rect 0 9914 15 9946
rect 47 9914 59 9946
rect 91 9914 103 9946
rect 135 9914 147 9946
rect 179 9941 19093 9946
rect 179 9940 2267 9941
rect 179 9914 765 9940
rect 0 9912 765 9914
rect 793 9912 812 9940
rect 840 9912 859 9940
rect 887 9912 2267 9940
rect 0 9901 2267 9912
rect 0 9869 15 9901
rect 47 9869 59 9901
rect 91 9869 103 9901
rect 135 9869 147 9901
rect 179 9893 2267 9901
rect 179 9869 765 9893
rect 0 9865 765 9869
rect 793 9865 812 9893
rect 840 9865 859 9893
rect 887 9865 2267 9893
rect 0 9856 2267 9865
rect 0 9824 15 9856
rect 47 9824 59 9856
rect 91 9824 103 9856
rect 135 9824 147 9856
rect 179 9846 2267 9856
rect 179 9824 765 9846
rect 0 9818 765 9824
rect 793 9818 812 9846
rect 840 9818 859 9846
rect 887 9819 2267 9846
rect 2430 9819 4267 9941
rect 4430 9819 6267 9941
rect 6430 9819 8267 9941
rect 8430 9819 10267 9941
rect 10430 9819 12267 9941
rect 12430 9819 14267 9941
rect 14430 9819 16267 9941
rect 16430 9819 18267 9941
rect 18430 9935 19093 9941
rect 18430 9907 18565 9935
rect 18593 9907 18612 9935
rect 18640 9907 18659 9935
rect 18687 9914 19093 9935
rect 19125 9914 19137 9946
rect 19169 9914 19181 9946
rect 19213 9914 19225 9946
rect 19257 9914 19272 9946
rect 18687 9907 19272 9914
rect 18430 9901 19272 9907
rect 18430 9888 19093 9901
rect 18430 9860 18565 9888
rect 18593 9860 18612 9888
rect 18640 9860 18659 9888
rect 18687 9869 19093 9888
rect 19125 9869 19137 9901
rect 19169 9869 19181 9901
rect 19213 9869 19225 9901
rect 19257 9869 19272 9901
rect 18687 9860 19272 9869
rect 18430 9856 19272 9860
rect 18430 9841 19093 9856
rect 18430 9819 18565 9841
rect 887 9818 18565 9819
rect 0 9813 18565 9818
rect 18593 9813 18612 9841
rect 18640 9813 18659 9841
rect 18687 9824 19093 9841
rect 19125 9824 19137 9856
rect 19169 9824 19181 9856
rect 19213 9824 19225 9856
rect 19257 9824 19272 9856
rect 18687 9813 19272 9824
rect 0 9810 19272 9813
rect 21346 9828 21762 9834
rect 18361 9805 18697 9810
rect 21346 9747 21637 9828
rect 21756 9747 21762 9828
rect 21346 9742 21762 9747
rect 238 9727 19272 9731
rect 238 9695 253 9727
rect 285 9695 297 9727
rect 329 9695 341 9727
rect 373 9695 385 9727
rect 417 9721 18855 9727
rect 417 9695 954 9721
rect 238 9693 954 9695
rect 982 9693 1001 9721
rect 1029 9693 1048 9721
rect 1076 9693 1497 9721
rect 1525 9693 1544 9721
rect 1572 9693 1591 9721
rect 1619 9693 1847 9721
rect 1875 9693 1894 9721
rect 1922 9693 1941 9721
rect 1969 9693 3061 9721
rect 3089 9693 3108 9721
rect 3136 9693 3155 9721
rect 3183 9693 3497 9721
rect 3525 9693 3544 9721
rect 3572 9693 3591 9721
rect 3619 9693 3847 9721
rect 3875 9693 3894 9721
rect 3922 9693 3941 9721
rect 3969 9693 5061 9721
rect 5089 9693 5108 9721
rect 5136 9693 5155 9721
rect 5183 9693 5497 9721
rect 5525 9693 5544 9721
rect 5572 9693 5591 9721
rect 5619 9693 5847 9721
rect 5875 9693 5894 9721
rect 5922 9693 5941 9721
rect 5969 9693 7061 9721
rect 7089 9693 7108 9721
rect 7136 9693 7155 9721
rect 7183 9693 7497 9721
rect 7525 9693 7544 9721
rect 7572 9693 7591 9721
rect 7619 9693 7847 9721
rect 7875 9693 7894 9721
rect 7922 9693 7941 9721
rect 7969 9693 9061 9721
rect 9089 9693 9108 9721
rect 9136 9693 9155 9721
rect 9183 9693 9497 9721
rect 9525 9693 9544 9721
rect 9572 9693 9591 9721
rect 9619 9693 9847 9721
rect 9875 9693 9894 9721
rect 9922 9693 9941 9721
rect 9969 9693 11061 9721
rect 11089 9693 11108 9721
rect 11136 9693 11155 9721
rect 11183 9693 11497 9721
rect 11525 9693 11544 9721
rect 11572 9693 11591 9721
rect 11619 9693 11847 9721
rect 11875 9693 11894 9721
rect 11922 9693 11941 9721
rect 11969 9693 13061 9721
rect 13089 9693 13108 9721
rect 13136 9693 13155 9721
rect 13183 9693 13497 9721
rect 13525 9693 13544 9721
rect 13572 9693 13591 9721
rect 13619 9693 13847 9721
rect 13875 9693 13894 9721
rect 13922 9693 13941 9721
rect 13969 9693 15061 9721
rect 15089 9693 15108 9721
rect 15136 9693 15155 9721
rect 15183 9693 15497 9721
rect 15525 9693 15544 9721
rect 15572 9693 15591 9721
rect 15619 9693 15847 9721
rect 15875 9693 15894 9721
rect 15922 9693 15941 9721
rect 15969 9693 17061 9721
rect 17089 9693 17108 9721
rect 17136 9693 17155 9721
rect 17183 9693 17497 9721
rect 17525 9693 17544 9721
rect 17572 9693 17591 9721
rect 17619 9693 17847 9721
rect 17875 9693 17894 9721
rect 17922 9693 17941 9721
rect 17969 9716 18855 9721
rect 17969 9693 18376 9716
rect 238 9688 18376 9693
rect 18404 9688 18423 9716
rect 18451 9688 18470 9716
rect 18498 9695 18855 9716
rect 18887 9695 18899 9727
rect 18931 9695 18943 9727
rect 18975 9695 18987 9727
rect 19019 9721 19272 9727
rect 19019 9695 19061 9721
rect 18498 9693 19061 9695
rect 19089 9693 19108 9721
rect 19136 9693 19155 9721
rect 19183 9693 19272 9721
rect 18498 9688 19272 9693
rect 238 9682 19272 9688
rect 238 9650 253 9682
rect 285 9650 297 9682
rect 329 9650 341 9682
rect 373 9650 385 9682
rect 417 9674 18855 9682
rect 417 9650 954 9674
rect 238 9646 954 9650
rect 982 9646 1001 9674
rect 1029 9646 1048 9674
rect 1076 9646 1497 9674
rect 1525 9646 1544 9674
rect 1572 9646 1591 9674
rect 1619 9646 1847 9674
rect 1875 9646 1894 9674
rect 1922 9646 1941 9674
rect 1969 9646 3061 9674
rect 3089 9646 3108 9674
rect 3136 9646 3155 9674
rect 3183 9646 3497 9674
rect 3525 9646 3544 9674
rect 3572 9646 3591 9674
rect 3619 9646 3847 9674
rect 3875 9646 3894 9674
rect 3922 9646 3941 9674
rect 3969 9646 5061 9674
rect 5089 9646 5108 9674
rect 5136 9646 5155 9674
rect 5183 9646 5497 9674
rect 5525 9646 5544 9674
rect 5572 9646 5591 9674
rect 5619 9646 5847 9674
rect 5875 9646 5894 9674
rect 5922 9646 5941 9674
rect 5969 9646 7061 9674
rect 7089 9646 7108 9674
rect 7136 9646 7155 9674
rect 7183 9646 7497 9674
rect 7525 9646 7544 9674
rect 7572 9646 7591 9674
rect 7619 9646 7847 9674
rect 7875 9646 7894 9674
rect 7922 9646 7941 9674
rect 7969 9646 9061 9674
rect 9089 9646 9108 9674
rect 9136 9646 9155 9674
rect 9183 9646 9497 9674
rect 9525 9646 9544 9674
rect 9572 9646 9591 9674
rect 9619 9646 9847 9674
rect 9875 9646 9894 9674
rect 9922 9646 9941 9674
rect 9969 9646 11061 9674
rect 11089 9646 11108 9674
rect 11136 9646 11155 9674
rect 11183 9646 11497 9674
rect 11525 9646 11544 9674
rect 11572 9646 11591 9674
rect 11619 9646 11847 9674
rect 11875 9646 11894 9674
rect 11922 9646 11941 9674
rect 11969 9646 13061 9674
rect 13089 9646 13108 9674
rect 13136 9646 13155 9674
rect 13183 9646 13497 9674
rect 13525 9646 13544 9674
rect 13572 9646 13591 9674
rect 13619 9646 13847 9674
rect 13875 9646 13894 9674
rect 13922 9646 13941 9674
rect 13969 9646 15061 9674
rect 15089 9646 15108 9674
rect 15136 9646 15155 9674
rect 15183 9646 15497 9674
rect 15525 9646 15544 9674
rect 15572 9646 15591 9674
rect 15619 9646 15847 9674
rect 15875 9646 15894 9674
rect 15922 9646 15941 9674
rect 15969 9646 17061 9674
rect 17089 9646 17108 9674
rect 17136 9646 17155 9674
rect 17183 9646 17497 9674
rect 17525 9646 17544 9674
rect 17572 9646 17591 9674
rect 17619 9646 17847 9674
rect 17875 9646 17894 9674
rect 17922 9646 17941 9674
rect 17969 9669 18855 9674
rect 17969 9646 18376 9669
rect 238 9641 18376 9646
rect 18404 9641 18423 9669
rect 18451 9641 18470 9669
rect 18498 9650 18855 9669
rect 18887 9650 18899 9682
rect 18931 9650 18943 9682
rect 18975 9650 18987 9682
rect 19019 9674 19272 9682
rect 19019 9650 19061 9674
rect 18498 9646 19061 9650
rect 19089 9646 19108 9674
rect 19136 9646 19155 9674
rect 19183 9646 19272 9674
rect 18498 9641 19272 9646
rect 238 9637 19272 9641
rect 238 9605 253 9637
rect 285 9605 297 9637
rect 329 9605 341 9637
rect 373 9605 385 9637
rect 417 9627 18855 9637
rect 417 9605 954 9627
rect 238 9599 954 9605
rect 982 9599 1001 9627
rect 1029 9599 1048 9627
rect 1076 9599 1497 9627
rect 1525 9599 1544 9627
rect 1572 9599 1591 9627
rect 1619 9599 1847 9627
rect 1875 9599 1894 9627
rect 1922 9599 1941 9627
rect 1969 9599 3061 9627
rect 3089 9599 3108 9627
rect 3136 9599 3155 9627
rect 3183 9599 3497 9627
rect 3525 9599 3544 9627
rect 3572 9599 3591 9627
rect 3619 9599 3847 9627
rect 3875 9599 3894 9627
rect 3922 9599 3941 9627
rect 3969 9599 5061 9627
rect 5089 9599 5108 9627
rect 5136 9599 5155 9627
rect 5183 9599 5497 9627
rect 5525 9599 5544 9627
rect 5572 9599 5591 9627
rect 5619 9599 5847 9627
rect 5875 9599 5894 9627
rect 5922 9599 5941 9627
rect 5969 9599 7061 9627
rect 7089 9599 7108 9627
rect 7136 9599 7155 9627
rect 7183 9599 7497 9627
rect 7525 9599 7544 9627
rect 7572 9599 7591 9627
rect 7619 9599 7847 9627
rect 7875 9599 7894 9627
rect 7922 9599 7941 9627
rect 7969 9599 9061 9627
rect 9089 9599 9108 9627
rect 9136 9599 9155 9627
rect 9183 9599 9497 9627
rect 9525 9599 9544 9627
rect 9572 9599 9591 9627
rect 9619 9599 9847 9627
rect 9875 9599 9894 9627
rect 9922 9599 9941 9627
rect 9969 9599 11061 9627
rect 11089 9599 11108 9627
rect 11136 9599 11155 9627
rect 11183 9599 11497 9627
rect 11525 9599 11544 9627
rect 11572 9599 11591 9627
rect 11619 9599 11847 9627
rect 11875 9599 11894 9627
rect 11922 9599 11941 9627
rect 11969 9599 13061 9627
rect 13089 9599 13108 9627
rect 13136 9599 13155 9627
rect 13183 9599 13497 9627
rect 13525 9599 13544 9627
rect 13572 9599 13591 9627
rect 13619 9599 13847 9627
rect 13875 9599 13894 9627
rect 13922 9599 13941 9627
rect 13969 9599 15061 9627
rect 15089 9599 15108 9627
rect 15136 9599 15155 9627
rect 15183 9599 15497 9627
rect 15525 9599 15544 9627
rect 15572 9599 15591 9627
rect 15619 9599 15847 9627
rect 15875 9599 15894 9627
rect 15922 9599 15941 9627
rect 15969 9599 17061 9627
rect 17089 9599 17108 9627
rect 17136 9599 17155 9627
rect 17183 9599 17497 9627
rect 17525 9599 17544 9627
rect 17572 9599 17591 9627
rect 17619 9599 17847 9627
rect 17875 9599 17894 9627
rect 17922 9599 17941 9627
rect 17969 9622 18855 9627
rect 17969 9599 18376 9622
rect 238 9594 18376 9599
rect 18404 9594 18423 9622
rect 18451 9594 18470 9622
rect 18498 9605 18855 9622
rect 18887 9605 18899 9637
rect 18931 9605 18943 9637
rect 18975 9605 18987 9637
rect 19019 9627 19272 9637
rect 19019 9605 19061 9627
rect 18498 9599 19061 9605
rect 19089 9599 19108 9627
rect 19136 9599 19155 9627
rect 19183 9599 19272 9627
rect 18498 9594 19272 9599
rect 238 9592 19272 9594
rect 239 9591 19272 9592
rect 21630 9625 21762 9638
rect 18361 9586 18697 9591
rect 21630 9419 21643 9625
rect 21749 9419 21762 9625
rect 755 9414 1195 9418
rect 755 9394 761 9414
rect 781 9394 800 9414
rect 820 9394 839 9414
rect 859 9394 878 9414
rect 898 9394 1195 9414
rect 755 9390 1195 9394
rect 18263 9414 18698 9418
rect 18263 9394 18554 9414
rect 18574 9394 18593 9414
rect 18613 9394 18632 9414
rect 18652 9394 18671 9414
rect 18691 9394 18698 9414
rect 21630 9407 21762 9419
rect 18263 9390 18698 9394
rect 21346 9394 21514 9403
rect 755 9372 1195 9376
rect 755 9352 761 9372
rect 781 9352 800 9372
rect 820 9352 839 9372
rect 859 9352 878 9372
rect 898 9362 1195 9372
rect 898 9352 904 9362
rect 755 9348 904 9352
rect 246 9305 252 9331
rect 427 9305 433 9331
rect 18839 9330 18845 9331
rect 18363 9322 18845 9330
rect 19020 9330 19026 9331
rect 19020 9329 19034 9330
rect 18363 9294 18377 9322
rect 18405 9294 18424 9322
rect 18452 9294 18471 9322
rect 18499 9305 18845 9322
rect 18499 9294 18856 9305
rect 18363 9284 18856 9294
rect 18888 9284 18900 9305
rect 18932 9284 18944 9305
rect 18976 9284 18988 9305
rect 19020 9284 19035 9329
rect 21346 9319 21397 9394
rect 21503 9319 21514 9394
rect 21346 9312 21514 9319
rect 18363 9275 19035 9284
rect 755 9247 1195 9261
rect 18363 9247 18377 9275
rect 18405 9247 18424 9275
rect 18452 9247 18471 9275
rect 18499 9271 19035 9275
rect 18499 9247 18856 9271
rect 755 9244 904 9247
rect 755 9224 761 9244
rect 781 9224 800 9244
rect 820 9224 839 9244
rect 859 9224 878 9244
rect 898 9224 904 9244
rect 755 9220 904 9224
rect 18363 9239 18856 9247
rect 18888 9239 18900 9271
rect 18932 9239 18944 9271
rect 18976 9239 18988 9271
rect 19020 9239 19035 9271
rect 18363 9228 19035 9239
rect 755 9206 1195 9220
rect 18363 9200 18377 9228
rect 18405 9200 18424 9228
rect 18452 9200 18471 9228
rect 18499 9226 19035 9228
rect 18499 9200 18856 9226
rect 18363 9194 18856 9200
rect 18888 9194 18900 9226
rect 18932 9194 18944 9226
rect 18976 9194 18988 9226
rect 19020 9194 19035 9226
rect 944 9188 1195 9192
rect 18363 9190 19035 9194
rect 944 9168 950 9188
rect 970 9168 989 9188
rect 1009 9168 1028 9188
rect 1048 9168 1067 9188
rect 1087 9178 1195 9188
rect 1087 9168 1093 9178
rect 944 9164 1093 9168
rect 21346 9123 21514 9132
rect 644 9118 730 9121
rect 644 9098 650 9118
rect 670 9098 689 9118
rect 709 9115 730 9118
rect 18722 9118 18808 9121
rect 18722 9115 18743 9118
rect 709 9101 1195 9115
rect 18263 9101 18743 9115
rect 709 9098 730 9101
rect 644 9095 730 9098
rect 18722 9098 18743 9101
rect 18763 9098 18782 9118
rect 18802 9098 18808 9118
rect 18722 9095 18808 9098
rect 944 9083 1195 9087
rect 944 9063 950 9083
rect 970 9063 989 9083
rect 1009 9063 1028 9083
rect 1048 9063 1067 9083
rect 1087 9063 1195 9083
rect 944 9059 1195 9063
rect 18263 9083 18508 9087
rect 18263 9063 18365 9083
rect 18385 9063 18404 9083
rect 18424 9063 18443 9083
rect 18463 9063 18482 9083
rect 18502 9063 18508 9083
rect 18263 9059 18508 9063
rect 21346 9048 21397 9123
rect 21503 9048 21514 9123
rect 21346 9041 21514 9048
rect 755 8912 1195 8916
rect 755 8892 761 8912
rect 781 8892 800 8912
rect 820 8892 839 8912
rect 859 8892 878 8912
rect 898 8892 1195 8912
rect 246 8865 252 8891
rect 427 8865 433 8891
rect 755 8888 1195 8892
rect 18263 8912 18698 8916
rect 18263 8892 18554 8912
rect 18574 8892 18593 8912
rect 18613 8892 18632 8912
rect 18652 8892 18671 8912
rect 18691 8892 18698 8912
rect 18263 8888 18698 8892
rect 536 8881 570 8884
rect 536 8864 544 8881
rect 561 8874 570 8881
rect 561 8864 1195 8874
rect 18839 8865 18845 8891
rect 19020 8865 19026 8891
rect 536 8860 1195 8864
rect 21346 8845 21514 8854
rect 18550 8837 18698 8838
rect 18550 8830 19272 8837
rect 18550 8802 18565 8830
rect 18593 8802 18612 8830
rect 18640 8802 18659 8830
rect 18687 8823 19272 8830
rect 18687 8802 19093 8823
rect 18550 8791 19093 8802
rect 19125 8791 19137 8823
rect 19169 8791 19181 8823
rect 19213 8791 19225 8823
rect 19257 8791 19272 8823
rect 18550 8783 19272 8791
rect 522 8745 1195 8759
rect 18550 8755 18565 8783
rect 18593 8755 18612 8783
rect 18640 8755 18659 8783
rect 18687 8778 19272 8783
rect 18687 8755 19093 8778
rect 18550 8746 19093 8755
rect 19125 8746 19137 8778
rect 19169 8746 19181 8778
rect 19213 8746 19225 8778
rect 19257 8746 19272 8778
rect 21346 8770 21397 8845
rect 21503 8770 21514 8845
rect 21346 8763 21514 8770
rect 18550 8736 19272 8746
rect 522 8704 1195 8718
rect 18550 8708 18565 8736
rect 18593 8708 18612 8736
rect 18640 8708 18659 8736
rect 18687 8733 19272 8736
rect 18687 8708 19093 8733
rect 18550 8701 19093 8708
rect 19125 8701 19137 8733
rect 19169 8701 19181 8733
rect 19213 8701 19225 8733
rect 19257 8701 19272 8733
rect 18550 8697 19272 8701
rect 21630 8746 21762 8759
rect 590 8687 1195 8690
rect 590 8670 598 8687
rect 615 8676 1195 8687
rect 615 8670 624 8676
rect 590 8666 624 8670
rect 644 8616 730 8619
rect 644 8596 650 8616
rect 670 8596 689 8616
rect 709 8613 730 8616
rect 18722 8616 18808 8619
rect 18722 8613 18743 8616
rect 709 8599 1195 8613
rect 18263 8599 18743 8613
rect 709 8596 730 8599
rect 644 8593 730 8596
rect 18722 8596 18743 8599
rect 18763 8596 18782 8616
rect 18802 8596 18808 8616
rect 18722 8593 18808 8596
rect 944 8581 1195 8585
rect 944 8561 950 8581
rect 970 8561 989 8581
rect 1009 8561 1028 8581
rect 1048 8561 1067 8581
rect 1087 8561 1195 8581
rect 944 8557 1195 8561
rect 18263 8581 18508 8585
rect 18263 8561 18365 8581
rect 18385 8561 18404 8581
rect 18424 8561 18443 8581
rect 18463 8561 18482 8581
rect 18502 8561 18508 8581
rect 18263 8557 18508 8561
rect 21630 8540 21643 8746
rect 21749 8540 21762 8746
rect 21630 8528 21762 8540
rect 246 8425 252 8451
rect 427 8425 433 8451
rect 18839 8425 18845 8451
rect 19020 8425 19026 8451
rect 755 8410 1195 8414
rect 755 8390 761 8410
rect 781 8390 800 8410
rect 820 8390 839 8410
rect 859 8390 878 8410
rect 898 8390 1195 8410
rect 755 8386 1195 8390
rect 18263 8410 18698 8414
rect 18263 8390 18554 8410
rect 18574 8390 18593 8410
rect 18613 8390 18632 8410
rect 18652 8390 18671 8410
rect 18691 8390 18698 8410
rect 18263 8386 18698 8390
rect 536 8379 570 8382
rect 536 8362 544 8379
rect 561 8372 570 8379
rect 561 8362 1195 8372
rect 536 8358 1195 8362
rect 18362 8321 19033 8322
rect 18362 8314 19034 8321
rect 18362 8286 18376 8314
rect 18404 8286 18423 8314
rect 18451 8286 18470 8314
rect 18498 8308 19034 8314
rect 18498 8286 18855 8308
rect 18362 8276 18855 8286
rect 18887 8276 18899 8308
rect 18931 8276 18943 8308
rect 18975 8276 18987 8308
rect 19019 8276 19034 8308
rect 18362 8267 19034 8276
rect 522 8243 1195 8257
rect 18362 8239 18376 8267
rect 18404 8239 18423 8267
rect 18451 8239 18470 8267
rect 18498 8263 19034 8267
rect 18498 8239 18855 8263
rect 18362 8231 18855 8239
rect 18887 8231 18899 8263
rect 18931 8231 18943 8263
rect 18975 8231 18987 8263
rect 19019 8231 19034 8263
rect 18362 8220 19034 8231
rect 522 8202 1195 8216
rect 18362 8192 18376 8220
rect 18404 8192 18423 8220
rect 18451 8192 18470 8220
rect 18498 8218 19034 8220
rect 18498 8192 18855 8218
rect 590 8185 1195 8188
rect 590 8168 598 8185
rect 615 8174 1195 8185
rect 18362 8186 18855 8192
rect 18887 8186 18899 8218
rect 18931 8186 18943 8218
rect 18975 8186 18987 8218
rect 19019 8186 19034 8218
rect 21346 8273 21762 8279
rect 21346 8192 21637 8273
rect 21756 8192 21762 8273
rect 21346 8187 21762 8192
rect 18362 8182 19034 8186
rect 615 8168 624 8174
rect 590 8164 624 8168
rect 644 8114 730 8117
rect 644 8094 650 8114
rect 670 8094 689 8114
rect 709 8111 730 8114
rect 18722 8114 18808 8117
rect 18722 8111 18743 8114
rect 709 8097 1195 8111
rect 18263 8097 18743 8111
rect 709 8094 730 8097
rect 644 8091 730 8094
rect 18722 8094 18743 8097
rect 18763 8094 18782 8114
rect 18802 8094 18808 8114
rect 18722 8091 18808 8094
rect 944 8079 1195 8083
rect 944 8059 950 8079
rect 970 8059 989 8079
rect 1009 8059 1028 8079
rect 1048 8059 1067 8079
rect 1087 8059 1195 8079
rect 944 8055 1195 8059
rect 18263 8079 18508 8083
rect 18263 8059 18365 8079
rect 18385 8059 18404 8079
rect 18424 8059 18443 8079
rect 18463 8059 18482 8079
rect 18502 8059 18508 8079
rect 18263 8055 18508 8059
rect 246 7985 252 8011
rect 427 7985 433 8011
rect 18839 7985 18845 8011
rect 19020 7985 19026 8011
rect 755 7908 1195 7912
rect 755 7888 761 7908
rect 781 7888 800 7908
rect 820 7888 839 7908
rect 859 7888 878 7908
rect 898 7888 1195 7908
rect 755 7884 1195 7888
rect 18263 7908 18698 7912
rect 18263 7888 18554 7908
rect 18574 7888 18593 7908
rect 18613 7888 18632 7908
rect 18652 7888 18671 7908
rect 18691 7888 18698 7908
rect 18263 7884 18698 7888
rect 536 7877 570 7880
rect 536 7860 544 7877
rect 561 7870 570 7877
rect 561 7860 1195 7870
rect 536 7856 1195 7860
rect 21346 7828 21762 7834
rect 18550 7776 19272 7783
rect 522 7741 1195 7755
rect 18550 7748 18565 7776
rect 18593 7748 18612 7776
rect 18640 7748 18659 7776
rect 18687 7769 19272 7776
rect 18687 7748 19093 7769
rect 18550 7737 19093 7748
rect 19125 7737 19137 7769
rect 19169 7737 19181 7769
rect 19213 7737 19225 7769
rect 19257 7737 19272 7769
rect 21346 7747 21637 7828
rect 21756 7747 21762 7828
rect 21346 7742 21762 7747
rect 18550 7729 19272 7737
rect 522 7700 1195 7714
rect 18550 7701 18565 7729
rect 18593 7701 18612 7729
rect 18640 7701 18659 7729
rect 18687 7724 19272 7729
rect 18687 7701 19093 7724
rect 18550 7692 19093 7701
rect 19125 7692 19137 7724
rect 19169 7692 19181 7724
rect 19213 7692 19225 7724
rect 19257 7692 19272 7724
rect 590 7683 1195 7686
rect 590 7666 598 7683
rect 615 7672 1195 7683
rect 18550 7682 19272 7692
rect 615 7666 624 7672
rect 590 7662 624 7666
rect 18550 7654 18565 7682
rect 18593 7654 18612 7682
rect 18640 7654 18659 7682
rect 18687 7679 19272 7682
rect 18687 7654 19093 7679
rect 18550 7647 19093 7654
rect 19125 7647 19137 7679
rect 19169 7647 19181 7679
rect 19213 7647 19225 7679
rect 19257 7647 19272 7679
rect 18550 7643 19272 7647
rect 21630 7625 21762 7638
rect 644 7612 730 7615
rect 644 7592 650 7612
rect 670 7592 689 7612
rect 709 7609 730 7612
rect 18722 7612 18808 7615
rect 18722 7609 18743 7612
rect 709 7595 1195 7609
rect 18263 7595 18743 7609
rect 709 7592 730 7595
rect 644 7589 730 7592
rect 18722 7592 18743 7595
rect 18763 7592 18782 7612
rect 18802 7592 18808 7612
rect 18722 7589 18808 7592
rect 944 7577 1195 7581
rect 246 7545 252 7571
rect 427 7545 433 7571
rect 944 7557 950 7577
rect 970 7557 989 7577
rect 1009 7557 1028 7577
rect 1048 7557 1067 7577
rect 1087 7557 1195 7577
rect 944 7553 1195 7557
rect 18263 7577 18508 7581
rect 18263 7557 18365 7577
rect 18385 7557 18404 7577
rect 18424 7557 18443 7577
rect 18463 7557 18482 7577
rect 18502 7557 18508 7577
rect 18263 7553 18508 7557
rect 18839 7545 18845 7571
rect 19020 7545 19026 7571
rect 21630 7419 21643 7625
rect 21749 7419 21762 7625
rect 755 7406 1195 7410
rect 755 7386 761 7406
rect 781 7386 800 7406
rect 820 7386 839 7406
rect 859 7386 878 7406
rect 898 7386 1195 7406
rect 755 7382 1195 7386
rect 18263 7406 18698 7410
rect 21630 7407 21762 7419
rect 18263 7386 18554 7406
rect 18574 7386 18593 7406
rect 18613 7386 18632 7406
rect 18652 7386 18671 7406
rect 18691 7386 18698 7406
rect 18263 7382 18698 7386
rect 21346 7394 21514 7403
rect 536 7375 570 7378
rect 536 7358 544 7375
rect 561 7368 570 7375
rect 561 7358 1195 7368
rect 536 7354 1195 7358
rect 18362 7321 19033 7322
rect 18362 7314 19034 7321
rect 18362 7286 18376 7314
rect 18404 7286 18423 7314
rect 18451 7286 18470 7314
rect 18498 7308 19034 7314
rect 21346 7319 21397 7394
rect 21503 7319 21514 7394
rect 21346 7312 21514 7319
rect 18498 7286 18855 7308
rect 18362 7276 18855 7286
rect 18887 7276 18899 7308
rect 18931 7276 18943 7308
rect 18975 7276 18987 7308
rect 19019 7276 19034 7308
rect 18362 7267 19034 7276
rect 522 7239 1195 7253
rect 18362 7239 18376 7267
rect 18404 7239 18423 7267
rect 18451 7239 18470 7267
rect 18498 7263 19034 7267
rect 18498 7239 18855 7263
rect 18362 7231 18855 7239
rect 18887 7231 18899 7263
rect 18931 7231 18943 7263
rect 18975 7231 18987 7263
rect 19019 7231 19034 7263
rect 18362 7220 19034 7231
rect 522 7198 1195 7212
rect 18362 7192 18376 7220
rect 18404 7192 18423 7220
rect 18451 7192 18470 7220
rect 18498 7218 19034 7220
rect 18498 7192 18855 7218
rect 18362 7186 18855 7192
rect 18887 7186 18899 7218
rect 18931 7186 18943 7218
rect 18975 7186 18987 7218
rect 19019 7186 19034 7218
rect 590 7181 1195 7184
rect 18362 7183 19034 7186
rect 590 7164 598 7181
rect 615 7170 1195 7181
rect 615 7164 624 7170
rect 590 7160 624 7164
rect 246 7105 252 7131
rect 427 7105 433 7131
rect 644 7110 730 7113
rect 644 7090 650 7110
rect 670 7090 689 7110
rect 709 7107 730 7110
rect 18722 7110 18808 7113
rect 18722 7107 18743 7110
rect 709 7093 1195 7107
rect 18263 7093 18743 7107
rect 709 7090 730 7093
rect 644 7087 730 7090
rect 18722 7090 18743 7093
rect 18763 7090 18782 7110
rect 18802 7090 18808 7110
rect 18839 7105 18845 7131
rect 19020 7105 19026 7131
rect 21346 7123 21514 7132
rect 18722 7087 18808 7090
rect 944 7075 1195 7079
rect 944 7055 950 7075
rect 970 7055 989 7075
rect 1009 7055 1028 7075
rect 1048 7055 1067 7075
rect 1087 7055 1195 7075
rect 944 7051 1195 7055
rect 18263 7075 18508 7079
rect 18263 7055 18365 7075
rect 18385 7055 18404 7075
rect 18424 7055 18443 7075
rect 18463 7055 18482 7075
rect 18502 7055 18508 7075
rect 18263 7051 18508 7055
rect 21346 7048 21397 7123
rect 21503 7048 21514 7123
rect 21346 7041 21514 7048
rect 755 6904 1195 6908
rect 755 6884 761 6904
rect 781 6884 800 6904
rect 820 6884 839 6904
rect 859 6884 878 6904
rect 898 6884 1195 6904
rect 755 6880 1195 6884
rect 18263 6904 18698 6908
rect 18263 6884 18554 6904
rect 18574 6884 18593 6904
rect 18613 6884 18632 6904
rect 18652 6884 18671 6904
rect 18691 6884 18698 6904
rect 18263 6880 18698 6884
rect 536 6873 570 6876
rect 536 6856 544 6873
rect 561 6866 570 6873
rect 561 6856 1195 6866
rect 536 6852 1195 6856
rect 21346 6845 21514 6854
rect 18549 6811 19271 6818
rect 18549 6783 18564 6811
rect 18592 6783 18611 6811
rect 18639 6783 18658 6811
rect 18686 6804 19271 6811
rect 18686 6783 19092 6804
rect 18549 6772 19092 6783
rect 19124 6772 19136 6804
rect 19168 6772 19180 6804
rect 19212 6772 19224 6804
rect 19256 6772 19271 6804
rect 18549 6764 19271 6772
rect 522 6737 1195 6751
rect 18549 6736 18564 6764
rect 18592 6736 18611 6764
rect 18639 6736 18658 6764
rect 18686 6759 19271 6764
rect 21346 6770 21397 6845
rect 21503 6770 21514 6845
rect 21346 6763 21514 6770
rect 18686 6736 19092 6759
rect 18549 6727 19092 6736
rect 19124 6727 19136 6759
rect 19168 6727 19180 6759
rect 19212 6727 19224 6759
rect 19256 6727 19271 6759
rect 18549 6717 19271 6727
rect 522 6696 1195 6710
rect 246 6665 252 6691
rect 427 6665 433 6691
rect 18549 6689 18564 6717
rect 18592 6689 18611 6717
rect 18639 6689 18658 6717
rect 18686 6714 19271 6717
rect 18686 6689 19092 6714
rect 18549 6682 19092 6689
rect 19124 6682 19136 6714
rect 19168 6682 19180 6714
rect 19212 6682 19224 6714
rect 19256 6682 19271 6714
rect 590 6679 1195 6682
rect 590 6662 598 6679
rect 615 6668 1195 6679
rect 18549 6678 19271 6682
rect 21630 6746 21762 6759
rect 615 6662 624 6668
rect 590 6658 624 6662
rect 644 6608 730 6611
rect 644 6588 650 6608
rect 670 6588 689 6608
rect 709 6605 730 6608
rect 18722 6608 18808 6611
rect 18722 6605 18743 6608
rect 709 6591 1195 6605
rect 18263 6591 18743 6605
rect 709 6588 730 6591
rect 644 6585 730 6588
rect 18722 6588 18743 6591
rect 18763 6588 18782 6608
rect 18802 6588 18808 6608
rect 18722 6585 18808 6588
rect 944 6573 1195 6577
rect 944 6553 950 6573
rect 970 6553 989 6573
rect 1009 6553 1028 6573
rect 1048 6553 1067 6573
rect 1087 6553 1195 6573
rect 944 6549 1195 6553
rect 18263 6573 18508 6577
rect 18263 6553 18365 6573
rect 18385 6553 18404 6573
rect 18424 6553 18443 6573
rect 18463 6553 18482 6573
rect 18502 6553 18508 6573
rect 18263 6549 18508 6553
rect 21630 6540 21643 6746
rect 21749 6540 21762 6746
rect 21630 6528 21762 6540
rect 755 6402 1195 6406
rect 755 6382 761 6402
rect 781 6382 800 6402
rect 820 6382 839 6402
rect 859 6382 878 6402
rect 898 6382 1195 6402
rect 755 6378 1195 6382
rect 18263 6402 18698 6406
rect 18263 6382 18554 6402
rect 18574 6382 18593 6402
rect 18613 6382 18632 6402
rect 18652 6382 18671 6402
rect 18691 6382 18698 6402
rect 18263 6378 18698 6382
rect 536 6371 570 6374
rect 536 6354 544 6371
rect 561 6364 570 6371
rect 561 6354 1195 6364
rect 536 6350 1195 6354
rect 18363 6359 19034 6360
rect 18363 6352 19035 6359
rect 18363 6324 18377 6352
rect 18405 6324 18424 6352
rect 18452 6324 18471 6352
rect 18499 6346 19035 6352
rect 18499 6324 18856 6346
rect 18363 6314 18856 6324
rect 18888 6314 18900 6346
rect 18932 6314 18944 6346
rect 18976 6314 18988 6346
rect 19020 6314 19035 6346
rect 18363 6305 19035 6314
rect 18363 6277 18377 6305
rect 18405 6277 18424 6305
rect 18452 6277 18471 6305
rect 18499 6301 19035 6305
rect 18499 6277 18856 6301
rect 18363 6269 18856 6277
rect 18888 6269 18900 6301
rect 18932 6269 18944 6301
rect 18976 6269 18988 6301
rect 19020 6269 19035 6301
rect 18363 6258 19035 6269
rect 246 6225 252 6251
rect 427 6225 433 6251
rect 522 6235 1195 6249
rect 18363 6230 18377 6258
rect 18405 6230 18424 6258
rect 18452 6230 18471 6258
rect 18499 6256 19035 6258
rect 18499 6251 18856 6256
rect 18888 6251 18900 6256
rect 18932 6251 18944 6256
rect 18976 6251 18988 6256
rect 18499 6230 18845 6251
rect 18363 6225 18845 6230
rect 18363 6224 18856 6225
rect 18888 6224 18900 6225
rect 18932 6224 18944 6225
rect 18976 6224 18988 6225
rect 19020 6224 19035 6256
rect 18363 6220 19035 6224
rect 21346 6273 21762 6279
rect 522 6194 1195 6208
rect 21346 6192 21637 6273
rect 21756 6192 21762 6273
rect 21346 6187 21762 6192
rect 590 6177 1195 6180
rect 590 6160 598 6177
rect 615 6166 1195 6177
rect 615 6160 624 6166
rect 590 6156 624 6160
rect 644 6106 730 6109
rect 644 6086 650 6106
rect 670 6086 689 6106
rect 709 6103 730 6106
rect 18722 6106 18808 6109
rect 18722 6103 18743 6106
rect 709 6089 1195 6103
rect 18263 6089 18743 6103
rect 709 6086 730 6089
rect 644 6083 730 6086
rect 18722 6086 18743 6089
rect 18763 6086 18782 6106
rect 18802 6086 18808 6106
rect 18722 6083 18808 6086
rect 944 6071 1195 6075
rect 944 6051 950 6071
rect 970 6051 989 6071
rect 1009 6051 1028 6071
rect 1048 6051 1067 6071
rect 1087 6051 1195 6071
rect 944 6047 1195 6051
rect 18263 6071 18508 6075
rect 18263 6051 18365 6071
rect 18385 6051 18404 6071
rect 18424 6051 18443 6071
rect 18463 6051 18482 6071
rect 18502 6051 18508 6071
rect 18263 6047 18508 6051
rect 755 5900 1195 5904
rect 755 5880 761 5900
rect 781 5880 800 5900
rect 820 5880 839 5900
rect 859 5880 878 5900
rect 898 5880 1195 5900
rect 755 5876 1195 5880
rect 18263 5900 18698 5904
rect 18263 5880 18554 5900
rect 18574 5880 18593 5900
rect 18613 5880 18632 5900
rect 18652 5880 18671 5900
rect 18691 5880 18698 5900
rect 18263 5876 18698 5880
rect 536 5869 570 5872
rect 536 5852 544 5869
rect 561 5862 570 5869
rect 561 5852 1195 5862
rect 536 5848 1195 5852
rect 21346 5828 21762 5834
rect 246 5785 252 5811
rect 427 5785 433 5811
rect 18550 5803 19272 5810
rect 18550 5775 18565 5803
rect 18593 5775 18612 5803
rect 18640 5775 18659 5803
rect 18687 5796 19272 5803
rect 18687 5775 19093 5796
rect 18550 5764 19093 5775
rect 19125 5764 19137 5796
rect 19169 5764 19181 5796
rect 19213 5764 19225 5796
rect 19257 5764 19272 5796
rect 18550 5756 19272 5764
rect 522 5733 1195 5747
rect 18550 5728 18565 5756
rect 18593 5728 18612 5756
rect 18640 5728 18659 5756
rect 18687 5751 19272 5756
rect 18687 5728 19093 5751
rect 18550 5719 19093 5728
rect 19125 5719 19137 5751
rect 19169 5719 19181 5751
rect 19213 5719 19225 5751
rect 19257 5719 19272 5751
rect 21346 5747 21637 5828
rect 21756 5747 21762 5828
rect 21346 5742 21762 5747
rect 18550 5709 19272 5719
rect 522 5692 1195 5706
rect 18550 5681 18565 5709
rect 18593 5681 18612 5709
rect 18640 5681 18659 5709
rect 18687 5706 19272 5709
rect 18687 5681 19093 5706
rect 590 5675 1195 5678
rect 590 5658 598 5675
rect 615 5664 1195 5675
rect 18550 5674 19093 5681
rect 19125 5674 19137 5706
rect 19169 5674 19181 5706
rect 19213 5674 19225 5706
rect 19257 5674 19272 5706
rect 18550 5670 19272 5674
rect 615 5658 624 5664
rect 590 5654 624 5658
rect 21630 5625 21762 5638
rect 644 5604 730 5607
rect 644 5584 650 5604
rect 670 5584 689 5604
rect 709 5601 730 5604
rect 18722 5604 18808 5607
rect 18722 5601 18743 5604
rect 709 5587 1195 5601
rect 18263 5587 18743 5601
rect 709 5584 730 5587
rect 644 5581 730 5584
rect 18722 5584 18743 5587
rect 18763 5584 18782 5604
rect 18802 5584 18808 5604
rect 18722 5581 18808 5584
rect 944 5569 1195 5573
rect 944 5549 950 5569
rect 970 5549 989 5569
rect 1009 5549 1028 5569
rect 1048 5549 1067 5569
rect 1087 5549 1195 5569
rect 944 5545 1195 5549
rect 18263 5569 18508 5573
rect 18263 5549 18365 5569
rect 18385 5549 18404 5569
rect 18424 5549 18443 5569
rect 18463 5549 18482 5569
rect 18502 5549 18508 5569
rect 18263 5545 18508 5549
rect 21630 5419 21643 5625
rect 21749 5419 21762 5625
rect 21630 5407 21762 5419
rect 755 5398 1195 5402
rect 755 5378 761 5398
rect 781 5378 800 5398
rect 820 5378 839 5398
rect 859 5378 878 5398
rect 898 5378 1195 5398
rect 755 5374 1195 5378
rect 18263 5398 18698 5402
rect 18263 5378 18554 5398
rect 18574 5378 18593 5398
rect 18613 5378 18632 5398
rect 18652 5378 18671 5398
rect 18691 5378 18698 5398
rect 18263 5374 18698 5378
rect 21346 5394 21514 5403
rect 246 5345 252 5371
rect 427 5345 433 5371
rect 536 5367 570 5370
rect 536 5350 544 5367
rect 561 5360 570 5367
rect 561 5350 1195 5360
rect 536 5346 1195 5350
rect 18839 5345 18845 5371
rect 19020 5345 19026 5371
rect 21346 5319 21397 5394
rect 21503 5319 21514 5394
rect 21346 5312 21514 5319
rect 18362 5296 19033 5297
rect 18362 5289 19034 5296
rect 18362 5261 18376 5289
rect 18404 5261 18423 5289
rect 18451 5261 18470 5289
rect 18498 5283 19034 5289
rect 18498 5261 18855 5283
rect 18362 5251 18855 5261
rect 18887 5251 18899 5283
rect 18931 5251 18943 5283
rect 18975 5251 18987 5283
rect 19019 5251 19034 5283
rect 522 5231 1195 5245
rect 18362 5242 19034 5251
rect 18362 5214 18376 5242
rect 18404 5214 18423 5242
rect 18451 5214 18470 5242
rect 18498 5238 19034 5242
rect 18498 5214 18855 5238
rect 18362 5206 18855 5214
rect 18887 5206 18899 5238
rect 18931 5206 18943 5238
rect 18975 5206 18987 5238
rect 19019 5206 19034 5238
rect 522 5190 1195 5204
rect 18362 5195 19034 5206
rect 590 5173 1195 5176
rect 590 5156 598 5173
rect 615 5162 1195 5173
rect 18362 5167 18376 5195
rect 18404 5167 18423 5195
rect 18451 5167 18470 5195
rect 18498 5193 19034 5195
rect 18498 5167 18855 5193
rect 615 5156 624 5162
rect 18362 5161 18855 5167
rect 18887 5161 18899 5193
rect 18931 5161 18943 5193
rect 18975 5161 18987 5193
rect 19019 5161 19034 5193
rect 18362 5157 19034 5161
rect 590 5152 624 5156
rect 21346 5123 21514 5132
rect 644 5102 730 5105
rect 644 5082 650 5102
rect 670 5082 689 5102
rect 709 5099 730 5102
rect 18722 5102 18808 5105
rect 18722 5099 18743 5102
rect 709 5085 1195 5099
rect 18263 5085 18743 5099
rect 709 5082 730 5085
rect 644 5079 730 5082
rect 18722 5082 18743 5085
rect 18763 5082 18782 5102
rect 18802 5082 18808 5102
rect 18722 5079 18808 5082
rect 944 5067 1195 5071
rect 944 5047 950 5067
rect 970 5047 989 5067
rect 1009 5047 1028 5067
rect 1048 5047 1067 5067
rect 1087 5047 1195 5067
rect 944 5043 1195 5047
rect 18263 5067 18508 5071
rect 18263 5047 18365 5067
rect 18385 5047 18404 5067
rect 18424 5047 18443 5067
rect 18463 5047 18482 5067
rect 18502 5047 18508 5067
rect 18263 5043 18508 5047
rect 21346 5048 21397 5123
rect 21503 5048 21514 5123
rect 21346 5041 21514 5048
rect 246 4905 252 4931
rect 427 4905 433 4931
rect 18839 4905 18845 4931
rect 19020 4905 19026 4931
rect 755 4896 1195 4900
rect 755 4876 761 4896
rect 781 4876 800 4896
rect 820 4876 839 4896
rect 859 4876 878 4896
rect 898 4876 1195 4896
rect 755 4872 1195 4876
rect 18263 4896 18698 4900
rect 18263 4876 18554 4896
rect 18574 4876 18593 4896
rect 18613 4876 18632 4896
rect 18652 4876 18671 4896
rect 18691 4876 18698 4896
rect 18263 4872 18698 4876
rect 536 4865 570 4868
rect 536 4848 544 4865
rect 561 4858 570 4865
rect 561 4848 1195 4858
rect 536 4844 1195 4848
rect 21346 4845 21514 4854
rect 18550 4802 19272 4809
rect 18550 4774 18565 4802
rect 18593 4774 18612 4802
rect 18640 4774 18659 4802
rect 18687 4795 19272 4802
rect 18687 4774 19093 4795
rect 18550 4763 19093 4774
rect 19125 4763 19137 4795
rect 19169 4763 19181 4795
rect 19213 4763 19225 4795
rect 19257 4763 19272 4795
rect 21346 4770 21397 4845
rect 21503 4770 21514 4845
rect 21346 4763 21514 4770
rect 18550 4755 19272 4763
rect 522 4729 1195 4743
rect 18550 4727 18565 4755
rect 18593 4727 18612 4755
rect 18640 4727 18659 4755
rect 18687 4750 19272 4755
rect 18687 4727 19093 4750
rect 18550 4718 19093 4727
rect 19125 4718 19137 4750
rect 19169 4718 19181 4750
rect 19213 4718 19225 4750
rect 19257 4718 19272 4750
rect 18550 4708 19272 4718
rect 522 4688 1195 4702
rect 18550 4680 18565 4708
rect 18593 4680 18612 4708
rect 18640 4680 18659 4708
rect 18687 4705 19272 4708
rect 18687 4680 19093 4705
rect 590 4671 1195 4674
rect 590 4654 598 4671
rect 615 4660 1195 4671
rect 18550 4673 19093 4680
rect 19125 4673 19137 4705
rect 19169 4673 19181 4705
rect 19213 4673 19225 4705
rect 19257 4673 19272 4705
rect 18550 4669 19272 4673
rect 21630 4746 21762 4759
rect 615 4654 624 4660
rect 590 4650 624 4654
rect 644 4600 730 4603
rect 644 4580 650 4600
rect 670 4580 689 4600
rect 709 4597 730 4600
rect 18722 4600 18808 4603
rect 18722 4597 18743 4600
rect 709 4583 1195 4597
rect 18263 4583 18743 4597
rect 709 4580 730 4583
rect 644 4577 730 4580
rect 18722 4580 18743 4583
rect 18763 4580 18782 4600
rect 18802 4580 18808 4600
rect 18722 4577 18808 4580
rect 944 4565 1195 4569
rect 944 4545 950 4565
rect 970 4545 989 4565
rect 1009 4545 1028 4565
rect 1048 4545 1067 4565
rect 1087 4545 1195 4565
rect 944 4541 1195 4545
rect 18263 4565 18508 4569
rect 18263 4545 18365 4565
rect 18385 4545 18404 4565
rect 18424 4545 18443 4565
rect 18463 4545 18482 4565
rect 18502 4545 18508 4565
rect 18263 4541 18508 4545
rect 21630 4540 21643 4746
rect 21749 4540 21762 4746
rect 21630 4528 21762 4540
rect 246 4465 252 4491
rect 427 4465 433 4491
rect 18839 4465 18845 4491
rect 19020 4465 19026 4491
rect 755 4394 1195 4398
rect 755 4374 761 4394
rect 781 4374 800 4394
rect 820 4374 839 4394
rect 859 4374 878 4394
rect 898 4374 1195 4394
rect 755 4370 1195 4374
rect 18263 4394 18698 4398
rect 18263 4374 18554 4394
rect 18574 4374 18593 4394
rect 18613 4374 18632 4394
rect 18652 4374 18671 4394
rect 18691 4374 18698 4394
rect 18263 4370 18698 4374
rect 536 4363 570 4366
rect 536 4346 544 4363
rect 561 4356 570 4363
rect 561 4346 1195 4356
rect 536 4342 1195 4346
rect 18363 4308 19034 4309
rect 18363 4301 19035 4308
rect 18363 4273 18377 4301
rect 18405 4273 18424 4301
rect 18452 4273 18471 4301
rect 18499 4295 19035 4301
rect 18499 4273 18856 4295
rect 18363 4263 18856 4273
rect 18888 4263 18900 4295
rect 18932 4263 18944 4295
rect 18976 4263 18988 4295
rect 19020 4263 19035 4295
rect 18363 4254 19035 4263
rect 522 4227 1195 4241
rect 18363 4226 18377 4254
rect 18405 4226 18424 4254
rect 18452 4226 18471 4254
rect 18499 4250 19035 4254
rect 18499 4226 18856 4250
rect 18363 4218 18856 4226
rect 18888 4218 18900 4250
rect 18932 4218 18944 4250
rect 18976 4218 18988 4250
rect 19020 4218 19035 4250
rect 18363 4207 19035 4218
rect 522 4186 1195 4200
rect 18363 4179 18377 4207
rect 18405 4179 18424 4207
rect 18452 4179 18471 4207
rect 18499 4205 19035 4207
rect 18499 4179 18856 4205
rect 18363 4173 18856 4179
rect 18888 4173 18900 4205
rect 18932 4173 18944 4205
rect 18976 4173 18988 4205
rect 19020 4173 19035 4205
rect 21346 4273 21762 4279
rect 21346 4192 21637 4273
rect 21756 4192 21762 4273
rect 21346 4187 21762 4192
rect 590 4169 1195 4172
rect 18363 4169 19035 4173
rect 590 4152 598 4169
rect 615 4158 1195 4169
rect 615 4152 624 4158
rect 590 4148 624 4152
rect 644 4098 730 4101
rect 644 4078 650 4098
rect 670 4078 689 4098
rect 709 4095 730 4098
rect 18722 4098 18808 4101
rect 18722 4095 18743 4098
rect 709 4081 1195 4095
rect 18263 4081 18743 4095
rect 709 4078 730 4081
rect 644 4075 730 4078
rect 18722 4078 18743 4081
rect 18763 4078 18782 4098
rect 18802 4078 18808 4098
rect 18722 4075 18808 4078
rect 944 4063 1195 4067
rect 246 4025 252 4051
rect 427 4025 433 4051
rect 944 4043 950 4063
rect 970 4043 989 4063
rect 1009 4043 1028 4063
rect 1048 4043 1067 4063
rect 1087 4043 1195 4063
rect 944 4039 1195 4043
rect 18263 4063 18508 4067
rect 18263 4043 18365 4063
rect 18385 4043 18404 4063
rect 18424 4043 18443 4063
rect 18463 4043 18482 4063
rect 18502 4043 18508 4063
rect 18263 4039 18508 4043
rect 18839 4025 18845 4051
rect 19020 4025 19026 4051
rect 755 3892 1195 3896
rect 755 3872 761 3892
rect 781 3872 800 3892
rect 820 3872 839 3892
rect 859 3872 878 3892
rect 898 3872 1195 3892
rect 755 3868 1195 3872
rect 18263 3892 18698 3896
rect 18263 3872 18554 3892
rect 18574 3872 18593 3892
rect 18613 3872 18632 3892
rect 18652 3872 18671 3892
rect 18691 3872 18698 3892
rect 18263 3868 18698 3872
rect 536 3861 570 3864
rect 536 3844 544 3861
rect 561 3854 570 3861
rect 561 3844 1195 3854
rect 536 3840 1195 3844
rect 21346 3828 21762 3834
rect 18549 3803 19271 3810
rect 18549 3775 18564 3803
rect 18592 3775 18611 3803
rect 18639 3775 18658 3803
rect 18686 3796 19271 3803
rect 18686 3775 19092 3796
rect 18549 3764 19092 3775
rect 19124 3764 19136 3796
rect 19168 3764 19180 3796
rect 19212 3764 19224 3796
rect 19256 3764 19271 3796
rect 18549 3756 19271 3764
rect 522 3725 1195 3739
rect 18549 3728 18564 3756
rect 18592 3728 18611 3756
rect 18639 3728 18658 3756
rect 18686 3751 19271 3756
rect 18686 3728 19092 3751
rect 18549 3719 19092 3728
rect 19124 3719 19136 3751
rect 19168 3719 19180 3751
rect 19212 3719 19224 3751
rect 19256 3719 19271 3751
rect 21346 3747 21637 3828
rect 21756 3747 21762 3828
rect 21346 3742 21762 3747
rect 18549 3709 19271 3719
rect 522 3684 1195 3698
rect 18549 3681 18564 3709
rect 18592 3681 18611 3709
rect 18639 3681 18658 3709
rect 18686 3706 19271 3709
rect 18686 3681 19092 3706
rect 18549 3674 19092 3681
rect 19124 3674 19136 3706
rect 19168 3674 19180 3706
rect 19212 3674 19224 3706
rect 19256 3674 19271 3706
rect 18549 3670 19271 3674
rect 590 3667 1195 3670
rect 590 3650 598 3667
rect 615 3656 1195 3667
rect 615 3650 624 3656
rect 590 3646 624 3650
rect 21630 3625 21762 3638
rect 246 3585 252 3611
rect 427 3585 433 3611
rect 644 3596 730 3599
rect 644 3576 650 3596
rect 670 3576 689 3596
rect 709 3593 730 3596
rect 18722 3596 18808 3599
rect 18722 3593 18743 3596
rect 709 3579 1195 3593
rect 18263 3579 18743 3593
rect 709 3576 730 3579
rect 644 3573 730 3576
rect 18722 3576 18743 3579
rect 18763 3576 18782 3596
rect 18802 3576 18808 3596
rect 18839 3585 18845 3611
rect 19020 3585 19026 3611
rect 18722 3573 18808 3576
rect 944 3561 1195 3565
rect 944 3541 950 3561
rect 970 3541 989 3561
rect 1009 3541 1028 3561
rect 1048 3541 1067 3561
rect 1087 3541 1195 3561
rect 944 3537 1195 3541
rect 18263 3561 18508 3565
rect 18263 3541 18365 3561
rect 18385 3541 18404 3561
rect 18424 3541 18443 3561
rect 18463 3541 18482 3561
rect 18502 3541 18508 3561
rect 18263 3537 18508 3541
rect 21630 3419 21643 3625
rect 21749 3419 21762 3625
rect 21630 3407 21762 3419
rect 21346 3394 21514 3403
rect 755 3390 1195 3394
rect 755 3370 761 3390
rect 781 3370 800 3390
rect 820 3370 839 3390
rect 859 3370 878 3390
rect 898 3370 1195 3390
rect 755 3366 1195 3370
rect 18263 3390 18698 3394
rect 18263 3370 18554 3390
rect 18574 3370 18593 3390
rect 18613 3370 18632 3390
rect 18652 3370 18671 3390
rect 18691 3370 18698 3390
rect 18263 3366 18698 3370
rect 536 3359 570 3362
rect 536 3342 544 3359
rect 561 3352 570 3359
rect 561 3342 1195 3352
rect 536 3338 1195 3342
rect 21346 3319 21397 3394
rect 21503 3319 21514 3394
rect 21346 3312 21514 3319
rect 18363 3286 19034 3287
rect 18363 3279 19035 3286
rect 18363 3251 18377 3279
rect 18405 3251 18424 3279
rect 18452 3251 18471 3279
rect 18499 3273 19035 3279
rect 18499 3251 18856 3273
rect 18363 3241 18856 3251
rect 18888 3241 18900 3273
rect 18932 3241 18944 3273
rect 18976 3241 18988 3273
rect 19020 3241 19035 3273
rect 522 3223 1195 3237
rect 18363 3232 19035 3241
rect 18363 3204 18377 3232
rect 18405 3204 18424 3232
rect 18452 3204 18471 3232
rect 18499 3228 19035 3232
rect 18499 3204 18856 3228
rect 18363 3196 18856 3204
rect 18888 3196 18900 3228
rect 18932 3196 18944 3228
rect 18976 3196 18988 3228
rect 19020 3196 19035 3228
rect 522 3182 1195 3196
rect 18363 3185 19035 3196
rect 246 3145 252 3171
rect 427 3145 433 3171
rect 590 3165 1195 3168
rect 590 3148 598 3165
rect 615 3154 1195 3165
rect 18363 3157 18377 3185
rect 18405 3157 18424 3185
rect 18452 3157 18471 3185
rect 18499 3183 19035 3185
rect 18499 3171 18856 3183
rect 18888 3171 18900 3183
rect 18932 3171 18944 3183
rect 18976 3171 18988 3183
rect 18499 3157 18845 3171
rect 615 3148 624 3154
rect 590 3144 624 3148
rect 18363 3147 18845 3157
rect 18839 3145 18845 3147
rect 19020 3147 19035 3183
rect 19020 3145 19026 3147
rect 21346 3123 21514 3132
rect 644 3094 730 3097
rect 644 3074 650 3094
rect 670 3074 689 3094
rect 709 3091 730 3094
rect 18722 3094 18808 3097
rect 18722 3091 18743 3094
rect 709 3077 1195 3091
rect 18263 3077 18743 3091
rect 709 3074 730 3077
rect 644 3071 730 3074
rect 18722 3074 18743 3077
rect 18763 3074 18782 3094
rect 18802 3074 18808 3094
rect 18722 3071 18808 3074
rect 944 3059 1195 3063
rect 944 3039 950 3059
rect 970 3039 989 3059
rect 1009 3039 1028 3059
rect 1048 3039 1067 3059
rect 1087 3039 1195 3059
rect 944 3035 1195 3039
rect 18263 3059 18508 3063
rect 18263 3039 18365 3059
rect 18385 3039 18404 3059
rect 18424 3039 18443 3059
rect 18463 3039 18482 3059
rect 18502 3039 18508 3059
rect 21346 3048 21397 3123
rect 21503 3048 21514 3123
rect 21346 3041 21514 3048
rect 18263 3035 18508 3039
rect 755 2888 1195 2892
rect 755 2868 761 2888
rect 781 2868 800 2888
rect 820 2868 839 2888
rect 859 2868 878 2888
rect 898 2868 1195 2888
rect 755 2864 1195 2868
rect 18263 2888 18698 2892
rect 18263 2868 18554 2888
rect 18574 2868 18593 2888
rect 18613 2868 18632 2888
rect 18652 2868 18671 2888
rect 18691 2868 18698 2888
rect 18263 2864 18698 2868
rect 536 2857 570 2860
rect 536 2840 544 2857
rect 561 2850 570 2857
rect 561 2840 1195 2850
rect 536 2836 1195 2840
rect 21346 2845 21514 2854
rect 18550 2769 19272 2776
rect 18550 2741 18565 2769
rect 18593 2741 18612 2769
rect 18640 2741 18659 2769
rect 18687 2762 19272 2769
rect 21346 2770 21397 2845
rect 21503 2770 21514 2845
rect 21346 2763 21514 2770
rect 18687 2741 19093 2762
rect 246 2705 252 2731
rect 427 2705 433 2731
rect 522 2721 1195 2735
rect 18550 2730 19093 2741
rect 19125 2730 19137 2762
rect 19169 2730 19181 2762
rect 19213 2730 19225 2762
rect 19257 2730 19272 2762
rect 18550 2722 19272 2730
rect 18550 2694 18565 2722
rect 18593 2694 18612 2722
rect 18640 2694 18659 2722
rect 18687 2717 19272 2722
rect 18687 2694 19093 2717
rect 522 2680 1195 2694
rect 18550 2685 19093 2694
rect 19125 2685 19137 2717
rect 19169 2685 19181 2717
rect 19213 2685 19225 2717
rect 19257 2685 19272 2717
rect 18550 2675 19272 2685
rect 590 2663 1195 2666
rect 590 2646 598 2663
rect 615 2652 1195 2663
rect 615 2646 624 2652
rect 590 2642 624 2646
rect 18550 2647 18565 2675
rect 18593 2647 18612 2675
rect 18640 2647 18659 2675
rect 18687 2672 19272 2675
rect 18687 2647 19093 2672
rect 18550 2640 19093 2647
rect 19125 2640 19137 2672
rect 19169 2640 19181 2672
rect 19213 2640 19225 2672
rect 19257 2640 19272 2672
rect 18550 2636 19272 2640
rect 21630 2746 21762 2759
rect 644 2592 730 2595
rect 644 2572 650 2592
rect 670 2572 689 2592
rect 709 2589 730 2592
rect 18722 2592 18808 2595
rect 18722 2589 18743 2592
rect 709 2575 1195 2589
rect 18263 2575 18743 2589
rect 709 2572 730 2575
rect 644 2569 730 2572
rect 18722 2572 18743 2575
rect 18763 2572 18782 2592
rect 18802 2572 18808 2592
rect 18722 2569 18808 2572
rect 944 2557 1195 2561
rect 944 2537 950 2557
rect 970 2537 989 2557
rect 1009 2537 1028 2557
rect 1048 2537 1067 2557
rect 1087 2537 1195 2557
rect 944 2533 1195 2537
rect 18263 2557 18508 2561
rect 18263 2537 18365 2557
rect 18385 2537 18404 2557
rect 18424 2537 18443 2557
rect 18463 2537 18482 2557
rect 18502 2537 18508 2557
rect 18263 2533 18508 2537
rect 21630 2540 21643 2746
rect 21749 2540 21762 2746
rect 21630 2528 21762 2540
rect 755 2386 1195 2390
rect 755 2366 761 2386
rect 781 2366 800 2386
rect 820 2366 839 2386
rect 859 2366 878 2386
rect 898 2366 1195 2386
rect 755 2362 1195 2366
rect 18263 2386 18698 2390
rect 18263 2366 18554 2386
rect 18574 2366 18593 2386
rect 18613 2366 18632 2386
rect 18652 2366 18671 2386
rect 18691 2366 18698 2386
rect 18263 2362 18698 2366
rect 536 2355 570 2358
rect 536 2338 544 2355
rect 561 2348 570 2355
rect 561 2338 1195 2348
rect 536 2334 1195 2338
rect 246 2265 252 2291
rect 427 2265 433 2291
rect 18839 2290 18845 2291
rect 18362 2282 18845 2290
rect 19020 2290 19026 2291
rect 18362 2254 18377 2282
rect 18405 2254 18424 2282
rect 18452 2254 18471 2282
rect 18499 2265 18845 2282
rect 18499 2254 18856 2265
rect 18362 2244 18856 2254
rect 18888 2244 18900 2265
rect 18932 2244 18944 2265
rect 18976 2244 18988 2265
rect 19020 2244 19034 2290
rect 18362 2235 19034 2244
rect 522 2219 1195 2233
rect 18362 2207 18377 2235
rect 18405 2207 18424 2235
rect 18452 2207 18471 2235
rect 18499 2231 19034 2235
rect 18499 2207 18856 2231
rect 18362 2199 18856 2207
rect 18888 2199 18900 2231
rect 18932 2199 18944 2231
rect 18976 2199 18988 2231
rect 19020 2199 19034 2231
rect 522 2178 1195 2192
rect 18362 2188 19034 2199
rect 590 2161 1195 2164
rect 590 2144 598 2161
rect 615 2150 1195 2161
rect 18362 2160 18377 2188
rect 18405 2160 18424 2188
rect 18452 2160 18471 2188
rect 18499 2186 19034 2188
rect 21346 2273 21762 2279
rect 21346 2192 21637 2273
rect 21756 2192 21762 2273
rect 21346 2187 21762 2192
rect 18499 2160 18856 2186
rect 18362 2154 18856 2160
rect 18888 2154 18900 2186
rect 18932 2154 18944 2186
rect 18976 2154 18988 2186
rect 19020 2154 19034 2186
rect 18362 2150 19034 2154
rect 615 2144 624 2150
rect 590 2140 624 2144
rect 644 2090 730 2093
rect 644 2070 650 2090
rect 670 2070 689 2090
rect 709 2087 730 2090
rect 18722 2090 18808 2093
rect 18722 2087 18743 2090
rect 709 2073 1195 2087
rect 18263 2073 18743 2087
rect 709 2070 730 2073
rect 644 2067 730 2070
rect 18722 2070 18743 2073
rect 18763 2070 18782 2090
rect 18802 2070 18808 2090
rect 18722 2067 18808 2070
rect 944 2055 1195 2059
rect 944 2035 950 2055
rect 970 2035 989 2055
rect 1009 2035 1028 2055
rect 1048 2035 1067 2055
rect 1087 2035 1195 2055
rect 944 2031 1195 2035
rect 18263 2055 18508 2059
rect 18263 2035 18365 2055
rect 18385 2035 18404 2055
rect 18424 2035 18443 2055
rect 18463 2035 18482 2055
rect 18502 2035 18508 2055
rect 18263 2031 18508 2035
rect 755 1884 1195 1888
rect 755 1864 761 1884
rect 781 1864 800 1884
rect 820 1864 839 1884
rect 859 1864 878 1884
rect 898 1864 1195 1884
rect 755 1860 1195 1864
rect 18263 1884 18698 1888
rect 18263 1864 18554 1884
rect 18574 1864 18593 1884
rect 18613 1864 18632 1884
rect 18652 1864 18671 1884
rect 18691 1864 18698 1884
rect 18263 1860 18698 1864
rect 536 1853 570 1856
rect 246 1825 252 1851
rect 427 1825 433 1851
rect 536 1836 544 1853
rect 561 1846 570 1853
rect 561 1836 1195 1846
rect 536 1832 1195 1836
rect 18839 1825 18845 1851
rect 19020 1825 19026 1851
rect 21346 1828 21762 1834
rect 18550 1767 19272 1774
rect 18550 1739 18565 1767
rect 18593 1739 18612 1767
rect 18640 1739 18659 1767
rect 18687 1760 19272 1767
rect 18687 1739 19093 1760
rect 522 1717 1195 1731
rect 18550 1728 19093 1739
rect 19125 1728 19137 1760
rect 19169 1728 19181 1760
rect 19213 1728 19225 1760
rect 19257 1728 19272 1760
rect 21346 1747 21637 1828
rect 21756 1747 21762 1828
rect 21346 1742 21762 1747
rect 18550 1720 19272 1728
rect 18550 1692 18565 1720
rect 18593 1692 18612 1720
rect 18640 1692 18659 1720
rect 18687 1715 19272 1720
rect 18687 1692 19093 1715
rect 522 1676 1195 1690
rect 18550 1683 19093 1692
rect 19125 1683 19137 1715
rect 19169 1683 19181 1715
rect 19213 1683 19225 1715
rect 19257 1683 19272 1715
rect 18550 1673 19272 1683
rect 590 1659 1195 1662
rect 590 1642 598 1659
rect 615 1648 1195 1659
rect 615 1642 624 1648
rect 590 1638 624 1642
rect 18550 1645 18565 1673
rect 18593 1645 18612 1673
rect 18640 1645 18659 1673
rect 18687 1670 19272 1673
rect 18687 1645 19093 1670
rect 18550 1638 19093 1645
rect 19125 1638 19137 1670
rect 19169 1638 19181 1670
rect 19213 1638 19225 1670
rect 19257 1638 19272 1670
rect 18550 1634 19272 1638
rect 21630 1625 21762 1638
rect 644 1588 730 1591
rect 644 1568 650 1588
rect 670 1568 689 1588
rect 709 1585 730 1588
rect 18722 1588 18808 1591
rect 18722 1585 18743 1588
rect 709 1571 1195 1585
rect 18263 1571 18743 1585
rect 709 1568 730 1571
rect 644 1565 730 1568
rect 18722 1568 18743 1571
rect 18763 1568 18782 1588
rect 18802 1568 18808 1588
rect 18722 1565 18808 1568
rect 944 1553 1195 1557
rect 944 1533 950 1553
rect 970 1533 989 1553
rect 1009 1533 1028 1553
rect 1048 1533 1067 1553
rect 1087 1533 1195 1553
rect 944 1529 1195 1533
rect 18263 1553 18508 1557
rect 18263 1533 18365 1553
rect 18385 1533 18404 1553
rect 18424 1533 18443 1553
rect 18463 1533 18482 1553
rect 18502 1533 18508 1553
rect 18263 1529 18508 1533
rect 21630 1419 21643 1625
rect 21749 1419 21762 1625
rect 246 1385 252 1411
rect 427 1385 433 1411
rect 755 1382 1195 1386
rect 755 1362 761 1382
rect 781 1362 800 1382
rect 820 1362 839 1382
rect 859 1362 878 1382
rect 898 1362 1195 1382
rect 755 1358 1195 1362
rect 18263 1382 18698 1386
rect 18839 1385 18845 1411
rect 19020 1385 19026 1411
rect 21630 1407 21762 1419
rect 21346 1394 21514 1403
rect 18263 1362 18554 1382
rect 18574 1362 18593 1382
rect 18613 1362 18632 1382
rect 18652 1362 18671 1382
rect 18691 1362 18698 1382
rect 18263 1358 18698 1362
rect 536 1351 570 1354
rect 536 1334 544 1351
rect 561 1344 570 1351
rect 561 1334 1195 1344
rect 536 1330 1195 1334
rect 21346 1319 21397 1394
rect 21503 1319 21514 1394
rect 21346 1312 21514 1319
rect 18361 1289 19032 1290
rect 18361 1282 19033 1289
rect 18361 1254 18375 1282
rect 18403 1254 18422 1282
rect 18450 1254 18469 1282
rect 18497 1276 19033 1282
rect 18497 1254 18854 1276
rect 18361 1244 18854 1254
rect 18886 1244 18898 1276
rect 18930 1244 18942 1276
rect 18974 1244 18986 1276
rect 19018 1244 19033 1276
rect 18361 1235 19033 1244
rect 522 1215 1195 1229
rect 18361 1207 18375 1235
rect 18403 1207 18422 1235
rect 18450 1207 18469 1235
rect 18497 1231 19033 1235
rect 18497 1207 18854 1231
rect 18361 1199 18854 1207
rect 18886 1199 18898 1231
rect 18930 1199 18942 1231
rect 18974 1199 18986 1231
rect 19018 1199 19033 1231
rect 18361 1188 19033 1199
rect 522 1174 1195 1188
rect 18361 1160 18375 1188
rect 18403 1160 18422 1188
rect 18450 1160 18469 1188
rect 18497 1186 19033 1188
rect 18497 1160 18854 1186
rect 590 1157 1195 1160
rect 590 1140 598 1157
rect 615 1146 1195 1157
rect 18361 1154 18854 1160
rect 18886 1154 18898 1186
rect 18930 1154 18942 1186
rect 18974 1154 18986 1186
rect 19018 1154 19033 1186
rect 18361 1150 19033 1154
rect 615 1140 624 1146
rect 590 1136 624 1140
rect 21346 1123 21514 1132
rect 644 1086 730 1089
rect 644 1066 650 1086
rect 670 1066 689 1086
rect 709 1083 730 1086
rect 18722 1086 18808 1089
rect 18722 1083 18743 1086
rect 709 1069 1195 1083
rect 18263 1069 18743 1083
rect 709 1066 730 1069
rect 644 1063 730 1066
rect 18722 1066 18743 1069
rect 18763 1066 18782 1086
rect 18802 1066 18808 1086
rect 18722 1063 18808 1066
rect 944 1051 1195 1055
rect 944 1031 950 1051
rect 970 1031 989 1051
rect 1009 1031 1028 1051
rect 1048 1031 1067 1051
rect 1087 1031 1195 1051
rect 944 1027 1195 1031
rect 18263 1051 18508 1055
rect 18263 1031 18365 1051
rect 18385 1031 18404 1051
rect 18424 1031 18443 1051
rect 18463 1031 18482 1051
rect 18502 1031 18508 1051
rect 21346 1048 21397 1123
rect 21503 1048 21514 1123
rect 21346 1041 21514 1048
rect 18263 1027 18508 1031
rect 246 945 252 971
rect 427 945 433 971
rect 18839 945 18845 971
rect 19020 945 19026 971
rect 755 880 1195 884
rect 755 860 761 880
rect 781 860 800 880
rect 820 860 839 880
rect 859 860 878 880
rect 898 860 1195 880
rect 755 856 1195 860
rect 18263 880 18698 884
rect 18263 860 18554 880
rect 18574 860 18593 880
rect 18613 860 18632 880
rect 18652 860 18671 880
rect 18691 860 18698 880
rect 18263 856 18698 860
rect 21346 845 21514 854
rect 755 838 1195 842
rect 755 818 761 838
rect 781 818 800 838
rect 820 818 839 838
rect 859 818 878 838
rect 898 828 1195 838
rect 898 818 904 828
rect 755 814 904 818
rect 18550 770 19272 777
rect 18550 742 18565 770
rect 18593 742 18612 770
rect 18640 742 18659 770
rect 18687 763 19272 770
rect 21346 770 21397 845
rect 21503 770 21514 845
rect 21346 763 21514 770
rect 18687 742 19093 763
rect 18550 731 19093 742
rect 19125 731 19137 763
rect 19169 731 19181 763
rect 19213 731 19225 763
rect 19257 731 19272 763
rect 944 713 1195 727
rect 18550 723 19272 731
rect 944 710 1093 713
rect 944 690 950 710
rect 970 690 989 710
rect 1009 690 1028 710
rect 1048 690 1067 710
rect 1087 690 1093 710
rect 944 686 1093 690
rect 18550 695 18565 723
rect 18593 695 18612 723
rect 18640 695 18659 723
rect 18687 718 19272 723
rect 18687 695 19093 718
rect 18550 686 19093 695
rect 19125 686 19137 718
rect 19169 686 19181 718
rect 19213 686 19225 718
rect 19257 686 19272 718
rect 944 672 1195 686
rect 18550 676 19272 686
rect 944 654 1195 658
rect 944 634 950 654
rect 970 634 989 654
rect 1009 634 1028 654
rect 1048 634 1067 654
rect 1087 644 1195 654
rect 18550 648 18565 676
rect 18593 648 18612 676
rect 18640 648 18659 676
rect 18687 673 19272 676
rect 18687 648 19093 673
rect 1087 634 1093 644
rect 18550 641 19093 648
rect 19125 641 19137 673
rect 19169 641 19181 673
rect 19213 641 19225 673
rect 19257 641 19272 673
rect 18550 637 19272 641
rect 21630 746 21762 759
rect 944 630 1093 634
rect 644 584 730 587
rect 644 564 650 584
rect 670 564 689 584
rect 709 581 730 584
rect 18722 584 18808 587
rect 18722 581 18743 584
rect 709 567 1195 581
rect 18263 567 18743 581
rect 709 564 730 567
rect 644 561 730 564
rect 18722 564 18743 567
rect 18763 564 18782 584
rect 18802 564 18808 584
rect 18722 561 18808 564
rect 944 549 1195 553
rect 246 505 252 531
rect 427 505 433 531
rect 944 529 950 549
rect 970 529 989 549
rect 1009 529 1028 549
rect 1048 529 1067 549
rect 1087 529 1195 549
rect 944 525 1195 529
rect 18263 549 18508 553
rect 18263 529 18365 549
rect 18385 529 18404 549
rect 18424 529 18443 549
rect 18463 529 18482 549
rect 18502 529 18508 549
rect 21630 540 21643 746
rect 21749 540 21762 746
rect 18263 525 18508 529
rect 18839 505 18845 531
rect 19020 505 19026 531
rect 21630 528 21762 540
rect 18341 444 19033 445
rect 18341 437 19034 444
rect 18341 409 18376 437
rect 18404 409 18423 437
rect 18451 409 18470 437
rect 18498 431 19034 437
rect 18498 409 18855 431
rect 18341 399 18855 409
rect 18887 399 18899 431
rect 18931 399 18943 431
rect 18975 399 18987 431
rect 19019 399 19034 431
rect 17293 393 17566 396
rect 239 379 445 380
rect 238 366 445 379
rect 238 334 253 366
rect 285 334 297 366
rect 329 334 341 366
rect 373 334 385 366
rect 417 334 445 366
rect 238 321 445 334
rect 238 289 253 321
rect 285 289 297 321
rect 329 289 341 321
rect 373 289 385 321
rect 417 289 445 321
rect 238 276 445 289
rect 238 244 253 276
rect 285 244 297 276
rect 329 244 341 276
rect 373 244 385 276
rect 417 244 445 276
rect 238 240 445 244
rect 922 372 1104 380
rect 17293 376 17299 393
rect 17316 376 17543 393
rect 17560 376 17566 393
rect 17293 372 17566 376
rect 18341 390 19034 399
rect 922 344 954 372
rect 982 344 1001 372
rect 1029 344 1048 372
rect 1076 344 1104 372
rect 922 325 1104 344
rect 922 297 954 325
rect 982 297 1001 325
rect 1029 297 1048 325
rect 1076 297 1104 325
rect 18341 362 18376 390
rect 18404 362 18423 390
rect 18451 362 18470 390
rect 18498 386 19034 390
rect 18498 362 18855 386
rect 18341 354 18855 362
rect 18887 354 18899 386
rect 18931 354 18943 386
rect 18975 354 18987 386
rect 19019 354 19034 386
rect 18341 343 19034 354
rect 14472 321 15701 324
rect 14472 304 14478 321
rect 14495 304 15678 321
rect 15695 304 15701 321
rect 18341 315 18376 343
rect 18404 315 18423 343
rect 18451 315 18470 343
rect 18498 341 19034 343
rect 18498 315 18855 341
rect 18341 309 18855 315
rect 18887 309 18899 341
rect 18931 309 18943 341
rect 18975 309 18987 341
rect 19019 309 19034 341
rect 18341 305 19034 309
rect 14472 300 15701 304
rect 922 278 1104 297
rect 922 250 954 278
rect 982 250 1001 278
rect 1029 250 1048 278
rect 1076 250 1104 278
rect 14574 282 16203 285
rect 14574 265 14580 282
rect 14597 265 16180 282
rect 16197 265 16203 282
rect 14574 261 16203 265
rect 21346 273 21762 279
rect 922 240 1104 250
rect 14676 244 16705 247
rect 14676 227 14682 244
rect 14699 227 16682 244
rect 16699 227 16705 244
rect 14676 223 16705 227
rect 18341 226 18698 227
rect 18341 219 19272 226
rect 14778 206 17207 209
rect 14778 189 14784 206
rect 14801 189 17184 206
rect 17201 189 17207 206
rect 14778 185 17207 189
rect 18341 191 18565 219
rect 18593 191 18612 219
rect 18640 191 18659 219
rect 18687 212 19272 219
rect 18687 191 19093 212
rect 18341 180 19093 191
rect 19125 180 19137 212
rect 19169 180 19181 212
rect 19213 180 19225 212
rect 19257 180 19272 212
rect 21346 192 21637 273
rect 21756 192 21762 273
rect 21346 187 21762 192
rect 18341 172 19272 180
rect 14880 168 17709 171
rect 1617 162 1643 165
rect 810 161 1620 162
rect 0 147 207 161
rect 0 115 15 147
rect 47 115 59 147
rect 91 115 103 147
rect 135 115 147 147
rect 179 115 207 147
rect 0 102 207 115
rect 0 70 15 102
rect 47 70 59 102
rect 91 70 103 102
rect 135 70 147 102
rect 179 70 207 102
rect 0 57 207 70
rect 0 25 15 57
rect 47 25 59 57
rect 91 25 103 57
rect 135 25 147 57
rect 179 25 207 57
rect 0 21 207 25
rect 733 153 1620 161
rect 733 125 765 153
rect 793 125 812 153
rect 840 125 859 153
rect 887 145 1620 153
rect 1637 145 1643 162
rect 14880 151 14886 168
rect 14903 151 17686 168
rect 17703 151 17709 168
rect 18341 162 18565 172
rect 14880 147 17709 151
rect 18184 159 18565 162
rect 887 141 1643 145
rect 18184 142 18190 159
rect 18207 144 18565 159
rect 18593 144 18612 172
rect 18640 144 18659 172
rect 18687 167 19272 172
rect 18687 144 19093 167
rect 18207 142 19093 144
rect 887 125 1104 141
rect 18184 138 19093 142
rect 733 106 1104 125
rect 733 78 765 106
rect 793 78 812 106
rect 840 78 859 106
rect 887 78 1104 106
rect 18341 135 19093 138
rect 19125 135 19137 167
rect 19169 135 19181 167
rect 19213 135 19225 167
rect 19257 135 19272 167
rect 18341 125 19272 135
rect 18341 97 18565 125
rect 18593 97 18612 125
rect 18640 97 18659 125
rect 18687 122 19272 125
rect 18687 97 19093 122
rect 18341 90 19093 97
rect 19125 90 19137 122
rect 19169 90 19181 122
rect 19213 90 19225 122
rect 19257 90 19272 122
rect 18341 86 19272 90
rect 733 59 1104 78
rect 733 31 765 59
rect 793 31 812 59
rect 840 31 859 59
rect 887 31 1104 59
rect 733 22 1104 31
rect 17590 25 19391 28
rect 733 21 915 22
rect 17590 8 17596 25
rect 17613 8 17632 25
rect 17649 8 19391 25
rect 17590 4 19391 8
<< via1 >>
rect 21637 11747 21756 11828
rect 21643 11419 21749 11625
rect 21397 11319 21503 11394
rect 21397 11048 21503 11123
rect 21397 10770 21503 10845
rect 21643 10540 21749 10746
rect 21637 10192 21756 10273
rect 1494 9973 1625 10052
rect 3058 9973 3189 10052
rect 3494 9973 3625 10052
rect 5058 9973 5189 10052
rect 5494 9973 5625 10052
rect 7058 9973 7189 10052
rect 7494 9973 7625 10052
rect 9058 9973 9189 10052
rect 9494 9973 9625 10052
rect 11058 9973 11189 10052
rect 11494 9973 11625 10052
rect 13058 9973 13189 10052
rect 13494 9973 13625 10052
rect 15058 9973 15189 10052
rect 15494 9973 15625 10052
rect 17058 9973 17189 10052
rect 17494 9973 17625 10052
rect 19058 9990 19189 10052
rect 15 9914 47 9946
rect 59 9914 91 9946
rect 103 9914 135 9946
rect 147 9914 179 9946
rect 15 9869 47 9901
rect 59 9869 91 9901
rect 103 9869 135 9901
rect 147 9869 179 9901
rect 15 9824 47 9856
rect 59 9824 91 9856
rect 103 9824 135 9856
rect 147 9824 179 9856
rect 2267 9819 2430 9941
rect 4267 9819 4430 9941
rect 6267 9819 6430 9941
rect 8267 9819 8430 9941
rect 10267 9819 10430 9941
rect 12267 9819 12430 9941
rect 14267 9819 14430 9941
rect 16267 9819 16430 9941
rect 18267 9819 18430 9941
rect 19093 9914 19125 9946
rect 19137 9914 19169 9946
rect 19181 9914 19213 9946
rect 19225 9914 19257 9946
rect 19093 9869 19125 9901
rect 19137 9869 19169 9901
rect 19181 9869 19213 9901
rect 19225 9869 19257 9901
rect 19093 9824 19125 9856
rect 19137 9824 19169 9856
rect 19181 9824 19213 9856
rect 19225 9824 19257 9856
rect 21637 9747 21756 9828
rect 253 9695 285 9727
rect 297 9695 329 9727
rect 341 9695 373 9727
rect 385 9695 417 9727
rect 18855 9695 18887 9727
rect 18899 9695 18931 9727
rect 18943 9695 18975 9727
rect 18987 9695 19019 9727
rect 253 9650 285 9682
rect 297 9650 329 9682
rect 341 9650 373 9682
rect 385 9650 417 9682
rect 18855 9650 18887 9682
rect 18899 9650 18931 9682
rect 18943 9650 18975 9682
rect 18987 9650 19019 9682
rect 253 9605 285 9637
rect 297 9605 329 9637
rect 341 9605 373 9637
rect 385 9605 417 9637
rect 18855 9605 18887 9637
rect 18899 9605 18931 9637
rect 18943 9605 18975 9637
rect 18987 9605 19019 9637
rect 21643 9419 21749 9625
rect 252 9327 427 9331
rect 252 9310 427 9327
rect 252 9305 427 9310
rect 18845 9327 19020 9331
rect 18845 9310 19020 9327
rect 18845 9305 19020 9310
rect 18856 9284 18888 9305
rect 18900 9284 18932 9305
rect 18944 9284 18976 9305
rect 18988 9284 19020 9305
rect 21397 9319 21503 9394
rect 18856 9239 18888 9271
rect 18900 9239 18932 9271
rect 18944 9239 18976 9271
rect 18988 9239 19020 9271
rect 18856 9194 18888 9226
rect 18900 9194 18932 9226
rect 18944 9194 18976 9226
rect 18988 9194 19020 9226
rect 21397 9048 21503 9123
rect 252 8887 427 8891
rect 252 8870 427 8887
rect 252 8865 427 8870
rect 18845 8887 19020 8891
rect 18845 8870 19020 8887
rect 18845 8865 19020 8870
rect 19093 8791 19125 8823
rect 19137 8791 19169 8823
rect 19181 8791 19213 8823
rect 19225 8791 19257 8823
rect 19093 8746 19125 8778
rect 19137 8746 19169 8778
rect 19181 8746 19213 8778
rect 19225 8746 19257 8778
rect 21397 8770 21503 8845
rect 19093 8701 19125 8733
rect 19137 8701 19169 8733
rect 19181 8701 19213 8733
rect 19225 8701 19257 8733
rect 21643 8540 21749 8746
rect 252 8447 427 8451
rect 252 8430 427 8447
rect 252 8425 427 8430
rect 18845 8447 19020 8451
rect 18845 8430 19020 8447
rect 18845 8425 19020 8430
rect 18855 8276 18887 8308
rect 18899 8276 18931 8308
rect 18943 8276 18975 8308
rect 18987 8276 19019 8308
rect 18855 8231 18887 8263
rect 18899 8231 18931 8263
rect 18943 8231 18975 8263
rect 18987 8231 19019 8263
rect 18855 8186 18887 8218
rect 18899 8186 18931 8218
rect 18943 8186 18975 8218
rect 18987 8186 19019 8218
rect 21637 8192 21756 8273
rect 252 8007 427 8011
rect 252 7990 427 8007
rect 252 7985 427 7990
rect 18845 8007 19020 8011
rect 18845 7990 19020 8007
rect 18845 7985 19020 7990
rect 19093 7737 19125 7769
rect 19137 7737 19169 7769
rect 19181 7737 19213 7769
rect 19225 7737 19257 7769
rect 21637 7747 21756 7828
rect 19093 7692 19125 7724
rect 19137 7692 19169 7724
rect 19181 7692 19213 7724
rect 19225 7692 19257 7724
rect 19093 7647 19125 7679
rect 19137 7647 19169 7679
rect 19181 7647 19213 7679
rect 19225 7647 19257 7679
rect 252 7567 427 7571
rect 252 7550 427 7567
rect 252 7545 427 7550
rect 18845 7567 19020 7571
rect 18845 7550 19020 7567
rect 18845 7545 19020 7550
rect 21643 7419 21749 7625
rect 21397 7319 21503 7394
rect 18855 7276 18887 7308
rect 18899 7276 18931 7308
rect 18943 7276 18975 7308
rect 18987 7276 19019 7308
rect 18855 7231 18887 7263
rect 18899 7231 18931 7263
rect 18943 7231 18975 7263
rect 18987 7231 19019 7263
rect 18855 7186 18887 7218
rect 18899 7186 18931 7218
rect 18943 7186 18975 7218
rect 18987 7186 19019 7218
rect 252 7127 427 7131
rect 252 7110 427 7127
rect 252 7105 427 7110
rect 18845 7127 19020 7131
rect 18845 7110 19020 7127
rect 18845 7105 19020 7110
rect 21397 7048 21503 7123
rect 19092 6772 19124 6804
rect 19136 6772 19168 6804
rect 19180 6772 19212 6804
rect 19224 6772 19256 6804
rect 21397 6770 21503 6845
rect 19092 6727 19124 6759
rect 19136 6727 19168 6759
rect 19180 6727 19212 6759
rect 19224 6727 19256 6759
rect 252 6687 427 6691
rect 252 6670 427 6687
rect 252 6665 427 6670
rect 19092 6682 19124 6714
rect 19136 6682 19168 6714
rect 19180 6682 19212 6714
rect 19224 6682 19256 6714
rect 21643 6540 21749 6746
rect 18856 6314 18888 6346
rect 18900 6314 18932 6346
rect 18944 6314 18976 6346
rect 18988 6314 19020 6346
rect 18856 6269 18888 6301
rect 18900 6269 18932 6301
rect 18944 6269 18976 6301
rect 18988 6269 19020 6301
rect 252 6247 427 6251
rect 252 6230 427 6247
rect 252 6225 427 6230
rect 18856 6251 18888 6256
rect 18900 6251 18932 6256
rect 18944 6251 18976 6256
rect 18988 6251 19020 6256
rect 18845 6247 19020 6251
rect 18845 6230 19020 6247
rect 18845 6225 19020 6230
rect 18856 6224 18888 6225
rect 18900 6224 18932 6225
rect 18944 6224 18976 6225
rect 18988 6224 19020 6225
rect 21637 6192 21756 6273
rect 252 5807 427 5811
rect 252 5790 427 5807
rect 252 5785 427 5790
rect 19093 5764 19125 5796
rect 19137 5764 19169 5796
rect 19181 5764 19213 5796
rect 19225 5764 19257 5796
rect 19093 5719 19125 5751
rect 19137 5719 19169 5751
rect 19181 5719 19213 5751
rect 19225 5719 19257 5751
rect 21637 5747 21756 5828
rect 19093 5674 19125 5706
rect 19137 5674 19169 5706
rect 19181 5674 19213 5706
rect 19225 5674 19257 5706
rect 21643 5419 21749 5625
rect 252 5367 427 5371
rect 252 5350 427 5367
rect 252 5345 427 5350
rect 18845 5367 19020 5371
rect 18845 5350 19020 5367
rect 18845 5345 19020 5350
rect 21397 5319 21503 5394
rect 18855 5251 18887 5283
rect 18899 5251 18931 5283
rect 18943 5251 18975 5283
rect 18987 5251 19019 5283
rect 18855 5206 18887 5238
rect 18899 5206 18931 5238
rect 18943 5206 18975 5238
rect 18987 5206 19019 5238
rect 18855 5161 18887 5193
rect 18899 5161 18931 5193
rect 18943 5161 18975 5193
rect 18987 5161 19019 5193
rect 21397 5048 21503 5123
rect 252 4927 427 4931
rect 252 4910 427 4927
rect 252 4905 427 4910
rect 18845 4927 19020 4931
rect 18845 4910 19020 4927
rect 18845 4905 19020 4910
rect 19093 4763 19125 4795
rect 19137 4763 19169 4795
rect 19181 4763 19213 4795
rect 19225 4763 19257 4795
rect 21397 4770 21503 4845
rect 19093 4718 19125 4750
rect 19137 4718 19169 4750
rect 19181 4718 19213 4750
rect 19225 4718 19257 4750
rect 19093 4673 19125 4705
rect 19137 4673 19169 4705
rect 19181 4673 19213 4705
rect 19225 4673 19257 4705
rect 21643 4540 21749 4746
rect 252 4487 427 4491
rect 252 4470 427 4487
rect 252 4465 427 4470
rect 18845 4487 19020 4491
rect 18845 4470 19020 4487
rect 18845 4465 19020 4470
rect 18856 4263 18888 4295
rect 18900 4263 18932 4295
rect 18944 4263 18976 4295
rect 18988 4263 19020 4295
rect 18856 4218 18888 4250
rect 18900 4218 18932 4250
rect 18944 4218 18976 4250
rect 18988 4218 19020 4250
rect 18856 4173 18888 4205
rect 18900 4173 18932 4205
rect 18944 4173 18976 4205
rect 18988 4173 19020 4205
rect 21637 4192 21756 4273
rect 252 4047 427 4051
rect 252 4030 427 4047
rect 252 4025 427 4030
rect 18845 4047 19020 4051
rect 18845 4030 19020 4047
rect 18845 4025 19020 4030
rect 19092 3764 19124 3796
rect 19136 3764 19168 3796
rect 19180 3764 19212 3796
rect 19224 3764 19256 3796
rect 19092 3719 19124 3751
rect 19136 3719 19168 3751
rect 19180 3719 19212 3751
rect 19224 3719 19256 3751
rect 21637 3747 21756 3828
rect 19092 3674 19124 3706
rect 19136 3674 19168 3706
rect 19180 3674 19212 3706
rect 19224 3674 19256 3706
rect 252 3607 427 3611
rect 252 3590 427 3607
rect 252 3585 427 3590
rect 18845 3607 19020 3611
rect 18845 3590 19020 3607
rect 18845 3585 19020 3590
rect 21643 3419 21749 3625
rect 21397 3319 21503 3394
rect 18856 3241 18888 3273
rect 18900 3241 18932 3273
rect 18944 3241 18976 3273
rect 18988 3241 19020 3273
rect 18856 3196 18888 3228
rect 18900 3196 18932 3228
rect 18944 3196 18976 3228
rect 18988 3196 19020 3228
rect 252 3167 427 3171
rect 252 3150 427 3167
rect 252 3145 427 3150
rect 18856 3171 18888 3183
rect 18900 3171 18932 3183
rect 18944 3171 18976 3183
rect 18988 3171 19020 3183
rect 18845 3167 19020 3171
rect 18845 3150 19020 3167
rect 18845 3145 19020 3150
rect 21397 3048 21503 3123
rect 21397 2770 21503 2845
rect 252 2727 427 2731
rect 252 2710 427 2727
rect 252 2705 427 2710
rect 19093 2730 19125 2762
rect 19137 2730 19169 2762
rect 19181 2730 19213 2762
rect 19225 2730 19257 2762
rect 19093 2685 19125 2717
rect 19137 2685 19169 2717
rect 19181 2685 19213 2717
rect 19225 2685 19257 2717
rect 19093 2640 19125 2672
rect 19137 2640 19169 2672
rect 19181 2640 19213 2672
rect 19225 2640 19257 2672
rect 21643 2540 21749 2746
rect 252 2287 427 2291
rect 252 2270 427 2287
rect 252 2265 427 2270
rect 18845 2287 19020 2291
rect 18845 2270 19020 2287
rect 18845 2265 19020 2270
rect 18856 2244 18888 2265
rect 18900 2244 18932 2265
rect 18944 2244 18976 2265
rect 18988 2244 19020 2265
rect 18856 2199 18888 2231
rect 18900 2199 18932 2231
rect 18944 2199 18976 2231
rect 18988 2199 19020 2231
rect 21637 2192 21756 2273
rect 18856 2154 18888 2186
rect 18900 2154 18932 2186
rect 18944 2154 18976 2186
rect 18988 2154 19020 2186
rect 252 1847 427 1851
rect 252 1830 427 1847
rect 252 1825 427 1830
rect 18845 1847 19020 1851
rect 18845 1830 19020 1847
rect 18845 1825 19020 1830
rect 19093 1728 19125 1760
rect 19137 1728 19169 1760
rect 19181 1728 19213 1760
rect 19225 1728 19257 1760
rect 21637 1747 21756 1828
rect 19093 1683 19125 1715
rect 19137 1683 19169 1715
rect 19181 1683 19213 1715
rect 19225 1683 19257 1715
rect 19093 1638 19125 1670
rect 19137 1638 19169 1670
rect 19181 1638 19213 1670
rect 19225 1638 19257 1670
rect 21643 1419 21749 1625
rect 252 1407 427 1411
rect 252 1390 427 1407
rect 252 1385 427 1390
rect 18845 1407 19020 1411
rect 18845 1390 19020 1407
rect 18845 1385 19020 1390
rect 21397 1319 21503 1394
rect 18854 1244 18886 1276
rect 18898 1244 18930 1276
rect 18942 1244 18974 1276
rect 18986 1244 19018 1276
rect 18854 1199 18886 1231
rect 18898 1199 18930 1231
rect 18942 1199 18974 1231
rect 18986 1199 19018 1231
rect 18854 1154 18886 1186
rect 18898 1154 18930 1186
rect 18942 1154 18974 1186
rect 18986 1154 19018 1186
rect 21397 1048 21503 1123
rect 252 967 427 971
rect 252 950 427 967
rect 252 945 427 950
rect 18845 967 19020 971
rect 18845 950 19020 967
rect 18845 945 19020 950
rect 21397 770 21503 845
rect 19093 731 19125 763
rect 19137 731 19169 763
rect 19181 731 19213 763
rect 19225 731 19257 763
rect 19093 686 19125 718
rect 19137 686 19169 718
rect 19181 686 19213 718
rect 19225 686 19257 718
rect 19093 641 19125 673
rect 19137 641 19169 673
rect 19181 641 19213 673
rect 19225 641 19257 673
rect 252 527 427 531
rect 252 510 427 527
rect 252 505 427 510
rect 21643 540 21749 746
rect 18845 527 19020 531
rect 18845 510 19020 527
rect 18845 505 19020 510
rect 18855 399 18887 431
rect 18899 399 18931 431
rect 18943 399 18975 431
rect 18987 399 19019 431
rect 253 334 285 366
rect 297 334 329 366
rect 341 334 373 366
rect 385 334 417 366
rect 253 289 285 321
rect 297 289 329 321
rect 341 289 373 321
rect 385 289 417 321
rect 253 244 285 276
rect 297 244 329 276
rect 341 244 373 276
rect 385 244 417 276
rect 954 344 982 372
rect 1001 344 1029 372
rect 1048 344 1076 372
rect 954 297 982 325
rect 1001 297 1029 325
rect 1048 297 1076 325
rect 18855 354 18887 386
rect 18899 354 18931 386
rect 18943 354 18975 386
rect 18987 354 19019 386
rect 18855 309 18887 341
rect 18899 309 18931 341
rect 18943 309 18975 341
rect 18987 309 19019 341
rect 954 250 982 278
rect 1001 250 1029 278
rect 1048 250 1076 278
rect 19093 180 19125 212
rect 19137 180 19169 212
rect 19181 180 19213 212
rect 19225 180 19257 212
rect 21637 192 21756 273
rect 15 115 47 147
rect 59 115 91 147
rect 103 115 135 147
rect 147 115 179 147
rect 15 70 47 102
rect 59 70 91 102
rect 103 70 135 102
rect 147 70 179 102
rect 15 25 47 57
rect 59 25 91 57
rect 103 25 135 57
rect 147 25 179 57
rect 765 125 793 153
rect 812 125 840 153
rect 859 125 887 153
rect 765 78 793 106
rect 812 78 840 106
rect 859 78 887 106
rect 19093 135 19125 167
rect 19137 135 19169 167
rect 19181 135 19213 167
rect 19225 135 19257 167
rect 19093 90 19125 122
rect 19137 90 19169 122
rect 19181 90 19213 122
rect 19225 90 19257 122
rect 765 31 793 59
rect 812 31 840 59
rect 859 31 887 59
<< metal2 >>
rect 21346 11828 21762 11834
rect 21346 11747 21637 11828
rect 21756 11747 21762 11828
rect 21346 11742 21762 11747
rect 21630 11625 21762 11638
rect 21630 11419 21643 11625
rect 21749 11419 21762 11625
rect 21630 11407 21762 11419
rect 21346 11394 21514 11403
rect 21346 11319 21397 11394
rect 21503 11319 21514 11394
rect 21346 11312 21514 11319
rect 21346 11123 21514 11132
rect 21346 11048 21397 11123
rect 21503 11048 21514 11123
rect 21346 11041 21514 11048
rect 21346 10845 21514 10854
rect 21346 10770 21397 10845
rect 21503 10770 21514 10845
rect 21346 10763 21514 10770
rect 21630 10746 21762 10759
rect 21630 10540 21643 10746
rect 21749 10540 21762 10746
rect 21630 10528 21762 10540
rect 21346 10273 21762 10279
rect 21346 10192 21637 10273
rect 21756 10192 21762 10273
rect 21346 10187 21762 10192
rect 1487 10052 1633 10060
rect 1487 9973 1494 10052
rect 1625 9973 1633 10052
rect 1487 9967 1633 9973
rect 3051 10052 3197 10060
rect 3051 9973 3058 10052
rect 3189 9973 3197 10052
rect 3051 9967 3197 9973
rect 3487 10052 3633 10060
rect 3487 9973 3494 10052
rect 3625 9973 3633 10052
rect 3487 9967 3633 9973
rect 5051 10052 5197 10060
rect 5051 9973 5058 10052
rect 5189 9973 5197 10052
rect 5051 9967 5197 9973
rect 5487 10052 5633 10060
rect 5487 9973 5494 10052
rect 5625 9973 5633 10052
rect 5487 9967 5633 9973
rect 7051 10052 7197 10060
rect 7051 9973 7058 10052
rect 7189 9973 7197 10052
rect 7051 9967 7197 9973
rect 7487 10052 7633 10060
rect 7487 9973 7494 10052
rect 7625 9973 7633 10052
rect 7487 9967 7633 9973
rect 9051 10052 9197 10060
rect 9051 9973 9058 10052
rect 9189 9973 9197 10052
rect 9051 9967 9197 9973
rect 9487 10052 9633 10060
rect 9487 9973 9494 10052
rect 9625 9973 9633 10052
rect 9487 9967 9633 9973
rect 11051 10052 11197 10060
rect 11051 9973 11058 10052
rect 11189 9973 11197 10052
rect 11051 9967 11197 9973
rect 11487 10052 11633 10060
rect 11487 9973 11494 10052
rect 11625 9973 11633 10052
rect 11487 9967 11633 9973
rect 13051 10052 13197 10060
rect 13051 9973 13058 10052
rect 13189 9973 13197 10052
rect 13051 9967 13197 9973
rect 13487 10052 13633 10060
rect 13487 9973 13494 10052
rect 13625 9973 13633 10052
rect 13487 9967 13633 9973
rect 15051 10052 15197 10060
rect 15051 9973 15058 10052
rect 15189 9973 15197 10052
rect 15051 9967 15197 9973
rect 15487 10052 15633 10060
rect 15487 9973 15494 10052
rect 15625 9973 15633 10052
rect 15487 9967 15633 9973
rect 17051 10052 17197 10060
rect 17051 9973 17058 10052
rect 17189 9973 17197 10052
rect 17051 9967 17197 9973
rect 17487 10052 17633 10060
rect 17487 9973 17494 10052
rect 17625 9973 17633 10052
rect 19051 10052 19197 10060
rect 19051 9990 19058 10052
rect 19189 9990 19197 10052
rect 19051 9984 19197 9990
rect 17487 9967 17633 9973
rect 0 9946 207 9950
rect 0 9914 15 9946
rect 47 9914 59 9946
rect 91 9914 103 9946
rect 135 9914 147 9946
rect 179 9914 207 9946
rect 0 9901 207 9914
rect 0 9869 15 9901
rect 47 9869 59 9901
rect 91 9869 103 9901
rect 135 9869 147 9901
rect 179 9869 207 9901
rect 0 9856 207 9869
rect 0 9824 15 9856
rect 47 9824 59 9856
rect 91 9824 103 9856
rect 135 9824 147 9856
rect 179 9824 207 9856
rect 0 9810 207 9824
rect 2255 9941 2440 9950
rect 2255 9819 2267 9941
rect 2430 9819 2440 9941
rect 2255 9810 2440 9819
rect 4255 9941 4440 9950
rect 4255 9819 4267 9941
rect 4430 9819 4440 9941
rect 4255 9810 4440 9819
rect 6255 9941 6440 9950
rect 6255 9819 6267 9941
rect 6430 9819 6440 9941
rect 6255 9810 6440 9819
rect 8255 9941 8440 9950
rect 8255 9819 8267 9941
rect 8430 9819 8440 9941
rect 8255 9810 8440 9819
rect 10255 9941 10440 9950
rect 10255 9819 10267 9941
rect 10430 9819 10440 9941
rect 10255 9810 10440 9819
rect 12255 9941 12440 9950
rect 12255 9819 12267 9941
rect 12430 9819 12440 9941
rect 12255 9810 12440 9819
rect 14255 9941 14440 9950
rect 14255 9819 14267 9941
rect 14430 9819 14440 9941
rect 14255 9810 14440 9819
rect 16255 9941 16440 9950
rect 16255 9819 16267 9941
rect 16430 9819 16440 9941
rect 16255 9810 16440 9819
rect 18255 9941 18440 9950
rect 18255 9819 18267 9941
rect 18430 9819 18440 9941
rect 18255 9810 18440 9819
rect 19065 9946 19272 9950
rect 19065 9914 19093 9946
rect 19125 9914 19137 9946
rect 19169 9914 19181 9946
rect 19213 9914 19225 9946
rect 19257 9914 19272 9946
rect 19065 9901 19272 9914
rect 19065 9869 19093 9901
rect 19125 9869 19137 9901
rect 19169 9869 19181 9901
rect 19213 9869 19225 9901
rect 19257 9869 19272 9901
rect 19065 9856 19272 9869
rect 19065 9824 19093 9856
rect 19125 9824 19137 9856
rect 19169 9824 19181 9856
rect 19213 9824 19225 9856
rect 19257 9824 19272 9856
rect 19065 9810 19272 9824
rect 21346 9828 21762 9834
rect 21346 9747 21637 9828
rect 21756 9747 21762 9828
rect 21346 9742 21762 9747
rect 238 9727 445 9731
rect 238 9695 253 9727
rect 285 9695 297 9727
rect 329 9695 341 9727
rect 373 9695 385 9727
rect 417 9695 445 9727
rect 238 9682 445 9695
rect 238 9650 253 9682
rect 285 9650 297 9682
rect 329 9650 341 9682
rect 373 9650 385 9682
rect 417 9650 445 9682
rect 238 9637 445 9650
rect 238 9605 253 9637
rect 285 9605 297 9637
rect 329 9605 341 9637
rect 373 9605 385 9637
rect 417 9605 445 9637
rect 238 9591 445 9605
rect 18827 9727 19346 9731
rect 18827 9695 18855 9727
rect 18887 9695 18899 9727
rect 18931 9695 18943 9727
rect 18975 9695 18987 9727
rect 19019 9695 19346 9727
rect 18827 9682 19346 9695
rect 18827 9650 18855 9682
rect 18887 9650 18899 9682
rect 18931 9650 18943 9682
rect 18975 9650 18987 9682
rect 19019 9650 19346 9682
rect 18827 9637 19346 9650
rect 18827 9605 18855 9637
rect 18887 9605 18899 9637
rect 18931 9605 18943 9637
rect 18975 9605 18987 9637
rect 19019 9605 19346 9637
rect 18827 9591 19346 9605
rect 21630 9625 21762 9638
rect 21630 9419 21643 9625
rect 21749 9419 21762 9625
rect 21630 9407 21762 9419
rect 21346 9394 21514 9403
rect 246 9304 252 9332
rect 427 9304 433 9332
rect 18839 9330 18845 9332
rect 18828 9304 18845 9330
rect 19020 9330 19026 9332
rect 18828 9284 18856 9304
rect 18888 9284 18900 9304
rect 18932 9284 18944 9304
rect 18976 9284 18988 9304
rect 19020 9284 19035 9330
rect 21346 9319 21397 9394
rect 21503 9319 21514 9394
rect 21346 9312 21514 9319
rect 18828 9271 19035 9284
rect 18828 9239 18856 9271
rect 18888 9239 18900 9271
rect 18932 9239 18944 9271
rect 18976 9239 18988 9271
rect 19020 9239 19035 9271
rect 18828 9226 19035 9239
rect 18828 9194 18856 9226
rect 18888 9194 18900 9226
rect 18932 9194 18944 9226
rect 18976 9194 18988 9226
rect 19020 9194 19035 9226
rect 18828 9190 19035 9194
rect 21346 9123 21514 9132
rect 21346 9048 21397 9123
rect 21503 9048 21514 9123
rect 21346 9041 21514 9048
rect 246 8864 252 8892
rect 427 8864 433 8892
rect 18839 8864 18845 8892
rect 19020 8864 19026 8892
rect 19065 8837 19346 8977
rect 21346 8845 21514 8854
rect 19065 8823 19272 8837
rect 19065 8791 19093 8823
rect 19125 8791 19137 8823
rect 19169 8791 19181 8823
rect 19213 8791 19225 8823
rect 19257 8791 19272 8823
rect 19065 8778 19272 8791
rect 19065 8746 19093 8778
rect 19125 8746 19137 8778
rect 19169 8746 19181 8778
rect 19213 8746 19225 8778
rect 19257 8746 19272 8778
rect 21346 8770 21397 8845
rect 21503 8770 21514 8845
rect 21346 8763 21514 8770
rect 19065 8733 19272 8746
rect 19065 8701 19093 8733
rect 19125 8701 19137 8733
rect 19169 8701 19181 8733
rect 19213 8701 19225 8733
rect 19257 8701 19272 8733
rect 19065 8697 19272 8701
rect 21630 8746 21762 8759
rect 21630 8540 21643 8746
rect 21749 8540 21762 8746
rect 21630 8528 21762 8540
rect 246 8424 252 8452
rect 427 8424 433 8452
rect 18839 8424 18845 8452
rect 19020 8424 19026 8452
rect 18827 8308 19346 8322
rect 18827 8276 18855 8308
rect 18887 8276 18899 8308
rect 18931 8276 18943 8308
rect 18975 8276 18987 8308
rect 19019 8276 19346 8308
rect 18827 8263 19346 8276
rect 18827 8231 18855 8263
rect 18887 8231 18899 8263
rect 18931 8231 18943 8263
rect 18975 8231 18987 8263
rect 19019 8231 19346 8263
rect 18827 8218 19346 8231
rect 18827 8186 18855 8218
rect 18887 8186 18899 8218
rect 18931 8186 18943 8218
rect 18975 8186 18987 8218
rect 19019 8186 19346 8218
rect 21346 8273 21762 8279
rect 21346 8192 21637 8273
rect 21756 8192 21762 8273
rect 21346 8187 21762 8192
rect 18827 8182 19346 8186
rect 246 7984 252 8012
rect 427 7984 433 8012
rect 18839 7984 18845 8012
rect 19020 7984 19026 8012
rect 21346 7828 21762 7834
rect 19065 7769 19272 7783
rect 19065 7737 19093 7769
rect 19125 7737 19137 7769
rect 19169 7737 19181 7769
rect 19213 7737 19225 7769
rect 19257 7737 19272 7769
rect 21346 7747 21637 7828
rect 21756 7747 21762 7828
rect 21346 7742 21762 7747
rect 19065 7724 19272 7737
rect 19065 7692 19093 7724
rect 19125 7692 19137 7724
rect 19169 7692 19181 7724
rect 19213 7692 19225 7724
rect 19257 7692 19272 7724
rect 19065 7679 19272 7692
rect 19065 7647 19093 7679
rect 19125 7647 19137 7679
rect 19169 7647 19181 7679
rect 19213 7647 19225 7679
rect 19257 7647 19272 7679
rect 19065 7643 19272 7647
rect 21630 7625 21762 7638
rect 246 7544 252 7572
rect 427 7544 433 7572
rect 18839 7544 18845 7572
rect 19020 7544 19026 7572
rect 21630 7419 21643 7625
rect 21749 7419 21762 7625
rect 21630 7407 21762 7419
rect 21346 7394 21514 7403
rect 18827 7308 19034 7322
rect 21346 7319 21397 7394
rect 21503 7319 21514 7394
rect 21346 7312 21514 7319
rect 18827 7276 18855 7308
rect 18887 7276 18899 7308
rect 18931 7276 18943 7308
rect 18975 7276 18987 7308
rect 19019 7276 19034 7308
rect 18827 7263 19034 7276
rect 18827 7231 18855 7263
rect 18887 7231 18899 7263
rect 18931 7231 18943 7263
rect 18975 7231 18987 7263
rect 19019 7231 19034 7263
rect 18827 7218 19034 7231
rect 18827 7186 18855 7218
rect 18887 7186 18899 7218
rect 18931 7186 18943 7218
rect 18975 7186 18987 7218
rect 19019 7186 19034 7218
rect 18827 7183 19034 7186
rect 246 7104 252 7132
rect 427 7104 433 7132
rect 18839 7104 18845 7132
rect 19020 7104 19026 7132
rect 21346 7123 21514 7132
rect 21346 7048 21397 7123
rect 21503 7048 21514 7123
rect 21346 7041 21514 7048
rect 19064 6818 19346 6959
rect 21346 6845 21514 6854
rect 19064 6804 19271 6818
rect 19064 6772 19092 6804
rect 19124 6772 19136 6804
rect 19168 6772 19180 6804
rect 19212 6772 19224 6804
rect 19256 6772 19271 6804
rect 19064 6759 19271 6772
rect 21346 6770 21397 6845
rect 21503 6770 21514 6845
rect 21346 6763 21514 6770
rect 19064 6727 19092 6759
rect 19124 6727 19136 6759
rect 19168 6727 19180 6759
rect 19212 6727 19224 6759
rect 19256 6727 19271 6759
rect 19064 6714 19271 6727
rect 246 6664 252 6692
rect 427 6664 433 6692
rect 19064 6682 19092 6714
rect 19124 6682 19136 6714
rect 19168 6682 19180 6714
rect 19212 6682 19224 6714
rect 19256 6682 19271 6714
rect 19064 6678 19271 6682
rect 21630 6746 21762 6759
rect 21630 6540 21643 6746
rect 21749 6540 21762 6746
rect 21630 6528 21762 6540
rect 19033 6360 19346 6361
rect 18828 6346 19346 6360
rect 18828 6314 18856 6346
rect 18888 6314 18900 6346
rect 18932 6314 18944 6346
rect 18976 6314 18988 6346
rect 19020 6314 19346 6346
rect 18828 6301 19346 6314
rect 18828 6269 18856 6301
rect 18888 6269 18900 6301
rect 18932 6269 18944 6301
rect 18976 6269 18988 6301
rect 19020 6269 19346 6301
rect 18828 6256 19346 6269
rect 18828 6252 18856 6256
rect 246 6224 252 6252
rect 427 6224 433 6252
rect 18828 6224 18845 6252
rect 18888 6252 18900 6256
rect 18932 6252 18944 6256
rect 18976 6252 18988 6256
rect 19020 6224 19346 6256
rect 18828 6220 19346 6224
rect 21346 6273 21762 6279
rect 21346 6192 21637 6273
rect 21756 6192 21762 6273
rect 21346 6187 21762 6192
rect 21346 5828 21762 5834
rect 246 5784 252 5812
rect 427 5784 433 5812
rect 19065 5796 19272 5810
rect 19065 5764 19093 5796
rect 19125 5764 19137 5796
rect 19169 5764 19181 5796
rect 19213 5764 19225 5796
rect 19257 5764 19272 5796
rect 19065 5751 19272 5764
rect 19065 5719 19093 5751
rect 19125 5719 19137 5751
rect 19169 5719 19181 5751
rect 19213 5719 19225 5751
rect 19257 5719 19272 5751
rect 21346 5747 21637 5828
rect 21756 5747 21762 5828
rect 21346 5742 21762 5747
rect 19065 5706 19272 5719
rect 19065 5674 19093 5706
rect 19125 5674 19137 5706
rect 19169 5674 19181 5706
rect 19213 5674 19225 5706
rect 19257 5674 19272 5706
rect 19065 5670 19272 5674
rect 21630 5625 21762 5638
rect 21630 5419 21643 5625
rect 21749 5419 21762 5625
rect 21630 5407 21762 5419
rect 21346 5394 21514 5403
rect 246 5344 252 5372
rect 427 5344 433 5372
rect 18839 5344 18845 5372
rect 19020 5344 19026 5372
rect 21346 5319 21397 5394
rect 21503 5319 21514 5394
rect 21346 5312 21514 5319
rect 18827 5283 19034 5297
rect 18827 5251 18855 5283
rect 18887 5251 18899 5283
rect 18931 5251 18943 5283
rect 18975 5251 18987 5283
rect 19019 5251 19034 5283
rect 18827 5238 19034 5251
rect 18827 5206 18855 5238
rect 18887 5206 18899 5238
rect 18931 5206 18943 5238
rect 18975 5206 18987 5238
rect 19019 5206 19034 5238
rect 18827 5193 19034 5206
rect 18827 5161 18855 5193
rect 18887 5161 18899 5193
rect 18931 5161 18943 5193
rect 18975 5161 18987 5193
rect 19019 5161 19034 5193
rect 18827 5157 19034 5161
rect 21346 5123 21514 5132
rect 21346 5048 21397 5123
rect 21503 5048 21514 5123
rect 21346 5041 21514 5048
rect 246 4904 252 4932
rect 427 4904 433 4932
rect 18839 4904 18845 4932
rect 19020 4904 19026 4932
rect 19065 4809 19346 4948
rect 21346 4845 21514 4854
rect 19065 4795 19272 4809
rect 19065 4763 19093 4795
rect 19125 4763 19137 4795
rect 19169 4763 19181 4795
rect 19213 4763 19225 4795
rect 19257 4763 19272 4795
rect 21346 4770 21397 4845
rect 21503 4770 21514 4845
rect 21346 4763 21514 4770
rect 19065 4750 19272 4763
rect 19065 4718 19093 4750
rect 19125 4718 19137 4750
rect 19169 4718 19181 4750
rect 19213 4718 19225 4750
rect 19257 4718 19272 4750
rect 19065 4705 19272 4718
rect 19065 4673 19093 4705
rect 19125 4673 19137 4705
rect 19169 4673 19181 4705
rect 19213 4673 19225 4705
rect 19257 4673 19272 4705
rect 19065 4669 19272 4673
rect 21630 4746 21762 4759
rect 21630 4540 21643 4746
rect 21749 4540 21762 4746
rect 21630 4528 21762 4540
rect 246 4464 252 4492
rect 427 4464 433 4492
rect 18839 4464 18845 4492
rect 19020 4464 19026 4492
rect 18828 4295 19346 4309
rect 18828 4263 18856 4295
rect 18888 4263 18900 4295
rect 18932 4263 18944 4295
rect 18976 4263 18988 4295
rect 19020 4263 19346 4295
rect 18828 4250 19346 4263
rect 18828 4218 18856 4250
rect 18888 4218 18900 4250
rect 18932 4218 18944 4250
rect 18976 4218 18988 4250
rect 19020 4218 19346 4250
rect 18828 4205 19346 4218
rect 18828 4173 18856 4205
rect 18888 4173 18900 4205
rect 18932 4173 18944 4205
rect 18976 4173 18988 4205
rect 19020 4173 19346 4205
rect 21346 4273 21762 4279
rect 21346 4192 21637 4273
rect 21756 4192 21762 4273
rect 21346 4187 21762 4192
rect 18828 4169 19346 4173
rect 246 4024 252 4052
rect 427 4024 433 4052
rect 18839 4024 18845 4052
rect 19020 4024 19026 4052
rect 21346 3828 21762 3834
rect 19064 3796 19271 3810
rect 19064 3764 19092 3796
rect 19124 3764 19136 3796
rect 19168 3764 19180 3796
rect 19212 3764 19224 3796
rect 19256 3764 19271 3796
rect 19064 3751 19271 3764
rect 19064 3719 19092 3751
rect 19124 3719 19136 3751
rect 19168 3719 19180 3751
rect 19212 3719 19224 3751
rect 19256 3719 19271 3751
rect 21346 3747 21637 3828
rect 21756 3747 21762 3828
rect 21346 3742 21762 3747
rect 19064 3706 19271 3719
rect 19064 3674 19092 3706
rect 19124 3674 19136 3706
rect 19168 3674 19180 3706
rect 19212 3674 19224 3706
rect 19256 3674 19271 3706
rect 19064 3670 19271 3674
rect 21630 3625 21762 3638
rect 246 3584 252 3612
rect 427 3584 433 3612
rect 18839 3584 18845 3612
rect 19020 3584 19026 3612
rect 21630 3419 21643 3625
rect 21749 3419 21762 3625
rect 21630 3407 21762 3419
rect 21346 3394 21514 3403
rect 21346 3319 21397 3394
rect 21503 3319 21514 3394
rect 21346 3312 21514 3319
rect 18828 3273 19035 3287
rect 18828 3241 18856 3273
rect 18888 3241 18900 3273
rect 18932 3241 18944 3273
rect 18976 3241 18988 3273
rect 19020 3241 19035 3273
rect 18828 3228 19035 3241
rect 18828 3196 18856 3228
rect 18888 3196 18900 3228
rect 18932 3196 18944 3228
rect 18976 3196 18988 3228
rect 19020 3196 19035 3228
rect 18828 3183 19035 3196
rect 18828 3172 18856 3183
rect 246 3144 252 3172
rect 427 3144 433 3172
rect 18828 3147 18845 3172
rect 18888 3172 18900 3183
rect 18932 3172 18944 3183
rect 18976 3172 18988 3183
rect 18839 3144 18845 3147
rect 19020 3147 19035 3183
rect 19020 3144 19026 3147
rect 21346 3123 21514 3132
rect 21346 3048 21397 3123
rect 21503 3048 21514 3123
rect 21346 3041 21514 3048
rect 19065 2776 19346 2915
rect 21346 2845 21514 2854
rect 19065 2762 19272 2776
rect 21346 2770 21397 2845
rect 21503 2770 21514 2845
rect 21346 2763 21514 2770
rect 246 2704 252 2732
rect 427 2704 433 2732
rect 19065 2730 19093 2762
rect 19125 2730 19137 2762
rect 19169 2730 19181 2762
rect 19213 2730 19225 2762
rect 19257 2730 19272 2762
rect 19065 2717 19272 2730
rect 19065 2685 19093 2717
rect 19125 2685 19137 2717
rect 19169 2685 19181 2717
rect 19213 2685 19225 2717
rect 19257 2685 19272 2717
rect 19065 2672 19272 2685
rect 19065 2640 19093 2672
rect 19125 2640 19137 2672
rect 19169 2640 19181 2672
rect 19213 2640 19225 2672
rect 19257 2640 19272 2672
rect 19065 2636 19272 2640
rect 21630 2746 21762 2759
rect 21630 2540 21643 2746
rect 21749 2540 21762 2746
rect 21630 2528 21762 2540
rect 246 2264 252 2292
rect 427 2264 433 2292
rect 18839 2290 18845 2292
rect 18828 2264 18845 2290
rect 19020 2290 19026 2292
rect 18828 2244 18856 2264
rect 18888 2244 18900 2264
rect 18932 2244 18944 2264
rect 18976 2244 18988 2264
rect 19020 2244 19346 2290
rect 18828 2231 19346 2244
rect 18828 2199 18856 2231
rect 18888 2199 18900 2231
rect 18932 2199 18944 2231
rect 18976 2199 18988 2231
rect 19020 2199 19346 2231
rect 18828 2186 19346 2199
rect 21346 2273 21762 2279
rect 21346 2192 21637 2273
rect 21756 2192 21762 2273
rect 21346 2187 21762 2192
rect 18828 2154 18856 2186
rect 18888 2154 18900 2186
rect 18932 2154 18944 2186
rect 18976 2154 18988 2186
rect 19020 2154 19346 2186
rect 18828 2150 19346 2154
rect 246 1824 252 1852
rect 427 1824 433 1852
rect 18839 1824 18845 1852
rect 19020 1824 19026 1852
rect 21346 1828 21762 1834
rect 19065 1760 19272 1774
rect 19065 1728 19093 1760
rect 19125 1728 19137 1760
rect 19169 1728 19181 1760
rect 19213 1728 19225 1760
rect 19257 1728 19272 1760
rect 21346 1747 21637 1828
rect 21756 1747 21762 1828
rect 21346 1742 21762 1747
rect 19065 1715 19272 1728
rect 19065 1683 19093 1715
rect 19125 1683 19137 1715
rect 19169 1683 19181 1715
rect 19213 1683 19225 1715
rect 19257 1683 19272 1715
rect 19065 1670 19272 1683
rect 19065 1638 19093 1670
rect 19125 1638 19137 1670
rect 19169 1638 19181 1670
rect 19213 1638 19225 1670
rect 19257 1638 19272 1670
rect 19065 1634 19272 1638
rect 21630 1625 21762 1638
rect 21630 1419 21643 1625
rect 21749 1419 21762 1625
rect 246 1384 252 1412
rect 427 1384 433 1412
rect 18839 1384 18845 1412
rect 19020 1384 19026 1412
rect 21630 1407 21762 1419
rect 21346 1394 21514 1403
rect 21346 1319 21397 1394
rect 21503 1319 21514 1394
rect 21346 1312 21514 1319
rect 18826 1276 19033 1290
rect 18826 1244 18854 1276
rect 18886 1244 18898 1276
rect 18930 1244 18942 1276
rect 18974 1244 18986 1276
rect 19018 1244 19033 1276
rect 18826 1231 19033 1244
rect 18826 1199 18854 1231
rect 18886 1199 18898 1231
rect 18930 1199 18942 1231
rect 18974 1199 18986 1231
rect 19018 1199 19033 1231
rect 18826 1186 19033 1199
rect 18826 1154 18854 1186
rect 18886 1154 18898 1186
rect 18930 1154 18942 1186
rect 18974 1154 18986 1186
rect 19018 1154 19033 1186
rect 18826 1150 19033 1154
rect 21346 1123 21514 1132
rect 21346 1048 21397 1123
rect 21503 1048 21514 1123
rect 21346 1041 21514 1048
rect 246 944 252 972
rect 427 944 433 972
rect 18839 944 18845 972
rect 19020 944 19026 972
rect 19065 776 19346 897
rect 21346 845 21514 854
rect 19065 763 19272 776
rect 21346 770 21397 845
rect 21503 770 21514 845
rect 21346 763 21514 770
rect 19065 731 19093 763
rect 19125 731 19137 763
rect 19169 731 19181 763
rect 19213 731 19225 763
rect 19257 731 19272 763
rect 19065 718 19272 731
rect 19065 686 19093 718
rect 19125 686 19137 718
rect 19169 686 19181 718
rect 19213 686 19225 718
rect 19257 686 19272 718
rect 19065 673 19272 686
rect 19065 641 19093 673
rect 19125 641 19137 673
rect 19169 641 19181 673
rect 19213 641 19225 673
rect 19257 641 19272 673
rect 19065 637 19272 641
rect 21630 746 21762 759
rect 21630 540 21643 746
rect 21749 540 21762 746
rect 246 504 252 532
rect 427 504 433 532
rect 18839 504 18845 532
rect 19020 504 19026 532
rect 21630 528 21762 540
rect 18827 431 19346 445
rect 18827 399 18855 431
rect 18887 399 18899 431
rect 18931 399 18943 431
rect 18975 399 18987 431
rect 19019 399 19346 431
rect 18827 386 19346 399
rect 238 366 445 380
rect 238 334 253 366
rect 285 334 297 366
rect 329 334 341 366
rect 373 334 385 366
rect 417 334 445 366
rect 238 321 445 334
rect 238 289 253 321
rect 285 289 297 321
rect 329 289 341 321
rect 373 289 385 321
rect 417 289 445 321
rect 238 276 445 289
rect 238 244 253 276
rect 285 244 297 276
rect 329 244 341 276
rect 373 244 385 276
rect 417 244 445 276
rect 238 240 445 244
rect 922 372 1104 381
rect 922 344 954 372
rect 982 344 1001 372
rect 1029 344 1048 372
rect 1076 344 1104 372
rect 922 325 1104 344
rect 922 297 954 325
rect 982 297 1001 325
rect 1029 297 1048 325
rect 1076 297 1104 325
rect 18827 354 18855 386
rect 18887 354 18899 386
rect 18931 354 18943 386
rect 18975 354 18987 386
rect 19019 354 19346 386
rect 18827 341 19346 354
rect 18827 309 18855 341
rect 18887 309 18899 341
rect 18931 309 18943 341
rect 18975 309 18987 341
rect 19019 309 19346 341
rect 18827 305 19346 309
rect 922 278 1104 297
rect 922 250 954 278
rect 982 250 1001 278
rect 1029 250 1048 278
rect 1076 250 1104 278
rect 922 240 1104 250
rect 21346 273 21762 279
rect 19065 212 19272 226
rect 19065 180 19093 212
rect 19125 180 19137 212
rect 19169 180 19181 212
rect 19213 180 19225 212
rect 19257 180 19272 212
rect 21346 192 21637 273
rect 21756 192 21762 273
rect 21346 187 21762 192
rect 19065 167 19272 180
rect 0 147 207 161
rect 0 115 15 147
rect 47 115 59 147
rect 91 115 103 147
rect 135 115 147 147
rect 179 115 207 147
rect 0 102 207 115
rect 0 70 15 102
rect 47 70 59 102
rect 91 70 103 102
rect 135 70 147 102
rect 179 70 207 102
rect 0 57 207 70
rect 0 25 15 57
rect 47 25 59 57
rect 91 25 103 57
rect 135 25 147 57
rect 179 25 207 57
rect 0 21 207 25
rect 733 153 915 162
rect 733 125 765 153
rect 793 125 812 153
rect 840 125 859 153
rect 887 125 915 153
rect 733 106 915 125
rect 733 78 765 106
rect 793 78 812 106
rect 840 78 859 106
rect 887 78 915 106
rect 19065 135 19093 167
rect 19125 135 19137 167
rect 19169 135 19181 167
rect 19213 135 19225 167
rect 19257 135 19272 167
rect 19065 122 19272 135
rect 19065 90 19093 122
rect 19125 90 19137 122
rect 19169 90 19181 122
rect 19213 90 19225 122
rect 19257 90 19272 122
rect 19065 86 19272 90
rect 733 59 915 78
rect 733 31 765 59
rect 793 31 812 59
rect 840 31 859 59
rect 887 31 915 59
rect 733 21 915 31
<< via2 >>
rect 21637 11747 21756 11828
rect 21643 11419 21749 11625
rect 21397 11319 21503 11394
rect 21397 11048 21503 11123
rect 21397 10770 21503 10845
rect 21643 10540 21749 10746
rect 21637 10192 21756 10273
rect 1494 9973 1625 10052
rect 3058 9973 3189 10052
rect 3494 9973 3625 10052
rect 5058 9973 5189 10052
rect 5494 9973 5625 10052
rect 7058 9973 7189 10052
rect 7494 9973 7625 10052
rect 9058 9973 9189 10052
rect 9494 9973 9625 10052
rect 11058 9973 11189 10052
rect 11494 9973 11625 10052
rect 13058 9973 13189 10052
rect 13494 9973 13625 10052
rect 15058 9973 15189 10052
rect 15494 9973 15625 10052
rect 17058 9973 17189 10052
rect 17494 9973 17625 10052
rect 19058 9990 19189 10052
rect 15 9914 47 9946
rect 59 9914 91 9946
rect 103 9914 135 9946
rect 147 9914 179 9946
rect 15 9869 47 9901
rect 59 9869 91 9901
rect 103 9869 135 9901
rect 147 9869 179 9901
rect 15 9824 47 9856
rect 59 9824 91 9856
rect 103 9824 135 9856
rect 147 9824 179 9856
rect 2267 9819 2430 9941
rect 4267 9819 4430 9941
rect 6267 9819 6430 9941
rect 8267 9819 8430 9941
rect 10267 9819 10430 9941
rect 12267 9819 12430 9941
rect 14267 9819 14430 9941
rect 16267 9819 16430 9941
rect 18267 9819 18430 9941
rect 19093 9914 19125 9946
rect 19137 9914 19169 9946
rect 19181 9914 19213 9946
rect 19225 9914 19257 9946
rect 19093 9869 19125 9901
rect 19137 9869 19169 9901
rect 19181 9869 19213 9901
rect 19225 9869 19257 9901
rect 19093 9824 19125 9856
rect 19137 9824 19169 9856
rect 19181 9824 19213 9856
rect 19225 9824 19257 9856
rect 21637 9747 21756 9828
rect 253 9695 285 9727
rect 297 9695 329 9727
rect 341 9695 373 9727
rect 385 9695 417 9727
rect 253 9650 285 9682
rect 297 9650 329 9682
rect 341 9650 373 9682
rect 385 9650 417 9682
rect 253 9605 285 9637
rect 297 9605 329 9637
rect 341 9605 373 9637
rect 385 9605 417 9637
rect 18855 9695 18887 9727
rect 18899 9695 18931 9727
rect 18943 9695 18975 9727
rect 18987 9695 19019 9727
rect 18855 9650 18887 9682
rect 18899 9650 18931 9682
rect 18943 9650 18975 9682
rect 18987 9650 19019 9682
rect 18855 9605 18887 9637
rect 18899 9605 18931 9637
rect 18943 9605 18975 9637
rect 18987 9605 19019 9637
rect 21643 9419 21749 9625
rect 252 9331 427 9332
rect 252 9305 427 9331
rect 252 9304 427 9305
rect 18845 9331 19020 9332
rect 18845 9305 19020 9331
rect 18845 9304 18856 9305
rect 18856 9284 18888 9305
rect 18888 9304 18900 9305
rect 18900 9284 18932 9305
rect 18932 9304 18944 9305
rect 18944 9284 18976 9305
rect 18976 9304 18988 9305
rect 18988 9284 19020 9305
rect 21397 9319 21503 9394
rect 18856 9239 18888 9271
rect 18900 9239 18932 9271
rect 18944 9239 18976 9271
rect 18988 9239 19020 9271
rect 18856 9194 18888 9226
rect 18900 9194 18932 9226
rect 18944 9194 18976 9226
rect 18988 9194 19020 9226
rect 21397 9048 21503 9123
rect 252 8891 427 8892
rect 252 8865 427 8891
rect 252 8864 427 8865
rect 18845 8891 19020 8892
rect 18845 8865 19020 8891
rect 18845 8864 19020 8865
rect 19093 8791 19125 8823
rect 19137 8791 19169 8823
rect 19181 8791 19213 8823
rect 19225 8791 19257 8823
rect 19093 8746 19125 8778
rect 19137 8746 19169 8778
rect 19181 8746 19213 8778
rect 19225 8746 19257 8778
rect 21397 8770 21503 8845
rect 19093 8701 19125 8733
rect 19137 8701 19169 8733
rect 19181 8701 19213 8733
rect 19225 8701 19257 8733
rect 21643 8540 21749 8746
rect 252 8451 427 8452
rect 252 8425 427 8451
rect 252 8424 427 8425
rect 18845 8451 19020 8452
rect 18845 8425 19020 8451
rect 18845 8424 19020 8425
rect 18855 8276 18887 8308
rect 18899 8276 18931 8308
rect 18943 8276 18975 8308
rect 18987 8276 19019 8308
rect 18855 8231 18887 8263
rect 18899 8231 18931 8263
rect 18943 8231 18975 8263
rect 18987 8231 19019 8263
rect 18855 8186 18887 8218
rect 18899 8186 18931 8218
rect 18943 8186 18975 8218
rect 18987 8186 19019 8218
rect 21637 8192 21756 8273
rect 252 8011 427 8012
rect 252 7985 427 8011
rect 252 7984 427 7985
rect 18845 8011 19020 8012
rect 18845 7985 19020 8011
rect 18845 7984 19020 7985
rect 19093 7737 19125 7769
rect 19137 7737 19169 7769
rect 19181 7737 19213 7769
rect 19225 7737 19257 7769
rect 21637 7747 21756 7828
rect 19093 7692 19125 7724
rect 19137 7692 19169 7724
rect 19181 7692 19213 7724
rect 19225 7692 19257 7724
rect 19093 7647 19125 7679
rect 19137 7647 19169 7679
rect 19181 7647 19213 7679
rect 19225 7647 19257 7679
rect 252 7571 427 7572
rect 252 7545 427 7571
rect 252 7544 427 7545
rect 18845 7571 19020 7572
rect 18845 7545 19020 7571
rect 18845 7544 19020 7545
rect 21643 7419 21749 7625
rect 21397 7319 21503 7394
rect 18855 7276 18887 7308
rect 18899 7276 18931 7308
rect 18943 7276 18975 7308
rect 18987 7276 19019 7308
rect 18855 7231 18887 7263
rect 18899 7231 18931 7263
rect 18943 7231 18975 7263
rect 18987 7231 19019 7263
rect 18855 7186 18887 7218
rect 18899 7186 18931 7218
rect 18943 7186 18975 7218
rect 18987 7186 19019 7218
rect 252 7131 427 7132
rect 252 7105 427 7131
rect 252 7104 427 7105
rect 18845 7131 19020 7132
rect 18845 7105 19020 7131
rect 18845 7104 19020 7105
rect 21397 7048 21503 7123
rect 19092 6772 19124 6804
rect 19136 6772 19168 6804
rect 19180 6772 19212 6804
rect 19224 6772 19256 6804
rect 21397 6770 21503 6845
rect 19092 6727 19124 6759
rect 19136 6727 19168 6759
rect 19180 6727 19212 6759
rect 19224 6727 19256 6759
rect 252 6691 427 6692
rect 252 6665 427 6691
rect 252 6664 427 6665
rect 19092 6682 19124 6714
rect 19136 6682 19168 6714
rect 19180 6682 19212 6714
rect 19224 6682 19256 6714
rect 21643 6540 21749 6746
rect 18856 6314 18888 6346
rect 18900 6314 18932 6346
rect 18944 6314 18976 6346
rect 18988 6314 19020 6346
rect 18856 6269 18888 6301
rect 18900 6269 18932 6301
rect 18944 6269 18976 6301
rect 18988 6269 19020 6301
rect 252 6251 427 6252
rect 252 6225 427 6251
rect 252 6224 427 6225
rect 18845 6251 18856 6252
rect 18856 6251 18888 6256
rect 18888 6251 18900 6252
rect 18900 6251 18932 6256
rect 18932 6251 18944 6252
rect 18944 6251 18976 6256
rect 18976 6251 18988 6252
rect 18988 6251 19020 6256
rect 18845 6225 19020 6251
rect 18845 6224 18856 6225
rect 18856 6224 18888 6225
rect 18888 6224 18900 6225
rect 18900 6224 18932 6225
rect 18932 6224 18944 6225
rect 18944 6224 18976 6225
rect 18976 6224 18988 6225
rect 18988 6224 19020 6225
rect 21637 6192 21756 6273
rect 252 5811 427 5812
rect 252 5785 427 5811
rect 252 5784 427 5785
rect 19093 5764 19125 5796
rect 19137 5764 19169 5796
rect 19181 5764 19213 5796
rect 19225 5764 19257 5796
rect 19093 5719 19125 5751
rect 19137 5719 19169 5751
rect 19181 5719 19213 5751
rect 19225 5719 19257 5751
rect 21637 5747 21756 5828
rect 19093 5674 19125 5706
rect 19137 5674 19169 5706
rect 19181 5674 19213 5706
rect 19225 5674 19257 5706
rect 21643 5419 21749 5625
rect 252 5371 427 5372
rect 252 5345 427 5371
rect 252 5344 427 5345
rect 18845 5371 19020 5372
rect 18845 5345 19020 5371
rect 18845 5344 19020 5345
rect 21397 5319 21503 5394
rect 18855 5251 18887 5283
rect 18899 5251 18931 5283
rect 18943 5251 18975 5283
rect 18987 5251 19019 5283
rect 18855 5206 18887 5238
rect 18899 5206 18931 5238
rect 18943 5206 18975 5238
rect 18987 5206 19019 5238
rect 18855 5161 18887 5193
rect 18899 5161 18931 5193
rect 18943 5161 18975 5193
rect 18987 5161 19019 5193
rect 21397 5048 21503 5123
rect 252 4931 427 4932
rect 252 4905 427 4931
rect 252 4904 427 4905
rect 18845 4931 19020 4932
rect 18845 4905 19020 4931
rect 18845 4904 19020 4905
rect 19093 4763 19125 4795
rect 19137 4763 19169 4795
rect 19181 4763 19213 4795
rect 19225 4763 19257 4795
rect 21397 4770 21503 4845
rect 19093 4718 19125 4750
rect 19137 4718 19169 4750
rect 19181 4718 19213 4750
rect 19225 4718 19257 4750
rect 19093 4673 19125 4705
rect 19137 4673 19169 4705
rect 19181 4673 19213 4705
rect 19225 4673 19257 4705
rect 21643 4540 21749 4746
rect 252 4491 427 4492
rect 252 4465 427 4491
rect 252 4464 427 4465
rect 18845 4491 19020 4492
rect 18845 4465 19020 4491
rect 18845 4464 19020 4465
rect 18856 4263 18888 4295
rect 18900 4263 18932 4295
rect 18944 4263 18976 4295
rect 18988 4263 19020 4295
rect 18856 4218 18888 4250
rect 18900 4218 18932 4250
rect 18944 4218 18976 4250
rect 18988 4218 19020 4250
rect 18856 4173 18888 4205
rect 18900 4173 18932 4205
rect 18944 4173 18976 4205
rect 18988 4173 19020 4205
rect 21637 4192 21756 4273
rect 252 4051 427 4052
rect 252 4025 427 4051
rect 252 4024 427 4025
rect 18845 4051 19020 4052
rect 18845 4025 19020 4051
rect 18845 4024 19020 4025
rect 19092 3764 19124 3796
rect 19136 3764 19168 3796
rect 19180 3764 19212 3796
rect 19224 3764 19256 3796
rect 19092 3719 19124 3751
rect 19136 3719 19168 3751
rect 19180 3719 19212 3751
rect 19224 3719 19256 3751
rect 21637 3747 21756 3828
rect 19092 3674 19124 3706
rect 19136 3674 19168 3706
rect 19180 3674 19212 3706
rect 19224 3674 19256 3706
rect 252 3611 427 3612
rect 252 3585 427 3611
rect 252 3584 427 3585
rect 18845 3611 19020 3612
rect 18845 3585 19020 3611
rect 18845 3584 19020 3585
rect 21643 3419 21749 3625
rect 21397 3319 21503 3394
rect 18856 3241 18888 3273
rect 18900 3241 18932 3273
rect 18944 3241 18976 3273
rect 18988 3241 19020 3273
rect 18856 3196 18888 3228
rect 18900 3196 18932 3228
rect 18944 3196 18976 3228
rect 18988 3196 19020 3228
rect 252 3171 427 3172
rect 252 3145 427 3171
rect 252 3144 427 3145
rect 18845 3171 18856 3172
rect 18856 3171 18888 3183
rect 18888 3171 18900 3172
rect 18900 3171 18932 3183
rect 18932 3171 18944 3172
rect 18944 3171 18976 3183
rect 18976 3171 18988 3172
rect 18988 3171 19020 3183
rect 18845 3145 19020 3171
rect 18845 3144 19020 3145
rect 21397 3048 21503 3123
rect 21397 2770 21503 2845
rect 252 2731 427 2732
rect 252 2705 427 2731
rect 252 2704 427 2705
rect 19093 2730 19125 2762
rect 19137 2730 19169 2762
rect 19181 2730 19213 2762
rect 19225 2730 19257 2762
rect 19093 2685 19125 2717
rect 19137 2685 19169 2717
rect 19181 2685 19213 2717
rect 19225 2685 19257 2717
rect 19093 2640 19125 2672
rect 19137 2640 19169 2672
rect 19181 2640 19213 2672
rect 19225 2640 19257 2672
rect 21643 2540 21749 2746
rect 252 2291 427 2292
rect 252 2265 427 2291
rect 252 2264 427 2265
rect 18845 2291 19020 2292
rect 18845 2265 19020 2291
rect 18845 2264 18856 2265
rect 18856 2244 18888 2265
rect 18888 2264 18900 2265
rect 18900 2244 18932 2265
rect 18932 2264 18944 2265
rect 18944 2244 18976 2265
rect 18976 2264 18988 2265
rect 18988 2244 19020 2265
rect 18856 2199 18888 2231
rect 18900 2199 18932 2231
rect 18944 2199 18976 2231
rect 18988 2199 19020 2231
rect 21637 2192 21756 2273
rect 18856 2154 18888 2186
rect 18900 2154 18932 2186
rect 18944 2154 18976 2186
rect 18988 2154 19020 2186
rect 252 1851 427 1852
rect 252 1825 427 1851
rect 252 1824 427 1825
rect 18845 1851 19020 1852
rect 18845 1825 19020 1851
rect 18845 1824 19020 1825
rect 19093 1728 19125 1760
rect 19137 1728 19169 1760
rect 19181 1728 19213 1760
rect 19225 1728 19257 1760
rect 21637 1747 21756 1828
rect 19093 1683 19125 1715
rect 19137 1683 19169 1715
rect 19181 1683 19213 1715
rect 19225 1683 19257 1715
rect 19093 1638 19125 1670
rect 19137 1638 19169 1670
rect 19181 1638 19213 1670
rect 19225 1638 19257 1670
rect 21643 1419 21749 1625
rect 252 1411 427 1412
rect 252 1385 427 1411
rect 252 1384 427 1385
rect 18845 1411 19020 1412
rect 18845 1385 19020 1411
rect 18845 1384 19020 1385
rect 21397 1319 21503 1394
rect 18854 1244 18886 1276
rect 18898 1244 18930 1276
rect 18942 1244 18974 1276
rect 18986 1244 19018 1276
rect 18854 1199 18886 1231
rect 18898 1199 18930 1231
rect 18942 1199 18974 1231
rect 18986 1199 19018 1231
rect 18854 1154 18886 1186
rect 18898 1154 18930 1186
rect 18942 1154 18974 1186
rect 18986 1154 19018 1186
rect 21397 1048 21503 1123
rect 252 971 427 972
rect 252 945 427 971
rect 252 944 427 945
rect 18845 971 19020 972
rect 18845 945 19020 971
rect 18845 944 19020 945
rect 21397 770 21503 845
rect 19093 731 19125 763
rect 19137 731 19169 763
rect 19181 731 19213 763
rect 19225 731 19257 763
rect 19093 686 19125 718
rect 19137 686 19169 718
rect 19181 686 19213 718
rect 19225 686 19257 718
rect 19093 641 19125 673
rect 19137 641 19169 673
rect 19181 641 19213 673
rect 19225 641 19257 673
rect 21643 540 21749 746
rect 252 531 427 532
rect 252 505 427 531
rect 252 504 427 505
rect 18845 531 19020 532
rect 18845 505 19020 531
rect 18845 504 19020 505
rect 18855 399 18887 431
rect 18899 399 18931 431
rect 18943 399 18975 431
rect 18987 399 19019 431
rect 253 334 285 366
rect 297 334 329 366
rect 341 334 373 366
rect 385 334 417 366
rect 253 289 285 321
rect 297 289 329 321
rect 341 289 373 321
rect 385 289 417 321
rect 253 244 285 276
rect 297 244 329 276
rect 341 244 373 276
rect 385 244 417 276
rect 954 344 982 372
rect 1001 344 1029 372
rect 1048 344 1076 372
rect 954 297 982 325
rect 1001 297 1029 325
rect 1048 297 1076 325
rect 18855 354 18887 386
rect 18899 354 18931 386
rect 18943 354 18975 386
rect 18987 354 19019 386
rect 18855 309 18887 341
rect 18899 309 18931 341
rect 18943 309 18975 341
rect 18987 309 19019 341
rect 954 250 982 278
rect 1001 250 1029 278
rect 1048 250 1076 278
rect 19093 180 19125 212
rect 19137 180 19169 212
rect 19181 180 19213 212
rect 19225 180 19257 212
rect 21637 192 21756 273
rect 15 115 47 147
rect 59 115 91 147
rect 103 115 135 147
rect 147 115 179 147
rect 15 70 47 102
rect 59 70 91 102
rect 103 70 135 102
rect 147 70 179 102
rect 15 25 47 57
rect 59 25 91 57
rect 103 25 135 57
rect 147 25 179 57
rect 765 125 793 153
rect 812 125 840 153
rect 859 125 887 153
rect 765 78 793 106
rect 812 78 840 106
rect 859 78 887 106
rect 19093 135 19125 167
rect 19137 135 19169 167
rect 19181 135 19213 167
rect 19225 135 19257 167
rect 19093 90 19125 122
rect 19137 90 19169 122
rect 19181 90 19213 122
rect 19225 90 19257 122
rect 765 31 793 59
rect 812 31 840 59
rect 859 31 887 59
<< metal3 >>
rect 21346 11828 21762 11834
rect 21346 11747 21637 11828
rect 21756 11747 21762 11828
rect 21346 11742 21762 11747
rect 21630 11625 21762 11638
rect 21630 11419 21643 11625
rect 21749 11419 21762 11625
rect 21630 11407 21762 11419
rect 21346 11394 21514 11403
rect 21346 11319 21397 11394
rect 21503 11319 21514 11394
rect 21346 11312 21514 11319
rect 21346 11123 21514 11132
rect 21346 11048 21397 11123
rect 21503 11048 21514 11123
rect 21346 11041 21514 11048
rect 21346 10845 21514 10854
rect 21346 10770 21397 10845
rect 21503 10770 21514 10845
rect 21346 10763 21514 10770
rect 21630 10746 21762 10759
rect 21630 10540 21643 10746
rect 21749 10540 21762 10746
rect 21630 10528 21762 10540
rect 21346 10273 21762 10279
rect 21346 10192 21637 10273
rect 21756 10192 21762 10273
rect 21346 10187 21762 10192
rect 1487 10052 1633 10084
rect 1487 9973 1494 10052
rect 1625 9973 1633 10052
rect 1487 9967 1633 9973
rect 3051 10052 3197 10083
rect 3051 9973 3058 10052
rect 3189 9973 3197 10052
rect 3051 9967 3197 9973
rect 3487 10052 3633 10083
rect 3487 9973 3494 10052
rect 3625 9973 3633 10052
rect 3487 9967 3633 9973
rect 5051 10052 5197 10083
rect 5051 9973 5058 10052
rect 5189 9973 5197 10052
rect 5051 9967 5197 9973
rect 5487 10052 5633 10083
rect 5487 9973 5494 10052
rect 5625 9973 5633 10052
rect 5487 9967 5633 9973
rect 7051 10052 7197 10083
rect 7051 9973 7058 10052
rect 7189 9973 7197 10052
rect 7051 9967 7197 9973
rect 7487 10052 7633 10083
rect 7487 9973 7494 10052
rect 7625 9973 7633 10052
rect 7487 9967 7633 9973
rect 9051 10052 9197 10083
rect 9051 9973 9058 10052
rect 9189 9973 9197 10052
rect 9051 9967 9197 9973
rect 9487 10052 9633 10083
rect 9487 9973 9494 10052
rect 9625 9973 9633 10052
rect 9487 9967 9633 9973
rect 11051 10052 11197 10083
rect 11051 9973 11058 10052
rect 11189 9973 11197 10052
rect 11051 9967 11197 9973
rect 11487 10052 11633 10083
rect 11487 9973 11494 10052
rect 11625 9973 11633 10052
rect 11487 9967 11633 9973
rect 13051 10052 13197 10083
rect 13051 9973 13058 10052
rect 13189 9973 13197 10052
rect 13051 9967 13197 9973
rect 13487 10052 13633 10083
rect 13487 9973 13494 10052
rect 13625 9973 13633 10052
rect 13487 9967 13633 9973
rect 15051 10052 15197 10083
rect 15051 9973 15058 10052
rect 15189 9973 15197 10052
rect 15051 9967 15197 9973
rect 15487 10052 15633 10083
rect 15487 9973 15494 10052
rect 15625 9973 15633 10052
rect 15487 9967 15633 9973
rect 17051 10052 17197 10083
rect 17051 9973 17058 10052
rect 17189 9973 17197 10052
rect 17051 9967 17197 9973
rect 17487 10052 17633 10083
rect 17487 9973 17494 10052
rect 17625 9973 17633 10052
rect 19051 10052 19197 10083
rect 19051 9990 19058 10052
rect 19189 9990 19197 10052
rect 19051 9984 19197 9990
rect 17487 9967 17633 9973
rect 0 9946 207 9950
rect 0 9914 15 9946
rect 47 9914 59 9946
rect 91 9914 103 9946
rect 135 9914 147 9946
rect 179 9914 207 9946
rect 0 9901 207 9914
rect 0 9869 15 9901
rect 47 9869 59 9901
rect 91 9869 103 9901
rect 135 9869 147 9901
rect 179 9869 207 9901
rect 0 9856 207 9869
rect 0 9824 15 9856
rect 47 9824 59 9856
rect 91 9824 103 9856
rect 135 9824 147 9856
rect 179 9824 207 9856
rect 0 9810 207 9824
rect 2255 9941 2440 9950
rect 2255 9819 2267 9941
rect 2430 9819 2440 9941
rect 2255 9810 2440 9819
rect 4255 9941 4440 9950
rect 4255 9819 4267 9941
rect 4430 9819 4440 9941
rect 4255 9810 4440 9819
rect 6255 9941 6440 9950
rect 6255 9819 6267 9941
rect 6430 9819 6440 9941
rect 6255 9810 6440 9819
rect 8255 9941 8440 9950
rect 8255 9819 8267 9941
rect 8430 9819 8440 9941
rect 8255 9810 8440 9819
rect 10255 9941 10440 9950
rect 10255 9819 10267 9941
rect 10430 9819 10440 9941
rect 10255 9810 10440 9819
rect 12255 9941 12440 9950
rect 12255 9819 12267 9941
rect 12430 9819 12440 9941
rect 12255 9810 12440 9819
rect 14255 9941 14440 9950
rect 14255 9819 14267 9941
rect 14430 9819 14440 9941
rect 14255 9810 14440 9819
rect 16255 9941 16440 9950
rect 16255 9819 16267 9941
rect 16430 9819 16440 9941
rect 16255 9810 16440 9819
rect 18255 9941 18440 9950
rect 18255 9819 18267 9941
rect 18430 9819 18440 9941
rect 18255 9810 18440 9819
rect 19065 9946 19272 9950
rect 19065 9914 19093 9946
rect 19125 9914 19137 9946
rect 19169 9914 19181 9946
rect 19213 9914 19225 9946
rect 19257 9914 19272 9946
rect 19065 9901 19272 9914
rect 19065 9869 19093 9901
rect 19125 9869 19137 9901
rect 19169 9869 19181 9901
rect 19213 9869 19225 9901
rect 19257 9869 19272 9901
rect 19065 9856 19272 9869
rect 19065 9824 19093 9856
rect 19125 9824 19137 9856
rect 19169 9824 19181 9856
rect 19213 9824 19225 9856
rect 19257 9824 19272 9856
rect 19065 9810 19272 9824
rect 21346 9828 21762 9834
rect 21346 9747 21637 9828
rect 21756 9747 21762 9828
rect 21346 9742 21762 9747
rect 238 9727 445 9731
rect 238 9695 253 9727
rect 285 9695 297 9727
rect 329 9695 341 9727
rect 373 9695 385 9727
rect 417 9695 445 9727
rect 238 9682 445 9695
rect 238 9650 253 9682
rect 285 9650 297 9682
rect 329 9650 341 9682
rect 373 9650 385 9682
rect 417 9650 445 9682
rect 238 9637 445 9650
rect 238 9605 253 9637
rect 285 9605 297 9637
rect 329 9605 341 9637
rect 373 9605 385 9637
rect 417 9605 445 9637
rect 238 9591 445 9605
rect 18827 9727 19034 9731
rect 18827 9695 18855 9727
rect 18887 9695 18899 9727
rect 18931 9695 18943 9727
rect 18975 9695 18987 9727
rect 19019 9695 19034 9727
rect 18827 9682 19034 9695
rect 18827 9650 18855 9682
rect 18887 9650 18899 9682
rect 18931 9650 18943 9682
rect 18975 9650 18987 9682
rect 19019 9650 19034 9682
rect 18827 9637 19034 9650
rect 18827 9605 18855 9637
rect 18887 9605 18899 9637
rect 18931 9605 18943 9637
rect 18975 9605 18987 9637
rect 19019 9605 19034 9637
rect 18827 9591 19034 9605
rect 21630 9625 21762 9638
rect 21630 9419 21643 9625
rect 21749 9419 21762 9625
rect 21630 9407 21762 9419
rect 21346 9394 21514 9403
rect 246 9334 433 9335
rect 246 9302 252 9334
rect 427 9302 433 9334
rect 18839 9334 19026 9335
rect 18839 9330 18845 9334
rect 246 9301 433 9302
rect 18828 9302 18845 9330
rect 19020 9330 19026 9334
rect 18828 9284 18856 9302
rect 18888 9284 18900 9302
rect 18932 9284 18944 9302
rect 18976 9284 18988 9302
rect 19020 9284 19035 9330
rect 21346 9319 21397 9394
rect 21503 9319 21514 9394
rect 21346 9312 21514 9319
rect 18828 9271 19035 9284
rect 18828 9239 18856 9271
rect 18888 9239 18900 9271
rect 18932 9239 18944 9271
rect 18976 9239 18988 9271
rect 19020 9239 19035 9271
rect 18828 9226 19035 9239
rect 18828 9194 18856 9226
rect 18888 9194 18900 9226
rect 18932 9194 18944 9226
rect 18976 9194 18988 9226
rect 19020 9194 19035 9226
rect 18828 9190 19035 9194
rect 21346 9123 21514 9132
rect 21346 9048 21397 9123
rect 21503 9048 21514 9123
rect 21346 9041 21514 9048
rect 246 8894 433 8895
rect 246 8862 252 8894
rect 427 8862 433 8894
rect 246 8861 433 8862
rect 18839 8894 19026 8895
rect 18839 8862 18845 8894
rect 19020 8862 19026 8894
rect 18839 8861 19026 8862
rect 21346 8845 21514 8854
rect 19065 8823 19272 8837
rect 19065 8791 19093 8823
rect 19125 8791 19137 8823
rect 19169 8791 19181 8823
rect 19213 8791 19225 8823
rect 19257 8791 19272 8823
rect 19065 8778 19272 8791
rect 19065 8746 19093 8778
rect 19125 8746 19137 8778
rect 19169 8746 19181 8778
rect 19213 8746 19225 8778
rect 19257 8746 19272 8778
rect 21346 8770 21397 8845
rect 21503 8770 21514 8845
rect 21346 8763 21514 8770
rect 19065 8733 19272 8746
rect 19065 8701 19093 8733
rect 19125 8701 19137 8733
rect 19169 8701 19181 8733
rect 19213 8701 19225 8733
rect 19257 8701 19272 8733
rect 19065 8697 19272 8701
rect 21630 8746 21762 8759
rect 21630 8540 21643 8746
rect 21749 8540 21762 8746
rect 21630 8528 21762 8540
rect 246 8454 433 8455
rect 246 8422 252 8454
rect 427 8422 433 8454
rect 246 8421 433 8422
rect 18839 8454 19026 8455
rect 18839 8422 18845 8454
rect 19020 8422 19026 8454
rect 18839 8421 19026 8422
rect 18827 8308 19346 8322
rect 18827 8276 18855 8308
rect 18887 8276 18899 8308
rect 18931 8276 18943 8308
rect 18975 8276 18987 8308
rect 19019 8276 19346 8308
rect 18827 8263 19346 8276
rect 18827 8231 18855 8263
rect 18887 8231 18899 8263
rect 18931 8231 18943 8263
rect 18975 8231 18987 8263
rect 19019 8231 19346 8263
rect 18827 8218 19346 8231
rect 18827 8186 18855 8218
rect 18887 8186 18899 8218
rect 18931 8186 18943 8218
rect 18975 8186 18987 8218
rect 19019 8186 19346 8218
rect 21346 8273 21762 8279
rect 21346 8192 21637 8273
rect 21756 8192 21762 8273
rect 21346 8187 21762 8192
rect 18827 8183 19346 8186
rect 18827 8182 19034 8183
rect 246 8014 433 8015
rect 246 7982 252 8014
rect 427 7982 433 8014
rect 246 7981 433 7982
rect 18839 8014 19026 8015
rect 18839 7982 18845 8014
rect 19020 7982 19026 8014
rect 18839 7981 19026 7982
rect 21346 7828 21762 7834
rect 19065 7769 19272 7783
rect 19065 7737 19093 7769
rect 19125 7737 19137 7769
rect 19169 7737 19181 7769
rect 19213 7737 19225 7769
rect 19257 7737 19272 7769
rect 21346 7747 21637 7828
rect 21756 7747 21762 7828
rect 21346 7742 21762 7747
rect 19065 7724 19272 7737
rect 19065 7692 19093 7724
rect 19125 7692 19137 7724
rect 19169 7692 19181 7724
rect 19213 7692 19225 7724
rect 19257 7692 19272 7724
rect 19065 7679 19272 7692
rect 19065 7647 19093 7679
rect 19125 7647 19137 7679
rect 19169 7647 19181 7679
rect 19213 7647 19225 7679
rect 19257 7647 19272 7679
rect 19065 7643 19272 7647
rect 21630 7625 21762 7638
rect 246 7574 433 7575
rect 246 7542 252 7574
rect 427 7542 433 7574
rect 246 7541 433 7542
rect 18839 7574 19026 7575
rect 18839 7542 18845 7574
rect 19020 7542 19026 7574
rect 18839 7541 19026 7542
rect 21630 7419 21643 7625
rect 21749 7419 21762 7625
rect 21630 7407 21762 7419
rect 21346 7394 21514 7403
rect 18827 7308 19034 7322
rect 21346 7319 21397 7394
rect 21503 7319 21514 7394
rect 21346 7312 21514 7319
rect 18827 7276 18855 7308
rect 18887 7276 18899 7308
rect 18931 7276 18943 7308
rect 18975 7276 18987 7308
rect 19019 7276 19034 7308
rect 18827 7263 19034 7276
rect 18827 7231 18855 7263
rect 18887 7231 18899 7263
rect 18931 7231 18943 7263
rect 18975 7231 18987 7263
rect 19019 7231 19034 7263
rect 18827 7218 19034 7231
rect 18827 7186 18855 7218
rect 18887 7186 18899 7218
rect 18931 7186 18943 7218
rect 18975 7186 18987 7218
rect 19019 7186 19034 7218
rect 18827 7183 19034 7186
rect 246 7134 433 7135
rect 246 7102 252 7134
rect 427 7102 433 7134
rect 246 7101 433 7102
rect 18839 7134 19026 7135
rect 18839 7102 18845 7134
rect 19020 7102 19026 7134
rect 18839 7101 19026 7102
rect 21346 7123 21514 7132
rect 21346 7048 21397 7123
rect 21503 7048 21514 7123
rect 21346 7041 21514 7048
rect 21346 6845 21514 6854
rect 19064 6804 19271 6818
rect 19064 6772 19092 6804
rect 19124 6772 19136 6804
rect 19168 6772 19180 6804
rect 19212 6772 19224 6804
rect 19256 6772 19271 6804
rect 19064 6759 19271 6772
rect 21346 6770 21397 6845
rect 21503 6770 21514 6845
rect 21346 6763 21514 6770
rect 19064 6727 19092 6759
rect 19124 6727 19136 6759
rect 19168 6727 19180 6759
rect 19212 6727 19224 6759
rect 19256 6727 19271 6759
rect 19064 6714 19271 6727
rect 246 6694 433 6695
rect 246 6662 252 6694
rect 427 6662 433 6694
rect 19064 6682 19092 6714
rect 19124 6682 19136 6714
rect 19168 6682 19180 6714
rect 19212 6682 19224 6714
rect 19256 6682 19271 6714
rect 19064 6678 19271 6682
rect 21630 6746 21762 6759
rect 246 6661 433 6662
rect 21630 6540 21643 6746
rect 21749 6540 21762 6746
rect 21630 6528 21762 6540
rect 18828 6359 19035 6360
rect 18828 6346 19346 6359
rect 18828 6314 18856 6346
rect 18888 6314 18900 6346
rect 18932 6314 18944 6346
rect 18976 6314 18988 6346
rect 19020 6314 19346 6346
rect 18828 6301 19346 6314
rect 18828 6269 18856 6301
rect 18888 6269 18900 6301
rect 18932 6269 18944 6301
rect 18976 6269 18988 6301
rect 19020 6269 19346 6301
rect 18828 6256 19346 6269
rect 246 6254 433 6255
rect 246 6222 252 6254
rect 427 6222 433 6254
rect 246 6221 433 6222
rect 18828 6254 18856 6256
rect 18828 6222 18845 6254
rect 18888 6254 18900 6256
rect 18932 6254 18944 6256
rect 18976 6254 18988 6256
rect 19020 6222 19346 6256
rect 18828 6220 19346 6222
rect 21346 6273 21762 6279
rect 21346 6192 21637 6273
rect 21756 6192 21762 6273
rect 21346 6187 21762 6192
rect 21346 5828 21762 5834
rect 246 5814 433 5815
rect 246 5782 252 5814
rect 427 5782 433 5814
rect 246 5781 433 5782
rect 19065 5796 19272 5810
rect 19065 5764 19093 5796
rect 19125 5764 19137 5796
rect 19169 5764 19181 5796
rect 19213 5764 19225 5796
rect 19257 5764 19272 5796
rect 19065 5751 19272 5764
rect 19065 5719 19093 5751
rect 19125 5719 19137 5751
rect 19169 5719 19181 5751
rect 19213 5719 19225 5751
rect 19257 5719 19272 5751
rect 21346 5747 21637 5828
rect 21756 5747 21762 5828
rect 21346 5742 21762 5747
rect 19065 5706 19272 5719
rect 19065 5674 19093 5706
rect 19125 5674 19137 5706
rect 19169 5674 19181 5706
rect 19213 5674 19225 5706
rect 19257 5674 19272 5706
rect 19065 5670 19272 5674
rect 21630 5625 21762 5638
rect 21630 5419 21643 5625
rect 21749 5419 21762 5625
rect 21630 5407 21762 5419
rect 21346 5394 21514 5403
rect 246 5374 433 5375
rect 246 5342 252 5374
rect 427 5342 433 5374
rect 246 5341 433 5342
rect 18839 5374 19026 5375
rect 18839 5342 18845 5374
rect 19020 5342 19026 5374
rect 18839 5341 19026 5342
rect 21346 5319 21397 5394
rect 21503 5319 21514 5394
rect 21346 5312 21514 5319
rect 18827 5283 19034 5297
rect 18827 5251 18855 5283
rect 18887 5251 18899 5283
rect 18931 5251 18943 5283
rect 18975 5251 18987 5283
rect 19019 5251 19034 5283
rect 18827 5238 19034 5251
rect 18827 5206 18855 5238
rect 18887 5206 18899 5238
rect 18931 5206 18943 5238
rect 18975 5206 18987 5238
rect 19019 5206 19034 5238
rect 18827 5193 19034 5206
rect 18827 5161 18855 5193
rect 18887 5161 18899 5193
rect 18931 5161 18943 5193
rect 18975 5161 18987 5193
rect 19019 5161 19034 5193
rect 18827 5157 19034 5161
rect 21346 5123 21514 5132
rect 21346 5048 21397 5123
rect 21503 5048 21514 5123
rect 21346 5041 21514 5048
rect 246 4934 433 4935
rect 246 4902 252 4934
rect 427 4902 433 4934
rect 246 4901 433 4902
rect 18839 4934 19026 4935
rect 18839 4902 18845 4934
rect 19020 4902 19026 4934
rect 18839 4901 19026 4902
rect 21346 4845 21514 4854
rect 19065 4795 19272 4809
rect 19065 4763 19093 4795
rect 19125 4763 19137 4795
rect 19169 4763 19181 4795
rect 19213 4763 19225 4795
rect 19257 4763 19272 4795
rect 21346 4770 21397 4845
rect 21503 4770 21514 4845
rect 21346 4763 21514 4770
rect 19065 4750 19272 4763
rect 19065 4718 19093 4750
rect 19125 4718 19137 4750
rect 19169 4718 19181 4750
rect 19213 4718 19225 4750
rect 19257 4718 19272 4750
rect 19065 4705 19272 4718
rect 19065 4673 19093 4705
rect 19125 4673 19137 4705
rect 19169 4673 19181 4705
rect 19213 4673 19225 4705
rect 19257 4673 19272 4705
rect 19065 4669 19272 4673
rect 21630 4746 21762 4759
rect 21630 4540 21643 4746
rect 21749 4540 21762 4746
rect 21630 4528 21762 4540
rect 246 4494 433 4495
rect 246 4462 252 4494
rect 427 4462 433 4494
rect 246 4461 433 4462
rect 18839 4494 19026 4495
rect 18839 4462 18845 4494
rect 19020 4462 19026 4494
rect 18839 4461 19026 4462
rect 18828 4308 19035 4309
rect 18828 4295 19346 4308
rect 18828 4263 18856 4295
rect 18888 4263 18900 4295
rect 18932 4263 18944 4295
rect 18976 4263 18988 4295
rect 19020 4263 19346 4295
rect 18828 4250 19346 4263
rect 18828 4218 18856 4250
rect 18888 4218 18900 4250
rect 18932 4218 18944 4250
rect 18976 4218 18988 4250
rect 19020 4218 19346 4250
rect 18828 4205 19346 4218
rect 18828 4173 18856 4205
rect 18888 4173 18900 4205
rect 18932 4173 18944 4205
rect 18976 4173 18988 4205
rect 19020 4173 19346 4205
rect 21346 4273 21762 4279
rect 21346 4192 21637 4273
rect 21756 4192 21762 4273
rect 21346 4187 21762 4192
rect 18828 4169 19346 4173
rect 246 4054 433 4055
rect 246 4022 252 4054
rect 427 4022 433 4054
rect 246 4021 433 4022
rect 18839 4054 19026 4055
rect 18839 4022 18845 4054
rect 19020 4022 19026 4054
rect 18839 4021 19026 4022
rect 21346 3828 21762 3834
rect 19064 3796 19271 3810
rect 19064 3764 19092 3796
rect 19124 3764 19136 3796
rect 19168 3764 19180 3796
rect 19212 3764 19224 3796
rect 19256 3764 19271 3796
rect 19064 3751 19271 3764
rect 19064 3719 19092 3751
rect 19124 3719 19136 3751
rect 19168 3719 19180 3751
rect 19212 3719 19224 3751
rect 19256 3719 19271 3751
rect 21346 3747 21637 3828
rect 21756 3747 21762 3828
rect 21346 3742 21762 3747
rect 19064 3706 19271 3719
rect 19064 3674 19092 3706
rect 19124 3674 19136 3706
rect 19168 3674 19180 3706
rect 19212 3674 19224 3706
rect 19256 3674 19271 3706
rect 19064 3670 19271 3674
rect 21630 3625 21762 3638
rect 246 3614 433 3615
rect 246 3582 252 3614
rect 427 3582 433 3614
rect 246 3581 433 3582
rect 18839 3614 19026 3615
rect 18839 3582 18845 3614
rect 19020 3582 19026 3614
rect 18839 3581 19026 3582
rect 21630 3419 21643 3625
rect 21749 3419 21762 3625
rect 21630 3407 21762 3419
rect 21346 3394 21514 3403
rect 21346 3319 21397 3394
rect 21503 3319 21514 3394
rect 21346 3312 21514 3319
rect 18828 3273 19035 3287
rect 18828 3241 18856 3273
rect 18888 3241 18900 3273
rect 18932 3241 18944 3273
rect 18976 3241 18988 3273
rect 19020 3241 19035 3273
rect 18828 3228 19035 3241
rect 18828 3196 18856 3228
rect 18888 3196 18900 3228
rect 18932 3196 18944 3228
rect 18976 3196 18988 3228
rect 19020 3196 19035 3228
rect 18828 3183 19035 3196
rect 246 3174 433 3175
rect 246 3142 252 3174
rect 427 3142 433 3174
rect 18828 3174 18856 3183
rect 18828 3147 18845 3174
rect 18888 3174 18900 3183
rect 18932 3174 18944 3183
rect 18976 3174 18988 3183
rect 246 3141 433 3142
rect 18839 3142 18845 3147
rect 19020 3147 19035 3183
rect 19020 3142 19026 3147
rect 18839 3141 19026 3142
rect 21346 3123 21514 3132
rect 21346 3048 21397 3123
rect 21503 3048 21514 3123
rect 21346 3041 21514 3048
rect 21346 2845 21514 2854
rect 19065 2762 19272 2776
rect 21346 2770 21397 2845
rect 21503 2770 21514 2845
rect 21346 2763 21514 2770
rect 246 2734 433 2735
rect 246 2702 252 2734
rect 427 2702 433 2734
rect 246 2701 433 2702
rect 19065 2730 19093 2762
rect 19125 2730 19137 2762
rect 19169 2730 19181 2762
rect 19213 2730 19225 2762
rect 19257 2730 19272 2762
rect 19065 2717 19272 2730
rect 19065 2685 19093 2717
rect 19125 2685 19137 2717
rect 19169 2685 19181 2717
rect 19213 2685 19225 2717
rect 19257 2685 19272 2717
rect 19065 2672 19272 2685
rect 19065 2640 19093 2672
rect 19125 2640 19137 2672
rect 19169 2640 19181 2672
rect 19213 2640 19225 2672
rect 19257 2640 19272 2672
rect 19065 2636 19272 2640
rect 21630 2746 21762 2759
rect 21630 2540 21643 2746
rect 21749 2540 21762 2746
rect 21630 2528 21762 2540
rect 246 2294 433 2295
rect 246 2262 252 2294
rect 427 2262 433 2294
rect 18839 2294 19026 2295
rect 18839 2290 18845 2294
rect 246 2261 433 2262
rect 18828 2262 18845 2290
rect 19020 2290 19026 2294
rect 18828 2244 18856 2262
rect 18888 2244 18900 2262
rect 18932 2244 18944 2262
rect 18976 2244 18988 2262
rect 19020 2244 19346 2290
rect 18828 2231 19346 2244
rect 18828 2199 18856 2231
rect 18888 2199 18900 2231
rect 18932 2199 18944 2231
rect 18976 2199 18988 2231
rect 19020 2199 19346 2231
rect 18828 2186 19346 2199
rect 21346 2273 21762 2279
rect 21346 2192 21637 2273
rect 21756 2192 21762 2273
rect 21346 2187 21762 2192
rect 18828 2154 18856 2186
rect 18888 2154 18900 2186
rect 18932 2154 18944 2186
rect 18976 2154 18988 2186
rect 19020 2154 19346 2186
rect 18828 2151 19346 2154
rect 18828 2150 19034 2151
rect 246 1854 433 1855
rect 246 1822 252 1854
rect 427 1822 433 1854
rect 246 1821 433 1822
rect 18839 1854 19026 1855
rect 18839 1822 18845 1854
rect 19020 1822 19026 1854
rect 18839 1821 19026 1822
rect 21346 1828 21762 1834
rect 19065 1760 19272 1774
rect 19065 1728 19093 1760
rect 19125 1728 19137 1760
rect 19169 1728 19181 1760
rect 19213 1728 19225 1760
rect 19257 1728 19272 1760
rect 21346 1747 21637 1828
rect 21756 1747 21762 1828
rect 21346 1742 21762 1747
rect 19065 1715 19272 1728
rect 19065 1683 19093 1715
rect 19125 1683 19137 1715
rect 19169 1683 19181 1715
rect 19213 1683 19225 1715
rect 19257 1683 19272 1715
rect 19065 1670 19272 1683
rect 19065 1638 19093 1670
rect 19125 1638 19137 1670
rect 19169 1638 19181 1670
rect 19213 1638 19225 1670
rect 19257 1638 19272 1670
rect 19065 1634 19272 1638
rect 21630 1625 21762 1638
rect 21630 1419 21643 1625
rect 21749 1419 21762 1625
rect 246 1414 433 1415
rect 246 1382 252 1414
rect 427 1382 433 1414
rect 246 1381 433 1382
rect 18839 1414 19026 1415
rect 18839 1382 18845 1414
rect 19020 1382 19026 1414
rect 21630 1407 21762 1419
rect 18839 1381 19026 1382
rect 21346 1394 21514 1403
rect 21346 1319 21397 1394
rect 21503 1319 21514 1394
rect 21346 1312 21514 1319
rect 18826 1276 19033 1290
rect 18826 1244 18854 1276
rect 18886 1244 18898 1276
rect 18930 1244 18942 1276
rect 18974 1244 18986 1276
rect 19018 1244 19033 1276
rect 18826 1231 19033 1244
rect 18826 1199 18854 1231
rect 18886 1199 18898 1231
rect 18930 1199 18942 1231
rect 18974 1199 18986 1231
rect 19018 1199 19033 1231
rect 18826 1186 19033 1199
rect 18826 1154 18854 1186
rect 18886 1154 18898 1186
rect 18930 1154 18942 1186
rect 18974 1154 18986 1186
rect 19018 1154 19033 1186
rect 18826 1150 19033 1154
rect 21346 1123 21514 1132
rect 21346 1048 21397 1123
rect 21503 1048 21514 1123
rect 21346 1041 21514 1048
rect 246 974 433 975
rect 246 942 252 974
rect 427 942 433 974
rect 246 941 433 942
rect 18839 974 19026 975
rect 18839 942 18845 974
rect 19020 942 19026 974
rect 18839 941 19026 942
rect 21346 845 21514 854
rect 19065 763 19272 777
rect 21346 770 21397 845
rect 21503 770 21514 845
rect 21346 763 21514 770
rect 19065 731 19093 763
rect 19125 731 19137 763
rect 19169 731 19181 763
rect 19213 731 19225 763
rect 19257 731 19272 763
rect 19065 718 19272 731
rect 19065 686 19093 718
rect 19125 686 19137 718
rect 19169 686 19181 718
rect 19213 686 19225 718
rect 19257 686 19272 718
rect 19065 673 19272 686
rect 19065 641 19093 673
rect 19125 641 19137 673
rect 19169 641 19181 673
rect 19213 641 19225 673
rect 19257 641 19272 673
rect 19065 637 19272 641
rect 21630 746 21762 759
rect 21630 540 21643 746
rect 21749 540 21762 746
rect 246 534 433 535
rect 246 502 252 534
rect 427 502 433 534
rect 246 501 433 502
rect 18839 534 19026 535
rect 18839 502 18845 534
rect 19020 502 19026 534
rect 21630 528 21762 540
rect 18839 501 19026 502
rect 18827 444 19034 445
rect 18827 431 19346 444
rect 18827 399 18855 431
rect 18887 399 18899 431
rect 18931 399 18943 431
rect 18975 399 18987 431
rect 19019 399 19346 431
rect 18827 386 19346 399
rect 237 372 1104 381
rect 237 366 954 372
rect 237 334 253 366
rect 285 334 297 366
rect 329 334 341 366
rect 373 334 385 366
rect 417 344 954 366
rect 982 344 1001 372
rect 1029 344 1048 372
rect 1076 344 1104 372
rect 417 334 1104 344
rect 237 325 1104 334
rect 237 321 954 325
rect 237 289 253 321
rect 285 289 297 321
rect 329 289 341 321
rect 373 289 385 321
rect 417 297 954 321
rect 982 297 1001 325
rect 1029 297 1048 325
rect 1076 297 1104 325
rect 18827 354 18855 386
rect 18887 354 18899 386
rect 18931 354 18943 386
rect 18975 354 18987 386
rect 19019 354 19346 386
rect 18827 341 19346 354
rect 18827 309 18855 341
rect 18887 309 18899 341
rect 18931 309 18943 341
rect 18975 309 18987 341
rect 19019 309 19346 341
rect 18827 305 19346 309
rect 417 289 1104 297
rect 237 278 1104 289
rect 237 276 954 278
rect 237 244 253 276
rect 285 244 297 276
rect 329 244 341 276
rect 373 244 385 276
rect 417 250 954 276
rect 982 250 1001 278
rect 1029 250 1048 278
rect 1076 250 1104 278
rect 417 244 1104 250
rect 237 240 1104 244
rect 21346 273 21762 279
rect 19065 212 19272 226
rect 19065 180 19093 212
rect 19125 180 19137 212
rect 19169 180 19181 212
rect 19213 180 19225 212
rect 19257 180 19272 212
rect 21346 192 21637 273
rect 21756 192 21762 273
rect 21346 187 21762 192
rect 19065 167 19272 180
rect 207 161 915 162
rect 0 153 915 161
rect 0 147 765 153
rect 0 115 15 147
rect 47 115 59 147
rect 91 115 103 147
rect 135 115 147 147
rect 179 125 765 147
rect 793 125 812 153
rect 840 125 859 153
rect 887 125 915 153
rect 179 115 915 125
rect 0 106 915 115
rect 0 102 765 106
rect 0 70 15 102
rect 47 70 59 102
rect 91 70 103 102
rect 135 70 147 102
rect 179 78 765 102
rect 793 78 812 106
rect 840 78 859 106
rect 887 78 915 106
rect 19065 135 19093 167
rect 19125 135 19137 167
rect 19169 135 19181 167
rect 19213 135 19225 167
rect 19257 135 19272 167
rect 19065 122 19272 135
rect 19065 90 19093 122
rect 19125 90 19137 122
rect 19169 90 19181 122
rect 19213 90 19225 122
rect 19257 90 19272 122
rect 19065 86 19272 90
rect 179 70 915 78
rect 0 59 915 70
rect 0 57 765 59
rect 0 25 15 57
rect 47 25 59 57
rect 91 25 103 57
rect 135 25 147 57
rect 179 31 765 57
rect 793 31 812 59
rect 840 31 859 59
rect 887 31 915 59
rect 179 25 915 31
rect 0 21 915 25
<< via3 >>
rect 21637 11747 21756 11828
rect 21643 11419 21749 11625
rect 21397 11319 21503 11394
rect 21397 11048 21503 11123
rect 21397 10770 21503 10845
rect 21643 10540 21749 10746
rect 21637 10192 21756 10273
rect 15 9914 47 9946
rect 59 9914 91 9946
rect 103 9914 135 9946
rect 147 9914 179 9946
rect 15 9869 47 9901
rect 59 9869 91 9901
rect 103 9869 135 9901
rect 147 9869 179 9901
rect 15 9824 47 9856
rect 59 9824 91 9856
rect 103 9824 135 9856
rect 147 9824 179 9856
rect 2267 9819 2430 9941
rect 4267 9819 4430 9941
rect 6267 9819 6430 9941
rect 8267 9819 8430 9941
rect 10267 9819 10430 9941
rect 12267 9819 12430 9941
rect 14267 9819 14430 9941
rect 16267 9819 16430 9941
rect 18267 9819 18430 9941
rect 19093 9914 19125 9946
rect 19137 9914 19169 9946
rect 19181 9914 19213 9946
rect 19225 9914 19257 9946
rect 19093 9869 19125 9901
rect 19137 9869 19169 9901
rect 19181 9869 19213 9901
rect 19225 9869 19257 9901
rect 19093 9824 19125 9856
rect 19137 9824 19169 9856
rect 19181 9824 19213 9856
rect 19225 9824 19257 9856
rect 21637 9747 21756 9828
rect 253 9695 285 9727
rect 297 9695 329 9727
rect 341 9695 373 9727
rect 385 9695 417 9727
rect 253 9650 285 9682
rect 297 9650 329 9682
rect 341 9650 373 9682
rect 385 9650 417 9682
rect 253 9605 285 9637
rect 297 9605 329 9637
rect 341 9605 373 9637
rect 385 9605 417 9637
rect 18855 9695 18887 9727
rect 18899 9695 18931 9727
rect 18943 9695 18975 9727
rect 18987 9695 19019 9727
rect 18855 9650 18887 9682
rect 18899 9650 18931 9682
rect 18943 9650 18975 9682
rect 18987 9650 19019 9682
rect 18855 9605 18887 9637
rect 18899 9605 18931 9637
rect 18943 9605 18975 9637
rect 18987 9605 19019 9637
rect 21643 9419 21749 9625
rect 252 9332 427 9334
rect 252 9304 427 9332
rect 252 9302 427 9304
rect 18845 9332 19020 9334
rect 18845 9304 19020 9332
rect 18845 9302 18856 9304
rect 18856 9284 18888 9304
rect 18888 9302 18900 9304
rect 18900 9284 18932 9304
rect 18932 9302 18944 9304
rect 18944 9284 18976 9304
rect 18976 9302 18988 9304
rect 18988 9284 19020 9304
rect 21397 9319 21503 9394
rect 18856 9239 18888 9271
rect 18900 9239 18932 9271
rect 18944 9239 18976 9271
rect 18988 9239 19020 9271
rect 18856 9194 18888 9226
rect 18900 9194 18932 9226
rect 18944 9194 18976 9226
rect 18988 9194 19020 9226
rect 21397 9048 21503 9123
rect 252 8892 427 8894
rect 252 8864 427 8892
rect 252 8862 427 8864
rect 18845 8892 19020 8894
rect 18845 8864 19020 8892
rect 18845 8862 19020 8864
rect 19093 8791 19125 8823
rect 19137 8791 19169 8823
rect 19181 8791 19213 8823
rect 19225 8791 19257 8823
rect 19093 8746 19125 8778
rect 19137 8746 19169 8778
rect 19181 8746 19213 8778
rect 19225 8746 19257 8778
rect 21397 8770 21503 8845
rect 19093 8701 19125 8733
rect 19137 8701 19169 8733
rect 19181 8701 19213 8733
rect 19225 8701 19257 8733
rect 21643 8540 21749 8746
rect 252 8452 427 8454
rect 252 8424 427 8452
rect 252 8422 427 8424
rect 18845 8452 19020 8454
rect 18845 8424 19020 8452
rect 18845 8422 19020 8424
rect 18855 8276 18887 8308
rect 18899 8276 18931 8308
rect 18943 8276 18975 8308
rect 18987 8276 19019 8308
rect 18855 8231 18887 8263
rect 18899 8231 18931 8263
rect 18943 8231 18975 8263
rect 18987 8231 19019 8263
rect 18855 8186 18887 8218
rect 18899 8186 18931 8218
rect 18943 8186 18975 8218
rect 18987 8186 19019 8218
rect 21637 8192 21756 8273
rect 252 8012 427 8014
rect 252 7984 427 8012
rect 252 7982 427 7984
rect 18845 8012 19020 8014
rect 18845 7984 19020 8012
rect 18845 7982 19020 7984
rect 19093 7737 19125 7769
rect 19137 7737 19169 7769
rect 19181 7737 19213 7769
rect 19225 7737 19257 7769
rect 21637 7747 21756 7828
rect 19093 7692 19125 7724
rect 19137 7692 19169 7724
rect 19181 7692 19213 7724
rect 19225 7692 19257 7724
rect 19093 7647 19125 7679
rect 19137 7647 19169 7679
rect 19181 7647 19213 7679
rect 19225 7647 19257 7679
rect 252 7572 427 7574
rect 252 7544 427 7572
rect 252 7542 427 7544
rect 18845 7572 19020 7574
rect 18845 7544 19020 7572
rect 18845 7542 19020 7544
rect 21643 7419 21749 7625
rect 21397 7319 21503 7394
rect 18855 7276 18887 7308
rect 18899 7276 18931 7308
rect 18943 7276 18975 7308
rect 18987 7276 19019 7308
rect 18855 7231 18887 7263
rect 18899 7231 18931 7263
rect 18943 7231 18975 7263
rect 18987 7231 19019 7263
rect 18855 7186 18887 7218
rect 18899 7186 18931 7218
rect 18943 7186 18975 7218
rect 18987 7186 19019 7218
rect 252 7132 427 7134
rect 252 7104 427 7132
rect 252 7102 427 7104
rect 18845 7132 19020 7134
rect 18845 7104 19020 7132
rect 18845 7102 19020 7104
rect 21397 7048 21503 7123
rect 19092 6772 19124 6804
rect 19136 6772 19168 6804
rect 19180 6772 19212 6804
rect 19224 6772 19256 6804
rect 21397 6770 21503 6845
rect 19092 6727 19124 6759
rect 19136 6727 19168 6759
rect 19180 6727 19212 6759
rect 19224 6727 19256 6759
rect 252 6692 427 6694
rect 252 6664 427 6692
rect 252 6662 427 6664
rect 19092 6682 19124 6714
rect 19136 6682 19168 6714
rect 19180 6682 19212 6714
rect 19224 6682 19256 6714
rect 21643 6540 21749 6746
rect 18856 6314 18888 6346
rect 18900 6314 18932 6346
rect 18944 6314 18976 6346
rect 18988 6314 19020 6346
rect 18856 6269 18888 6301
rect 18900 6269 18932 6301
rect 18944 6269 18976 6301
rect 18988 6269 19020 6301
rect 252 6252 427 6254
rect 252 6224 427 6252
rect 252 6222 427 6224
rect 18845 6252 18856 6254
rect 18856 6252 18888 6256
rect 18888 6252 18900 6254
rect 18900 6252 18932 6256
rect 18932 6252 18944 6254
rect 18944 6252 18976 6256
rect 18976 6252 18988 6254
rect 18988 6252 19020 6256
rect 18845 6224 19020 6252
rect 18845 6222 19020 6224
rect 21637 6192 21756 6273
rect 252 5812 427 5814
rect 252 5784 427 5812
rect 252 5782 427 5784
rect 19093 5764 19125 5796
rect 19137 5764 19169 5796
rect 19181 5764 19213 5796
rect 19225 5764 19257 5796
rect 19093 5719 19125 5751
rect 19137 5719 19169 5751
rect 19181 5719 19213 5751
rect 19225 5719 19257 5751
rect 21637 5747 21756 5828
rect 19093 5674 19125 5706
rect 19137 5674 19169 5706
rect 19181 5674 19213 5706
rect 19225 5674 19257 5706
rect 21643 5419 21749 5625
rect 252 5372 427 5374
rect 252 5344 427 5372
rect 252 5342 427 5344
rect 18845 5372 19020 5374
rect 18845 5344 19020 5372
rect 18845 5342 19020 5344
rect 21397 5319 21503 5394
rect 18855 5251 18887 5283
rect 18899 5251 18931 5283
rect 18943 5251 18975 5283
rect 18987 5251 19019 5283
rect 18855 5206 18887 5238
rect 18899 5206 18931 5238
rect 18943 5206 18975 5238
rect 18987 5206 19019 5238
rect 18855 5161 18887 5193
rect 18899 5161 18931 5193
rect 18943 5161 18975 5193
rect 18987 5161 19019 5193
rect 21397 5048 21503 5123
rect 252 4932 427 4934
rect 252 4904 427 4932
rect 252 4902 427 4904
rect 18845 4932 19020 4934
rect 18845 4904 19020 4932
rect 18845 4902 19020 4904
rect 19093 4763 19125 4795
rect 19137 4763 19169 4795
rect 19181 4763 19213 4795
rect 19225 4763 19257 4795
rect 21397 4770 21503 4845
rect 19093 4718 19125 4750
rect 19137 4718 19169 4750
rect 19181 4718 19213 4750
rect 19225 4718 19257 4750
rect 19093 4673 19125 4705
rect 19137 4673 19169 4705
rect 19181 4673 19213 4705
rect 19225 4673 19257 4705
rect 21643 4540 21749 4746
rect 252 4492 427 4494
rect 252 4464 427 4492
rect 252 4462 427 4464
rect 18845 4492 19020 4494
rect 18845 4464 19020 4492
rect 18845 4462 19020 4464
rect 18856 4263 18888 4295
rect 18900 4263 18932 4295
rect 18944 4263 18976 4295
rect 18988 4263 19020 4295
rect 18856 4218 18888 4250
rect 18900 4218 18932 4250
rect 18944 4218 18976 4250
rect 18988 4218 19020 4250
rect 18856 4173 18888 4205
rect 18900 4173 18932 4205
rect 18944 4173 18976 4205
rect 18988 4173 19020 4205
rect 21637 4192 21756 4273
rect 252 4052 427 4054
rect 252 4024 427 4052
rect 252 4022 427 4024
rect 18845 4052 19020 4054
rect 18845 4024 19020 4052
rect 18845 4022 19020 4024
rect 19092 3764 19124 3796
rect 19136 3764 19168 3796
rect 19180 3764 19212 3796
rect 19224 3764 19256 3796
rect 19092 3719 19124 3751
rect 19136 3719 19168 3751
rect 19180 3719 19212 3751
rect 19224 3719 19256 3751
rect 21637 3747 21756 3828
rect 19092 3674 19124 3706
rect 19136 3674 19168 3706
rect 19180 3674 19212 3706
rect 19224 3674 19256 3706
rect 252 3612 427 3614
rect 252 3584 427 3612
rect 252 3582 427 3584
rect 18845 3612 19020 3614
rect 18845 3584 19020 3612
rect 18845 3582 19020 3584
rect 21643 3419 21749 3625
rect 21397 3319 21503 3394
rect 18856 3241 18888 3273
rect 18900 3241 18932 3273
rect 18944 3241 18976 3273
rect 18988 3241 19020 3273
rect 18856 3196 18888 3228
rect 18900 3196 18932 3228
rect 18944 3196 18976 3228
rect 18988 3196 19020 3228
rect 252 3172 427 3174
rect 252 3144 427 3172
rect 252 3142 427 3144
rect 18845 3172 18856 3174
rect 18856 3172 18888 3183
rect 18888 3172 18900 3174
rect 18900 3172 18932 3183
rect 18932 3172 18944 3174
rect 18944 3172 18976 3183
rect 18976 3172 18988 3174
rect 18988 3172 19020 3183
rect 18845 3144 19020 3172
rect 18845 3142 19020 3144
rect 21397 3048 21503 3123
rect 21397 2770 21503 2845
rect 252 2732 427 2734
rect 252 2704 427 2732
rect 252 2702 427 2704
rect 19093 2730 19125 2762
rect 19137 2730 19169 2762
rect 19181 2730 19213 2762
rect 19225 2730 19257 2762
rect 19093 2685 19125 2717
rect 19137 2685 19169 2717
rect 19181 2685 19213 2717
rect 19225 2685 19257 2717
rect 19093 2640 19125 2672
rect 19137 2640 19169 2672
rect 19181 2640 19213 2672
rect 19225 2640 19257 2672
rect 21643 2540 21749 2746
rect 252 2292 427 2294
rect 252 2264 427 2292
rect 252 2262 427 2264
rect 18845 2292 19020 2294
rect 18845 2264 19020 2292
rect 18845 2262 18856 2264
rect 18856 2244 18888 2264
rect 18888 2262 18900 2264
rect 18900 2244 18932 2264
rect 18932 2262 18944 2264
rect 18944 2244 18976 2264
rect 18976 2262 18988 2264
rect 18988 2244 19020 2264
rect 18856 2199 18888 2231
rect 18900 2199 18932 2231
rect 18944 2199 18976 2231
rect 18988 2199 19020 2231
rect 21637 2192 21756 2273
rect 18856 2154 18888 2186
rect 18900 2154 18932 2186
rect 18944 2154 18976 2186
rect 18988 2154 19020 2186
rect 252 1852 427 1854
rect 252 1824 427 1852
rect 252 1822 427 1824
rect 18845 1852 19020 1854
rect 18845 1824 19020 1852
rect 18845 1822 19020 1824
rect 19093 1728 19125 1760
rect 19137 1728 19169 1760
rect 19181 1728 19213 1760
rect 19225 1728 19257 1760
rect 21637 1747 21756 1828
rect 19093 1683 19125 1715
rect 19137 1683 19169 1715
rect 19181 1683 19213 1715
rect 19225 1683 19257 1715
rect 19093 1638 19125 1670
rect 19137 1638 19169 1670
rect 19181 1638 19213 1670
rect 19225 1638 19257 1670
rect 21643 1419 21749 1625
rect 252 1412 427 1414
rect 252 1384 427 1412
rect 252 1382 427 1384
rect 18845 1412 19020 1414
rect 18845 1384 19020 1412
rect 18845 1382 19020 1384
rect 21397 1319 21503 1394
rect 18854 1244 18886 1276
rect 18898 1244 18930 1276
rect 18942 1244 18974 1276
rect 18986 1244 19018 1276
rect 18854 1199 18886 1231
rect 18898 1199 18930 1231
rect 18942 1199 18974 1231
rect 18986 1199 19018 1231
rect 18854 1154 18886 1186
rect 18898 1154 18930 1186
rect 18942 1154 18974 1186
rect 18986 1154 19018 1186
rect 21397 1048 21503 1123
rect 252 972 427 974
rect 252 944 427 972
rect 252 942 427 944
rect 18845 972 19020 974
rect 18845 944 19020 972
rect 18845 942 19020 944
rect 21397 770 21503 845
rect 19093 731 19125 763
rect 19137 731 19169 763
rect 19181 731 19213 763
rect 19225 731 19257 763
rect 19093 686 19125 718
rect 19137 686 19169 718
rect 19181 686 19213 718
rect 19225 686 19257 718
rect 19093 641 19125 673
rect 19137 641 19169 673
rect 19181 641 19213 673
rect 19225 641 19257 673
rect 21643 540 21749 746
rect 252 532 427 534
rect 252 504 427 532
rect 252 502 427 504
rect 18845 532 19020 534
rect 18845 504 19020 532
rect 18845 502 19020 504
rect 18855 399 18887 431
rect 18899 399 18931 431
rect 18943 399 18975 431
rect 18987 399 19019 431
rect 253 334 285 366
rect 297 334 329 366
rect 341 334 373 366
rect 385 334 417 366
rect 253 289 285 321
rect 297 289 329 321
rect 341 289 373 321
rect 385 289 417 321
rect 18855 354 18887 386
rect 18899 354 18931 386
rect 18943 354 18975 386
rect 18987 354 19019 386
rect 18855 309 18887 341
rect 18899 309 18931 341
rect 18943 309 18975 341
rect 18987 309 19019 341
rect 253 244 285 276
rect 297 244 329 276
rect 341 244 373 276
rect 385 244 417 276
rect 19093 180 19125 212
rect 19137 180 19169 212
rect 19181 180 19213 212
rect 19225 180 19257 212
rect 21637 192 21756 273
rect 15 115 47 147
rect 59 115 91 147
rect 103 115 135 147
rect 147 115 179 147
rect 15 70 47 102
rect 59 70 91 102
rect 103 70 135 102
rect 147 70 179 102
rect 19093 135 19125 167
rect 19137 135 19169 167
rect 19181 135 19213 167
rect 19225 135 19257 167
rect 19093 90 19125 122
rect 19137 90 19169 122
rect 19181 90 19213 122
rect 19225 90 19257 122
rect 15 25 47 57
rect 59 25 91 57
rect 103 25 135 57
rect 147 25 179 57
<< metal4 >>
rect 0 9946 207 12083
rect 0 9914 15 9946
rect 47 9914 59 9946
rect 91 9914 103 9946
rect 135 9914 147 9946
rect 179 9914 207 9946
rect 0 9901 207 9914
rect 0 9869 15 9901
rect 47 9869 59 9901
rect 91 9869 103 9901
rect 135 9869 147 9901
rect 179 9869 207 9901
rect 0 9856 207 9869
rect 0 9824 15 9856
rect 47 9824 59 9856
rect 91 9824 103 9856
rect 135 9824 147 9856
rect 179 9824 207 9856
rect 0 147 207 9824
rect 0 115 15 147
rect 47 115 59 147
rect 91 115 103 147
rect 135 115 147 147
rect 179 115 207 147
rect 0 102 207 115
rect 0 70 15 102
rect 47 70 59 102
rect 91 70 103 102
rect 135 70 147 102
rect 179 70 207 102
rect 0 57 207 70
rect 0 25 15 57
rect 47 25 59 57
rect 91 25 103 57
rect 135 25 147 57
rect 179 25 207 57
rect 0 21 207 25
rect 238 9727 445 12083
rect 21386 11403 21593 12083
rect 21346 11394 21593 11403
rect 21346 11319 21397 11394
rect 21503 11319 21593 11394
rect 21346 11312 21593 11319
rect 21386 11132 21593 11312
rect 21346 11123 21593 11132
rect 21346 11048 21397 11123
rect 21503 11048 21593 11123
rect 21346 11041 21593 11048
rect 21386 10854 21593 11041
rect 21346 10845 21593 10854
rect 21346 10770 21397 10845
rect 21503 10770 21593 10845
rect 21346 10763 21593 10770
rect 2255 9941 2440 10083
rect 2255 9819 2267 9941
rect 2430 9819 2440 9941
rect 2255 9810 2440 9819
rect 4255 9941 4440 10083
rect 4255 9819 4267 9941
rect 4430 9819 4440 9941
rect 4255 9810 4440 9819
rect 6255 9941 6440 10083
rect 6255 9819 6267 9941
rect 6430 9819 6440 9941
rect 6255 9810 6440 9819
rect 8255 9941 8440 10083
rect 8255 9819 8267 9941
rect 8430 9819 8440 9941
rect 8255 9810 8440 9819
rect 10255 9941 10440 10083
rect 10255 9819 10267 9941
rect 10430 9819 10440 9941
rect 10255 9810 10440 9819
rect 12255 9941 12440 10083
rect 12255 9819 12267 9941
rect 12430 9819 12440 9941
rect 12255 9810 12440 9819
rect 14255 9941 14440 10083
rect 14255 9819 14267 9941
rect 14430 9819 14440 9941
rect 14255 9810 14440 9819
rect 16255 9941 16440 10083
rect 16255 9819 16267 9941
rect 16430 9819 16440 9941
rect 16255 9810 16440 9819
rect 18255 9941 18440 10083
rect 18255 9819 18267 9941
rect 18430 9819 18440 9941
rect 18255 9810 18440 9819
rect 238 9695 253 9727
rect 285 9695 297 9727
rect 329 9695 341 9727
rect 373 9695 385 9727
rect 417 9695 445 9727
rect 238 9682 445 9695
rect 238 9650 253 9682
rect 285 9650 297 9682
rect 329 9650 341 9682
rect 373 9650 385 9682
rect 417 9650 445 9682
rect 238 9637 445 9650
rect 238 9605 253 9637
rect 285 9605 297 9637
rect 329 9605 341 9637
rect 373 9605 385 9637
rect 417 9605 445 9637
rect 238 9334 445 9605
rect 238 9302 252 9334
rect 427 9302 445 9334
rect 238 8894 445 9302
rect 18827 9727 19034 9951
rect 18827 9695 18855 9727
rect 18887 9695 18899 9727
rect 18931 9695 18943 9727
rect 18975 9695 18987 9727
rect 19019 9695 19034 9727
rect 18827 9682 19034 9695
rect 18827 9650 18855 9682
rect 18887 9650 18899 9682
rect 18931 9650 18943 9682
rect 18975 9650 18987 9682
rect 19019 9650 19034 9682
rect 18827 9637 19034 9650
rect 18827 9605 18855 9637
rect 18887 9605 18899 9637
rect 18931 9605 18943 9637
rect 18975 9605 18987 9637
rect 19019 9605 19034 9637
rect 18827 9334 19034 9605
rect 18827 9302 18845 9334
rect 19020 9331 19034 9334
rect 19065 9946 19272 9951
rect 19065 9914 19093 9946
rect 19125 9914 19137 9946
rect 19169 9914 19181 9946
rect 19213 9914 19225 9946
rect 19257 9914 19272 9946
rect 19065 9901 19272 9914
rect 19065 9869 19093 9901
rect 19125 9869 19137 9901
rect 19169 9869 19181 9901
rect 19213 9869 19225 9901
rect 19257 9869 19272 9901
rect 19065 9856 19272 9869
rect 19065 9824 19093 9856
rect 19125 9824 19137 9856
rect 19169 9824 19181 9856
rect 19213 9824 19225 9856
rect 19257 9824 19272 9856
rect 18827 9284 18856 9302
rect 18888 9284 18900 9302
rect 18932 9284 18944 9302
rect 18976 9284 18988 9302
rect 19020 9284 19035 9331
rect 18827 9271 19035 9284
rect 18827 9239 18856 9271
rect 18888 9239 18900 9271
rect 18932 9239 18944 9271
rect 18976 9239 18988 9271
rect 19020 9239 19035 9271
rect 18827 9226 19035 9239
rect 18827 9194 18856 9226
rect 18888 9194 18900 9226
rect 18932 9194 18944 9226
rect 18976 9194 18988 9226
rect 19020 9194 19035 9226
rect 18827 9190 19035 9194
rect 238 8862 252 8894
rect 427 8862 445 8894
rect 2164 8869 2234 8899
rect 2666 8869 2736 8899
rect 3168 8869 3238 8899
rect 3670 8869 3740 8899
rect 4172 8869 4242 8899
rect 4674 8869 4744 8899
rect 5176 8869 5246 8899
rect 5678 8869 5748 8899
rect 6180 8869 6250 8899
rect 6682 8869 6752 8899
rect 7184 8869 7254 8899
rect 7686 8869 7756 8899
rect 8188 8869 8258 8899
rect 8690 8869 8760 8899
rect 9192 8869 9262 8899
rect 9694 8869 9764 8899
rect 10196 8869 10266 8899
rect 10698 8869 10768 8899
rect 11200 8869 11270 8899
rect 11702 8869 11772 8899
rect 12204 8869 12274 8899
rect 12706 8869 12776 8899
rect 13208 8869 13278 8899
rect 13710 8869 13780 8899
rect 14212 8869 14282 8899
rect 14714 8869 14784 8899
rect 15216 8869 15286 8899
rect 15718 8869 15788 8899
rect 16220 8869 16290 8899
rect 16722 8869 16792 8899
rect 17224 8869 17294 8899
rect 18827 8894 19034 9190
rect 238 8454 445 8862
rect 18827 8862 18845 8894
rect 19020 8862 19034 8894
rect 2164 8581 2234 8611
rect 2666 8581 2736 8611
rect 3168 8581 3238 8611
rect 3670 8581 3740 8611
rect 4172 8581 4242 8611
rect 4674 8581 4744 8611
rect 5176 8581 5246 8611
rect 5678 8581 5748 8611
rect 6180 8581 6250 8611
rect 6682 8581 6752 8611
rect 7184 8581 7254 8611
rect 7686 8581 7756 8611
rect 8188 8581 8258 8611
rect 8690 8581 8760 8611
rect 9192 8581 9262 8611
rect 9694 8581 9764 8611
rect 10196 8581 10266 8611
rect 10698 8581 10768 8611
rect 11200 8581 11270 8611
rect 11702 8581 11772 8611
rect 12204 8581 12274 8611
rect 12706 8581 12776 8611
rect 13208 8581 13278 8611
rect 13710 8581 13780 8611
rect 14212 8581 14282 8611
rect 14714 8581 14784 8611
rect 15216 8581 15286 8611
rect 15718 8581 15788 8611
rect 16220 8581 16290 8611
rect 16722 8581 16792 8611
rect 17224 8581 17294 8611
rect 1789 8454 1819 8524
rect 2077 8454 2107 8524
rect 2291 8454 2321 8524
rect 2579 8454 2609 8524
rect 2793 8454 2823 8524
rect 3081 8454 3111 8524
rect 3295 8454 3325 8524
rect 3583 8454 3613 8524
rect 3797 8454 3827 8524
rect 4085 8454 4115 8524
rect 4299 8454 4329 8524
rect 4587 8454 4617 8524
rect 4801 8454 4831 8524
rect 5089 8454 5119 8524
rect 5303 8454 5333 8524
rect 5591 8454 5621 8524
rect 5805 8454 5835 8524
rect 6093 8454 6123 8524
rect 6307 8454 6337 8524
rect 6595 8454 6625 8524
rect 6809 8454 6839 8524
rect 7097 8454 7127 8524
rect 7311 8454 7341 8524
rect 7599 8454 7629 8524
rect 7813 8454 7843 8524
rect 8101 8454 8131 8524
rect 8315 8454 8345 8524
rect 8603 8454 8633 8524
rect 8817 8454 8847 8524
rect 9105 8454 9135 8524
rect 9319 8454 9349 8524
rect 9607 8454 9637 8524
rect 9821 8454 9851 8524
rect 10109 8454 10139 8524
rect 10323 8454 10353 8524
rect 10611 8454 10641 8524
rect 10825 8454 10855 8524
rect 11113 8454 11143 8524
rect 11327 8454 11357 8524
rect 11615 8454 11645 8524
rect 11829 8454 11859 8524
rect 12117 8454 12147 8524
rect 12331 8454 12361 8524
rect 12619 8454 12649 8524
rect 12833 8454 12863 8524
rect 13121 8454 13151 8524
rect 13335 8454 13365 8524
rect 13623 8454 13653 8524
rect 13837 8454 13867 8524
rect 14125 8454 14155 8524
rect 14339 8454 14369 8524
rect 14627 8454 14657 8524
rect 14841 8454 14871 8524
rect 15129 8454 15159 8524
rect 15343 8454 15373 8524
rect 15631 8454 15661 8524
rect 15845 8454 15875 8524
rect 16133 8454 16163 8524
rect 16347 8454 16377 8524
rect 16635 8454 16665 8524
rect 16849 8454 16879 8524
rect 17137 8454 17167 8524
rect 17351 8454 17381 8524
rect 17639 8454 17669 8524
rect 18827 8454 19034 8862
rect 238 8422 252 8454
rect 427 8422 445 8454
rect 238 8014 445 8422
rect 18827 8422 18845 8454
rect 19020 8422 19034 8454
rect 2164 8367 2234 8397
rect 2666 8367 2736 8397
rect 3168 8367 3238 8397
rect 3670 8367 3740 8397
rect 4172 8367 4242 8397
rect 4674 8367 4744 8397
rect 5176 8367 5246 8397
rect 5678 8367 5748 8397
rect 6180 8367 6250 8397
rect 6682 8367 6752 8397
rect 7184 8367 7254 8397
rect 7686 8367 7756 8397
rect 8188 8367 8258 8397
rect 8690 8367 8760 8397
rect 9192 8367 9262 8397
rect 9694 8367 9764 8397
rect 10196 8367 10266 8397
rect 10698 8367 10768 8397
rect 11200 8367 11270 8397
rect 11702 8367 11772 8397
rect 12204 8367 12274 8397
rect 12706 8367 12776 8397
rect 13208 8367 13278 8397
rect 13710 8367 13780 8397
rect 14212 8367 14282 8397
rect 14714 8367 14784 8397
rect 15216 8367 15286 8397
rect 15718 8367 15788 8397
rect 16220 8367 16290 8397
rect 16722 8367 16792 8397
rect 17224 8367 17294 8397
rect 18827 8308 19034 8422
rect 18827 8276 18855 8308
rect 18887 8276 18899 8308
rect 18931 8276 18943 8308
rect 18975 8276 18987 8308
rect 19019 8276 19034 8308
rect 18827 8263 19034 8276
rect 18827 8231 18855 8263
rect 18887 8231 18899 8263
rect 18931 8231 18943 8263
rect 18975 8231 18987 8263
rect 19019 8231 19034 8263
rect 18827 8218 19034 8231
rect 18827 8186 18855 8218
rect 18887 8186 18899 8218
rect 18931 8186 18943 8218
rect 18975 8186 18987 8218
rect 19019 8186 19034 8218
rect 2164 8079 2234 8109
rect 2666 8079 2736 8109
rect 3168 8079 3238 8109
rect 3670 8079 3740 8109
rect 4172 8079 4242 8109
rect 4674 8079 4744 8109
rect 5176 8079 5246 8109
rect 5678 8079 5748 8109
rect 6180 8079 6250 8109
rect 6682 8079 6752 8109
rect 7184 8079 7254 8109
rect 7686 8079 7756 8109
rect 8188 8079 8258 8109
rect 8690 8079 8760 8109
rect 9192 8079 9262 8109
rect 9694 8079 9764 8109
rect 10196 8079 10266 8109
rect 10698 8079 10768 8109
rect 11200 8079 11270 8109
rect 11702 8079 11772 8109
rect 12204 8079 12274 8109
rect 12706 8079 12776 8109
rect 13208 8079 13278 8109
rect 13710 8079 13780 8109
rect 14212 8079 14282 8109
rect 14714 8079 14784 8109
rect 15216 8079 15286 8109
rect 15718 8079 15788 8109
rect 16220 8079 16290 8109
rect 16722 8079 16792 8109
rect 17224 8079 17294 8109
rect 238 7982 252 8014
rect 427 7982 445 8014
rect 238 7574 445 7982
rect 1789 7952 1819 8022
rect 2077 7952 2107 8022
rect 2291 7952 2321 8022
rect 2579 7952 2609 8022
rect 2793 7952 2823 8022
rect 3081 7952 3111 8022
rect 3295 7952 3325 8022
rect 3583 7952 3613 8022
rect 3797 7952 3827 8022
rect 4085 7952 4115 8022
rect 4299 7952 4329 8022
rect 4587 7952 4617 8022
rect 4801 7952 4831 8022
rect 5089 7952 5119 8022
rect 5303 7952 5333 8022
rect 5591 7952 5621 8022
rect 5805 7952 5835 8022
rect 6093 7952 6123 8022
rect 6307 7952 6337 8022
rect 6595 7952 6625 8022
rect 6809 7952 6839 8022
rect 7097 7952 7127 8022
rect 7311 7952 7341 8022
rect 7599 7952 7629 8022
rect 7813 7952 7843 8022
rect 8101 7952 8131 8022
rect 8315 7952 8345 8022
rect 8603 7952 8633 8022
rect 8817 7952 8847 8022
rect 9105 7952 9135 8022
rect 9319 7952 9349 8022
rect 9607 7952 9637 8022
rect 9821 7952 9851 8022
rect 10109 7952 10139 8022
rect 10323 7952 10353 8022
rect 10611 7952 10641 8022
rect 10825 7952 10855 8022
rect 11113 7952 11143 8022
rect 11327 7952 11357 8022
rect 11615 7952 11645 8022
rect 11829 7952 11859 8022
rect 12117 7952 12147 8022
rect 12331 7952 12361 8022
rect 12619 7952 12649 8022
rect 12833 7952 12863 8022
rect 13121 7952 13151 8022
rect 13335 7952 13365 8022
rect 13623 7952 13653 8022
rect 13837 7952 13867 8022
rect 14125 7952 14155 8022
rect 14339 7952 14369 8022
rect 14627 7952 14657 8022
rect 14841 7952 14871 8022
rect 15129 7952 15159 8022
rect 15343 7952 15373 8022
rect 15631 7952 15661 8022
rect 15845 7952 15875 8022
rect 16133 7952 16163 8022
rect 16347 7952 16377 8022
rect 16635 7952 16665 8022
rect 16849 7952 16879 8022
rect 17137 7952 17167 8022
rect 17351 7952 17381 8022
rect 17639 7952 17669 8022
rect 18827 8014 19034 8186
rect 18827 7982 18845 8014
rect 19020 7982 19034 8014
rect 2164 7865 2234 7895
rect 2666 7865 2736 7895
rect 3168 7865 3238 7895
rect 3670 7865 3740 7895
rect 4172 7865 4242 7895
rect 4674 7865 4744 7895
rect 5176 7865 5246 7895
rect 5678 7865 5748 7895
rect 6180 7865 6250 7895
rect 6682 7865 6752 7895
rect 7184 7865 7254 7895
rect 7686 7865 7756 7895
rect 8188 7865 8258 7895
rect 8690 7865 8760 7895
rect 9192 7865 9262 7895
rect 9694 7865 9764 7895
rect 10196 7865 10266 7895
rect 10698 7865 10768 7895
rect 11200 7865 11270 7895
rect 11702 7865 11772 7895
rect 12204 7865 12274 7895
rect 12706 7865 12776 7895
rect 13208 7865 13278 7895
rect 13710 7865 13780 7895
rect 14212 7865 14282 7895
rect 14714 7865 14784 7895
rect 15216 7865 15286 7895
rect 15718 7865 15788 7895
rect 16220 7865 16290 7895
rect 16722 7865 16792 7895
rect 17224 7865 17294 7895
rect 2164 7577 2234 7607
rect 2666 7577 2736 7607
rect 3168 7577 3238 7607
rect 3670 7577 3740 7607
rect 4172 7577 4242 7607
rect 4674 7577 4744 7607
rect 5176 7577 5246 7607
rect 5678 7577 5748 7607
rect 6180 7577 6250 7607
rect 6682 7577 6752 7607
rect 7184 7577 7254 7607
rect 7686 7577 7756 7607
rect 8188 7577 8258 7607
rect 8690 7577 8760 7607
rect 9192 7577 9262 7607
rect 9694 7577 9764 7607
rect 10196 7577 10266 7607
rect 10698 7577 10768 7607
rect 11200 7577 11270 7607
rect 11702 7577 11772 7607
rect 12204 7577 12274 7607
rect 12706 7577 12776 7607
rect 13208 7577 13278 7607
rect 13710 7577 13780 7607
rect 14212 7577 14282 7607
rect 14714 7577 14784 7607
rect 15216 7577 15286 7607
rect 15718 7577 15788 7607
rect 16220 7577 16290 7607
rect 16722 7577 16792 7607
rect 17224 7577 17294 7607
rect 238 7542 252 7574
rect 427 7542 445 7574
rect 238 7134 445 7542
rect 18827 7574 19034 7982
rect 18827 7542 18845 7574
rect 19020 7542 19034 7574
rect 1789 7450 1819 7520
rect 2077 7450 2107 7520
rect 2291 7450 2321 7520
rect 2579 7450 2609 7520
rect 2793 7450 2823 7520
rect 3081 7450 3111 7520
rect 3295 7450 3325 7520
rect 3583 7450 3613 7520
rect 3797 7450 3827 7520
rect 4085 7450 4115 7520
rect 4299 7450 4329 7520
rect 4587 7450 4617 7520
rect 4801 7450 4831 7520
rect 5089 7450 5119 7520
rect 5303 7450 5333 7520
rect 5591 7450 5621 7520
rect 5805 7450 5835 7520
rect 6093 7450 6123 7520
rect 6307 7450 6337 7520
rect 6595 7450 6625 7520
rect 6809 7450 6839 7520
rect 7097 7450 7127 7520
rect 7311 7450 7341 7520
rect 7599 7450 7629 7520
rect 7813 7450 7843 7520
rect 8101 7450 8131 7520
rect 8315 7450 8345 7520
rect 8603 7450 8633 7520
rect 8817 7450 8847 7520
rect 9105 7450 9135 7520
rect 9319 7450 9349 7520
rect 9607 7450 9637 7520
rect 9821 7450 9851 7520
rect 10109 7450 10139 7520
rect 10323 7450 10353 7520
rect 10611 7450 10641 7520
rect 10825 7450 10855 7520
rect 11113 7450 11143 7520
rect 11327 7450 11357 7520
rect 11615 7450 11645 7520
rect 11829 7450 11859 7520
rect 12117 7450 12147 7520
rect 12331 7450 12361 7520
rect 12619 7450 12649 7520
rect 12833 7450 12863 7520
rect 13121 7450 13151 7520
rect 13335 7450 13365 7520
rect 13623 7450 13653 7520
rect 13837 7450 13867 7520
rect 14125 7450 14155 7520
rect 14339 7450 14369 7520
rect 14627 7450 14657 7520
rect 14841 7450 14871 7520
rect 15129 7450 15159 7520
rect 15343 7450 15373 7520
rect 15631 7450 15661 7520
rect 15845 7450 15875 7520
rect 16133 7450 16163 7520
rect 16347 7450 16377 7520
rect 16635 7450 16665 7520
rect 16849 7450 16879 7520
rect 17137 7450 17167 7520
rect 17351 7450 17381 7520
rect 17639 7450 17669 7520
rect 2164 7363 2234 7393
rect 2666 7363 2736 7393
rect 3168 7363 3238 7393
rect 3670 7363 3740 7393
rect 4172 7363 4242 7393
rect 4674 7363 4744 7393
rect 5176 7363 5246 7393
rect 5678 7363 5748 7393
rect 6180 7363 6250 7393
rect 6682 7363 6752 7393
rect 7184 7363 7254 7393
rect 7686 7363 7756 7393
rect 8188 7363 8258 7393
rect 8690 7363 8760 7393
rect 9192 7363 9262 7393
rect 9694 7363 9764 7393
rect 10196 7363 10266 7393
rect 10698 7363 10768 7393
rect 11200 7363 11270 7393
rect 11702 7363 11772 7393
rect 12204 7363 12274 7393
rect 12706 7363 12776 7393
rect 13208 7363 13278 7393
rect 13710 7363 13780 7393
rect 14212 7363 14282 7393
rect 14714 7363 14784 7393
rect 15216 7363 15286 7393
rect 15718 7363 15788 7393
rect 16220 7363 16290 7393
rect 16722 7363 16792 7393
rect 17224 7363 17294 7393
rect 238 7102 252 7134
rect 427 7102 445 7134
rect 18827 7308 19034 7542
rect 18827 7276 18855 7308
rect 18887 7276 18899 7308
rect 18931 7276 18943 7308
rect 18975 7276 18987 7308
rect 19019 7276 19034 7308
rect 18827 7263 19034 7276
rect 18827 7231 18855 7263
rect 18887 7231 18899 7263
rect 18931 7231 18943 7263
rect 18975 7231 18987 7263
rect 19019 7231 19034 7263
rect 18827 7218 19034 7231
rect 18827 7186 18855 7218
rect 18887 7186 18899 7218
rect 18931 7186 18943 7218
rect 18975 7186 18987 7218
rect 19019 7186 19034 7218
rect 18827 7134 19034 7186
rect 238 6694 445 7102
rect 2164 7075 2234 7105
rect 2666 7075 2736 7105
rect 3168 7075 3238 7105
rect 3670 7075 3740 7105
rect 4172 7075 4242 7105
rect 4674 7075 4744 7105
rect 5176 7075 5246 7105
rect 5678 7075 5748 7105
rect 6180 7075 6250 7105
rect 6682 7075 6752 7105
rect 7184 7075 7254 7105
rect 7686 7075 7756 7105
rect 8188 7075 8258 7105
rect 8690 7075 8760 7105
rect 9192 7075 9262 7105
rect 9694 7075 9764 7105
rect 10196 7075 10266 7105
rect 10698 7075 10768 7105
rect 11200 7075 11270 7105
rect 11702 7075 11772 7105
rect 12204 7075 12274 7105
rect 12706 7075 12776 7105
rect 13208 7075 13278 7105
rect 13710 7075 13780 7105
rect 14212 7075 14282 7105
rect 14714 7075 14784 7105
rect 15216 7075 15286 7105
rect 15718 7075 15788 7105
rect 16220 7075 16290 7105
rect 16722 7075 16792 7105
rect 17224 7075 17294 7105
rect 18827 7102 18845 7134
rect 19020 7102 19034 7134
rect 1789 6948 1819 7018
rect 2077 6948 2107 7018
rect 2291 6948 2321 7018
rect 2579 6948 2609 7018
rect 2793 6948 2823 7018
rect 3081 6948 3111 7018
rect 3295 6948 3325 7018
rect 3583 6948 3613 7018
rect 3797 6948 3827 7018
rect 4085 6948 4115 7018
rect 4299 6948 4329 7018
rect 4587 6948 4617 7018
rect 4801 6948 4831 7018
rect 5089 6948 5119 7018
rect 5303 6948 5333 7018
rect 5591 6948 5621 7018
rect 5805 6948 5835 7018
rect 6093 6948 6123 7018
rect 6307 6948 6337 7018
rect 6595 6948 6625 7018
rect 6809 6948 6839 7018
rect 7097 6948 7127 7018
rect 7311 6948 7341 7018
rect 7599 6948 7629 7018
rect 7813 6948 7843 7018
rect 8101 6948 8131 7018
rect 8315 6948 8345 7018
rect 8603 6948 8633 7018
rect 8817 6948 8847 7018
rect 9105 6948 9135 7018
rect 9319 6948 9349 7018
rect 9607 6948 9637 7018
rect 9821 6948 9851 7018
rect 10109 6948 10139 7018
rect 10323 6948 10353 7018
rect 10611 6948 10641 7018
rect 10825 6948 10855 7018
rect 11113 6948 11143 7018
rect 11327 6948 11357 7018
rect 11615 6948 11645 7018
rect 11829 6948 11859 7018
rect 12117 6948 12147 7018
rect 12331 6948 12361 7018
rect 12619 6948 12649 7018
rect 12833 6948 12863 7018
rect 13121 6948 13151 7018
rect 13335 6948 13365 7018
rect 13623 6948 13653 7018
rect 13837 6948 13867 7018
rect 14125 6948 14155 7018
rect 14339 6948 14369 7018
rect 14627 6948 14657 7018
rect 14841 6948 14871 7018
rect 15129 6948 15159 7018
rect 15343 6948 15373 7018
rect 15631 6948 15661 7018
rect 15845 6948 15875 7018
rect 16133 6948 16163 7018
rect 16347 6948 16377 7018
rect 16635 6948 16665 7018
rect 16849 6948 16879 7018
rect 17137 6948 17167 7018
rect 17351 6948 17381 7018
rect 17639 6948 17669 7018
rect 2164 6861 2234 6891
rect 2666 6861 2736 6891
rect 3168 6861 3238 6891
rect 3670 6861 3740 6891
rect 4172 6861 4242 6891
rect 4674 6861 4744 6891
rect 5176 6861 5246 6891
rect 5678 6861 5748 6891
rect 6180 6861 6250 6891
rect 6682 6861 6752 6891
rect 7184 6861 7254 6891
rect 7686 6861 7756 6891
rect 8188 6861 8258 6891
rect 8690 6861 8760 6891
rect 9192 6861 9262 6891
rect 9694 6861 9764 6891
rect 10196 6861 10266 6891
rect 10698 6861 10768 6891
rect 11200 6861 11270 6891
rect 11702 6861 11772 6891
rect 12204 6861 12274 6891
rect 12706 6861 12776 6891
rect 13208 6861 13278 6891
rect 13710 6861 13780 6891
rect 14212 6861 14282 6891
rect 14714 6861 14784 6891
rect 15216 6861 15286 6891
rect 15718 6861 15788 6891
rect 16220 6861 16290 6891
rect 16722 6861 16792 6891
rect 17224 6861 17294 6891
rect 238 6662 252 6694
rect 427 6662 445 6694
rect 238 6254 445 6662
rect 2164 6573 2234 6603
rect 2666 6573 2736 6603
rect 3168 6573 3238 6603
rect 3670 6573 3740 6603
rect 4172 6573 4242 6603
rect 4674 6573 4744 6603
rect 5176 6573 5246 6603
rect 5678 6573 5748 6603
rect 6180 6573 6250 6603
rect 6682 6573 6752 6603
rect 7184 6573 7254 6603
rect 7686 6573 7756 6603
rect 8188 6573 8258 6603
rect 8690 6573 8760 6603
rect 9192 6573 9262 6603
rect 9694 6573 9764 6603
rect 10196 6573 10266 6603
rect 10698 6573 10768 6603
rect 11200 6573 11270 6603
rect 11702 6573 11772 6603
rect 12204 6573 12274 6603
rect 12706 6573 12776 6603
rect 13208 6573 13278 6603
rect 13710 6573 13780 6603
rect 14212 6573 14282 6603
rect 14714 6573 14784 6603
rect 15216 6573 15286 6603
rect 15718 6573 15788 6603
rect 16220 6573 16290 6603
rect 16722 6573 16792 6603
rect 17224 6573 17294 6603
rect 1789 6446 1819 6516
rect 2077 6446 2107 6516
rect 2291 6446 2321 6516
rect 2579 6446 2609 6516
rect 2793 6446 2823 6516
rect 3081 6446 3111 6516
rect 3295 6446 3325 6516
rect 3583 6446 3613 6516
rect 3797 6446 3827 6516
rect 4085 6446 4115 6516
rect 4299 6446 4329 6516
rect 4587 6446 4617 6516
rect 4801 6446 4831 6516
rect 5089 6446 5119 6516
rect 5303 6446 5333 6516
rect 5591 6446 5621 6516
rect 5805 6446 5835 6516
rect 6093 6446 6123 6516
rect 6307 6446 6337 6516
rect 6595 6446 6625 6516
rect 6809 6446 6839 6516
rect 7097 6446 7127 6516
rect 7311 6446 7341 6516
rect 7599 6446 7629 6516
rect 7813 6446 7843 6516
rect 8101 6446 8131 6516
rect 8315 6446 8345 6516
rect 8603 6446 8633 6516
rect 8817 6446 8847 6516
rect 9105 6446 9135 6516
rect 9319 6446 9349 6516
rect 9607 6446 9637 6516
rect 9821 6446 9851 6516
rect 10109 6446 10139 6516
rect 10323 6446 10353 6516
rect 10611 6446 10641 6516
rect 10825 6446 10855 6516
rect 11113 6446 11143 6516
rect 11327 6446 11357 6516
rect 11615 6446 11645 6516
rect 11829 6446 11859 6516
rect 12117 6446 12147 6516
rect 12331 6446 12361 6516
rect 12619 6446 12649 6516
rect 12833 6446 12863 6516
rect 13121 6446 13151 6516
rect 13335 6446 13365 6516
rect 13623 6446 13653 6516
rect 13837 6446 13867 6516
rect 14125 6446 14155 6516
rect 14339 6446 14369 6516
rect 14627 6446 14657 6516
rect 14841 6446 14871 6516
rect 15129 6446 15159 6516
rect 15343 6446 15373 6516
rect 15631 6446 15661 6516
rect 15845 6446 15875 6516
rect 16133 6446 16163 6516
rect 16347 6446 16377 6516
rect 16635 6446 16665 6516
rect 16849 6446 16879 6516
rect 17137 6446 17167 6516
rect 17351 6446 17381 6516
rect 17639 6446 17669 6516
rect 2164 6359 2234 6389
rect 2666 6359 2736 6389
rect 3168 6359 3238 6389
rect 3670 6359 3740 6389
rect 4172 6359 4242 6389
rect 4674 6359 4744 6389
rect 5176 6359 5246 6389
rect 5678 6359 5748 6389
rect 6180 6359 6250 6389
rect 6682 6359 6752 6389
rect 7184 6359 7254 6389
rect 7686 6359 7756 6389
rect 8188 6359 8258 6389
rect 8690 6359 8760 6389
rect 9192 6359 9262 6389
rect 9694 6359 9764 6389
rect 10196 6359 10266 6389
rect 10698 6359 10768 6389
rect 11200 6359 11270 6389
rect 11702 6359 11772 6389
rect 12204 6359 12274 6389
rect 12706 6359 12776 6389
rect 13208 6359 13278 6389
rect 13710 6359 13780 6389
rect 14212 6359 14282 6389
rect 14714 6359 14784 6389
rect 15216 6359 15286 6389
rect 15718 6359 15788 6389
rect 16220 6359 16290 6389
rect 16722 6359 16792 6389
rect 17224 6359 17294 6389
rect 18827 6361 19034 7102
rect 19065 9166 19272 9824
rect 21386 9403 21593 10763
rect 21346 9394 21593 9403
rect 21346 9319 21397 9394
rect 21503 9319 21593 9394
rect 21346 9312 21593 9319
rect 19065 8994 19346 9166
rect 21386 9132 21593 9312
rect 21346 9123 21593 9132
rect 21346 9048 21397 9123
rect 21503 9048 21593 9123
rect 21346 9041 21593 9048
rect 19065 8823 19272 8994
rect 21386 8854 21593 9041
rect 19065 8791 19093 8823
rect 19125 8791 19137 8823
rect 19169 8791 19181 8823
rect 19213 8791 19225 8823
rect 19257 8791 19272 8823
rect 19065 8778 19272 8791
rect 19065 8746 19093 8778
rect 19125 8746 19137 8778
rect 19169 8746 19181 8778
rect 19213 8746 19225 8778
rect 19257 8746 19272 8778
rect 21346 8845 21593 8854
rect 21346 8770 21397 8845
rect 21503 8770 21593 8845
rect 21346 8763 21593 8770
rect 19065 8733 19272 8746
rect 19065 8701 19093 8733
rect 19125 8701 19137 8733
rect 19169 8701 19181 8733
rect 19213 8701 19225 8733
rect 19257 8701 19272 8733
rect 19065 7769 19272 8701
rect 19065 7737 19093 7769
rect 19125 7737 19137 7769
rect 19169 7737 19181 7769
rect 19213 7737 19225 7769
rect 19257 7737 19272 7769
rect 19065 7724 19272 7737
rect 19065 7692 19093 7724
rect 19125 7692 19137 7724
rect 19169 7692 19181 7724
rect 19213 7692 19225 7724
rect 19257 7692 19272 7724
rect 19065 7679 19272 7692
rect 19065 7647 19093 7679
rect 19125 7647 19137 7679
rect 19169 7647 19181 7679
rect 19213 7647 19225 7679
rect 19257 7647 19272 7679
rect 19065 7166 19272 7647
rect 21386 7403 21593 8763
rect 21346 7394 21593 7403
rect 21346 7319 21397 7394
rect 21503 7319 21593 7394
rect 21346 7312 21593 7319
rect 19065 6994 19346 7166
rect 21386 7132 21593 7312
rect 21346 7123 21593 7132
rect 21346 7048 21397 7123
rect 21503 7048 21593 7123
rect 21346 7041 21593 7048
rect 19065 6818 19272 6994
rect 21386 6854 21593 7041
rect 19064 6804 19272 6818
rect 19064 6772 19092 6804
rect 19124 6772 19136 6804
rect 19168 6772 19180 6804
rect 19212 6772 19224 6804
rect 19256 6772 19272 6804
rect 19064 6759 19272 6772
rect 21346 6845 21593 6854
rect 21346 6770 21397 6845
rect 21503 6770 21593 6845
rect 21346 6763 21593 6770
rect 19064 6727 19092 6759
rect 19124 6727 19136 6759
rect 19168 6727 19180 6759
rect 19212 6727 19224 6759
rect 19256 6727 19272 6759
rect 19064 6714 19272 6727
rect 19064 6682 19092 6714
rect 19124 6682 19136 6714
rect 19168 6682 19180 6714
rect 19212 6682 19224 6714
rect 19256 6682 19272 6714
rect 19064 6678 19272 6682
rect 238 6222 252 6254
rect 427 6222 445 6254
rect 238 5814 445 6222
rect 18827 6346 19035 6361
rect 18827 6314 18856 6346
rect 18888 6314 18900 6346
rect 18932 6314 18944 6346
rect 18976 6314 18988 6346
rect 19020 6314 19035 6346
rect 18827 6301 19035 6314
rect 18827 6269 18856 6301
rect 18888 6269 18900 6301
rect 18932 6269 18944 6301
rect 18976 6269 18988 6301
rect 19020 6269 19035 6301
rect 18827 6256 19035 6269
rect 18827 6254 18856 6256
rect 18888 6254 18900 6256
rect 18932 6254 18944 6256
rect 18976 6254 18988 6256
rect 18827 6222 18845 6254
rect 19020 6222 19035 6256
rect 18827 6220 19035 6222
rect 2164 6071 2234 6101
rect 2666 6071 2736 6101
rect 3168 6071 3238 6101
rect 3670 6071 3740 6101
rect 4172 6071 4242 6101
rect 4674 6071 4744 6101
rect 5176 6071 5246 6101
rect 5678 6071 5748 6101
rect 6180 6071 6250 6101
rect 6682 6071 6752 6101
rect 7184 6071 7254 6101
rect 7686 6071 7756 6101
rect 8188 6071 8258 6101
rect 8690 6071 8760 6101
rect 9192 6071 9262 6101
rect 9694 6071 9764 6101
rect 10196 6071 10266 6101
rect 10698 6071 10768 6101
rect 11200 6071 11270 6101
rect 11702 6071 11772 6101
rect 12204 6071 12274 6101
rect 12706 6071 12776 6101
rect 13208 6071 13278 6101
rect 13710 6071 13780 6101
rect 14212 6071 14282 6101
rect 14714 6071 14784 6101
rect 15216 6071 15286 6101
rect 15718 6071 15788 6101
rect 16220 6071 16290 6101
rect 16722 6071 16792 6101
rect 17224 6071 17294 6101
rect 1789 5944 1819 6014
rect 2077 5944 2107 6014
rect 2291 5944 2321 6014
rect 2579 5944 2609 6014
rect 2793 5944 2823 6014
rect 3081 5944 3111 6014
rect 3295 5944 3325 6014
rect 3583 5944 3613 6014
rect 3797 5944 3827 6014
rect 4085 5944 4115 6014
rect 4299 5944 4329 6014
rect 4587 5944 4617 6014
rect 4801 5944 4831 6014
rect 5089 5944 5119 6014
rect 5303 5944 5333 6014
rect 5591 5944 5621 6014
rect 5805 5944 5835 6014
rect 6093 5944 6123 6014
rect 6307 5944 6337 6014
rect 6595 5944 6625 6014
rect 6809 5944 6839 6014
rect 7097 5944 7127 6014
rect 7311 5944 7341 6014
rect 7599 5944 7629 6014
rect 7813 5944 7843 6014
rect 8101 5944 8131 6014
rect 8315 5944 8345 6014
rect 8603 5944 8633 6014
rect 8817 5944 8847 6014
rect 9105 5944 9135 6014
rect 9319 5944 9349 6014
rect 9607 5944 9637 6014
rect 9821 5944 9851 6014
rect 10109 5944 10139 6014
rect 10323 5944 10353 6014
rect 10611 5944 10641 6014
rect 10825 5944 10855 6014
rect 11113 5944 11143 6014
rect 11327 5944 11357 6014
rect 11615 5944 11645 6014
rect 11829 5944 11859 6014
rect 12117 5944 12147 6014
rect 12331 5944 12361 6014
rect 12619 5944 12649 6014
rect 12833 5944 12863 6014
rect 13121 5944 13151 6014
rect 13335 5944 13365 6014
rect 13623 5944 13653 6014
rect 13837 5944 13867 6014
rect 14125 5944 14155 6014
rect 14339 5944 14369 6014
rect 14627 5944 14657 6014
rect 14841 5944 14871 6014
rect 15129 5944 15159 6014
rect 15343 5944 15373 6014
rect 15631 5944 15661 6014
rect 15845 5944 15875 6014
rect 16133 5944 16163 6014
rect 16347 5944 16377 6014
rect 16635 5944 16665 6014
rect 16849 5944 16879 6014
rect 17137 5944 17167 6014
rect 17351 5944 17381 6014
rect 17639 5944 17669 6014
rect 2164 5857 2234 5887
rect 2666 5857 2736 5887
rect 3168 5857 3238 5887
rect 3670 5857 3740 5887
rect 4172 5857 4242 5887
rect 4674 5857 4744 5887
rect 5176 5857 5246 5887
rect 5678 5857 5748 5887
rect 6180 5857 6250 5887
rect 6682 5857 6752 5887
rect 7184 5857 7254 5887
rect 7686 5857 7756 5887
rect 8188 5857 8258 5887
rect 8690 5857 8760 5887
rect 9192 5857 9262 5887
rect 9694 5857 9764 5887
rect 10196 5857 10266 5887
rect 10698 5857 10768 5887
rect 11200 5857 11270 5887
rect 11702 5857 11772 5887
rect 12204 5857 12274 5887
rect 12706 5857 12776 5887
rect 13208 5857 13278 5887
rect 13710 5857 13780 5887
rect 14212 5857 14282 5887
rect 14714 5857 14784 5887
rect 15216 5857 15286 5887
rect 15718 5857 15788 5887
rect 16220 5857 16290 5887
rect 16722 5857 16792 5887
rect 17224 5857 17294 5887
rect 238 5782 252 5814
rect 427 5782 445 5814
rect 238 5374 445 5782
rect 2164 5569 2234 5599
rect 2666 5569 2736 5599
rect 3168 5569 3238 5599
rect 3670 5569 3740 5599
rect 4172 5569 4242 5599
rect 4674 5569 4744 5599
rect 5176 5569 5246 5599
rect 5678 5569 5748 5599
rect 6180 5569 6250 5599
rect 6682 5569 6752 5599
rect 7184 5569 7254 5599
rect 7686 5569 7756 5599
rect 8188 5569 8258 5599
rect 8690 5569 8760 5599
rect 9192 5569 9262 5599
rect 9694 5569 9764 5599
rect 10196 5569 10266 5599
rect 10698 5569 10768 5599
rect 11200 5569 11270 5599
rect 11702 5569 11772 5599
rect 12204 5569 12274 5599
rect 12706 5569 12776 5599
rect 13208 5569 13278 5599
rect 13710 5569 13780 5599
rect 14212 5569 14282 5599
rect 14714 5569 14784 5599
rect 15216 5569 15286 5599
rect 15718 5569 15788 5599
rect 16220 5569 16290 5599
rect 16722 5569 16792 5599
rect 17224 5569 17294 5599
rect 1789 5442 1819 5512
rect 2077 5442 2107 5512
rect 2291 5442 2321 5512
rect 2579 5442 2609 5512
rect 2793 5442 2823 5512
rect 3081 5442 3111 5512
rect 3295 5442 3325 5512
rect 3583 5442 3613 5512
rect 3797 5442 3827 5512
rect 4085 5442 4115 5512
rect 4299 5442 4329 5512
rect 4587 5442 4617 5512
rect 4801 5442 4831 5512
rect 5089 5442 5119 5512
rect 5303 5442 5333 5512
rect 5591 5442 5621 5512
rect 5805 5442 5835 5512
rect 6093 5442 6123 5512
rect 6307 5442 6337 5512
rect 6595 5442 6625 5512
rect 6809 5442 6839 5512
rect 7097 5442 7127 5512
rect 7311 5442 7341 5512
rect 7599 5442 7629 5512
rect 7813 5442 7843 5512
rect 8101 5442 8131 5512
rect 8315 5442 8345 5512
rect 8603 5442 8633 5512
rect 8817 5442 8847 5512
rect 9105 5442 9135 5512
rect 9319 5442 9349 5512
rect 9607 5442 9637 5512
rect 9821 5442 9851 5512
rect 10109 5442 10139 5512
rect 10323 5442 10353 5512
rect 10611 5442 10641 5512
rect 10825 5442 10855 5512
rect 11113 5442 11143 5512
rect 11327 5442 11357 5512
rect 11615 5442 11645 5512
rect 11829 5442 11859 5512
rect 12117 5442 12147 5512
rect 12331 5442 12361 5512
rect 12619 5442 12649 5512
rect 12833 5442 12863 5512
rect 13121 5442 13151 5512
rect 13335 5442 13365 5512
rect 13623 5442 13653 5512
rect 13837 5442 13867 5512
rect 14125 5442 14155 5512
rect 14339 5442 14369 5512
rect 14627 5442 14657 5512
rect 14841 5442 14871 5512
rect 15129 5442 15159 5512
rect 15343 5442 15373 5512
rect 15631 5442 15661 5512
rect 15845 5442 15875 5512
rect 16133 5442 16163 5512
rect 16347 5442 16377 5512
rect 16635 5442 16665 5512
rect 16849 5442 16879 5512
rect 17137 5442 17167 5512
rect 17351 5442 17381 5512
rect 17639 5442 17669 5512
rect 238 5342 252 5374
rect 427 5342 445 5374
rect 2164 5355 2234 5385
rect 2666 5355 2736 5385
rect 3168 5355 3238 5385
rect 3670 5355 3740 5385
rect 4172 5355 4242 5385
rect 4674 5355 4744 5385
rect 5176 5355 5246 5385
rect 5678 5355 5748 5385
rect 6180 5355 6250 5385
rect 6682 5355 6752 5385
rect 7184 5355 7254 5385
rect 7686 5355 7756 5385
rect 8188 5355 8258 5385
rect 8690 5355 8760 5385
rect 9192 5355 9262 5385
rect 9694 5355 9764 5385
rect 10196 5355 10266 5385
rect 10698 5355 10768 5385
rect 11200 5355 11270 5385
rect 11702 5355 11772 5385
rect 12204 5355 12274 5385
rect 12706 5355 12776 5385
rect 13208 5355 13278 5385
rect 13710 5355 13780 5385
rect 14212 5355 14282 5385
rect 14714 5355 14784 5385
rect 15216 5355 15286 5385
rect 15718 5355 15788 5385
rect 16220 5355 16290 5385
rect 16722 5355 16792 5385
rect 17224 5355 17294 5385
rect 18827 5374 19034 6220
rect 238 4934 445 5342
rect 18827 5342 18845 5374
rect 19020 5342 19034 5374
rect 18827 5283 19034 5342
rect 18827 5251 18855 5283
rect 18887 5251 18899 5283
rect 18931 5251 18943 5283
rect 18975 5251 18987 5283
rect 19019 5251 19034 5283
rect 18827 5238 19034 5251
rect 18827 5206 18855 5238
rect 18887 5206 18899 5238
rect 18931 5206 18943 5238
rect 18975 5206 18987 5238
rect 19019 5206 19034 5238
rect 18827 5193 19034 5206
rect 18827 5161 18855 5193
rect 18887 5161 18899 5193
rect 18931 5161 18943 5193
rect 18975 5161 18987 5193
rect 19019 5161 19034 5193
rect 2164 5067 2234 5097
rect 2666 5067 2736 5097
rect 3168 5067 3238 5097
rect 3670 5067 3740 5097
rect 4172 5067 4242 5097
rect 4674 5067 4744 5097
rect 5176 5067 5246 5097
rect 5678 5067 5748 5097
rect 6180 5067 6250 5097
rect 6682 5067 6752 5097
rect 7184 5067 7254 5097
rect 7686 5067 7756 5097
rect 8188 5067 8258 5097
rect 8690 5067 8760 5097
rect 9192 5067 9262 5097
rect 9694 5067 9764 5097
rect 10196 5067 10266 5097
rect 10698 5067 10768 5097
rect 11200 5067 11270 5097
rect 11702 5067 11772 5097
rect 12204 5067 12274 5097
rect 12706 5067 12776 5097
rect 13208 5067 13278 5097
rect 13710 5067 13780 5097
rect 14212 5067 14282 5097
rect 14714 5067 14784 5097
rect 15216 5067 15286 5097
rect 15718 5067 15788 5097
rect 16220 5067 16290 5097
rect 16722 5067 16792 5097
rect 17224 5067 17294 5097
rect 1789 4940 1819 5010
rect 2077 4940 2107 5010
rect 2291 4940 2321 5010
rect 2579 4940 2609 5010
rect 2793 4940 2823 5010
rect 3081 4940 3111 5010
rect 3295 4940 3325 5010
rect 3583 4940 3613 5010
rect 3797 4940 3827 5010
rect 4085 4940 4115 5010
rect 4299 4940 4329 5010
rect 4587 4940 4617 5010
rect 4801 4940 4831 5010
rect 5089 4940 5119 5010
rect 5303 4940 5333 5010
rect 5591 4940 5621 5010
rect 5805 4940 5835 5010
rect 6093 4940 6123 5010
rect 6307 4940 6337 5010
rect 6595 4940 6625 5010
rect 6809 4940 6839 5010
rect 7097 4940 7127 5010
rect 7311 4940 7341 5010
rect 7599 4940 7629 5010
rect 7813 4940 7843 5010
rect 8101 4940 8131 5010
rect 8315 4940 8345 5010
rect 8603 4940 8633 5010
rect 8817 4940 8847 5010
rect 9105 4940 9135 5010
rect 9319 4940 9349 5010
rect 9607 4940 9637 5010
rect 9821 4940 9851 5010
rect 10109 4940 10139 5010
rect 10323 4940 10353 5010
rect 10611 4940 10641 5010
rect 10825 4940 10855 5010
rect 11113 4940 11143 5010
rect 11327 4940 11357 5010
rect 11615 4940 11645 5010
rect 11829 4940 11859 5010
rect 12117 4940 12147 5010
rect 12331 4940 12361 5010
rect 12619 4940 12649 5010
rect 12833 4940 12863 5010
rect 13121 4940 13151 5010
rect 13335 4940 13365 5010
rect 13623 4940 13653 5010
rect 13837 4940 13867 5010
rect 14125 4940 14155 5010
rect 14339 4940 14369 5010
rect 14627 4940 14657 5010
rect 14841 4940 14871 5010
rect 15129 4940 15159 5010
rect 15343 4940 15373 5010
rect 15631 4940 15661 5010
rect 15845 4940 15875 5010
rect 16133 4940 16163 5010
rect 16347 4940 16377 5010
rect 16635 4940 16665 5010
rect 16849 4940 16879 5010
rect 17137 4940 17167 5010
rect 17351 4940 17381 5010
rect 17639 4940 17669 5010
rect 238 4902 252 4934
rect 427 4902 445 4934
rect 238 4494 445 4902
rect 18827 4934 19034 5161
rect 18827 4902 18845 4934
rect 19020 4902 19034 4934
rect 2164 4853 2234 4883
rect 2666 4853 2736 4883
rect 3168 4853 3238 4883
rect 3670 4853 3740 4883
rect 4172 4853 4242 4883
rect 4674 4853 4744 4883
rect 5176 4853 5246 4883
rect 5678 4853 5748 4883
rect 6180 4853 6250 4883
rect 6682 4853 6752 4883
rect 7184 4853 7254 4883
rect 7686 4853 7756 4883
rect 8188 4853 8258 4883
rect 8690 4853 8760 4883
rect 9192 4853 9262 4883
rect 9694 4853 9764 4883
rect 10196 4853 10266 4883
rect 10698 4853 10768 4883
rect 11200 4853 11270 4883
rect 11702 4853 11772 4883
rect 12204 4853 12274 4883
rect 12706 4853 12776 4883
rect 13208 4853 13278 4883
rect 13710 4853 13780 4883
rect 14212 4853 14282 4883
rect 14714 4853 14784 4883
rect 15216 4853 15286 4883
rect 15718 4853 15788 4883
rect 16220 4853 16290 4883
rect 16722 4853 16792 4883
rect 17224 4853 17294 4883
rect 2164 4565 2234 4595
rect 2666 4565 2736 4595
rect 3168 4565 3238 4595
rect 3670 4565 3740 4595
rect 4172 4565 4242 4595
rect 4674 4565 4744 4595
rect 5176 4565 5246 4595
rect 5678 4565 5748 4595
rect 6180 4565 6250 4595
rect 6682 4565 6752 4595
rect 7184 4565 7254 4595
rect 7686 4565 7756 4595
rect 8188 4565 8258 4595
rect 8690 4565 8760 4595
rect 9192 4565 9262 4595
rect 9694 4565 9764 4595
rect 10196 4565 10266 4595
rect 10698 4565 10768 4595
rect 11200 4565 11270 4595
rect 11702 4565 11772 4595
rect 12204 4565 12274 4595
rect 12706 4565 12776 4595
rect 13208 4565 13278 4595
rect 13710 4565 13780 4595
rect 14212 4565 14282 4595
rect 14714 4565 14784 4595
rect 15216 4565 15286 4595
rect 15718 4565 15788 4595
rect 16220 4565 16290 4595
rect 16722 4565 16792 4595
rect 17224 4565 17294 4595
rect 238 4462 252 4494
rect 427 4462 445 4494
rect 238 4054 445 4462
rect 1789 4438 1819 4508
rect 2077 4438 2107 4508
rect 2291 4438 2321 4508
rect 2579 4438 2609 4508
rect 2793 4438 2823 4508
rect 3081 4438 3111 4508
rect 3295 4438 3325 4508
rect 3583 4438 3613 4508
rect 3797 4438 3827 4508
rect 4085 4438 4115 4508
rect 4299 4438 4329 4508
rect 4587 4438 4617 4508
rect 4801 4438 4831 4508
rect 5089 4438 5119 4508
rect 5303 4438 5333 4508
rect 5591 4438 5621 4508
rect 5805 4438 5835 4508
rect 6093 4438 6123 4508
rect 6307 4438 6337 4508
rect 6595 4438 6625 4508
rect 6809 4438 6839 4508
rect 7097 4438 7127 4508
rect 7311 4438 7341 4508
rect 7599 4438 7629 4508
rect 7813 4438 7843 4508
rect 8101 4438 8131 4508
rect 8315 4438 8345 4508
rect 8603 4438 8633 4508
rect 8817 4438 8847 4508
rect 9105 4438 9135 4508
rect 9319 4438 9349 4508
rect 9607 4438 9637 4508
rect 9821 4438 9851 4508
rect 10109 4438 10139 4508
rect 10323 4438 10353 4508
rect 10611 4438 10641 4508
rect 10825 4438 10855 4508
rect 11113 4438 11143 4508
rect 11327 4438 11357 4508
rect 11615 4438 11645 4508
rect 11829 4438 11859 4508
rect 12117 4438 12147 4508
rect 12331 4438 12361 4508
rect 12619 4438 12649 4508
rect 12833 4438 12863 4508
rect 13121 4438 13151 4508
rect 13335 4438 13365 4508
rect 13623 4438 13653 4508
rect 13837 4438 13867 4508
rect 14125 4438 14155 4508
rect 14339 4438 14369 4508
rect 14627 4438 14657 4508
rect 14841 4438 14871 4508
rect 15129 4438 15159 4508
rect 15343 4438 15373 4508
rect 15631 4438 15661 4508
rect 15845 4438 15875 4508
rect 16133 4438 16163 4508
rect 16347 4438 16377 4508
rect 16635 4438 16665 4508
rect 16849 4438 16879 4508
rect 17137 4438 17167 4508
rect 17351 4438 17381 4508
rect 17639 4438 17669 4508
rect 18827 4494 19034 4902
rect 18827 4462 18845 4494
rect 19020 4462 19034 4494
rect 2164 4351 2234 4381
rect 2666 4351 2736 4381
rect 3168 4351 3238 4381
rect 3670 4351 3740 4381
rect 4172 4351 4242 4381
rect 4674 4351 4744 4381
rect 5176 4351 5246 4381
rect 5678 4351 5748 4381
rect 6180 4351 6250 4381
rect 6682 4351 6752 4381
rect 7184 4351 7254 4381
rect 7686 4351 7756 4381
rect 8188 4351 8258 4381
rect 8690 4351 8760 4381
rect 9192 4351 9262 4381
rect 9694 4351 9764 4381
rect 10196 4351 10266 4381
rect 10698 4351 10768 4381
rect 11200 4351 11270 4381
rect 11702 4351 11772 4381
rect 12204 4351 12274 4381
rect 12706 4351 12776 4381
rect 13208 4351 13278 4381
rect 13710 4351 13780 4381
rect 14212 4351 14282 4381
rect 14714 4351 14784 4381
rect 15216 4351 15286 4381
rect 15718 4351 15788 4381
rect 16220 4351 16290 4381
rect 16722 4351 16792 4381
rect 17224 4351 17294 4381
rect 18827 4310 19034 4462
rect 19065 5796 19272 6678
rect 19065 5764 19093 5796
rect 19125 5764 19137 5796
rect 19169 5764 19181 5796
rect 19213 5764 19225 5796
rect 19257 5764 19272 5796
rect 19065 5751 19272 5764
rect 19065 5719 19093 5751
rect 19125 5719 19137 5751
rect 19169 5719 19181 5751
rect 19213 5719 19225 5751
rect 19257 5719 19272 5751
rect 19065 5706 19272 5719
rect 19065 5674 19093 5706
rect 19125 5674 19137 5706
rect 19169 5674 19181 5706
rect 19213 5674 19225 5706
rect 19257 5674 19272 5706
rect 19065 5166 19272 5674
rect 21386 5403 21593 6763
rect 21346 5394 21593 5403
rect 21346 5319 21397 5394
rect 21503 5319 21593 5394
rect 21346 5312 21593 5319
rect 19065 4994 19346 5166
rect 21386 5132 21593 5312
rect 21346 5123 21593 5132
rect 21346 5048 21397 5123
rect 21503 5048 21593 5123
rect 21346 5041 21593 5048
rect 19065 4795 19272 4994
rect 21386 4854 21593 5041
rect 19065 4763 19093 4795
rect 19125 4763 19137 4795
rect 19169 4763 19181 4795
rect 19213 4763 19225 4795
rect 19257 4763 19272 4795
rect 21346 4845 21593 4854
rect 21346 4770 21397 4845
rect 21503 4770 21593 4845
rect 21346 4763 21593 4770
rect 19065 4750 19272 4763
rect 19065 4718 19093 4750
rect 19125 4718 19137 4750
rect 19169 4718 19181 4750
rect 19213 4718 19225 4750
rect 19257 4718 19272 4750
rect 19065 4705 19272 4718
rect 19065 4673 19093 4705
rect 19125 4673 19137 4705
rect 19169 4673 19181 4705
rect 19213 4673 19225 4705
rect 19257 4673 19272 4705
rect 18827 4295 19035 4310
rect 18827 4263 18856 4295
rect 18888 4263 18900 4295
rect 18932 4263 18944 4295
rect 18976 4263 18988 4295
rect 19020 4263 19035 4295
rect 18827 4250 19035 4263
rect 18827 4218 18856 4250
rect 18888 4218 18900 4250
rect 18932 4218 18944 4250
rect 18976 4218 18988 4250
rect 19020 4218 19035 4250
rect 18827 4205 19035 4218
rect 18827 4173 18856 4205
rect 18888 4173 18900 4205
rect 18932 4173 18944 4205
rect 18976 4173 18988 4205
rect 19020 4173 19035 4205
rect 18827 4169 19035 4173
rect 2164 4063 2234 4093
rect 2666 4063 2736 4093
rect 3168 4063 3238 4093
rect 3670 4063 3740 4093
rect 4172 4063 4242 4093
rect 4674 4063 4744 4093
rect 5176 4063 5246 4093
rect 5678 4063 5748 4093
rect 6180 4063 6250 4093
rect 6682 4063 6752 4093
rect 7184 4063 7254 4093
rect 7686 4063 7756 4093
rect 8188 4063 8258 4093
rect 8690 4063 8760 4093
rect 9192 4063 9262 4093
rect 9694 4063 9764 4093
rect 10196 4063 10266 4093
rect 10698 4063 10768 4093
rect 11200 4063 11270 4093
rect 11702 4063 11772 4093
rect 12204 4063 12274 4093
rect 12706 4063 12776 4093
rect 13208 4063 13278 4093
rect 13710 4063 13780 4093
rect 14212 4063 14282 4093
rect 14714 4063 14784 4093
rect 15216 4063 15286 4093
rect 15718 4063 15788 4093
rect 16220 4063 16290 4093
rect 16722 4063 16792 4093
rect 17224 4063 17294 4093
rect 238 4022 252 4054
rect 427 4022 445 4054
rect 238 3614 445 4022
rect 18827 4054 19034 4169
rect 18827 4022 18845 4054
rect 19020 4022 19034 4054
rect 1789 3936 1819 4006
rect 2077 3936 2107 4006
rect 2291 3936 2321 4006
rect 2579 3936 2609 4006
rect 2793 3936 2823 4006
rect 3081 3936 3111 4006
rect 3295 3936 3325 4006
rect 3583 3936 3613 4006
rect 3797 3936 3827 4006
rect 4085 3936 4115 4006
rect 4299 3936 4329 4006
rect 4587 3936 4617 4006
rect 4801 3936 4831 4006
rect 5089 3936 5119 4006
rect 5303 3936 5333 4006
rect 5591 3936 5621 4006
rect 5805 3936 5835 4006
rect 6093 3936 6123 4006
rect 6307 3936 6337 4006
rect 6595 3936 6625 4006
rect 6809 3936 6839 4006
rect 7097 3936 7127 4006
rect 7311 3936 7341 4006
rect 7599 3936 7629 4006
rect 7813 3936 7843 4006
rect 8101 3936 8131 4006
rect 8315 3936 8345 4006
rect 8603 3936 8633 4006
rect 8817 3936 8847 4006
rect 9105 3936 9135 4006
rect 9319 3936 9349 4006
rect 9607 3936 9637 4006
rect 9821 3936 9851 4006
rect 10109 3936 10139 4006
rect 10323 3936 10353 4006
rect 10611 3936 10641 4006
rect 10825 3936 10855 4006
rect 11113 3936 11143 4006
rect 11327 3936 11357 4006
rect 11615 3936 11645 4006
rect 11829 3936 11859 4006
rect 12117 3936 12147 4006
rect 12331 3936 12361 4006
rect 12619 3936 12649 4006
rect 12833 3936 12863 4006
rect 13121 3936 13151 4006
rect 13335 3936 13365 4006
rect 13623 3936 13653 4006
rect 13837 3936 13867 4006
rect 14125 3936 14155 4006
rect 14339 3936 14369 4006
rect 14627 3936 14657 4006
rect 14841 3936 14871 4006
rect 15129 3936 15159 4006
rect 15343 3936 15373 4006
rect 15631 3936 15661 4006
rect 15845 3936 15875 4006
rect 16133 3936 16163 4006
rect 16347 3936 16377 4006
rect 16635 3936 16665 4006
rect 16849 3936 16879 4006
rect 17137 3936 17167 4006
rect 17351 3936 17381 4006
rect 17639 3936 17669 4006
rect 2164 3849 2234 3879
rect 2666 3849 2736 3879
rect 3168 3849 3238 3879
rect 3670 3849 3740 3879
rect 4172 3849 4242 3879
rect 4674 3849 4744 3879
rect 5176 3849 5246 3879
rect 5678 3849 5748 3879
rect 6180 3849 6250 3879
rect 6682 3849 6752 3879
rect 7184 3849 7254 3879
rect 7686 3849 7756 3879
rect 8188 3849 8258 3879
rect 8690 3849 8760 3879
rect 9192 3849 9262 3879
rect 9694 3849 9764 3879
rect 10196 3849 10266 3879
rect 10698 3849 10768 3879
rect 11200 3849 11270 3879
rect 11702 3849 11772 3879
rect 12204 3849 12274 3879
rect 12706 3849 12776 3879
rect 13208 3849 13278 3879
rect 13710 3849 13780 3879
rect 14212 3849 14282 3879
rect 14714 3849 14784 3879
rect 15216 3849 15286 3879
rect 15718 3849 15788 3879
rect 16220 3849 16290 3879
rect 16722 3849 16792 3879
rect 17224 3849 17294 3879
rect 238 3582 252 3614
rect 427 3582 445 3614
rect 18827 3614 19034 4022
rect 19065 3810 19272 4673
rect 19064 3796 19272 3810
rect 19064 3764 19092 3796
rect 19124 3764 19136 3796
rect 19168 3764 19180 3796
rect 19212 3764 19224 3796
rect 19256 3764 19272 3796
rect 19064 3751 19272 3764
rect 19064 3719 19092 3751
rect 19124 3719 19136 3751
rect 19168 3719 19180 3751
rect 19212 3719 19224 3751
rect 19256 3719 19272 3751
rect 19064 3706 19272 3719
rect 19064 3674 19092 3706
rect 19124 3674 19136 3706
rect 19168 3674 19180 3706
rect 19212 3674 19224 3706
rect 19256 3674 19272 3706
rect 19064 3670 19272 3674
rect 238 3174 445 3582
rect 2164 3561 2234 3591
rect 2666 3561 2736 3591
rect 3168 3561 3238 3591
rect 3670 3561 3740 3591
rect 4172 3561 4242 3591
rect 4674 3561 4744 3591
rect 5176 3561 5246 3591
rect 5678 3561 5748 3591
rect 6180 3561 6250 3591
rect 6682 3561 6752 3591
rect 7184 3561 7254 3591
rect 7686 3561 7756 3591
rect 8188 3561 8258 3591
rect 8690 3561 8760 3591
rect 9192 3561 9262 3591
rect 9694 3561 9764 3591
rect 10196 3561 10266 3591
rect 10698 3561 10768 3591
rect 11200 3561 11270 3591
rect 11702 3561 11772 3591
rect 12204 3561 12274 3591
rect 12706 3561 12776 3591
rect 13208 3561 13278 3591
rect 13710 3561 13780 3591
rect 14212 3561 14282 3591
rect 14714 3561 14784 3591
rect 15216 3561 15286 3591
rect 15718 3561 15788 3591
rect 16220 3561 16290 3591
rect 16722 3561 16792 3591
rect 17224 3561 17294 3591
rect 18827 3582 18845 3614
rect 19020 3582 19034 3614
rect 1789 3434 1819 3504
rect 2077 3434 2107 3504
rect 2291 3434 2321 3504
rect 2579 3434 2609 3504
rect 2793 3434 2823 3504
rect 3081 3434 3111 3504
rect 3295 3434 3325 3504
rect 3583 3434 3613 3504
rect 3797 3434 3827 3504
rect 4085 3434 4115 3504
rect 4299 3434 4329 3504
rect 4587 3434 4617 3504
rect 4801 3434 4831 3504
rect 5089 3434 5119 3504
rect 5303 3434 5333 3504
rect 5591 3434 5621 3504
rect 5805 3434 5835 3504
rect 6093 3434 6123 3504
rect 6307 3434 6337 3504
rect 6595 3434 6625 3504
rect 6809 3434 6839 3504
rect 7097 3434 7127 3504
rect 7311 3434 7341 3504
rect 7599 3434 7629 3504
rect 7813 3434 7843 3504
rect 8101 3434 8131 3504
rect 8315 3434 8345 3504
rect 8603 3434 8633 3504
rect 8817 3434 8847 3504
rect 9105 3434 9135 3504
rect 9319 3434 9349 3504
rect 9607 3434 9637 3504
rect 9821 3434 9851 3504
rect 10109 3434 10139 3504
rect 10323 3434 10353 3504
rect 10611 3434 10641 3504
rect 10825 3434 10855 3504
rect 11113 3434 11143 3504
rect 11327 3434 11357 3504
rect 11615 3434 11645 3504
rect 11829 3434 11859 3504
rect 12117 3434 12147 3504
rect 12331 3434 12361 3504
rect 12619 3434 12649 3504
rect 12833 3434 12863 3504
rect 13121 3434 13151 3504
rect 13335 3434 13365 3504
rect 13623 3434 13653 3504
rect 13837 3434 13867 3504
rect 14125 3434 14155 3504
rect 14339 3434 14369 3504
rect 14627 3434 14657 3504
rect 14841 3434 14871 3504
rect 15129 3434 15159 3504
rect 15343 3434 15373 3504
rect 15631 3434 15661 3504
rect 15845 3434 15875 3504
rect 16133 3434 16163 3504
rect 16347 3434 16377 3504
rect 16635 3434 16665 3504
rect 16849 3434 16879 3504
rect 17137 3434 17167 3504
rect 17351 3434 17381 3504
rect 17639 3434 17669 3504
rect 2164 3347 2234 3377
rect 2666 3347 2736 3377
rect 3168 3347 3238 3377
rect 3670 3347 3740 3377
rect 4172 3347 4242 3377
rect 4674 3347 4744 3377
rect 5176 3347 5246 3377
rect 5678 3347 5748 3377
rect 6180 3347 6250 3377
rect 6682 3347 6752 3377
rect 7184 3347 7254 3377
rect 7686 3347 7756 3377
rect 8188 3347 8258 3377
rect 8690 3347 8760 3377
rect 9192 3347 9262 3377
rect 9694 3347 9764 3377
rect 10196 3347 10266 3377
rect 10698 3347 10768 3377
rect 11200 3347 11270 3377
rect 11702 3347 11772 3377
rect 12204 3347 12274 3377
rect 12706 3347 12776 3377
rect 13208 3347 13278 3377
rect 13710 3347 13780 3377
rect 14212 3347 14282 3377
rect 14714 3347 14784 3377
rect 15216 3347 15286 3377
rect 15718 3347 15788 3377
rect 16220 3347 16290 3377
rect 16722 3347 16792 3377
rect 17224 3347 17294 3377
rect 238 3142 252 3174
rect 427 3142 445 3174
rect 238 2734 445 3142
rect 18827 3288 19034 3582
rect 18827 3273 19035 3288
rect 18827 3241 18856 3273
rect 18888 3241 18900 3273
rect 18932 3241 18944 3273
rect 18976 3241 18988 3273
rect 19020 3241 19035 3273
rect 18827 3228 19035 3241
rect 18827 3196 18856 3228
rect 18888 3196 18900 3228
rect 18932 3196 18944 3228
rect 18976 3196 18988 3228
rect 19020 3196 19035 3228
rect 18827 3183 19035 3196
rect 18827 3174 18856 3183
rect 18888 3174 18900 3183
rect 18932 3174 18944 3183
rect 18976 3174 18988 3183
rect 18827 3142 18845 3174
rect 19020 3147 19035 3183
rect 19065 3165 19272 3670
rect 21386 3403 21593 4763
rect 21346 3394 21593 3403
rect 21346 3319 21397 3394
rect 21503 3319 21593 3394
rect 21346 3312 21593 3319
rect 19020 3142 19034 3147
rect 2164 3059 2234 3089
rect 2666 3059 2736 3089
rect 3168 3059 3238 3089
rect 3670 3059 3740 3089
rect 4172 3059 4242 3089
rect 4674 3059 4744 3089
rect 5176 3059 5246 3089
rect 5678 3059 5748 3089
rect 6180 3059 6250 3089
rect 6682 3059 6752 3089
rect 7184 3059 7254 3089
rect 7686 3059 7756 3089
rect 8188 3059 8258 3089
rect 8690 3059 8760 3089
rect 9192 3059 9262 3089
rect 9694 3059 9764 3089
rect 10196 3059 10266 3089
rect 10698 3059 10768 3089
rect 11200 3059 11270 3089
rect 11702 3059 11772 3089
rect 12204 3059 12274 3089
rect 12706 3059 12776 3089
rect 13208 3059 13278 3089
rect 13710 3059 13780 3089
rect 14212 3059 14282 3089
rect 14714 3059 14784 3089
rect 15216 3059 15286 3089
rect 15718 3059 15788 3089
rect 16220 3059 16290 3089
rect 16722 3059 16792 3089
rect 17224 3059 17294 3089
rect 1789 2932 1819 3002
rect 2077 2932 2107 3002
rect 2291 2932 2321 3002
rect 2579 2932 2609 3002
rect 2793 2932 2823 3002
rect 3081 2932 3111 3002
rect 3295 2932 3325 3002
rect 3583 2932 3613 3002
rect 3797 2932 3827 3002
rect 4085 2932 4115 3002
rect 4299 2932 4329 3002
rect 4587 2932 4617 3002
rect 4801 2932 4831 3002
rect 5089 2932 5119 3002
rect 5303 2932 5333 3002
rect 5591 2932 5621 3002
rect 5805 2932 5835 3002
rect 6093 2932 6123 3002
rect 6307 2932 6337 3002
rect 6595 2932 6625 3002
rect 6809 2932 6839 3002
rect 7097 2932 7127 3002
rect 7311 2932 7341 3002
rect 7599 2932 7629 3002
rect 7813 2932 7843 3002
rect 8101 2932 8131 3002
rect 8315 2932 8345 3002
rect 8603 2932 8633 3002
rect 8817 2932 8847 3002
rect 9105 2932 9135 3002
rect 9319 2932 9349 3002
rect 9607 2932 9637 3002
rect 9821 2932 9851 3002
rect 10109 2932 10139 3002
rect 10323 2932 10353 3002
rect 10611 2932 10641 3002
rect 10825 2932 10855 3002
rect 11113 2932 11143 3002
rect 11327 2932 11357 3002
rect 11615 2932 11645 3002
rect 11829 2932 11859 3002
rect 12117 2932 12147 3002
rect 12331 2932 12361 3002
rect 12619 2932 12649 3002
rect 12833 2932 12863 3002
rect 13121 2932 13151 3002
rect 13335 2932 13365 3002
rect 13623 2932 13653 3002
rect 13837 2932 13867 3002
rect 14125 2932 14155 3002
rect 14339 2932 14369 3002
rect 14627 2932 14657 3002
rect 14841 2932 14871 3002
rect 15129 2932 15159 3002
rect 15343 2932 15373 3002
rect 15631 2932 15661 3002
rect 15845 2932 15875 3002
rect 16133 2932 16163 3002
rect 16347 2932 16377 3002
rect 16635 2932 16665 3002
rect 16849 2932 16879 3002
rect 17137 2932 17167 3002
rect 17351 2932 17381 3002
rect 17639 2932 17669 3002
rect 2164 2845 2234 2875
rect 2666 2845 2736 2875
rect 3168 2845 3238 2875
rect 3670 2845 3740 2875
rect 4172 2845 4242 2875
rect 4674 2845 4744 2875
rect 5176 2845 5246 2875
rect 5678 2845 5748 2875
rect 6180 2845 6250 2875
rect 6682 2845 6752 2875
rect 7184 2845 7254 2875
rect 7686 2845 7756 2875
rect 8188 2845 8258 2875
rect 8690 2845 8760 2875
rect 9192 2845 9262 2875
rect 9694 2845 9764 2875
rect 10196 2845 10266 2875
rect 10698 2845 10768 2875
rect 11200 2845 11270 2875
rect 11702 2845 11772 2875
rect 12204 2845 12274 2875
rect 12706 2845 12776 2875
rect 13208 2845 13278 2875
rect 13710 2845 13780 2875
rect 14212 2845 14282 2875
rect 14714 2845 14784 2875
rect 15216 2845 15286 2875
rect 15718 2845 15788 2875
rect 16220 2845 16290 2875
rect 16722 2845 16792 2875
rect 17224 2845 17294 2875
rect 238 2702 252 2734
rect 427 2702 445 2734
rect 238 2294 445 2702
rect 2164 2557 2234 2587
rect 2666 2557 2736 2587
rect 3168 2557 3238 2587
rect 3670 2557 3740 2587
rect 4172 2557 4242 2587
rect 4674 2557 4744 2587
rect 5176 2557 5246 2587
rect 5678 2557 5748 2587
rect 6180 2557 6250 2587
rect 6682 2557 6752 2587
rect 7184 2557 7254 2587
rect 7686 2557 7756 2587
rect 8188 2557 8258 2587
rect 8690 2557 8760 2587
rect 9192 2557 9262 2587
rect 9694 2557 9764 2587
rect 10196 2557 10266 2587
rect 10698 2557 10768 2587
rect 11200 2557 11270 2587
rect 11702 2557 11772 2587
rect 12204 2557 12274 2587
rect 12706 2557 12776 2587
rect 13208 2557 13278 2587
rect 13710 2557 13780 2587
rect 14212 2557 14282 2587
rect 14714 2557 14784 2587
rect 15216 2557 15286 2587
rect 15718 2557 15788 2587
rect 16220 2557 16290 2587
rect 16722 2557 16792 2587
rect 17224 2557 17294 2587
rect 1789 2430 1819 2500
rect 2077 2430 2107 2500
rect 2291 2430 2321 2500
rect 2579 2430 2609 2500
rect 2793 2430 2823 2500
rect 3081 2430 3111 2500
rect 3295 2430 3325 2500
rect 3583 2430 3613 2500
rect 3797 2430 3827 2500
rect 4085 2430 4115 2500
rect 4299 2430 4329 2500
rect 4587 2430 4617 2500
rect 4801 2430 4831 2500
rect 5089 2430 5119 2500
rect 5303 2430 5333 2500
rect 5591 2430 5621 2500
rect 5805 2430 5835 2500
rect 6093 2430 6123 2500
rect 6307 2430 6337 2500
rect 6595 2430 6625 2500
rect 6809 2430 6839 2500
rect 7097 2430 7127 2500
rect 7311 2430 7341 2500
rect 7599 2430 7629 2500
rect 7813 2430 7843 2500
rect 8101 2430 8131 2500
rect 8315 2430 8345 2500
rect 8603 2430 8633 2500
rect 8817 2430 8847 2500
rect 9105 2430 9135 2500
rect 9319 2430 9349 2500
rect 9607 2430 9637 2500
rect 9821 2430 9851 2500
rect 10109 2430 10139 2500
rect 10323 2430 10353 2500
rect 10611 2430 10641 2500
rect 10825 2430 10855 2500
rect 11113 2430 11143 2500
rect 11327 2430 11357 2500
rect 11615 2430 11645 2500
rect 11829 2430 11859 2500
rect 12117 2430 12147 2500
rect 12331 2430 12361 2500
rect 12619 2430 12649 2500
rect 12833 2430 12863 2500
rect 13121 2430 13151 2500
rect 13335 2430 13365 2500
rect 13623 2430 13653 2500
rect 13837 2430 13867 2500
rect 14125 2430 14155 2500
rect 14339 2430 14369 2500
rect 14627 2430 14657 2500
rect 14841 2430 14871 2500
rect 15129 2430 15159 2500
rect 15343 2430 15373 2500
rect 15631 2430 15661 2500
rect 15845 2430 15875 2500
rect 16133 2430 16163 2500
rect 16347 2430 16377 2500
rect 16635 2430 16665 2500
rect 16849 2430 16879 2500
rect 17137 2430 17167 2500
rect 17351 2430 17381 2500
rect 17639 2430 17669 2500
rect 2164 2343 2234 2373
rect 2666 2343 2736 2373
rect 3168 2343 3238 2373
rect 3670 2343 3740 2373
rect 4172 2343 4242 2373
rect 4674 2343 4744 2373
rect 5176 2343 5246 2373
rect 5678 2343 5748 2373
rect 6180 2343 6250 2373
rect 6682 2343 6752 2373
rect 7184 2343 7254 2373
rect 7686 2343 7756 2373
rect 8188 2343 8258 2373
rect 8690 2343 8760 2373
rect 9192 2343 9262 2373
rect 9694 2343 9764 2373
rect 10196 2343 10266 2373
rect 10698 2343 10768 2373
rect 11200 2343 11270 2373
rect 11702 2343 11772 2373
rect 12204 2343 12274 2373
rect 12706 2343 12776 2373
rect 13208 2343 13278 2373
rect 13710 2343 13780 2373
rect 14212 2343 14282 2373
rect 14714 2343 14784 2373
rect 15216 2343 15286 2373
rect 15718 2343 15788 2373
rect 16220 2343 16290 2373
rect 16722 2343 16792 2373
rect 17224 2343 17294 2373
rect 238 2262 252 2294
rect 427 2262 445 2294
rect 238 1854 445 2262
rect 18827 2294 19034 3142
rect 18827 2262 18845 2294
rect 18827 2244 18856 2262
rect 18888 2244 18900 2262
rect 18932 2244 18944 2262
rect 18976 2244 18988 2262
rect 19020 2244 19034 2294
rect 18827 2231 19034 2244
rect 18827 2199 18856 2231
rect 18888 2199 18900 2231
rect 18932 2199 18944 2231
rect 18976 2199 18988 2231
rect 19020 2199 19034 2231
rect 18827 2186 19034 2199
rect 18827 2154 18856 2186
rect 18888 2154 18900 2186
rect 18932 2154 18944 2186
rect 18976 2154 18988 2186
rect 19020 2154 19034 2186
rect 2164 2055 2234 2085
rect 2666 2055 2736 2085
rect 3168 2055 3238 2085
rect 3670 2055 3740 2085
rect 4172 2055 4242 2085
rect 4674 2055 4744 2085
rect 5176 2055 5246 2085
rect 5678 2055 5748 2085
rect 6180 2055 6250 2085
rect 6682 2055 6752 2085
rect 7184 2055 7254 2085
rect 7686 2055 7756 2085
rect 8188 2055 8258 2085
rect 8690 2055 8760 2085
rect 9192 2055 9262 2085
rect 9694 2055 9764 2085
rect 10196 2055 10266 2085
rect 10698 2055 10768 2085
rect 11200 2055 11270 2085
rect 11702 2055 11772 2085
rect 12204 2055 12274 2085
rect 12706 2055 12776 2085
rect 13208 2055 13278 2085
rect 13710 2055 13780 2085
rect 14212 2055 14282 2085
rect 14714 2055 14784 2085
rect 15216 2055 15286 2085
rect 15718 2055 15788 2085
rect 16220 2055 16290 2085
rect 16722 2055 16792 2085
rect 17224 2055 17294 2085
rect 1789 1928 1819 1998
rect 2077 1928 2107 1998
rect 2291 1928 2321 1998
rect 2579 1928 2609 1998
rect 2793 1928 2823 1998
rect 3081 1928 3111 1998
rect 3295 1928 3325 1998
rect 3583 1928 3613 1998
rect 3797 1928 3827 1998
rect 4085 1928 4115 1998
rect 4299 1928 4329 1998
rect 4587 1928 4617 1998
rect 4801 1928 4831 1998
rect 5089 1928 5119 1998
rect 5303 1928 5333 1998
rect 5591 1928 5621 1998
rect 5805 1928 5835 1998
rect 6093 1928 6123 1998
rect 6307 1928 6337 1998
rect 6595 1928 6625 1998
rect 6809 1928 6839 1998
rect 7097 1928 7127 1998
rect 7311 1928 7341 1998
rect 7599 1928 7629 1998
rect 7813 1928 7843 1998
rect 8101 1928 8131 1998
rect 8315 1928 8345 1998
rect 8603 1928 8633 1998
rect 8817 1928 8847 1998
rect 9105 1928 9135 1998
rect 9319 1928 9349 1998
rect 9607 1928 9637 1998
rect 9821 1928 9851 1998
rect 10109 1928 10139 1998
rect 10323 1928 10353 1998
rect 10611 1928 10641 1998
rect 10825 1928 10855 1998
rect 11113 1928 11143 1998
rect 11327 1928 11357 1998
rect 11615 1928 11645 1998
rect 11829 1928 11859 1998
rect 12117 1928 12147 1998
rect 12331 1928 12361 1998
rect 12619 1928 12649 1998
rect 12833 1928 12863 1998
rect 13121 1928 13151 1998
rect 13335 1928 13365 1998
rect 13623 1928 13653 1998
rect 13837 1928 13867 1998
rect 14125 1928 14155 1998
rect 14339 1928 14369 1998
rect 14627 1928 14657 1998
rect 14841 1928 14871 1998
rect 15129 1928 15159 1998
rect 15343 1928 15373 1998
rect 15631 1928 15661 1998
rect 15845 1928 15875 1998
rect 16133 1928 16163 1998
rect 16347 1928 16377 1998
rect 16635 1928 16665 1998
rect 16849 1928 16879 1998
rect 17137 1928 17167 1998
rect 17351 1928 17381 1998
rect 17639 1928 17669 1998
rect 238 1822 252 1854
rect 427 1822 445 1854
rect 2164 1841 2234 1871
rect 2666 1841 2736 1871
rect 3168 1841 3238 1871
rect 3670 1841 3740 1871
rect 4172 1841 4242 1871
rect 4674 1841 4744 1871
rect 5176 1841 5246 1871
rect 5678 1841 5748 1871
rect 6180 1841 6250 1871
rect 6682 1841 6752 1871
rect 7184 1841 7254 1871
rect 7686 1841 7756 1871
rect 8188 1841 8258 1871
rect 8690 1841 8760 1871
rect 9192 1841 9262 1871
rect 9694 1841 9764 1871
rect 10196 1841 10266 1871
rect 10698 1841 10768 1871
rect 11200 1841 11270 1871
rect 11702 1841 11772 1871
rect 12204 1841 12274 1871
rect 12706 1841 12776 1871
rect 13208 1841 13278 1871
rect 13710 1841 13780 1871
rect 14212 1841 14282 1871
rect 14714 1841 14784 1871
rect 15216 1841 15286 1871
rect 15718 1841 15788 1871
rect 16220 1841 16290 1871
rect 16722 1841 16792 1871
rect 17224 1841 17294 1871
rect 18827 1854 19034 2154
rect 238 1414 445 1822
rect 18827 1822 18845 1854
rect 19020 1822 19034 1854
rect 2164 1553 2234 1583
rect 2666 1553 2736 1583
rect 3168 1553 3238 1583
rect 3670 1553 3740 1583
rect 4172 1553 4242 1583
rect 4674 1553 4744 1583
rect 5176 1553 5246 1583
rect 5678 1553 5748 1583
rect 6180 1553 6250 1583
rect 6682 1553 6752 1583
rect 7184 1553 7254 1583
rect 7686 1553 7756 1583
rect 8188 1553 8258 1583
rect 8690 1553 8760 1583
rect 9192 1553 9262 1583
rect 9694 1553 9764 1583
rect 10196 1553 10266 1583
rect 10698 1553 10768 1583
rect 11200 1553 11270 1583
rect 11702 1553 11772 1583
rect 12204 1553 12274 1583
rect 12706 1553 12776 1583
rect 13208 1553 13278 1583
rect 13710 1553 13780 1583
rect 14212 1553 14282 1583
rect 14714 1553 14784 1583
rect 15216 1553 15286 1583
rect 15718 1553 15788 1583
rect 16220 1553 16290 1583
rect 16722 1553 16792 1583
rect 17224 1553 17294 1583
rect 1789 1426 1819 1496
rect 2077 1426 2107 1496
rect 2291 1426 2321 1496
rect 2579 1426 2609 1496
rect 2793 1426 2823 1496
rect 3081 1426 3111 1496
rect 3295 1426 3325 1496
rect 3583 1426 3613 1496
rect 3797 1426 3827 1496
rect 4085 1426 4115 1496
rect 4299 1426 4329 1496
rect 4587 1426 4617 1496
rect 4801 1426 4831 1496
rect 5089 1426 5119 1496
rect 5303 1426 5333 1496
rect 5591 1426 5621 1496
rect 5805 1426 5835 1496
rect 6093 1426 6123 1496
rect 6307 1426 6337 1496
rect 6595 1426 6625 1496
rect 6809 1426 6839 1496
rect 7097 1426 7127 1496
rect 7311 1426 7341 1496
rect 7599 1426 7629 1496
rect 7813 1426 7843 1496
rect 8101 1426 8131 1496
rect 8315 1426 8345 1496
rect 8603 1426 8633 1496
rect 8817 1426 8847 1496
rect 9105 1426 9135 1496
rect 9319 1426 9349 1496
rect 9607 1426 9637 1496
rect 9821 1426 9851 1496
rect 10109 1426 10139 1496
rect 10323 1426 10353 1496
rect 10611 1426 10641 1496
rect 10825 1426 10855 1496
rect 11113 1426 11143 1496
rect 11327 1426 11357 1496
rect 11615 1426 11645 1496
rect 11829 1426 11859 1496
rect 12117 1426 12147 1496
rect 12331 1426 12361 1496
rect 12619 1426 12649 1496
rect 12833 1426 12863 1496
rect 13121 1426 13151 1496
rect 13335 1426 13365 1496
rect 13623 1426 13653 1496
rect 13837 1426 13867 1496
rect 14125 1426 14155 1496
rect 14339 1426 14369 1496
rect 14627 1426 14657 1496
rect 14841 1426 14871 1496
rect 15129 1426 15159 1496
rect 15343 1426 15373 1496
rect 15631 1426 15661 1496
rect 15845 1426 15875 1496
rect 16133 1426 16163 1496
rect 16347 1426 16377 1496
rect 16635 1426 16665 1496
rect 16849 1426 16879 1496
rect 17137 1426 17167 1496
rect 17351 1426 17381 1496
rect 17639 1426 17669 1496
rect 238 1382 252 1414
rect 427 1382 445 1414
rect 238 974 445 1382
rect 18827 1414 19034 1822
rect 18827 1382 18845 1414
rect 19020 1382 19034 1414
rect 2164 1339 2234 1369
rect 2666 1339 2736 1369
rect 3168 1339 3238 1369
rect 3670 1339 3740 1369
rect 4172 1339 4242 1369
rect 4674 1339 4744 1369
rect 5176 1339 5246 1369
rect 5678 1339 5748 1369
rect 6180 1339 6250 1369
rect 6682 1339 6752 1369
rect 7184 1339 7254 1369
rect 7686 1339 7756 1369
rect 8188 1339 8258 1369
rect 8690 1339 8760 1369
rect 9192 1339 9262 1369
rect 9694 1339 9764 1369
rect 10196 1339 10266 1369
rect 10698 1339 10768 1369
rect 11200 1339 11270 1369
rect 11702 1339 11772 1369
rect 12204 1339 12274 1369
rect 12706 1339 12776 1369
rect 13208 1339 13278 1369
rect 13710 1339 13780 1369
rect 14212 1339 14282 1369
rect 14714 1339 14784 1369
rect 15216 1339 15286 1369
rect 15718 1339 15788 1369
rect 16220 1339 16290 1369
rect 16722 1339 16792 1369
rect 17224 1339 17294 1369
rect 18827 1291 19034 1382
rect 18826 1276 19034 1291
rect 18826 1244 18854 1276
rect 18886 1244 18898 1276
rect 18930 1244 18942 1276
rect 18974 1244 18986 1276
rect 19018 1244 19034 1276
rect 18826 1231 19034 1244
rect 18826 1199 18854 1231
rect 18886 1199 18898 1231
rect 18930 1199 18942 1231
rect 18974 1199 18986 1231
rect 19018 1199 19034 1231
rect 18826 1186 19034 1199
rect 18826 1154 18854 1186
rect 18886 1154 18898 1186
rect 18930 1154 18942 1186
rect 18974 1154 18986 1186
rect 19018 1154 19034 1186
rect 18826 1150 19034 1154
rect 2164 1051 2234 1081
rect 2666 1051 2736 1081
rect 3168 1051 3238 1081
rect 3670 1051 3740 1081
rect 4172 1051 4242 1081
rect 4674 1051 4744 1081
rect 5176 1051 5246 1081
rect 5678 1051 5748 1081
rect 6180 1051 6250 1081
rect 6682 1051 6752 1081
rect 7184 1051 7254 1081
rect 7686 1051 7756 1081
rect 8188 1051 8258 1081
rect 8690 1051 8760 1081
rect 9192 1051 9262 1081
rect 9694 1051 9764 1081
rect 10196 1051 10266 1081
rect 10698 1051 10768 1081
rect 11200 1051 11270 1081
rect 11702 1051 11772 1081
rect 12204 1051 12274 1081
rect 12706 1051 12776 1081
rect 13208 1051 13278 1081
rect 13710 1051 13780 1081
rect 14212 1051 14282 1081
rect 14714 1051 14784 1081
rect 15216 1051 15286 1081
rect 15718 1051 15788 1081
rect 16220 1051 16290 1081
rect 16722 1051 16792 1081
rect 17224 1051 17294 1081
rect 238 942 252 974
rect 427 942 445 974
rect 238 534 445 942
rect 5805 924 5835 994
rect 6093 924 6123 994
rect 7957 924 7987 994
rect 9821 924 9851 994
rect 9965 924 9995 994
rect 13837 924 13867 994
rect 15487 924 15517 994
rect 17495 924 17525 994
rect 18827 974 19034 1150
rect 18827 942 18845 974
rect 19020 942 19034 974
rect 5713 837 5748 867
rect 6180 837 6215 867
rect 238 502 252 534
rect 427 502 445 534
rect 238 366 445 502
rect 18827 534 19034 942
rect 18827 502 18845 534
rect 19020 502 19034 534
rect 238 334 253 366
rect 285 334 297 366
rect 329 334 341 366
rect 373 334 385 366
rect 417 334 445 366
rect 238 321 445 334
rect 238 289 253 321
rect 285 289 297 321
rect 329 289 341 321
rect 373 289 385 321
rect 417 289 445 321
rect 238 276 445 289
rect 238 244 253 276
rect 285 244 297 276
rect 329 244 341 276
rect 373 244 385 276
rect 417 244 445 276
rect 238 21 445 244
rect 17495 1 17525 457
rect 18827 431 19034 502
rect 18827 399 18855 431
rect 18887 399 18899 431
rect 18931 399 18943 431
rect 18975 399 18987 431
rect 19019 399 19034 431
rect 18827 386 19034 399
rect 18827 354 18855 386
rect 18887 354 18899 386
rect 18931 354 18943 386
rect 18975 354 18987 386
rect 19019 354 19034 386
rect 18827 341 19034 354
rect 18827 309 18855 341
rect 18887 309 18899 341
rect 18931 309 18943 341
rect 18975 309 18987 341
rect 19019 309 19034 341
rect 18827 86 19034 309
rect 19065 2993 19346 3165
rect 21386 3132 21593 3312
rect 21346 3123 21593 3132
rect 21346 3048 21397 3123
rect 21503 3048 21593 3123
rect 21346 3041 21593 3048
rect 19065 2762 19272 2993
rect 21386 2854 21593 3041
rect 21346 2845 21593 2854
rect 21346 2770 21397 2845
rect 21503 2770 21593 2845
rect 21346 2763 21593 2770
rect 19065 2730 19093 2762
rect 19125 2730 19137 2762
rect 19169 2730 19181 2762
rect 19213 2730 19225 2762
rect 19257 2730 19272 2762
rect 19065 2717 19272 2730
rect 19065 2685 19093 2717
rect 19125 2685 19137 2717
rect 19169 2685 19181 2717
rect 19213 2685 19225 2717
rect 19257 2685 19272 2717
rect 19065 2672 19272 2685
rect 19065 2640 19093 2672
rect 19125 2640 19137 2672
rect 19169 2640 19181 2672
rect 19213 2640 19225 2672
rect 19257 2640 19272 2672
rect 19065 1760 19272 2640
rect 19065 1728 19093 1760
rect 19125 1728 19137 1760
rect 19169 1728 19181 1760
rect 19213 1728 19225 1760
rect 19257 1728 19272 1760
rect 19065 1715 19272 1728
rect 19065 1683 19093 1715
rect 19125 1683 19137 1715
rect 19169 1683 19181 1715
rect 19213 1683 19225 1715
rect 19257 1683 19272 1715
rect 19065 1670 19272 1683
rect 19065 1638 19093 1670
rect 19125 1638 19137 1670
rect 19169 1638 19181 1670
rect 19213 1638 19225 1670
rect 19257 1638 19272 1670
rect 19065 1168 19272 1638
rect 21386 1403 21593 2763
rect 21346 1394 21593 1403
rect 21346 1319 21397 1394
rect 21503 1319 21593 1394
rect 21346 1312 21593 1319
rect 19065 996 19346 1168
rect 21386 1132 21593 1312
rect 21346 1123 21593 1132
rect 21346 1048 21397 1123
rect 21503 1048 21593 1123
rect 21346 1041 21593 1048
rect 19065 763 19272 996
rect 21386 854 21593 1041
rect 21346 845 21593 854
rect 21346 770 21397 845
rect 21503 770 21593 845
rect 21346 763 21593 770
rect 19065 731 19093 763
rect 19125 731 19137 763
rect 19169 731 19181 763
rect 19213 731 19225 763
rect 19257 731 19272 763
rect 19065 718 19272 731
rect 19065 686 19093 718
rect 19125 686 19137 718
rect 19169 686 19181 718
rect 19213 686 19225 718
rect 19257 686 19272 718
rect 19065 673 19272 686
rect 19065 641 19093 673
rect 19125 641 19137 673
rect 19169 641 19181 673
rect 19213 641 19225 673
rect 19257 641 19272 673
rect 19065 212 19272 641
rect 19065 180 19093 212
rect 19125 180 19137 212
rect 19169 180 19181 212
rect 19213 180 19225 212
rect 19257 180 19272 212
rect 19065 167 19272 180
rect 19065 135 19093 167
rect 19125 135 19137 167
rect 19169 135 19181 167
rect 19213 135 19225 167
rect 19257 135 19272 167
rect 19065 122 19272 135
rect 19065 90 19093 122
rect 19125 90 19137 122
rect 19169 90 19181 122
rect 19213 90 19225 122
rect 19257 90 19272 122
rect 19065 86 19272 90
rect 21386 83 21593 763
rect 21630 11828 21837 12084
rect 21630 11747 21637 11828
rect 21756 11747 21837 11828
rect 21630 11625 21837 11747
rect 21630 11419 21643 11625
rect 21749 11419 21837 11625
rect 21630 10746 21837 11419
rect 21630 10540 21643 10746
rect 21749 10540 21837 10746
rect 21630 10273 21837 10540
rect 21630 10192 21637 10273
rect 21756 10192 21837 10273
rect 21630 9828 21837 10192
rect 21630 9747 21637 9828
rect 21756 9747 21837 9828
rect 21630 9625 21837 9747
rect 21630 9419 21643 9625
rect 21749 9419 21837 9625
rect 21630 8746 21837 9419
rect 21630 8540 21643 8746
rect 21749 8540 21837 8746
rect 21630 8273 21837 8540
rect 21630 8192 21637 8273
rect 21756 8192 21837 8273
rect 21630 7828 21837 8192
rect 21630 7747 21637 7828
rect 21756 7747 21837 7828
rect 21630 7625 21837 7747
rect 21630 7419 21643 7625
rect 21749 7419 21837 7625
rect 21630 6746 21837 7419
rect 21630 6540 21643 6746
rect 21749 6540 21837 6746
rect 21630 6273 21837 6540
rect 21630 6192 21637 6273
rect 21756 6192 21837 6273
rect 21630 5828 21837 6192
rect 21630 5747 21637 5828
rect 21756 5747 21837 5828
rect 21630 5625 21837 5747
rect 21630 5419 21643 5625
rect 21749 5419 21837 5625
rect 21630 4746 21837 5419
rect 21630 4540 21643 4746
rect 21749 4540 21837 4746
rect 21630 4273 21837 4540
rect 21630 4192 21637 4273
rect 21756 4192 21837 4273
rect 21630 3828 21837 4192
rect 21630 3747 21637 3828
rect 21756 3747 21837 3828
rect 21630 3625 21837 3747
rect 21630 3419 21643 3625
rect 21749 3419 21837 3625
rect 21630 2746 21837 3419
rect 21630 2540 21643 2746
rect 21749 2540 21837 2746
rect 21630 2273 21837 2540
rect 21630 2192 21637 2273
rect 21756 2192 21837 2273
rect 21630 1828 21837 2192
rect 21630 1747 21637 1828
rect 21756 1747 21837 1828
rect 21630 1625 21837 1747
rect 21630 1419 21643 1625
rect 21749 1419 21837 1625
rect 21630 746 21837 1419
rect 21630 540 21643 746
rect 21749 540 21837 746
rect 21630 273 21837 540
rect 21630 192 21637 273
rect 21756 192 21837 273
rect 21630 84 21837 192
use adc_array_wafflecap_8_1  adc_array_wafflecap_8_1_0 ../adc_array_cap
timestamp 1662987872
transform 1 0 13745 0 1 457
box 0 0 502 502
use adc_array_wafflecap_8_2  adc_array_wafflecap_8_2_0 ../adc_array_cap
timestamp 1662983799
transform 1 0 9729 0 1 457
box 0 0 502 502
use adc_array_wafflecap_8_4  adc_array_wafflecap_8_4_0 ../adc_array_cap
timestamp 1662985026
transform 1 0 5713 0 1 457
box 0 0 502 502
use adc_array_wafflecap_8_8  adc_array_wafflecap_8_8_0 ../adc_array_cap
array 0 31 502 0 15 502
timestamp 1662984960
transform 1 0 1697 0 1 959
box 0 0 502 502
use adc_array_wafflecap_8_Drv  adc_array_wafflecap_8_Drv_0 ../adc_array_cap
array 0 0 502 0 15 502
timestamp 1663932020
transform 1 0 1195 0 1 959
box 0 0 502 502
use adc_array_wafflecap_8_Dummy  adc_array_wafflecap_8_Dummy_0 ../adc_array_cap
array 0 8 502 0 0 502
timestamp 1663073688
transform 1 0 1195 0 1 457
box 0 0 502 502
use adc_array_wafflecap_8_Dummy  adc_array_wafflecap_8_Dummy_1
array 0 6 502 0 0 502
timestamp 1663073688
transform 1 0 6215 0 1 457
box 0 0 502 502
use adc_array_wafflecap_8_Dummy  adc_array_wafflecap_8_Dummy_2
array 0 6 502 0 0 502
timestamp 1663073688
transform 1 0 10231 0 1 457
box 0 0 502 502
use adc_array_wafflecap_8_Dummy  adc_array_wafflecap_8_Dummy_3
array 0 5 502 0 0 502
timestamp 1663073688
transform 1 0 14247 0 1 457
box 0 0 502 502
use adc_array_wafflecap_8_Dummy  adc_array_wafflecap_8_Dummy_4
array 0 33 502 0 0 502
timestamp 1663073688
transform 1 0 1195 0 1 8991
box 0 0 502 502
use adc_array_wafflecap_8_Dummy  adc_array_wafflecap_8_Dummy_5
array 0 0 502 0 15 502
timestamp 1663073688
transform 1 0 17761 0 1 959
box 0 0 502 502
use adc_array_wafflecap_8_Dummy  adc_array_wafflecap_8_Dummy_6
timestamp 1663073688
transform 1 0 17761 0 1 457
box 0 0 502 502
use adc_array_wafflecap_8_Gate  adc_array_wafflecap_8_Gate_0 ../adc_array_cap
timestamp 1663061126
transform 1 0 17259 0 1 457
box 0 0 502 502
use adc_noise_decoup_cell1  adc_noise_decoup_cell1_0 ../adc_noise_decoup_cell
array 0 0 2000 0 5 2000
timestamp 1663849571
transform 1 0 19346 0 1 83
box 0 0 2000 2000
use adc_noise_decoup_cell1  adc_noise_decoup_cell1_1
array 0 8 2000 0 0 2000
timestamp 1663849571
transform 1 0 1346 0 1 10083
box 0 0 2000 2000
<< labels >>
flabel locali s 536 0 570 21 5 FreeSans 40 0 0 0 sample_n
port 7 s signal input
flabel locali s 590 0 624 21 5 FreeSans 40 0 0 0 sample
port 6 s signal input
flabel locali s 644 0 712 21 5 FreeSans 40 0 0 0 vcm
port 3 s analog input
flabel locali s 755 0 901 21 5 FreeSans 40 0 0 0 VDD
port 1 s power bidirectional
flabel locali s 944 0 1090 21 5 FreeSans 40 0 0 0 VSS
port 2 s power bidirectional
flabel locali s 2124 0 2141 21 5 FreeSans 80 0 0 0 row_n[0]
port 70 s signal input
flabel locali s 2626 0 2643 21 5 FreeSans 80 0 0 0 row_n[1]
port 71 s signal input
flabel locali s 3128 0 3145 21 5 FreeSans 80 0 0 0 row_n[2]
port 72 s signal input
flabel locali s 3630 0 3647 21 5 FreeSans 80 0 0 0 row_n[3]
port 73 s signal input
flabel locali s 4132 0 4149 21 5 FreeSans 80 0 0 0 row_n[4]
port 74 s signal input
flabel locali s 4634 0 4651 21 5 FreeSans 80 0 0 0 row_n[5]
port 75 s signal input
flabel locali s 5136 0 5153 21 5 FreeSans 80 0 0 0 row_n[6]
port 76 s signal input
flabel locali s 5638 0 5655 21 5 FreeSans 80 0 0 0 row_n[7]
port 77 s signal input
flabel locali s 6140 0 6157 21 5 FreeSans 80 0 0 0 row_n[8]
port 78 s signal input
flabel locali s 6642 0 6659 21 5 FreeSans 80 0 0 0 row_n[9]
port 79 s signal input
flabel locali s 7144 0 7161 21 5 FreeSans 80 0 0 0 row_n[10]
port 80 s signal input
flabel locali s 7646 0 7663 21 5 FreeSans 80 0 0 0 row_n[11]
port 81 s signal input
flabel locali s 8148 0 8165 21 5 FreeSans 80 0 0 0 row_n[12]
port 82 s signal input
flabel locali s 8650 0 8667 21 5 FreeSans 80 0 0 0 row_n[13]
port 83 s signal input
flabel locali s 9152 0 9169 21 5 FreeSans 80 0 0 0 row_n[14]
port 84 s signal input
flabel locali s 9654 0 9671 21 5 FreeSans 80 0 0 0 row_n[15]
port 85 s signal input
flabel locali s 10156 0 10173 21 5 FreeSans 80 0 0 0 row_n[16]
port 86 s signal input
flabel locali s 10658 0 10675 21 5 FreeSans 80 0 0 0 row_n[17]
port 87 s signal input
flabel locali s 11160 0 11177 21 5 FreeSans 80 0 0 0 row_n[18]
port 88 s signal input
flabel locali s 11662 0 11679 21 5 FreeSans 80 0 0 0 row_n[19]
port 89 s signal input
flabel locali s 12164 0 12181 21 5 FreeSans 80 0 0 0 row_n[20]
port 90 s signal input
flabel locali s 12666 0 12683 21 5 FreeSans 80 0 0 0 row_n[21]
port 91 s signal input
flabel locali s 13168 0 13185 21 5 FreeSans 80 0 0 0 row_n[22]
port 92 s signal input
flabel locali s 13670 0 13687 21 5 FreeSans 80 0 0 0 row_n[23]
port 93 s signal input
flabel locali s 14172 0 14189 21 5 FreeSans 80 0 0 0 row_n[24]
port 94 s signal input
flabel locali s 5974 0 5991 21 5 FreeSans 80 0 0 0 en_n_bit[2]
port 102 s signal input
flabel locali s 9990 0 10007 21 5 FreeSans 80 0 0 0 en_n_bit[1]
port 103 s signal input
flabel locali s 14006 0 14023 21 5 FreeSans 80 0 0 0 en_n_bit[0]
port 104 s signal input
flabel locali s 14274 0 14291 21 5 FreeSans 80 0 0 0 row_n[25]
port 95 s signal input
flabel locali s 14376 0 14393 21 5 FreeSans 80 0 0 0 row_n[26]
port 96 s signal input
flabel locali s 14478 0 14495 21 5 FreeSans 80 0 0 0 row_n[27]
port 97 s signal input
flabel locali s 14580 0 14597 21 5 FreeSans 80 0 0 0 row_n[28]
port 98 s signal input
flabel locali s 14682 0 14699 21 5 FreeSans 80 0 0 0 row_n[29]
port 99 s signal input
flabel locali s 14784 0 14801 21 5 FreeSans 80 0 0 0 row_n[30]
port 100 s signal input
flabel locali s 14886 0 14903 21 5 FreeSans 80 0 0 0 row_n[31]
port 101 s signal input
flabel locali s 17238 1 17255 22 5 FreeSans 80 90 0 0 sw_n
port 9 s signal input
flabel locali s 17299 1 17316 22 5 FreeSans 80 90 0 0 sw
port 8 s signal input
flabel metal4 s 17495 1 17525 30 5 FreeSans 80 0 0 0 ctop
port 4 s analog output
flabel metal1 s 19297 4 19391 28 0 FreeSans 80 0 0 0 analog_in
port 5 nsew analog input
flabel metal1 s 522 1174 575 1188 7 FreeSans 80 0 0 0 col_n[0]
port 123 w signal input
flabel metal1 s 522 1676 575 1690 7 FreeSans 80 0 0 0 col_n[1]
port 124 w signal input
flabel metal1 s 522 2178 575 2192 7 FreeSans 80 0 0 0 col_n[2]
port 125 w signal input
flabel metal1 s 522 2680 575 2694 7 FreeSans 80 0 0 0 col_n[3]
port 126 w signal input
flabel metal1 s 522 3182 575 3196 7 FreeSans 80 0 0 0 col_n[4]
port 127 w signal input
flabel metal1 s 522 3684 575 3698 7 FreeSans 80 0 0 0 col_n[5]
port 128 w signal input
flabel metal1 s 522 4186 575 4200 7 FreeSans 80 0 0 0 col_n[6]
port 129 w signal input
flabel metal1 s 522 4688 575 4702 7 FreeSans 80 0 0 0 col_n[7]
port 130 w signal input
flabel metal1 s 522 5190 575 5204 7 FreeSans 80 0 0 0 col_n[8]
port 131 w signal input
flabel metal1 s 522 5692 575 5706 7 FreeSans 80 0 0 0 col_n[9]
port 132 w signal input
flabel metal1 s 522 6194 575 6208 7 FreeSans 80 0 0 0 col_n[10]
port 133 w signal input
flabel metal1 s 522 6696 575 6710 7 FreeSans 80 0 0 0 col_n[11]
port 134 w signal input
flabel metal1 s 522 7198 575 7212 7 FreeSans 80 0 0 0 col_n[12]
port 135 w signal input
flabel metal1 s 522 7700 575 7714 7 FreeSans 80 0 0 0 col_n[13]
port 136 w signal input
flabel metal1 s 522 8202 575 8216 7 FreeSans 80 0 0 0 col_n[14]
port 137 w signal input
flabel metal1 s 522 8704 575 8718 7 FreeSans 80 0 0 0 col_n[15]
port 138 w signal input
flabel metal1 s 522 1215 575 1229 7 FreeSans 80 0 0 0 colon_n[0]
port 139 w signal input
flabel metal1 s 522 1717 575 1731 7 FreeSans 80 0 0 0 colon_n[1]
port 140 w signal input
flabel metal1 s 522 2219 575 2233 7 FreeSans 80 0 0 0 colon_n[2]
port 141 w signal input
flabel metal1 s 522 2721 575 2735 7 FreeSans 80 0 0 0 colon_n[3]
port 142 w signal input
flabel metal1 s 521 3223 574 3237 7 FreeSans 80 0 0 0 colon_n[4]
port 143 w signal input
flabel metal1 s 522 3725 575 3739 7 FreeSans 80 0 0 0 colon_n[5]
port 144 w signal input
flabel metal1 s 522 4227 575 4241 7 FreeSans 80 0 0 0 colon_n[6]
port 145 w signal input
flabel metal1 s 522 4729 575 4743 7 FreeSans 80 0 0 0 colon_n[7]
port 146 w signal input
flabel metal1 s 522 5231 575 5245 7 FreeSans 80 0 0 0 colon_n[8]
port 147 w signal input
flabel metal1 s 522 5733 575 5747 7 FreeSans 80 0 0 0 colon_n[9]
port 148 w signal input
flabel metal1 s 522 6235 575 6249 7 FreeSans 80 0 0 0 colon_n[10]
port 149 w signal input
flabel metal1 s 522 6737 575 6751 7 FreeSans 80 0 0 0 colon_n[11]
port 150 w signal input
flabel metal1 s 522 7239 575 7253 7 FreeSans 80 0 0 0 colon_n[12]
port 151 w signal input
flabel metal1 s 522 7741 575 7755 7 FreeSans 80 0 0 0 colon_n[13]
port 152 w signal input
flabel metal1 s 522 8243 575 8257 7 FreeSans 80 0 0 0 colon_n[14]
port 153 w signal input
flabel metal1 s 522 8745 575 8759 7 FreeSans 80 0 0 0 colon_n[15]
port 154 w signal input
flabel metal4 s 0 21 207 12083 0 FreeSans 800 90 0 0 VDD
port 1 nsew power bidirectional
flabel metal4 s 238 21 445 12083 0 FreeSans 800 90 0 0 VSS
port 2 nsew power bidirectional
flabel metal4 s 18827 86 19034 9951 0 FreeSans 800 90 0 0 VSS
port 2 nsew power bidirectional
flabel metal4 s 19065 86 19272 9951 0 FreeSans 800 90 0 0 VDD
port 1 nsew power bidirectional
flabel metal4 s 21386 83 21593 12083 0 FreeSans 800 90 0 0 VDD
port 1 nsew power bidirectional
flabel metal4 s 21630 84 21837 12084 0 FreeSans 800 90 0 0 VSS
port 2 nsew power bidirectional
<< properties >>
string LEFclass CORE
string LEForigin 0 0
string LEFsource USER
<< end >>
